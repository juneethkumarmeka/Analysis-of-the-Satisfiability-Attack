module basic_500_3000_500_3_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_474,In_357);
and U1 (N_1,In_452,In_151);
nor U2 (N_2,In_310,In_197);
nor U3 (N_3,In_392,In_380);
xnor U4 (N_4,In_388,In_248);
xor U5 (N_5,In_98,In_202);
nand U6 (N_6,In_221,In_43);
xnor U7 (N_7,In_1,In_31);
nor U8 (N_8,In_445,In_231);
or U9 (N_9,In_130,In_264);
and U10 (N_10,In_378,In_29);
nand U11 (N_11,In_425,In_210);
xnor U12 (N_12,In_230,In_118);
and U13 (N_13,In_68,In_471);
or U14 (N_14,In_184,In_147);
nor U15 (N_15,In_244,In_363);
xnor U16 (N_16,In_482,In_191);
and U17 (N_17,In_195,In_290);
and U18 (N_18,In_389,In_106);
nor U19 (N_19,In_24,In_259);
xor U20 (N_20,In_490,In_278);
nand U21 (N_21,In_369,In_235);
and U22 (N_22,In_214,In_496);
and U23 (N_23,In_205,In_252);
or U24 (N_24,In_405,In_428);
or U25 (N_25,In_477,In_193);
xnor U26 (N_26,In_125,In_322);
or U27 (N_27,In_261,In_254);
nand U28 (N_28,In_132,In_181);
nor U29 (N_29,In_101,In_343);
or U30 (N_30,In_103,In_3);
or U31 (N_31,In_417,In_71);
or U32 (N_32,In_470,In_263);
or U33 (N_33,In_79,In_422);
xor U34 (N_34,In_274,In_346);
xor U35 (N_35,In_88,In_207);
and U36 (N_36,In_58,In_59);
nand U37 (N_37,In_485,In_134);
and U38 (N_38,In_86,In_149);
or U39 (N_39,In_367,In_267);
nand U40 (N_40,In_273,In_450);
and U41 (N_41,In_298,In_92);
xnor U42 (N_42,In_379,In_321);
nand U43 (N_43,In_69,In_228);
xnor U44 (N_44,In_393,In_413);
xnor U45 (N_45,In_365,In_277);
and U46 (N_46,In_176,In_443);
xnor U47 (N_47,In_352,In_319);
or U48 (N_48,In_497,In_345);
nor U49 (N_49,In_11,In_441);
xor U50 (N_50,In_61,In_240);
and U51 (N_51,In_74,In_476);
nand U52 (N_52,In_136,In_338);
and U53 (N_53,In_382,In_328);
nand U54 (N_54,In_279,In_62);
nor U55 (N_55,In_241,In_87);
and U56 (N_56,In_339,In_177);
nand U57 (N_57,In_289,In_494);
xnor U58 (N_58,In_186,In_459);
or U59 (N_59,In_311,In_187);
nor U60 (N_60,In_131,In_448);
nor U61 (N_61,In_233,In_342);
nor U62 (N_62,In_7,In_15);
xnor U63 (N_63,In_188,In_386);
nand U64 (N_64,In_9,In_46);
nor U65 (N_65,In_190,In_359);
nor U66 (N_66,In_371,In_461);
xor U67 (N_67,In_32,In_94);
nand U68 (N_68,In_66,In_280);
or U69 (N_69,In_312,In_418);
and U70 (N_70,In_8,In_314);
xnor U71 (N_71,In_141,In_407);
xor U72 (N_72,In_291,In_156);
xor U73 (N_73,In_242,In_324);
xnor U74 (N_74,In_377,In_238);
nand U75 (N_75,In_372,In_168);
nor U76 (N_76,In_415,In_18);
nor U77 (N_77,In_96,In_6);
or U78 (N_78,In_286,In_316);
xor U79 (N_79,In_148,In_257);
xor U80 (N_80,In_330,In_292);
or U81 (N_81,In_218,In_410);
nand U82 (N_82,In_198,In_276);
xnor U83 (N_83,In_26,In_137);
or U84 (N_84,In_196,In_424);
and U85 (N_85,In_299,In_281);
and U86 (N_86,In_271,In_348);
or U87 (N_87,In_374,In_127);
and U88 (N_88,In_111,In_262);
or U89 (N_89,In_329,In_206);
and U90 (N_90,In_323,In_126);
nand U91 (N_91,In_394,In_104);
and U92 (N_92,In_473,In_60);
xor U93 (N_93,In_27,In_483);
xor U94 (N_94,In_170,In_282);
nor U95 (N_95,In_347,In_436);
and U96 (N_96,In_128,In_462);
nor U97 (N_97,In_28,In_294);
nor U98 (N_98,In_307,In_385);
nand U99 (N_99,In_57,In_250);
nand U100 (N_100,In_56,In_399);
xnor U101 (N_101,In_301,In_303);
xor U102 (N_102,In_52,In_285);
nor U103 (N_103,In_150,In_437);
or U104 (N_104,In_107,In_256);
and U105 (N_105,In_491,In_460);
and U106 (N_106,In_463,In_90);
nor U107 (N_107,In_295,In_229);
and U108 (N_108,In_199,In_114);
nand U109 (N_109,In_91,In_213);
or U110 (N_110,In_2,In_397);
nand U111 (N_111,In_70,In_383);
or U112 (N_112,In_495,In_110);
nor U113 (N_113,In_78,In_48);
xor U114 (N_114,In_192,In_30);
and U115 (N_115,In_469,In_227);
nand U116 (N_116,In_67,In_159);
and U117 (N_117,In_19,In_161);
nor U118 (N_118,In_270,In_340);
xnor U119 (N_119,In_488,In_75);
and U120 (N_120,In_97,In_376);
xor U121 (N_121,In_166,In_456);
and U122 (N_122,In_284,In_412);
and U123 (N_123,In_430,In_396);
and U124 (N_124,In_366,In_423);
and U125 (N_125,In_245,In_480);
nand U126 (N_126,In_370,In_487);
nand U127 (N_127,In_465,In_403);
nand U128 (N_128,In_454,In_390);
or U129 (N_129,In_287,In_163);
and U130 (N_130,In_255,In_432);
and U131 (N_131,In_85,In_246);
xnor U132 (N_132,In_47,In_302);
or U133 (N_133,In_269,In_53);
or U134 (N_134,In_113,In_236);
and U135 (N_135,In_427,In_162);
or U136 (N_136,In_265,In_171);
or U137 (N_137,In_475,In_16);
nand U138 (N_138,In_309,In_100);
or U139 (N_139,In_344,In_120);
or U140 (N_140,In_395,In_249);
xor U141 (N_141,In_457,In_498);
xnor U142 (N_142,In_55,In_216);
nand U143 (N_143,In_408,In_447);
xor U144 (N_144,In_449,In_375);
nor U145 (N_145,In_440,In_51);
nand U146 (N_146,In_37,In_336);
nor U147 (N_147,In_65,In_121);
xnor U148 (N_148,In_325,In_160);
xor U149 (N_149,In_486,In_76);
or U150 (N_150,In_115,In_173);
xor U151 (N_151,In_93,In_73);
xnor U152 (N_152,In_212,In_154);
xnor U153 (N_153,In_401,In_38);
nand U154 (N_154,In_349,In_489);
nand U155 (N_155,In_182,In_327);
xnor U156 (N_156,In_81,In_466);
or U157 (N_157,In_217,In_350);
nand U158 (N_158,In_315,In_158);
nor U159 (N_159,In_165,In_409);
nand U160 (N_160,In_174,In_384);
nor U161 (N_161,In_124,In_49);
xnor U162 (N_162,In_167,In_80);
nand U163 (N_163,In_119,In_153);
nor U164 (N_164,In_332,In_260);
xor U165 (N_165,In_109,In_4);
or U166 (N_166,In_431,In_398);
or U167 (N_167,In_313,In_41);
nand U168 (N_168,In_499,In_203);
nor U169 (N_169,In_211,In_222);
nor U170 (N_170,In_155,In_36);
xor U171 (N_171,In_435,In_320);
xnor U172 (N_172,In_337,In_308);
nand U173 (N_173,In_142,In_39);
nor U174 (N_174,In_416,In_253);
nor U175 (N_175,In_224,In_183);
and U176 (N_176,In_364,In_306);
xnor U177 (N_177,In_25,In_44);
xnor U178 (N_178,In_391,In_63);
or U179 (N_179,In_362,In_34);
nand U180 (N_180,In_122,In_82);
and U181 (N_181,In_381,In_10);
and U182 (N_182,In_133,In_45);
or U183 (N_183,In_117,In_442);
xnor U184 (N_184,In_402,In_493);
nor U185 (N_185,In_411,In_185);
nor U186 (N_186,In_17,In_135);
nand U187 (N_187,In_84,In_108);
xnor U188 (N_188,In_208,In_50);
or U189 (N_189,In_200,In_464);
nand U190 (N_190,In_180,In_318);
nand U191 (N_191,In_215,In_258);
nor U192 (N_192,In_360,In_334);
xor U193 (N_193,In_144,In_478);
nand U194 (N_194,In_243,In_455);
xnor U195 (N_195,In_426,In_35);
or U196 (N_196,In_351,In_102);
or U197 (N_197,In_237,In_178);
and U198 (N_198,In_420,In_326);
or U199 (N_199,In_5,In_157);
xor U200 (N_200,In_438,In_226);
xor U201 (N_201,In_204,In_22);
and U202 (N_202,In_472,In_232);
and U203 (N_203,In_251,In_77);
xnor U204 (N_204,In_112,In_283);
or U205 (N_205,In_140,In_83);
nand U206 (N_206,In_201,In_54);
nor U207 (N_207,In_164,In_421);
xor U208 (N_208,In_139,In_444);
or U209 (N_209,In_481,In_219);
and U210 (N_210,In_239,In_468);
and U211 (N_211,In_341,In_123);
or U212 (N_212,In_368,In_20);
nor U213 (N_213,In_404,In_247);
or U214 (N_214,In_189,In_304);
or U215 (N_215,In_446,In_143);
nand U216 (N_216,In_116,In_429);
or U217 (N_217,In_297,In_272);
nor U218 (N_218,In_358,In_458);
nand U219 (N_219,In_400,In_172);
nand U220 (N_220,In_89,In_152);
xnor U221 (N_221,In_433,In_266);
nor U222 (N_222,In_317,In_220);
nor U223 (N_223,In_331,In_288);
and U224 (N_224,In_145,In_169);
nor U225 (N_225,In_234,In_296);
and U226 (N_226,In_72,In_387);
or U227 (N_227,In_419,In_439);
nor U228 (N_228,In_138,In_467);
nor U229 (N_229,In_305,In_268);
xnor U230 (N_230,In_225,In_209);
nor U231 (N_231,In_12,In_179);
or U232 (N_232,In_99,In_40);
nor U233 (N_233,In_492,In_175);
and U234 (N_234,In_406,In_21);
or U235 (N_235,In_293,In_33);
nor U236 (N_236,In_105,In_275);
or U237 (N_237,In_354,In_13);
and U238 (N_238,In_95,In_353);
xor U239 (N_239,In_355,In_434);
xnor U240 (N_240,In_335,In_484);
nor U241 (N_241,In_453,In_194);
or U242 (N_242,In_64,In_129);
xnor U243 (N_243,In_23,In_42);
nor U244 (N_244,In_356,In_333);
nor U245 (N_245,In_479,In_0);
nor U246 (N_246,In_373,In_361);
nand U247 (N_247,In_146,In_14);
or U248 (N_248,In_414,In_451);
nor U249 (N_249,In_223,In_300);
or U250 (N_250,In_184,In_482);
nand U251 (N_251,In_154,In_142);
xor U252 (N_252,In_231,In_202);
nand U253 (N_253,In_108,In_254);
xor U254 (N_254,In_444,In_328);
or U255 (N_255,In_450,In_473);
or U256 (N_256,In_275,In_15);
nand U257 (N_257,In_418,In_162);
or U258 (N_258,In_110,In_383);
and U259 (N_259,In_172,In_105);
nand U260 (N_260,In_134,In_210);
and U261 (N_261,In_140,In_21);
and U262 (N_262,In_204,In_334);
nor U263 (N_263,In_391,In_462);
and U264 (N_264,In_116,In_337);
or U265 (N_265,In_321,In_251);
nand U266 (N_266,In_193,In_186);
nor U267 (N_267,In_53,In_183);
nor U268 (N_268,In_22,In_341);
and U269 (N_269,In_210,In_137);
nand U270 (N_270,In_112,In_282);
nand U271 (N_271,In_300,In_25);
nand U272 (N_272,In_286,In_42);
nand U273 (N_273,In_105,In_371);
nand U274 (N_274,In_272,In_453);
or U275 (N_275,In_105,In_490);
or U276 (N_276,In_66,In_9);
and U277 (N_277,In_74,In_136);
or U278 (N_278,In_300,In_0);
nor U279 (N_279,In_362,In_214);
nand U280 (N_280,In_170,In_301);
and U281 (N_281,In_380,In_14);
and U282 (N_282,In_0,In_6);
nand U283 (N_283,In_103,In_394);
nand U284 (N_284,In_19,In_354);
nand U285 (N_285,In_282,In_305);
nor U286 (N_286,In_105,In_404);
or U287 (N_287,In_296,In_363);
xor U288 (N_288,In_99,In_190);
or U289 (N_289,In_86,In_167);
or U290 (N_290,In_197,In_421);
and U291 (N_291,In_280,In_468);
nand U292 (N_292,In_216,In_219);
nor U293 (N_293,In_460,In_255);
nand U294 (N_294,In_150,In_357);
nand U295 (N_295,In_71,In_27);
or U296 (N_296,In_327,In_274);
xor U297 (N_297,In_388,In_109);
or U298 (N_298,In_148,In_132);
nor U299 (N_299,In_48,In_412);
nor U300 (N_300,In_194,In_32);
and U301 (N_301,In_151,In_31);
nor U302 (N_302,In_247,In_356);
xnor U303 (N_303,In_234,In_92);
nor U304 (N_304,In_118,In_226);
xnor U305 (N_305,In_471,In_216);
and U306 (N_306,In_150,In_44);
or U307 (N_307,In_308,In_477);
and U308 (N_308,In_106,In_402);
or U309 (N_309,In_185,In_404);
xnor U310 (N_310,In_365,In_497);
nand U311 (N_311,In_21,In_86);
or U312 (N_312,In_363,In_412);
xor U313 (N_313,In_320,In_59);
xor U314 (N_314,In_319,In_385);
and U315 (N_315,In_214,In_145);
and U316 (N_316,In_116,In_425);
or U317 (N_317,In_97,In_34);
nand U318 (N_318,In_490,In_62);
xor U319 (N_319,In_397,In_361);
or U320 (N_320,In_106,In_243);
nand U321 (N_321,In_281,In_441);
and U322 (N_322,In_29,In_461);
nor U323 (N_323,In_91,In_469);
and U324 (N_324,In_203,In_108);
xnor U325 (N_325,In_175,In_222);
nand U326 (N_326,In_320,In_3);
or U327 (N_327,In_479,In_70);
or U328 (N_328,In_492,In_22);
nand U329 (N_329,In_192,In_208);
nand U330 (N_330,In_51,In_35);
nand U331 (N_331,In_455,In_326);
xor U332 (N_332,In_379,In_360);
nor U333 (N_333,In_50,In_229);
and U334 (N_334,In_359,In_177);
nand U335 (N_335,In_348,In_103);
nand U336 (N_336,In_440,In_307);
and U337 (N_337,In_27,In_160);
nand U338 (N_338,In_121,In_393);
nor U339 (N_339,In_481,In_305);
or U340 (N_340,In_401,In_334);
nand U341 (N_341,In_375,In_2);
xnor U342 (N_342,In_228,In_60);
and U343 (N_343,In_30,In_113);
nand U344 (N_344,In_223,In_266);
xor U345 (N_345,In_50,In_29);
and U346 (N_346,In_371,In_493);
or U347 (N_347,In_109,In_444);
or U348 (N_348,In_103,In_14);
or U349 (N_349,In_209,In_116);
nor U350 (N_350,In_379,In_346);
or U351 (N_351,In_349,In_149);
and U352 (N_352,In_144,In_425);
nor U353 (N_353,In_79,In_105);
xnor U354 (N_354,In_396,In_189);
or U355 (N_355,In_310,In_249);
nand U356 (N_356,In_381,In_384);
nor U357 (N_357,In_493,In_487);
or U358 (N_358,In_157,In_170);
xnor U359 (N_359,In_326,In_453);
nor U360 (N_360,In_62,In_263);
nand U361 (N_361,In_470,In_443);
and U362 (N_362,In_171,In_481);
nor U363 (N_363,In_337,In_100);
and U364 (N_364,In_150,In_424);
and U365 (N_365,In_349,In_377);
or U366 (N_366,In_238,In_460);
xnor U367 (N_367,In_447,In_434);
xor U368 (N_368,In_118,In_445);
xnor U369 (N_369,In_250,In_187);
and U370 (N_370,In_423,In_244);
nor U371 (N_371,In_270,In_19);
nand U372 (N_372,In_294,In_489);
and U373 (N_373,In_319,In_235);
xnor U374 (N_374,In_487,In_26);
nor U375 (N_375,In_193,In_397);
nand U376 (N_376,In_16,In_315);
nand U377 (N_377,In_34,In_329);
xor U378 (N_378,In_45,In_348);
nor U379 (N_379,In_248,In_422);
nand U380 (N_380,In_328,In_156);
xnor U381 (N_381,In_240,In_221);
nand U382 (N_382,In_392,In_8);
nand U383 (N_383,In_467,In_227);
nand U384 (N_384,In_136,In_346);
or U385 (N_385,In_229,In_38);
nand U386 (N_386,In_195,In_137);
nand U387 (N_387,In_445,In_455);
and U388 (N_388,In_84,In_126);
nand U389 (N_389,In_19,In_91);
nand U390 (N_390,In_447,In_61);
nor U391 (N_391,In_167,In_289);
or U392 (N_392,In_244,In_255);
and U393 (N_393,In_127,In_143);
and U394 (N_394,In_411,In_202);
nor U395 (N_395,In_415,In_234);
xor U396 (N_396,In_71,In_491);
nand U397 (N_397,In_235,In_164);
nand U398 (N_398,In_234,In_492);
or U399 (N_399,In_321,In_23);
nand U400 (N_400,In_441,In_398);
xnor U401 (N_401,In_177,In_489);
nor U402 (N_402,In_357,In_77);
and U403 (N_403,In_418,In_241);
nor U404 (N_404,In_193,In_496);
nor U405 (N_405,In_428,In_252);
xor U406 (N_406,In_224,In_302);
and U407 (N_407,In_327,In_464);
xor U408 (N_408,In_66,In_162);
or U409 (N_409,In_455,In_371);
xnor U410 (N_410,In_310,In_287);
nand U411 (N_411,In_407,In_408);
or U412 (N_412,In_129,In_173);
nor U413 (N_413,In_18,In_406);
xnor U414 (N_414,In_289,In_468);
xnor U415 (N_415,In_0,In_195);
nand U416 (N_416,In_469,In_115);
and U417 (N_417,In_84,In_282);
nand U418 (N_418,In_462,In_275);
or U419 (N_419,In_207,In_336);
and U420 (N_420,In_344,In_420);
nand U421 (N_421,In_426,In_149);
and U422 (N_422,In_237,In_462);
nand U423 (N_423,In_401,In_383);
and U424 (N_424,In_481,In_264);
and U425 (N_425,In_447,In_142);
xor U426 (N_426,In_88,In_335);
or U427 (N_427,In_66,In_33);
or U428 (N_428,In_342,In_53);
or U429 (N_429,In_314,In_255);
and U430 (N_430,In_353,In_50);
and U431 (N_431,In_15,In_218);
nor U432 (N_432,In_460,In_49);
xor U433 (N_433,In_311,In_341);
or U434 (N_434,In_453,In_118);
or U435 (N_435,In_325,In_405);
nand U436 (N_436,In_329,In_108);
nand U437 (N_437,In_281,In_258);
nor U438 (N_438,In_54,In_155);
or U439 (N_439,In_493,In_252);
nor U440 (N_440,In_196,In_256);
and U441 (N_441,In_0,In_430);
nand U442 (N_442,In_486,In_232);
nor U443 (N_443,In_302,In_42);
nor U444 (N_444,In_27,In_462);
and U445 (N_445,In_215,In_333);
or U446 (N_446,In_40,In_319);
xnor U447 (N_447,In_112,In_26);
xor U448 (N_448,In_58,In_457);
nand U449 (N_449,In_135,In_247);
and U450 (N_450,In_359,In_114);
nand U451 (N_451,In_228,In_315);
and U452 (N_452,In_71,In_313);
nor U453 (N_453,In_363,In_82);
nand U454 (N_454,In_262,In_91);
nor U455 (N_455,In_148,In_331);
xnor U456 (N_456,In_490,In_203);
and U457 (N_457,In_308,In_247);
or U458 (N_458,In_456,In_479);
and U459 (N_459,In_212,In_204);
nor U460 (N_460,In_128,In_351);
nand U461 (N_461,In_458,In_154);
xor U462 (N_462,In_231,In_110);
nor U463 (N_463,In_343,In_427);
xor U464 (N_464,In_442,In_438);
or U465 (N_465,In_269,In_419);
and U466 (N_466,In_499,In_411);
xnor U467 (N_467,In_301,In_229);
and U468 (N_468,In_351,In_265);
nand U469 (N_469,In_254,In_481);
nand U470 (N_470,In_141,In_209);
nand U471 (N_471,In_20,In_416);
and U472 (N_472,In_43,In_423);
or U473 (N_473,In_355,In_81);
nand U474 (N_474,In_218,In_105);
xor U475 (N_475,In_477,In_49);
nor U476 (N_476,In_130,In_487);
xnor U477 (N_477,In_401,In_129);
nor U478 (N_478,In_326,In_306);
nor U479 (N_479,In_115,In_151);
nand U480 (N_480,In_149,In_376);
xor U481 (N_481,In_359,In_492);
or U482 (N_482,In_354,In_186);
and U483 (N_483,In_59,In_256);
nor U484 (N_484,In_24,In_57);
nand U485 (N_485,In_76,In_299);
nand U486 (N_486,In_27,In_350);
and U487 (N_487,In_238,In_83);
or U488 (N_488,In_384,In_366);
or U489 (N_489,In_117,In_307);
nor U490 (N_490,In_390,In_401);
or U491 (N_491,In_247,In_160);
or U492 (N_492,In_67,In_466);
or U493 (N_493,In_352,In_71);
and U494 (N_494,In_403,In_324);
or U495 (N_495,In_187,In_288);
xnor U496 (N_496,In_492,In_283);
nor U497 (N_497,In_132,In_326);
and U498 (N_498,In_437,In_424);
and U499 (N_499,In_491,In_193);
nor U500 (N_500,In_296,In_431);
nor U501 (N_501,In_261,In_485);
or U502 (N_502,In_3,In_458);
nand U503 (N_503,In_191,In_230);
and U504 (N_504,In_114,In_338);
nand U505 (N_505,In_234,In_147);
nand U506 (N_506,In_161,In_236);
nand U507 (N_507,In_151,In_328);
and U508 (N_508,In_85,In_33);
nor U509 (N_509,In_469,In_73);
and U510 (N_510,In_4,In_147);
xnor U511 (N_511,In_412,In_123);
nand U512 (N_512,In_230,In_256);
and U513 (N_513,In_398,In_380);
xnor U514 (N_514,In_367,In_379);
and U515 (N_515,In_153,In_427);
nand U516 (N_516,In_198,In_323);
and U517 (N_517,In_305,In_224);
and U518 (N_518,In_330,In_293);
or U519 (N_519,In_155,In_288);
and U520 (N_520,In_67,In_365);
xor U521 (N_521,In_179,In_167);
or U522 (N_522,In_414,In_289);
xnor U523 (N_523,In_87,In_78);
nand U524 (N_524,In_265,In_266);
xor U525 (N_525,In_122,In_115);
or U526 (N_526,In_139,In_312);
or U527 (N_527,In_307,In_180);
or U528 (N_528,In_14,In_396);
nor U529 (N_529,In_288,In_453);
or U530 (N_530,In_7,In_335);
nand U531 (N_531,In_466,In_285);
and U532 (N_532,In_389,In_21);
and U533 (N_533,In_50,In_184);
xnor U534 (N_534,In_303,In_287);
or U535 (N_535,In_338,In_395);
nand U536 (N_536,In_139,In_174);
nor U537 (N_537,In_447,In_150);
nor U538 (N_538,In_344,In_201);
nand U539 (N_539,In_462,In_72);
nand U540 (N_540,In_343,In_460);
nand U541 (N_541,In_166,In_358);
nor U542 (N_542,In_301,In_68);
nor U543 (N_543,In_491,In_115);
or U544 (N_544,In_229,In_387);
nor U545 (N_545,In_382,In_403);
and U546 (N_546,In_7,In_338);
or U547 (N_547,In_399,In_227);
nand U548 (N_548,In_334,In_18);
nor U549 (N_549,In_303,In_355);
or U550 (N_550,In_14,In_46);
xor U551 (N_551,In_431,In_230);
or U552 (N_552,In_136,In_12);
xor U553 (N_553,In_310,In_489);
xnor U554 (N_554,In_0,In_97);
nor U555 (N_555,In_443,In_179);
and U556 (N_556,In_445,In_39);
or U557 (N_557,In_321,In_56);
xnor U558 (N_558,In_245,In_268);
nor U559 (N_559,In_60,In_226);
or U560 (N_560,In_124,In_198);
nand U561 (N_561,In_365,In_442);
or U562 (N_562,In_158,In_81);
nor U563 (N_563,In_167,In_186);
xor U564 (N_564,In_0,In_7);
or U565 (N_565,In_15,In_170);
nand U566 (N_566,In_24,In_417);
xnor U567 (N_567,In_272,In_2);
and U568 (N_568,In_52,In_451);
nor U569 (N_569,In_289,In_51);
xor U570 (N_570,In_64,In_372);
nand U571 (N_571,In_106,In_135);
and U572 (N_572,In_279,In_43);
nand U573 (N_573,In_497,In_417);
xor U574 (N_574,In_108,In_81);
nor U575 (N_575,In_13,In_415);
and U576 (N_576,In_130,In_118);
nor U577 (N_577,In_310,In_399);
or U578 (N_578,In_371,In_116);
nor U579 (N_579,In_355,In_271);
or U580 (N_580,In_484,In_175);
nor U581 (N_581,In_394,In_115);
and U582 (N_582,In_38,In_134);
nor U583 (N_583,In_226,In_94);
or U584 (N_584,In_145,In_107);
nand U585 (N_585,In_156,In_425);
nand U586 (N_586,In_33,In_52);
nand U587 (N_587,In_241,In_177);
and U588 (N_588,In_247,In_459);
xnor U589 (N_589,In_498,In_308);
nor U590 (N_590,In_265,In_381);
or U591 (N_591,In_229,In_257);
or U592 (N_592,In_35,In_346);
and U593 (N_593,In_30,In_288);
nand U594 (N_594,In_372,In_292);
xnor U595 (N_595,In_132,In_65);
nand U596 (N_596,In_274,In_99);
nand U597 (N_597,In_389,In_231);
or U598 (N_598,In_415,In_291);
nand U599 (N_599,In_171,In_21);
nand U600 (N_600,In_341,In_223);
nor U601 (N_601,In_180,In_371);
nand U602 (N_602,In_17,In_380);
and U603 (N_603,In_16,In_286);
and U604 (N_604,In_426,In_258);
nand U605 (N_605,In_41,In_318);
and U606 (N_606,In_347,In_351);
xor U607 (N_607,In_230,In_490);
xnor U608 (N_608,In_96,In_401);
xnor U609 (N_609,In_107,In_243);
nor U610 (N_610,In_29,In_293);
nand U611 (N_611,In_192,In_411);
xnor U612 (N_612,In_118,In_229);
nor U613 (N_613,In_384,In_413);
and U614 (N_614,In_21,In_189);
nand U615 (N_615,In_481,In_112);
and U616 (N_616,In_261,In_392);
or U617 (N_617,In_434,In_348);
and U618 (N_618,In_14,In_312);
or U619 (N_619,In_310,In_106);
and U620 (N_620,In_140,In_439);
or U621 (N_621,In_230,In_254);
nor U622 (N_622,In_413,In_15);
xnor U623 (N_623,In_339,In_42);
and U624 (N_624,In_89,In_225);
and U625 (N_625,In_474,In_483);
nor U626 (N_626,In_240,In_470);
nand U627 (N_627,In_18,In_132);
and U628 (N_628,In_140,In_218);
xnor U629 (N_629,In_140,In_166);
and U630 (N_630,In_461,In_493);
or U631 (N_631,In_110,In_59);
nor U632 (N_632,In_128,In_66);
and U633 (N_633,In_201,In_3);
xor U634 (N_634,In_469,In_289);
nand U635 (N_635,In_30,In_195);
xnor U636 (N_636,In_334,In_125);
nor U637 (N_637,In_200,In_398);
and U638 (N_638,In_463,In_356);
nor U639 (N_639,In_290,In_481);
xnor U640 (N_640,In_100,In_111);
xor U641 (N_641,In_23,In_202);
nand U642 (N_642,In_266,In_399);
xnor U643 (N_643,In_131,In_372);
nand U644 (N_644,In_488,In_405);
and U645 (N_645,In_405,In_370);
nand U646 (N_646,In_61,In_341);
nor U647 (N_647,In_474,In_187);
or U648 (N_648,In_222,In_391);
xor U649 (N_649,In_60,In_195);
or U650 (N_650,In_399,In_410);
xnor U651 (N_651,In_228,In_316);
and U652 (N_652,In_405,In_102);
nor U653 (N_653,In_240,In_38);
and U654 (N_654,In_445,In_203);
nand U655 (N_655,In_411,In_214);
xor U656 (N_656,In_498,In_426);
and U657 (N_657,In_162,In_455);
nor U658 (N_658,In_27,In_492);
nand U659 (N_659,In_394,In_397);
nor U660 (N_660,In_390,In_403);
nor U661 (N_661,In_322,In_263);
nor U662 (N_662,In_33,In_332);
and U663 (N_663,In_122,In_35);
or U664 (N_664,In_211,In_139);
nand U665 (N_665,In_129,In_415);
nand U666 (N_666,In_393,In_180);
nor U667 (N_667,In_222,In_313);
and U668 (N_668,In_97,In_28);
nand U669 (N_669,In_336,In_354);
nor U670 (N_670,In_412,In_433);
and U671 (N_671,In_124,In_105);
xnor U672 (N_672,In_372,In_407);
and U673 (N_673,In_336,In_27);
nor U674 (N_674,In_232,In_46);
and U675 (N_675,In_39,In_456);
nor U676 (N_676,In_330,In_235);
nand U677 (N_677,In_230,In_49);
nor U678 (N_678,In_94,In_17);
nand U679 (N_679,In_298,In_71);
nor U680 (N_680,In_78,In_137);
nand U681 (N_681,In_285,In_485);
nand U682 (N_682,In_337,In_140);
or U683 (N_683,In_249,In_142);
and U684 (N_684,In_216,In_22);
or U685 (N_685,In_27,In_56);
and U686 (N_686,In_261,In_462);
or U687 (N_687,In_349,In_485);
and U688 (N_688,In_169,In_422);
nor U689 (N_689,In_82,In_315);
or U690 (N_690,In_466,In_107);
nor U691 (N_691,In_465,In_205);
xnor U692 (N_692,In_192,In_107);
and U693 (N_693,In_177,In_398);
nor U694 (N_694,In_283,In_52);
xnor U695 (N_695,In_416,In_395);
nor U696 (N_696,In_477,In_346);
xor U697 (N_697,In_179,In_124);
nand U698 (N_698,In_186,In_267);
or U699 (N_699,In_272,In_474);
nand U700 (N_700,In_210,In_126);
xor U701 (N_701,In_192,In_217);
nand U702 (N_702,In_307,In_233);
xor U703 (N_703,In_383,In_78);
or U704 (N_704,In_383,In_261);
and U705 (N_705,In_419,In_354);
nand U706 (N_706,In_498,In_26);
or U707 (N_707,In_297,In_281);
and U708 (N_708,In_369,In_120);
nand U709 (N_709,In_255,In_419);
and U710 (N_710,In_374,In_299);
nor U711 (N_711,In_484,In_248);
xor U712 (N_712,In_254,In_363);
nand U713 (N_713,In_259,In_65);
xnor U714 (N_714,In_98,In_224);
nand U715 (N_715,In_158,In_290);
and U716 (N_716,In_433,In_109);
nand U717 (N_717,In_431,In_175);
nand U718 (N_718,In_389,In_432);
nand U719 (N_719,In_497,In_485);
xnor U720 (N_720,In_435,In_53);
nand U721 (N_721,In_291,In_69);
and U722 (N_722,In_131,In_241);
xor U723 (N_723,In_331,In_421);
xor U724 (N_724,In_272,In_361);
nor U725 (N_725,In_264,In_406);
or U726 (N_726,In_486,In_44);
nand U727 (N_727,In_397,In_313);
or U728 (N_728,In_390,In_423);
nor U729 (N_729,In_278,In_399);
xnor U730 (N_730,In_360,In_169);
xor U731 (N_731,In_365,In_297);
and U732 (N_732,In_43,In_482);
or U733 (N_733,In_27,In_213);
nand U734 (N_734,In_142,In_153);
nor U735 (N_735,In_305,In_419);
and U736 (N_736,In_100,In_248);
and U737 (N_737,In_301,In_6);
or U738 (N_738,In_72,In_335);
xor U739 (N_739,In_269,In_56);
or U740 (N_740,In_153,In_185);
nor U741 (N_741,In_395,In_104);
xnor U742 (N_742,In_225,In_46);
xnor U743 (N_743,In_147,In_401);
nand U744 (N_744,In_323,In_122);
xnor U745 (N_745,In_370,In_448);
xor U746 (N_746,In_40,In_5);
and U747 (N_747,In_348,In_91);
nor U748 (N_748,In_407,In_186);
nor U749 (N_749,In_475,In_5);
or U750 (N_750,In_19,In_96);
nor U751 (N_751,In_7,In_190);
nor U752 (N_752,In_50,In_472);
and U753 (N_753,In_198,In_34);
and U754 (N_754,In_277,In_243);
nor U755 (N_755,In_364,In_276);
or U756 (N_756,In_18,In_150);
nor U757 (N_757,In_220,In_74);
xor U758 (N_758,In_302,In_102);
nor U759 (N_759,In_363,In_253);
xnor U760 (N_760,In_343,In_285);
nor U761 (N_761,In_272,In_382);
nand U762 (N_762,In_364,In_482);
xnor U763 (N_763,In_81,In_403);
and U764 (N_764,In_320,In_298);
nand U765 (N_765,In_347,In_154);
and U766 (N_766,In_490,In_232);
xnor U767 (N_767,In_185,In_302);
nand U768 (N_768,In_341,In_403);
and U769 (N_769,In_137,In_312);
or U770 (N_770,In_201,In_422);
nor U771 (N_771,In_49,In_22);
xnor U772 (N_772,In_183,In_24);
or U773 (N_773,In_230,In_28);
nor U774 (N_774,In_193,In_471);
nor U775 (N_775,In_370,In_275);
nor U776 (N_776,In_457,In_436);
nand U777 (N_777,In_86,In_171);
nor U778 (N_778,In_285,In_298);
or U779 (N_779,In_118,In_63);
and U780 (N_780,In_34,In_255);
xor U781 (N_781,In_252,In_256);
nand U782 (N_782,In_88,In_489);
xnor U783 (N_783,In_6,In_127);
and U784 (N_784,In_133,In_467);
nor U785 (N_785,In_55,In_228);
nand U786 (N_786,In_417,In_169);
nor U787 (N_787,In_424,In_65);
and U788 (N_788,In_154,In_19);
and U789 (N_789,In_4,In_227);
nor U790 (N_790,In_58,In_96);
nand U791 (N_791,In_10,In_11);
or U792 (N_792,In_233,In_356);
nand U793 (N_793,In_234,In_399);
xnor U794 (N_794,In_195,In_352);
nor U795 (N_795,In_379,In_218);
nand U796 (N_796,In_263,In_16);
and U797 (N_797,In_17,In_483);
or U798 (N_798,In_318,In_390);
nand U799 (N_799,In_233,In_408);
nand U800 (N_800,In_485,In_113);
nor U801 (N_801,In_474,In_254);
and U802 (N_802,In_432,In_263);
nor U803 (N_803,In_462,In_243);
and U804 (N_804,In_315,In_166);
and U805 (N_805,In_404,In_8);
nand U806 (N_806,In_243,In_411);
nor U807 (N_807,In_466,In_233);
and U808 (N_808,In_150,In_52);
or U809 (N_809,In_346,In_397);
nand U810 (N_810,In_294,In_491);
and U811 (N_811,In_50,In_198);
and U812 (N_812,In_314,In_341);
or U813 (N_813,In_109,In_473);
xor U814 (N_814,In_199,In_463);
and U815 (N_815,In_203,In_50);
or U816 (N_816,In_345,In_433);
or U817 (N_817,In_95,In_55);
xnor U818 (N_818,In_355,In_298);
xor U819 (N_819,In_187,In_55);
or U820 (N_820,In_2,In_419);
and U821 (N_821,In_264,In_376);
or U822 (N_822,In_361,In_283);
xnor U823 (N_823,In_184,In_356);
or U824 (N_824,In_23,In_71);
xor U825 (N_825,In_177,In_243);
and U826 (N_826,In_307,In_174);
nor U827 (N_827,In_162,In_374);
xor U828 (N_828,In_148,In_150);
nand U829 (N_829,In_284,In_293);
xnor U830 (N_830,In_428,In_452);
nand U831 (N_831,In_90,In_238);
nand U832 (N_832,In_463,In_146);
or U833 (N_833,In_24,In_325);
nor U834 (N_834,In_427,In_430);
nor U835 (N_835,In_127,In_14);
xor U836 (N_836,In_143,In_168);
nand U837 (N_837,In_415,In_191);
or U838 (N_838,In_149,In_363);
or U839 (N_839,In_72,In_385);
xor U840 (N_840,In_326,In_330);
xor U841 (N_841,In_54,In_178);
nand U842 (N_842,In_352,In_404);
nor U843 (N_843,In_346,In_467);
nor U844 (N_844,In_146,In_311);
or U845 (N_845,In_157,In_299);
xor U846 (N_846,In_357,In_65);
nand U847 (N_847,In_291,In_73);
nand U848 (N_848,In_233,In_411);
xnor U849 (N_849,In_381,In_18);
or U850 (N_850,In_95,In_57);
xnor U851 (N_851,In_325,In_224);
nand U852 (N_852,In_354,In_450);
xor U853 (N_853,In_338,In_349);
or U854 (N_854,In_53,In_433);
nand U855 (N_855,In_201,In_25);
nand U856 (N_856,In_30,In_286);
nor U857 (N_857,In_315,In_156);
and U858 (N_858,In_430,In_234);
and U859 (N_859,In_107,In_379);
nand U860 (N_860,In_339,In_345);
xnor U861 (N_861,In_259,In_309);
and U862 (N_862,In_192,In_237);
nand U863 (N_863,In_100,In_204);
xnor U864 (N_864,In_418,In_240);
nand U865 (N_865,In_198,In_176);
and U866 (N_866,In_384,In_61);
nand U867 (N_867,In_395,In_478);
xor U868 (N_868,In_355,In_407);
nand U869 (N_869,In_2,In_333);
and U870 (N_870,In_54,In_151);
and U871 (N_871,In_471,In_305);
and U872 (N_872,In_311,In_174);
nor U873 (N_873,In_157,In_46);
or U874 (N_874,In_493,In_394);
and U875 (N_875,In_257,In_454);
nor U876 (N_876,In_497,In_257);
xor U877 (N_877,In_361,In_72);
nand U878 (N_878,In_214,In_281);
nor U879 (N_879,In_241,In_469);
nand U880 (N_880,In_391,In_343);
xor U881 (N_881,In_5,In_221);
and U882 (N_882,In_303,In_74);
or U883 (N_883,In_487,In_469);
or U884 (N_884,In_109,In_456);
nand U885 (N_885,In_141,In_192);
nor U886 (N_886,In_410,In_302);
or U887 (N_887,In_42,In_418);
or U888 (N_888,In_69,In_423);
and U889 (N_889,In_87,In_474);
nor U890 (N_890,In_69,In_232);
or U891 (N_891,In_138,In_461);
or U892 (N_892,In_345,In_86);
nor U893 (N_893,In_95,In_320);
nor U894 (N_894,In_228,In_492);
nand U895 (N_895,In_352,In_156);
and U896 (N_896,In_364,In_63);
and U897 (N_897,In_38,In_458);
nor U898 (N_898,In_241,In_45);
and U899 (N_899,In_313,In_307);
or U900 (N_900,In_222,In_280);
nand U901 (N_901,In_488,In_103);
and U902 (N_902,In_422,In_272);
xnor U903 (N_903,In_262,In_378);
nor U904 (N_904,In_293,In_471);
or U905 (N_905,In_197,In_493);
and U906 (N_906,In_190,In_124);
xor U907 (N_907,In_72,In_132);
or U908 (N_908,In_90,In_227);
or U909 (N_909,In_190,In_305);
or U910 (N_910,In_282,In_369);
nor U911 (N_911,In_373,In_95);
xnor U912 (N_912,In_464,In_398);
nand U913 (N_913,In_203,In_96);
or U914 (N_914,In_405,In_313);
and U915 (N_915,In_23,In_453);
and U916 (N_916,In_11,In_195);
and U917 (N_917,In_149,In_145);
and U918 (N_918,In_486,In_420);
and U919 (N_919,In_232,In_384);
or U920 (N_920,In_187,In_425);
or U921 (N_921,In_343,In_90);
or U922 (N_922,In_492,In_372);
nand U923 (N_923,In_102,In_200);
xnor U924 (N_924,In_286,In_360);
nand U925 (N_925,In_330,In_238);
xor U926 (N_926,In_170,In_478);
and U927 (N_927,In_66,In_24);
or U928 (N_928,In_198,In_110);
nand U929 (N_929,In_308,In_211);
nor U930 (N_930,In_138,In_253);
xnor U931 (N_931,In_381,In_178);
or U932 (N_932,In_133,In_124);
and U933 (N_933,In_357,In_61);
nand U934 (N_934,In_442,In_338);
nor U935 (N_935,In_8,In_67);
xor U936 (N_936,In_397,In_202);
nor U937 (N_937,In_397,In_485);
nor U938 (N_938,In_177,In_47);
and U939 (N_939,In_311,In_264);
nor U940 (N_940,In_353,In_362);
xnor U941 (N_941,In_297,In_318);
and U942 (N_942,In_100,In_378);
nor U943 (N_943,In_261,In_332);
xor U944 (N_944,In_290,In_225);
nand U945 (N_945,In_181,In_13);
xor U946 (N_946,In_469,In_280);
xnor U947 (N_947,In_261,In_88);
nor U948 (N_948,In_38,In_440);
or U949 (N_949,In_382,In_208);
nand U950 (N_950,In_494,In_284);
or U951 (N_951,In_172,In_345);
nand U952 (N_952,In_204,In_110);
nand U953 (N_953,In_354,In_6);
nor U954 (N_954,In_320,In_381);
nand U955 (N_955,In_132,In_294);
nand U956 (N_956,In_30,In_145);
xnor U957 (N_957,In_294,In_146);
and U958 (N_958,In_106,In_79);
xor U959 (N_959,In_46,In_422);
nand U960 (N_960,In_185,In_128);
nand U961 (N_961,In_181,In_58);
nor U962 (N_962,In_266,In_13);
or U963 (N_963,In_206,In_434);
xnor U964 (N_964,In_479,In_31);
nor U965 (N_965,In_13,In_20);
and U966 (N_966,In_1,In_132);
or U967 (N_967,In_183,In_124);
xor U968 (N_968,In_366,In_57);
and U969 (N_969,In_119,In_234);
nand U970 (N_970,In_211,In_34);
or U971 (N_971,In_13,In_121);
or U972 (N_972,In_471,In_218);
or U973 (N_973,In_96,In_229);
xnor U974 (N_974,In_188,In_142);
nand U975 (N_975,In_208,In_360);
or U976 (N_976,In_389,In_140);
nand U977 (N_977,In_92,In_286);
or U978 (N_978,In_341,In_161);
and U979 (N_979,In_40,In_324);
nand U980 (N_980,In_100,In_51);
xor U981 (N_981,In_55,In_89);
nor U982 (N_982,In_105,In_459);
nor U983 (N_983,In_104,In_216);
and U984 (N_984,In_314,In_15);
or U985 (N_985,In_48,In_368);
and U986 (N_986,In_412,In_120);
and U987 (N_987,In_316,In_468);
or U988 (N_988,In_449,In_335);
and U989 (N_989,In_432,In_32);
and U990 (N_990,In_393,In_38);
or U991 (N_991,In_153,In_422);
xnor U992 (N_992,In_190,In_301);
nor U993 (N_993,In_229,In_307);
xor U994 (N_994,In_343,In_303);
and U995 (N_995,In_296,In_171);
nor U996 (N_996,In_228,In_374);
xor U997 (N_997,In_360,In_195);
nor U998 (N_998,In_159,In_439);
and U999 (N_999,In_256,In_62);
nand U1000 (N_1000,N_691,N_955);
nor U1001 (N_1001,N_522,N_899);
nand U1002 (N_1002,N_352,N_905);
nand U1003 (N_1003,N_976,N_279);
nand U1004 (N_1004,N_659,N_934);
xnor U1005 (N_1005,N_668,N_344);
xnor U1006 (N_1006,N_540,N_918);
and U1007 (N_1007,N_386,N_680);
nand U1008 (N_1008,N_846,N_779);
nand U1009 (N_1009,N_327,N_852);
xor U1010 (N_1010,N_463,N_994);
or U1011 (N_1011,N_656,N_325);
or U1012 (N_1012,N_458,N_376);
or U1013 (N_1013,N_818,N_618);
and U1014 (N_1014,N_840,N_699);
xor U1015 (N_1015,N_917,N_484);
nand U1016 (N_1016,N_22,N_52);
or U1017 (N_1017,N_152,N_929);
nor U1018 (N_1018,N_294,N_998);
xnor U1019 (N_1019,N_438,N_639);
or U1020 (N_1020,N_729,N_483);
or U1021 (N_1021,N_206,N_742);
or U1022 (N_1022,N_837,N_684);
nor U1023 (N_1023,N_941,N_339);
xnor U1024 (N_1024,N_577,N_855);
and U1025 (N_1025,N_243,N_209);
and U1026 (N_1026,N_222,N_317);
and U1027 (N_1027,N_628,N_395);
or U1028 (N_1028,N_488,N_663);
or U1029 (N_1029,N_687,N_696);
nor U1030 (N_1030,N_58,N_298);
and U1031 (N_1031,N_417,N_419);
and U1032 (N_1032,N_297,N_290);
nand U1033 (N_1033,N_17,N_482);
xnor U1034 (N_1034,N_246,N_521);
xnor U1035 (N_1035,N_567,N_160);
nor U1036 (N_1036,N_553,N_295);
or U1037 (N_1037,N_153,N_786);
or U1038 (N_1038,N_373,N_812);
and U1039 (N_1039,N_235,N_194);
nor U1040 (N_1040,N_452,N_219);
or U1041 (N_1041,N_996,N_375);
nor U1042 (N_1042,N_861,N_203);
nand U1043 (N_1043,N_774,N_108);
xor U1044 (N_1044,N_581,N_563);
and U1045 (N_1045,N_435,N_45);
xor U1046 (N_1046,N_823,N_928);
nand U1047 (N_1047,N_971,N_888);
or U1048 (N_1048,N_670,N_42);
and U1049 (N_1049,N_806,N_586);
xnor U1050 (N_1050,N_371,N_20);
nor U1051 (N_1051,N_636,N_314);
and U1052 (N_1052,N_308,N_346);
nor U1053 (N_1053,N_141,N_7);
or U1054 (N_1054,N_236,N_651);
or U1055 (N_1055,N_804,N_936);
nand U1056 (N_1056,N_606,N_394);
xnor U1057 (N_1057,N_296,N_448);
nor U1058 (N_1058,N_843,N_5);
or U1059 (N_1059,N_410,N_772);
xnor U1060 (N_1060,N_103,N_213);
nand U1061 (N_1061,N_493,N_72);
and U1062 (N_1062,N_437,N_131);
and U1063 (N_1063,N_377,N_661);
and U1064 (N_1064,N_690,N_873);
nand U1065 (N_1065,N_220,N_902);
nand U1066 (N_1066,N_358,N_145);
nand U1067 (N_1067,N_285,N_24);
nand U1068 (N_1068,N_359,N_198);
and U1069 (N_1069,N_393,N_867);
nand U1070 (N_1070,N_286,N_939);
and U1071 (N_1071,N_431,N_723);
xor U1072 (N_1072,N_333,N_367);
or U1073 (N_1073,N_480,N_190);
and U1074 (N_1074,N_554,N_953);
nand U1075 (N_1075,N_626,N_890);
or U1076 (N_1076,N_43,N_114);
or U1077 (N_1077,N_60,N_519);
and U1078 (N_1078,N_37,N_865);
nor U1079 (N_1079,N_75,N_430);
xor U1080 (N_1080,N_698,N_368);
nand U1081 (N_1081,N_106,N_912);
and U1082 (N_1082,N_854,N_291);
nor U1083 (N_1083,N_559,N_65);
nand U1084 (N_1084,N_311,N_501);
nand U1085 (N_1085,N_151,N_543);
xnor U1086 (N_1086,N_113,N_514);
xnor U1087 (N_1087,N_879,N_859);
or U1088 (N_1088,N_566,N_172);
and U1089 (N_1089,N_218,N_138);
nand U1090 (N_1090,N_267,N_247);
xnor U1091 (N_1091,N_433,N_762);
nor U1092 (N_1092,N_557,N_84);
or U1093 (N_1093,N_157,N_616);
or U1094 (N_1094,N_401,N_582);
xor U1095 (N_1095,N_221,N_679);
nor U1096 (N_1096,N_797,N_895);
nor U1097 (N_1097,N_133,N_199);
xor U1098 (N_1098,N_984,N_569);
and U1099 (N_1099,N_730,N_316);
xor U1100 (N_1100,N_693,N_231);
and U1101 (N_1101,N_217,N_497);
and U1102 (N_1102,N_789,N_425);
xnor U1103 (N_1103,N_851,N_249);
nor U1104 (N_1104,N_966,N_946);
xnor U1105 (N_1105,N_301,N_92);
xnor U1106 (N_1106,N_261,N_86);
and U1107 (N_1107,N_332,N_183);
or U1108 (N_1108,N_340,N_214);
and U1109 (N_1109,N_364,N_594);
or U1110 (N_1110,N_348,N_838);
or U1111 (N_1111,N_755,N_26);
and U1112 (N_1112,N_624,N_83);
or U1113 (N_1113,N_461,N_695);
nor U1114 (N_1114,N_105,N_592);
nand U1115 (N_1115,N_828,N_983);
or U1116 (N_1116,N_657,N_671);
or U1117 (N_1117,N_385,N_252);
nand U1118 (N_1118,N_737,N_591);
and U1119 (N_1119,N_547,N_82);
xor U1120 (N_1120,N_415,N_293);
xor U1121 (N_1121,N_533,N_307);
and U1122 (N_1122,N_41,N_525);
nor U1123 (N_1123,N_354,N_305);
or U1124 (N_1124,N_485,N_253);
xor U1125 (N_1125,N_795,N_449);
or U1126 (N_1126,N_869,N_613);
xnor U1127 (N_1127,N_520,N_817);
or U1128 (N_1128,N_523,N_602);
or U1129 (N_1129,N_446,N_676);
nand U1130 (N_1130,N_334,N_617);
nand U1131 (N_1131,N_389,N_876);
or U1132 (N_1132,N_927,N_139);
nand U1133 (N_1133,N_977,N_539);
or U1134 (N_1134,N_842,N_940);
xnor U1135 (N_1135,N_724,N_502);
or U1136 (N_1136,N_787,N_426);
nor U1137 (N_1137,N_821,N_564);
or U1138 (N_1138,N_232,N_802);
nor U1139 (N_1139,N_109,N_406);
or U1140 (N_1140,N_732,N_248);
xor U1141 (N_1141,N_125,N_226);
nor U1142 (N_1142,N_825,N_632);
or U1143 (N_1143,N_791,N_185);
or U1144 (N_1144,N_622,N_726);
xnor U1145 (N_1145,N_465,N_712);
xor U1146 (N_1146,N_181,N_808);
or U1147 (N_1147,N_549,N_137);
xor U1148 (N_1148,N_643,N_49);
xnor U1149 (N_1149,N_749,N_748);
nor U1150 (N_1150,N_90,N_761);
and U1151 (N_1151,N_957,N_481);
or U1152 (N_1152,N_408,N_756);
xor U1153 (N_1153,N_120,N_140);
or U1154 (N_1154,N_829,N_949);
xnor U1155 (N_1155,N_439,N_738);
xnor U1156 (N_1156,N_973,N_504);
or U1157 (N_1157,N_926,N_441);
xor U1158 (N_1158,N_965,N_215);
or U1159 (N_1159,N_640,N_625);
nor U1160 (N_1160,N_132,N_413);
xnor U1161 (N_1161,N_440,N_173);
xor U1162 (N_1162,N_714,N_470);
xnor U1163 (N_1163,N_353,N_306);
nor U1164 (N_1164,N_149,N_341);
nor U1165 (N_1165,N_281,N_931);
and U1166 (N_1166,N_653,N_411);
xor U1167 (N_1167,N_831,N_605);
xor U1168 (N_1168,N_303,N_54);
and U1169 (N_1169,N_588,N_596);
nor U1170 (N_1170,N_604,N_323);
or U1171 (N_1171,N_127,N_526);
or U1172 (N_1172,N_897,N_416);
or U1173 (N_1173,N_79,N_558);
nor U1174 (N_1174,N_708,N_642);
nor U1175 (N_1175,N_8,N_369);
xor U1176 (N_1176,N_350,N_122);
xnor U1177 (N_1177,N_975,N_688);
nor U1178 (N_1178,N_981,N_943);
and U1179 (N_1179,N_74,N_302);
nor U1180 (N_1180,N_801,N_509);
and U1181 (N_1181,N_877,N_365);
and U1182 (N_1182,N_23,N_67);
or U1183 (N_1183,N_740,N_805);
and U1184 (N_1184,N_770,N_16);
and U1185 (N_1185,N_362,N_870);
nand U1186 (N_1186,N_678,N_283);
nand U1187 (N_1187,N_98,N_169);
and U1188 (N_1188,N_193,N_300);
or U1189 (N_1189,N_322,N_357);
xnor U1190 (N_1190,N_259,N_104);
and U1191 (N_1191,N_107,N_299);
nand U1192 (N_1192,N_675,N_278);
or U1193 (N_1193,N_950,N_562);
nand U1194 (N_1194,N_811,N_487);
or U1195 (N_1195,N_116,N_150);
xnor U1196 (N_1196,N_736,N_129);
or U1197 (N_1197,N_598,N_397);
nand U1198 (N_1198,N_32,N_46);
nand U1199 (N_1199,N_907,N_197);
nand U1200 (N_1200,N_318,N_719);
nor U1201 (N_1201,N_402,N_179);
or U1202 (N_1202,N_986,N_615);
nor U1203 (N_1203,N_987,N_508);
xnor U1204 (N_1204,N_398,N_570);
nand U1205 (N_1205,N_711,N_466);
nor U1206 (N_1206,N_478,N_399);
and U1207 (N_1207,N_100,N_768);
xor U1208 (N_1208,N_506,N_572);
nand U1209 (N_1209,N_701,N_421);
and U1210 (N_1210,N_263,N_383);
or U1211 (N_1211,N_400,N_94);
or U1212 (N_1212,N_621,N_979);
nor U1213 (N_1213,N_495,N_228);
nor U1214 (N_1214,N_930,N_21);
nand U1215 (N_1215,N_390,N_810);
nand U1216 (N_1216,N_27,N_324);
or U1217 (N_1217,N_524,N_993);
nor U1218 (N_1218,N_575,N_18);
xor U1219 (N_1219,N_351,N_257);
nand U1220 (N_1220,N_991,N_48);
nor U1221 (N_1221,N_99,N_937);
xnor U1222 (N_1222,N_2,N_64);
or U1223 (N_1223,N_40,N_757);
nor U1224 (N_1224,N_168,N_277);
nand U1225 (N_1225,N_967,N_775);
and U1226 (N_1226,N_595,N_326);
xnor U1227 (N_1227,N_610,N_118);
or U1228 (N_1228,N_959,N_744);
nor U1229 (N_1229,N_31,N_781);
xnor U1230 (N_1230,N_734,N_370);
and U1231 (N_1231,N_672,N_180);
or U1232 (N_1232,N_778,N_89);
nand U1233 (N_1233,N_689,N_240);
or U1234 (N_1234,N_492,N_751);
xnor U1235 (N_1235,N_208,N_538);
nand U1236 (N_1236,N_608,N_453);
nor U1237 (N_1237,N_637,N_382);
and U1238 (N_1238,N_391,N_469);
nor U1239 (N_1239,N_459,N_515);
nor U1240 (N_1240,N_360,N_735);
xor U1241 (N_1241,N_705,N_165);
nor U1242 (N_1242,N_251,N_664);
and U1243 (N_1243,N_134,N_55);
nand U1244 (N_1244,N_848,N_147);
or U1245 (N_1245,N_773,N_124);
xor U1246 (N_1246,N_420,N_312);
nand U1247 (N_1247,N_174,N_442);
nand U1248 (N_1248,N_913,N_503);
xor U1249 (N_1249,N_793,N_527);
nor U1250 (N_1250,N_310,N_710);
and U1251 (N_1251,N_537,N_479);
or U1252 (N_1252,N_677,N_143);
xor U1253 (N_1253,N_694,N_335);
or U1254 (N_1254,N_707,N_597);
or U1255 (N_1255,N_685,N_863);
and U1256 (N_1256,N_951,N_634);
nand U1257 (N_1257,N_355,N_667);
and U1258 (N_1258,N_916,N_552);
xnor U1259 (N_1259,N_780,N_91);
and U1260 (N_1260,N_704,N_836);
and U1261 (N_1261,N_891,N_792);
xor U1262 (N_1262,N_111,N_534);
nor U1263 (N_1263,N_952,N_414);
nand U1264 (N_1264,N_227,N_717);
or U1265 (N_1265,N_96,N_102);
and U1266 (N_1266,N_803,N_655);
nor U1267 (N_1267,N_702,N_337);
and U1268 (N_1268,N_250,N_654);
and U1269 (N_1269,N_56,N_545);
nand U1270 (N_1270,N_392,N_809);
xnor U1271 (N_1271,N_682,N_914);
nor U1272 (N_1272,N_573,N_212);
xor U1273 (N_1273,N_119,N_706);
and U1274 (N_1274,N_834,N_813);
nor U1275 (N_1275,N_990,N_130);
and U1276 (N_1276,N_343,N_258);
and U1277 (N_1277,N_532,N_182);
nor U1278 (N_1278,N_860,N_462);
and U1279 (N_1279,N_167,N_571);
nand U1280 (N_1280,N_210,N_234);
or U1281 (N_1281,N_600,N_404);
and U1282 (N_1282,N_450,N_839);
xor U1283 (N_1283,N_841,N_12);
or U1284 (N_1284,N_544,N_758);
and U1285 (N_1285,N_565,N_321);
nor U1286 (N_1286,N_901,N_171);
nand U1287 (N_1287,N_345,N_73);
xnor U1288 (N_1288,N_292,N_908);
nor U1289 (N_1289,N_882,N_342);
nor U1290 (N_1290,N_731,N_857);
or U1291 (N_1291,N_764,N_423);
nand U1292 (N_1292,N_578,N_403);
xnor U1293 (N_1293,N_126,N_239);
nand U1294 (N_1294,N_57,N_980);
xnor U1295 (N_1295,N_388,N_674);
nor U1296 (N_1296,N_530,N_555);
and U1297 (N_1297,N_510,N_507);
nor U1298 (N_1298,N_476,N_893);
nor U1299 (N_1299,N_170,N_436);
and U1300 (N_1300,N_999,N_464);
and U1301 (N_1301,N_760,N_911);
nand U1302 (N_1302,N_78,N_224);
nor U1303 (N_1303,N_904,N_785);
or U1304 (N_1304,N_319,N_216);
nor U1305 (N_1305,N_336,N_95);
or U1306 (N_1306,N_799,N_412);
xnor U1307 (N_1307,N_188,N_356);
nand U1308 (N_1308,N_826,N_948);
xor U1309 (N_1309,N_579,N_424);
nor U1310 (N_1310,N_255,N_783);
nor U1311 (N_1311,N_798,N_513);
or U1312 (N_1312,N_700,N_36);
xor U1313 (N_1313,N_472,N_517);
or U1314 (N_1314,N_874,N_242);
nor U1315 (N_1315,N_276,N_202);
nand U1316 (N_1316,N_87,N_518);
nor U1317 (N_1317,N_338,N_13);
nor U1318 (N_1318,N_123,N_593);
nand U1319 (N_1319,N_178,N_614);
or U1320 (N_1320,N_892,N_896);
xnor U1321 (N_1321,N_271,N_381);
xor U1322 (N_1322,N_611,N_71);
nand U1323 (N_1323,N_192,N_434);
and U1324 (N_1324,N_33,N_516);
nor U1325 (N_1325,N_175,N_101);
nand U1326 (N_1326,N_363,N_739);
nand U1327 (N_1327,N_752,N_405);
nand U1328 (N_1328,N_112,N_788);
xor U1329 (N_1329,N_496,N_641);
nor U1330 (N_1330,N_759,N_313);
xor U1331 (N_1331,N_697,N_238);
or U1332 (N_1332,N_128,N_275);
nor U1333 (N_1333,N_282,N_528);
xor U1334 (N_1334,N_885,N_945);
nor U1335 (N_1335,N_451,N_988);
and U1336 (N_1336,N_587,N_989);
and U1337 (N_1337,N_6,N_455);
nand U1338 (N_1338,N_796,N_568);
nand U1339 (N_1339,N_769,N_28);
nor U1340 (N_1340,N_328,N_163);
nand U1341 (N_1341,N_330,N_262);
or U1342 (N_1342,N_703,N_474);
or U1343 (N_1343,N_561,N_716);
nand U1344 (N_1344,N_919,N_771);
and U1345 (N_1345,N_824,N_14);
nor U1346 (N_1346,N_146,N_807);
nand U1347 (N_1347,N_747,N_947);
nor U1348 (N_1348,N_268,N_280);
xnor U1349 (N_1349,N_121,N_862);
and U1350 (N_1350,N_686,N_443);
nor U1351 (N_1351,N_230,N_550);
or U1352 (N_1352,N_548,N_47);
xnor U1353 (N_1353,N_864,N_347);
and U1354 (N_1354,N_254,N_871);
xor U1355 (N_1355,N_938,N_205);
nor U1356 (N_1356,N_794,N_601);
nand U1357 (N_1357,N_256,N_15);
nand U1358 (N_1358,N_50,N_471);
nor U1359 (N_1359,N_727,N_447);
nand U1360 (N_1360,N_883,N_673);
and U1361 (N_1361,N_144,N_407);
nand U1362 (N_1362,N_633,N_361);
and U1363 (N_1363,N_241,N_576);
and U1364 (N_1364,N_887,N_349);
and U1365 (N_1365,N_880,N_491);
nor U1366 (N_1366,N_709,N_427);
nand U1367 (N_1367,N_159,N_287);
xor U1368 (N_1368,N_894,N_962);
nor U1369 (N_1369,N_154,N_189);
nand U1370 (N_1370,N_884,N_142);
and U1371 (N_1371,N_162,N_148);
nor U1372 (N_1372,N_396,N_903);
and U1373 (N_1373,N_767,N_969);
nor U1374 (N_1374,N_827,N_832);
nand U1375 (N_1375,N_460,N_274);
or U1376 (N_1376,N_211,N_790);
xnor U1377 (N_1377,N_923,N_229);
and U1378 (N_1378,N_881,N_765);
xnor U1379 (N_1379,N_844,N_384);
or U1380 (N_1380,N_875,N_782);
or U1381 (N_1381,N_898,N_647);
nand U1382 (N_1382,N_847,N_68);
nand U1383 (N_1383,N_304,N_660);
and U1384 (N_1384,N_81,N_835);
xnor U1385 (N_1385,N_974,N_531);
nand U1386 (N_1386,N_623,N_260);
xnor U1387 (N_1387,N_814,N_590);
or U1388 (N_1388,N_535,N_117);
nor U1389 (N_1389,N_176,N_166);
nand U1390 (N_1390,N_720,N_646);
nor U1391 (N_1391,N_766,N_444);
nand U1392 (N_1392,N_428,N_186);
nand U1393 (N_1393,N_19,N_665);
and U1394 (N_1394,N_776,N_872);
xnor U1395 (N_1395,N_909,N_53);
nand U1396 (N_1396,N_777,N_387);
and U1397 (N_1397,N_85,N_63);
nor U1398 (N_1398,N_631,N_269);
nor U1399 (N_1399,N_754,N_379);
nand U1400 (N_1400,N_956,N_833);
and U1401 (N_1401,N_753,N_195);
xnor U1402 (N_1402,N_820,N_284);
and U1403 (N_1403,N_77,N_331);
nor U1404 (N_1404,N_76,N_191);
xnor U1405 (N_1405,N_978,N_29);
or U1406 (N_1406,N_652,N_932);
nor U1407 (N_1407,N_473,N_196);
nor U1408 (N_1408,N_609,N_910);
nand U1409 (N_1409,N_546,N_746);
nor U1410 (N_1410,N_589,N_964);
nand U1411 (N_1411,N_9,N_627);
xor U1412 (N_1412,N_264,N_156);
xnor U1413 (N_1413,N_995,N_816);
nand U1414 (N_1414,N_512,N_320);
nor U1415 (N_1415,N_970,N_915);
nand U1416 (N_1416,N_741,N_418);
xor U1417 (N_1417,N_972,N_868);
and U1418 (N_1418,N_66,N_61);
and U1419 (N_1419,N_457,N_886);
or U1420 (N_1420,N_635,N_982);
nor U1421 (N_1421,N_850,N_683);
or U1422 (N_1422,N_486,N_997);
nor U1423 (N_1423,N_0,N_135);
and U1424 (N_1424,N_830,N_273);
nor U1425 (N_1425,N_207,N_245);
and U1426 (N_1426,N_629,N_505);
or U1427 (N_1427,N_968,N_3);
nor U1428 (N_1428,N_620,N_244);
xnor U1429 (N_1429,N_960,N_815);
or U1430 (N_1430,N_529,N_648);
and U1431 (N_1431,N_11,N_422);
or U1432 (N_1432,N_511,N_374);
or U1433 (N_1433,N_88,N_658);
and U1434 (N_1434,N_542,N_201);
and U1435 (N_1435,N_136,N_763);
xor U1436 (N_1436,N_25,N_499);
xor U1437 (N_1437,N_681,N_432);
nand U1438 (N_1438,N_110,N_177);
nand U1439 (N_1439,N_498,N_266);
nor U1440 (N_1440,N_200,N_288);
or U1441 (N_1441,N_574,N_750);
xnor U1442 (N_1442,N_70,N_467);
or U1443 (N_1443,N_187,N_265);
or U1444 (N_1444,N_992,N_958);
and U1445 (N_1445,N_272,N_733);
nor U1446 (N_1446,N_963,N_942);
and U1447 (N_1447,N_35,N_644);
nor U1448 (N_1448,N_666,N_477);
and U1449 (N_1449,N_560,N_619);
or U1450 (N_1450,N_556,N_662);
nand U1451 (N_1451,N_184,N_580);
nor U1452 (N_1452,N_944,N_728);
nor U1453 (N_1453,N_489,N_409);
and U1454 (N_1454,N_289,N_961);
or U1455 (N_1455,N_158,N_4);
nor U1456 (N_1456,N_225,N_315);
xnor U1457 (N_1457,N_164,N_924);
xor U1458 (N_1458,N_722,N_603);
nor U1459 (N_1459,N_985,N_51);
or U1460 (N_1460,N_38,N_161);
nor U1461 (N_1461,N_309,N_541);
or U1462 (N_1462,N_233,N_630);
nor U1463 (N_1463,N_607,N_933);
and U1464 (N_1464,N_900,N_44);
nand U1465 (N_1465,N_429,N_743);
or U1466 (N_1466,N_490,N_649);
and U1467 (N_1467,N_819,N_853);
or U1468 (N_1468,N_925,N_650);
xor U1469 (N_1469,N_721,N_784);
nor U1470 (N_1470,N_1,N_454);
and U1471 (N_1471,N_59,N_270);
xor U1472 (N_1472,N_380,N_906);
nand U1473 (N_1473,N_93,N_878);
and U1474 (N_1474,N_858,N_39);
or U1475 (N_1475,N_866,N_366);
nand U1476 (N_1476,N_80,N_599);
or U1477 (N_1477,N_475,N_725);
xnor U1478 (N_1478,N_645,N_822);
and U1479 (N_1479,N_718,N_921);
nand U1480 (N_1480,N_329,N_583);
nor U1481 (N_1481,N_372,N_456);
xor U1482 (N_1482,N_584,N_856);
and U1483 (N_1483,N_500,N_713);
xor U1484 (N_1484,N_97,N_585);
xnor U1485 (N_1485,N_115,N_30);
and U1486 (N_1486,N_638,N_715);
nor U1487 (N_1487,N_669,N_10);
nand U1488 (N_1488,N_889,N_849);
nand U1489 (N_1489,N_69,N_745);
or U1490 (N_1490,N_378,N_692);
or U1491 (N_1491,N_612,N_494);
nor U1492 (N_1492,N_536,N_237);
and U1493 (N_1493,N_155,N_445);
xnor U1494 (N_1494,N_34,N_551);
and U1495 (N_1495,N_922,N_845);
nand U1496 (N_1496,N_935,N_468);
nand U1497 (N_1497,N_223,N_204);
or U1498 (N_1498,N_920,N_954);
nor U1499 (N_1499,N_62,N_800);
nand U1500 (N_1500,N_458,N_907);
xnor U1501 (N_1501,N_276,N_634);
nor U1502 (N_1502,N_587,N_904);
nor U1503 (N_1503,N_210,N_10);
and U1504 (N_1504,N_228,N_976);
and U1505 (N_1505,N_525,N_301);
xor U1506 (N_1506,N_150,N_51);
and U1507 (N_1507,N_891,N_713);
nand U1508 (N_1508,N_884,N_86);
and U1509 (N_1509,N_295,N_396);
or U1510 (N_1510,N_470,N_468);
xor U1511 (N_1511,N_873,N_649);
or U1512 (N_1512,N_707,N_507);
xnor U1513 (N_1513,N_805,N_940);
nor U1514 (N_1514,N_959,N_507);
nor U1515 (N_1515,N_107,N_199);
xnor U1516 (N_1516,N_625,N_626);
xnor U1517 (N_1517,N_268,N_474);
nor U1518 (N_1518,N_649,N_228);
nor U1519 (N_1519,N_754,N_355);
xor U1520 (N_1520,N_19,N_596);
and U1521 (N_1521,N_107,N_828);
nor U1522 (N_1522,N_215,N_538);
nand U1523 (N_1523,N_132,N_798);
or U1524 (N_1524,N_389,N_207);
xor U1525 (N_1525,N_427,N_938);
nor U1526 (N_1526,N_341,N_309);
xor U1527 (N_1527,N_976,N_799);
and U1528 (N_1528,N_927,N_392);
and U1529 (N_1529,N_78,N_175);
or U1530 (N_1530,N_756,N_951);
or U1531 (N_1531,N_76,N_671);
and U1532 (N_1532,N_621,N_368);
xnor U1533 (N_1533,N_77,N_504);
or U1534 (N_1534,N_862,N_197);
or U1535 (N_1535,N_222,N_570);
or U1536 (N_1536,N_236,N_616);
and U1537 (N_1537,N_106,N_556);
or U1538 (N_1538,N_94,N_322);
nand U1539 (N_1539,N_600,N_961);
nor U1540 (N_1540,N_394,N_34);
nand U1541 (N_1541,N_918,N_213);
nand U1542 (N_1542,N_127,N_892);
or U1543 (N_1543,N_371,N_840);
nand U1544 (N_1544,N_299,N_720);
or U1545 (N_1545,N_525,N_145);
nand U1546 (N_1546,N_109,N_215);
nand U1547 (N_1547,N_62,N_197);
nor U1548 (N_1548,N_696,N_686);
nand U1549 (N_1549,N_495,N_952);
and U1550 (N_1550,N_260,N_690);
xnor U1551 (N_1551,N_313,N_171);
nor U1552 (N_1552,N_658,N_181);
xnor U1553 (N_1553,N_323,N_85);
or U1554 (N_1554,N_708,N_42);
and U1555 (N_1555,N_552,N_231);
and U1556 (N_1556,N_911,N_384);
and U1557 (N_1557,N_777,N_147);
xnor U1558 (N_1558,N_753,N_308);
nand U1559 (N_1559,N_85,N_696);
and U1560 (N_1560,N_458,N_878);
and U1561 (N_1561,N_760,N_219);
xor U1562 (N_1562,N_632,N_912);
nor U1563 (N_1563,N_810,N_102);
xor U1564 (N_1564,N_889,N_715);
nor U1565 (N_1565,N_858,N_769);
or U1566 (N_1566,N_770,N_92);
xor U1567 (N_1567,N_876,N_699);
nor U1568 (N_1568,N_959,N_760);
nand U1569 (N_1569,N_865,N_121);
nor U1570 (N_1570,N_679,N_598);
nor U1571 (N_1571,N_177,N_896);
and U1572 (N_1572,N_460,N_47);
or U1573 (N_1573,N_367,N_13);
and U1574 (N_1574,N_8,N_933);
and U1575 (N_1575,N_101,N_335);
nor U1576 (N_1576,N_396,N_194);
or U1577 (N_1577,N_229,N_307);
and U1578 (N_1578,N_379,N_492);
xor U1579 (N_1579,N_200,N_409);
and U1580 (N_1580,N_480,N_411);
nand U1581 (N_1581,N_676,N_637);
or U1582 (N_1582,N_937,N_94);
or U1583 (N_1583,N_104,N_228);
and U1584 (N_1584,N_43,N_215);
nand U1585 (N_1585,N_457,N_685);
or U1586 (N_1586,N_972,N_688);
nand U1587 (N_1587,N_53,N_558);
nor U1588 (N_1588,N_410,N_119);
and U1589 (N_1589,N_554,N_949);
nor U1590 (N_1590,N_574,N_547);
xor U1591 (N_1591,N_386,N_343);
nor U1592 (N_1592,N_702,N_364);
nor U1593 (N_1593,N_107,N_89);
and U1594 (N_1594,N_507,N_77);
or U1595 (N_1595,N_504,N_139);
or U1596 (N_1596,N_858,N_556);
and U1597 (N_1597,N_94,N_876);
nor U1598 (N_1598,N_499,N_221);
or U1599 (N_1599,N_739,N_339);
and U1600 (N_1600,N_537,N_344);
nor U1601 (N_1601,N_829,N_572);
or U1602 (N_1602,N_16,N_342);
xnor U1603 (N_1603,N_752,N_707);
nand U1604 (N_1604,N_723,N_577);
nor U1605 (N_1605,N_47,N_969);
nand U1606 (N_1606,N_289,N_336);
and U1607 (N_1607,N_324,N_606);
and U1608 (N_1608,N_16,N_527);
nor U1609 (N_1609,N_32,N_560);
nand U1610 (N_1610,N_932,N_880);
nand U1611 (N_1611,N_225,N_541);
or U1612 (N_1612,N_544,N_978);
nor U1613 (N_1613,N_872,N_775);
nor U1614 (N_1614,N_376,N_786);
and U1615 (N_1615,N_94,N_629);
xnor U1616 (N_1616,N_168,N_264);
xor U1617 (N_1617,N_603,N_542);
xnor U1618 (N_1618,N_970,N_164);
nor U1619 (N_1619,N_954,N_820);
xor U1620 (N_1620,N_873,N_652);
or U1621 (N_1621,N_841,N_265);
nand U1622 (N_1622,N_963,N_116);
or U1623 (N_1623,N_852,N_412);
nor U1624 (N_1624,N_966,N_396);
or U1625 (N_1625,N_888,N_180);
nor U1626 (N_1626,N_696,N_578);
nor U1627 (N_1627,N_922,N_96);
and U1628 (N_1628,N_63,N_157);
xnor U1629 (N_1629,N_170,N_863);
nor U1630 (N_1630,N_121,N_821);
nand U1631 (N_1631,N_830,N_560);
or U1632 (N_1632,N_268,N_718);
and U1633 (N_1633,N_10,N_674);
or U1634 (N_1634,N_101,N_223);
xnor U1635 (N_1635,N_905,N_249);
nor U1636 (N_1636,N_552,N_472);
or U1637 (N_1637,N_615,N_159);
or U1638 (N_1638,N_823,N_931);
and U1639 (N_1639,N_839,N_133);
xnor U1640 (N_1640,N_153,N_185);
or U1641 (N_1641,N_523,N_985);
and U1642 (N_1642,N_16,N_435);
nor U1643 (N_1643,N_198,N_300);
nor U1644 (N_1644,N_729,N_604);
nor U1645 (N_1645,N_456,N_95);
and U1646 (N_1646,N_598,N_964);
nand U1647 (N_1647,N_32,N_122);
or U1648 (N_1648,N_375,N_755);
xnor U1649 (N_1649,N_684,N_165);
or U1650 (N_1650,N_32,N_496);
and U1651 (N_1651,N_618,N_45);
or U1652 (N_1652,N_277,N_628);
and U1653 (N_1653,N_466,N_423);
xor U1654 (N_1654,N_776,N_390);
nand U1655 (N_1655,N_100,N_701);
nor U1656 (N_1656,N_790,N_347);
or U1657 (N_1657,N_483,N_505);
and U1658 (N_1658,N_765,N_690);
nand U1659 (N_1659,N_788,N_57);
nand U1660 (N_1660,N_586,N_711);
xor U1661 (N_1661,N_47,N_386);
nand U1662 (N_1662,N_965,N_848);
nor U1663 (N_1663,N_287,N_293);
nand U1664 (N_1664,N_106,N_718);
xnor U1665 (N_1665,N_527,N_865);
nor U1666 (N_1666,N_640,N_705);
nor U1667 (N_1667,N_993,N_553);
and U1668 (N_1668,N_216,N_134);
nand U1669 (N_1669,N_606,N_989);
xnor U1670 (N_1670,N_910,N_423);
nor U1671 (N_1671,N_721,N_239);
and U1672 (N_1672,N_616,N_61);
and U1673 (N_1673,N_523,N_711);
and U1674 (N_1674,N_796,N_367);
xnor U1675 (N_1675,N_649,N_909);
xor U1676 (N_1676,N_710,N_617);
nor U1677 (N_1677,N_812,N_792);
or U1678 (N_1678,N_991,N_845);
nand U1679 (N_1679,N_733,N_215);
nand U1680 (N_1680,N_319,N_18);
or U1681 (N_1681,N_791,N_788);
and U1682 (N_1682,N_315,N_431);
and U1683 (N_1683,N_643,N_666);
or U1684 (N_1684,N_230,N_236);
nand U1685 (N_1685,N_896,N_862);
nor U1686 (N_1686,N_724,N_927);
and U1687 (N_1687,N_490,N_372);
or U1688 (N_1688,N_780,N_514);
nor U1689 (N_1689,N_699,N_796);
and U1690 (N_1690,N_410,N_859);
nand U1691 (N_1691,N_734,N_706);
nand U1692 (N_1692,N_470,N_249);
or U1693 (N_1693,N_522,N_736);
nor U1694 (N_1694,N_537,N_956);
or U1695 (N_1695,N_223,N_105);
or U1696 (N_1696,N_246,N_948);
nor U1697 (N_1697,N_438,N_560);
nor U1698 (N_1698,N_99,N_617);
nand U1699 (N_1699,N_394,N_527);
xnor U1700 (N_1700,N_91,N_960);
and U1701 (N_1701,N_991,N_859);
xnor U1702 (N_1702,N_481,N_488);
nand U1703 (N_1703,N_319,N_895);
nor U1704 (N_1704,N_722,N_792);
or U1705 (N_1705,N_169,N_833);
nor U1706 (N_1706,N_837,N_756);
nor U1707 (N_1707,N_418,N_619);
or U1708 (N_1708,N_659,N_813);
or U1709 (N_1709,N_805,N_381);
and U1710 (N_1710,N_923,N_616);
and U1711 (N_1711,N_326,N_93);
and U1712 (N_1712,N_595,N_469);
xnor U1713 (N_1713,N_907,N_898);
nor U1714 (N_1714,N_697,N_852);
or U1715 (N_1715,N_272,N_794);
or U1716 (N_1716,N_622,N_645);
xnor U1717 (N_1717,N_277,N_930);
nor U1718 (N_1718,N_912,N_520);
nor U1719 (N_1719,N_830,N_49);
nor U1720 (N_1720,N_933,N_206);
nor U1721 (N_1721,N_949,N_220);
nand U1722 (N_1722,N_117,N_159);
xnor U1723 (N_1723,N_795,N_75);
nor U1724 (N_1724,N_953,N_383);
nor U1725 (N_1725,N_607,N_223);
xor U1726 (N_1726,N_528,N_23);
xor U1727 (N_1727,N_819,N_716);
nand U1728 (N_1728,N_396,N_180);
and U1729 (N_1729,N_40,N_973);
nor U1730 (N_1730,N_17,N_600);
nand U1731 (N_1731,N_996,N_523);
nand U1732 (N_1732,N_223,N_509);
xor U1733 (N_1733,N_415,N_261);
nor U1734 (N_1734,N_408,N_725);
nor U1735 (N_1735,N_360,N_623);
nand U1736 (N_1736,N_423,N_957);
nor U1737 (N_1737,N_270,N_868);
and U1738 (N_1738,N_669,N_656);
and U1739 (N_1739,N_935,N_928);
or U1740 (N_1740,N_892,N_68);
and U1741 (N_1741,N_856,N_307);
nand U1742 (N_1742,N_513,N_455);
nand U1743 (N_1743,N_323,N_117);
nand U1744 (N_1744,N_348,N_642);
nand U1745 (N_1745,N_289,N_933);
or U1746 (N_1746,N_406,N_312);
or U1747 (N_1747,N_825,N_820);
nand U1748 (N_1748,N_384,N_794);
nor U1749 (N_1749,N_791,N_290);
and U1750 (N_1750,N_628,N_792);
nor U1751 (N_1751,N_716,N_145);
and U1752 (N_1752,N_556,N_971);
or U1753 (N_1753,N_212,N_594);
and U1754 (N_1754,N_614,N_783);
or U1755 (N_1755,N_398,N_702);
and U1756 (N_1756,N_290,N_186);
nor U1757 (N_1757,N_928,N_302);
nand U1758 (N_1758,N_133,N_80);
and U1759 (N_1759,N_747,N_229);
or U1760 (N_1760,N_343,N_881);
nor U1761 (N_1761,N_220,N_667);
xnor U1762 (N_1762,N_131,N_787);
nand U1763 (N_1763,N_123,N_557);
or U1764 (N_1764,N_83,N_325);
and U1765 (N_1765,N_405,N_111);
nand U1766 (N_1766,N_713,N_947);
and U1767 (N_1767,N_995,N_743);
and U1768 (N_1768,N_475,N_769);
xnor U1769 (N_1769,N_57,N_100);
xor U1770 (N_1770,N_869,N_616);
nand U1771 (N_1771,N_86,N_241);
and U1772 (N_1772,N_482,N_921);
or U1773 (N_1773,N_623,N_482);
nor U1774 (N_1774,N_588,N_237);
nand U1775 (N_1775,N_901,N_388);
xnor U1776 (N_1776,N_847,N_777);
or U1777 (N_1777,N_516,N_383);
and U1778 (N_1778,N_663,N_131);
nand U1779 (N_1779,N_498,N_509);
nor U1780 (N_1780,N_805,N_497);
or U1781 (N_1781,N_943,N_244);
nor U1782 (N_1782,N_482,N_542);
nor U1783 (N_1783,N_357,N_414);
or U1784 (N_1784,N_228,N_217);
or U1785 (N_1785,N_911,N_994);
and U1786 (N_1786,N_206,N_686);
and U1787 (N_1787,N_718,N_220);
or U1788 (N_1788,N_802,N_139);
and U1789 (N_1789,N_804,N_436);
and U1790 (N_1790,N_706,N_61);
or U1791 (N_1791,N_564,N_134);
nand U1792 (N_1792,N_279,N_702);
xnor U1793 (N_1793,N_937,N_208);
xnor U1794 (N_1794,N_640,N_469);
xnor U1795 (N_1795,N_307,N_339);
or U1796 (N_1796,N_765,N_216);
or U1797 (N_1797,N_827,N_456);
and U1798 (N_1798,N_903,N_927);
or U1799 (N_1799,N_424,N_361);
or U1800 (N_1800,N_526,N_737);
xor U1801 (N_1801,N_187,N_213);
xor U1802 (N_1802,N_200,N_12);
nand U1803 (N_1803,N_440,N_589);
nor U1804 (N_1804,N_583,N_296);
and U1805 (N_1805,N_686,N_838);
xor U1806 (N_1806,N_298,N_271);
nor U1807 (N_1807,N_52,N_343);
xor U1808 (N_1808,N_134,N_377);
and U1809 (N_1809,N_995,N_87);
or U1810 (N_1810,N_121,N_536);
nand U1811 (N_1811,N_383,N_67);
and U1812 (N_1812,N_372,N_287);
nor U1813 (N_1813,N_868,N_295);
nor U1814 (N_1814,N_942,N_204);
nand U1815 (N_1815,N_384,N_682);
xor U1816 (N_1816,N_363,N_570);
xor U1817 (N_1817,N_219,N_382);
nor U1818 (N_1818,N_515,N_982);
or U1819 (N_1819,N_157,N_111);
and U1820 (N_1820,N_102,N_821);
xor U1821 (N_1821,N_327,N_521);
xnor U1822 (N_1822,N_80,N_72);
nand U1823 (N_1823,N_380,N_917);
and U1824 (N_1824,N_259,N_185);
or U1825 (N_1825,N_998,N_490);
and U1826 (N_1826,N_292,N_14);
xnor U1827 (N_1827,N_746,N_276);
xnor U1828 (N_1828,N_570,N_370);
nand U1829 (N_1829,N_286,N_407);
nand U1830 (N_1830,N_660,N_151);
nor U1831 (N_1831,N_495,N_522);
nor U1832 (N_1832,N_904,N_656);
and U1833 (N_1833,N_493,N_535);
or U1834 (N_1834,N_911,N_702);
or U1835 (N_1835,N_653,N_721);
xnor U1836 (N_1836,N_910,N_480);
nand U1837 (N_1837,N_243,N_162);
nor U1838 (N_1838,N_300,N_133);
xnor U1839 (N_1839,N_446,N_828);
or U1840 (N_1840,N_782,N_18);
xnor U1841 (N_1841,N_748,N_573);
xnor U1842 (N_1842,N_215,N_620);
and U1843 (N_1843,N_612,N_11);
xor U1844 (N_1844,N_212,N_506);
xnor U1845 (N_1845,N_330,N_192);
nor U1846 (N_1846,N_565,N_796);
xnor U1847 (N_1847,N_778,N_967);
nand U1848 (N_1848,N_322,N_777);
and U1849 (N_1849,N_340,N_284);
nand U1850 (N_1850,N_737,N_434);
or U1851 (N_1851,N_305,N_5);
nor U1852 (N_1852,N_810,N_584);
and U1853 (N_1853,N_851,N_556);
nor U1854 (N_1854,N_64,N_882);
or U1855 (N_1855,N_27,N_345);
nand U1856 (N_1856,N_686,N_866);
and U1857 (N_1857,N_775,N_884);
and U1858 (N_1858,N_64,N_735);
nor U1859 (N_1859,N_216,N_430);
or U1860 (N_1860,N_478,N_284);
nor U1861 (N_1861,N_494,N_357);
or U1862 (N_1862,N_965,N_224);
xnor U1863 (N_1863,N_413,N_948);
and U1864 (N_1864,N_213,N_52);
nand U1865 (N_1865,N_80,N_749);
nand U1866 (N_1866,N_489,N_355);
nand U1867 (N_1867,N_851,N_734);
xor U1868 (N_1868,N_418,N_268);
and U1869 (N_1869,N_637,N_959);
xnor U1870 (N_1870,N_7,N_876);
nand U1871 (N_1871,N_936,N_898);
xor U1872 (N_1872,N_503,N_163);
xnor U1873 (N_1873,N_629,N_935);
and U1874 (N_1874,N_114,N_854);
xor U1875 (N_1875,N_655,N_12);
and U1876 (N_1876,N_200,N_923);
or U1877 (N_1877,N_265,N_549);
nand U1878 (N_1878,N_976,N_467);
xor U1879 (N_1879,N_501,N_957);
and U1880 (N_1880,N_208,N_787);
and U1881 (N_1881,N_993,N_112);
or U1882 (N_1882,N_231,N_114);
xnor U1883 (N_1883,N_0,N_376);
nor U1884 (N_1884,N_901,N_338);
and U1885 (N_1885,N_355,N_308);
and U1886 (N_1886,N_532,N_588);
xnor U1887 (N_1887,N_788,N_310);
nand U1888 (N_1888,N_357,N_928);
and U1889 (N_1889,N_622,N_828);
nand U1890 (N_1890,N_707,N_526);
nand U1891 (N_1891,N_769,N_797);
nand U1892 (N_1892,N_786,N_982);
and U1893 (N_1893,N_491,N_188);
nand U1894 (N_1894,N_767,N_470);
xor U1895 (N_1895,N_991,N_211);
xnor U1896 (N_1896,N_206,N_379);
nor U1897 (N_1897,N_295,N_490);
nand U1898 (N_1898,N_427,N_258);
nand U1899 (N_1899,N_107,N_180);
nor U1900 (N_1900,N_294,N_479);
xnor U1901 (N_1901,N_874,N_786);
xnor U1902 (N_1902,N_739,N_415);
xor U1903 (N_1903,N_993,N_829);
or U1904 (N_1904,N_884,N_429);
nand U1905 (N_1905,N_358,N_194);
nor U1906 (N_1906,N_560,N_713);
xor U1907 (N_1907,N_228,N_632);
nand U1908 (N_1908,N_700,N_800);
and U1909 (N_1909,N_439,N_45);
or U1910 (N_1910,N_811,N_760);
or U1911 (N_1911,N_466,N_896);
xor U1912 (N_1912,N_860,N_523);
and U1913 (N_1913,N_388,N_258);
xnor U1914 (N_1914,N_580,N_239);
and U1915 (N_1915,N_331,N_295);
or U1916 (N_1916,N_198,N_188);
xnor U1917 (N_1917,N_905,N_535);
xor U1918 (N_1918,N_6,N_879);
nor U1919 (N_1919,N_405,N_836);
or U1920 (N_1920,N_757,N_474);
and U1921 (N_1921,N_823,N_510);
or U1922 (N_1922,N_637,N_592);
or U1923 (N_1923,N_976,N_172);
and U1924 (N_1924,N_124,N_84);
or U1925 (N_1925,N_22,N_178);
nor U1926 (N_1926,N_126,N_423);
nand U1927 (N_1927,N_281,N_231);
nor U1928 (N_1928,N_542,N_193);
xnor U1929 (N_1929,N_254,N_36);
or U1930 (N_1930,N_881,N_404);
xnor U1931 (N_1931,N_133,N_236);
nor U1932 (N_1932,N_510,N_584);
or U1933 (N_1933,N_845,N_165);
or U1934 (N_1934,N_638,N_321);
xnor U1935 (N_1935,N_113,N_219);
or U1936 (N_1936,N_748,N_326);
and U1937 (N_1937,N_721,N_996);
xnor U1938 (N_1938,N_8,N_259);
xor U1939 (N_1939,N_221,N_984);
nor U1940 (N_1940,N_952,N_637);
or U1941 (N_1941,N_0,N_137);
nor U1942 (N_1942,N_408,N_33);
nand U1943 (N_1943,N_682,N_745);
or U1944 (N_1944,N_761,N_278);
xor U1945 (N_1945,N_237,N_687);
nand U1946 (N_1946,N_278,N_544);
and U1947 (N_1947,N_820,N_44);
and U1948 (N_1948,N_667,N_371);
and U1949 (N_1949,N_503,N_573);
and U1950 (N_1950,N_938,N_367);
xnor U1951 (N_1951,N_162,N_104);
nor U1952 (N_1952,N_988,N_208);
nor U1953 (N_1953,N_139,N_193);
and U1954 (N_1954,N_617,N_995);
xnor U1955 (N_1955,N_829,N_580);
and U1956 (N_1956,N_145,N_886);
xnor U1957 (N_1957,N_732,N_99);
or U1958 (N_1958,N_557,N_855);
nand U1959 (N_1959,N_670,N_77);
or U1960 (N_1960,N_380,N_12);
xor U1961 (N_1961,N_254,N_949);
or U1962 (N_1962,N_5,N_457);
and U1963 (N_1963,N_658,N_368);
or U1964 (N_1964,N_297,N_938);
nor U1965 (N_1965,N_518,N_65);
nand U1966 (N_1966,N_205,N_980);
xor U1967 (N_1967,N_680,N_137);
and U1968 (N_1968,N_93,N_521);
and U1969 (N_1969,N_879,N_477);
nor U1970 (N_1970,N_388,N_594);
nand U1971 (N_1971,N_968,N_204);
nand U1972 (N_1972,N_83,N_449);
or U1973 (N_1973,N_993,N_709);
nand U1974 (N_1974,N_370,N_913);
xor U1975 (N_1975,N_869,N_331);
or U1976 (N_1976,N_410,N_200);
or U1977 (N_1977,N_256,N_986);
nand U1978 (N_1978,N_5,N_918);
xnor U1979 (N_1979,N_301,N_147);
xnor U1980 (N_1980,N_318,N_396);
xnor U1981 (N_1981,N_294,N_951);
and U1982 (N_1982,N_96,N_407);
and U1983 (N_1983,N_218,N_580);
xor U1984 (N_1984,N_887,N_560);
or U1985 (N_1985,N_398,N_872);
and U1986 (N_1986,N_361,N_717);
nor U1987 (N_1987,N_577,N_433);
nor U1988 (N_1988,N_273,N_215);
or U1989 (N_1989,N_711,N_374);
nor U1990 (N_1990,N_582,N_386);
and U1991 (N_1991,N_481,N_592);
or U1992 (N_1992,N_374,N_97);
nor U1993 (N_1993,N_152,N_308);
and U1994 (N_1994,N_431,N_94);
xor U1995 (N_1995,N_213,N_281);
nor U1996 (N_1996,N_165,N_153);
nand U1997 (N_1997,N_282,N_795);
or U1998 (N_1998,N_614,N_79);
and U1999 (N_1999,N_303,N_544);
nand U2000 (N_2000,N_1819,N_1493);
and U2001 (N_2001,N_1628,N_1383);
xnor U2002 (N_2002,N_1990,N_1419);
nor U2003 (N_2003,N_1901,N_1980);
nor U2004 (N_2004,N_1597,N_1194);
nor U2005 (N_2005,N_1580,N_1035);
and U2006 (N_2006,N_1467,N_1827);
nand U2007 (N_2007,N_1171,N_1009);
xor U2008 (N_2008,N_1655,N_1535);
or U2009 (N_2009,N_1245,N_1501);
or U2010 (N_2010,N_1020,N_1301);
xnor U2011 (N_2011,N_1999,N_1998);
or U2012 (N_2012,N_1526,N_1500);
or U2013 (N_2013,N_1168,N_1314);
nor U2014 (N_2014,N_1831,N_1908);
and U2015 (N_2015,N_1636,N_1802);
nand U2016 (N_2016,N_1511,N_1460);
nand U2017 (N_2017,N_1991,N_1134);
and U2018 (N_2018,N_1119,N_1088);
or U2019 (N_2019,N_1400,N_1272);
nor U2020 (N_2020,N_1654,N_1611);
or U2021 (N_2021,N_1659,N_1118);
and U2022 (N_2022,N_1624,N_1914);
xnor U2023 (N_2023,N_1179,N_1974);
nand U2024 (N_2024,N_1239,N_1300);
nor U2025 (N_2025,N_1533,N_1102);
nor U2026 (N_2026,N_1787,N_1401);
nand U2027 (N_2027,N_1249,N_1713);
and U2028 (N_2028,N_1455,N_1421);
or U2029 (N_2029,N_1860,N_1283);
nand U2030 (N_2030,N_1108,N_1570);
nor U2031 (N_2031,N_1041,N_1717);
nand U2032 (N_2032,N_1862,N_1534);
and U2033 (N_2033,N_1374,N_1276);
or U2034 (N_2034,N_1917,N_1071);
nor U2035 (N_2035,N_1915,N_1816);
nand U2036 (N_2036,N_1855,N_1987);
and U2037 (N_2037,N_1191,N_1904);
nor U2038 (N_2038,N_1432,N_1122);
nand U2039 (N_2039,N_1721,N_1739);
and U2040 (N_2040,N_1436,N_1306);
nand U2041 (N_2041,N_1304,N_1696);
xnor U2042 (N_2042,N_1921,N_1403);
and U2043 (N_2043,N_1516,N_1858);
nor U2044 (N_2044,N_1656,N_1478);
xor U2045 (N_2045,N_1952,N_1155);
and U2046 (N_2046,N_1748,N_1657);
xnor U2047 (N_2047,N_1984,N_1641);
or U2048 (N_2048,N_1532,N_1172);
nand U2049 (N_2049,N_1658,N_1902);
nand U2050 (N_2050,N_1551,N_1878);
xor U2051 (N_2051,N_1224,N_1623);
and U2052 (N_2052,N_1277,N_1107);
xor U2053 (N_2053,N_1390,N_1817);
and U2054 (N_2054,N_1530,N_1664);
or U2055 (N_2055,N_1409,N_1520);
and U2056 (N_2056,N_1602,N_1142);
xnor U2057 (N_2057,N_1617,N_1517);
and U2058 (N_2058,N_1682,N_1295);
nand U2059 (N_2059,N_1693,N_1714);
nand U2060 (N_2060,N_1121,N_1826);
xnor U2061 (N_2061,N_1483,N_1269);
nand U2062 (N_2062,N_1210,N_1268);
nor U2063 (N_2063,N_1413,N_1583);
nand U2064 (N_2064,N_1913,N_1556);
nand U2065 (N_2065,N_1124,N_1876);
and U2066 (N_2066,N_1905,N_1446);
or U2067 (N_2067,N_1979,N_1968);
xor U2068 (N_2068,N_1285,N_1079);
and U2069 (N_2069,N_1680,N_1969);
nand U2070 (N_2070,N_1555,N_1289);
nand U2071 (N_2071,N_1476,N_1547);
or U2072 (N_2072,N_1491,N_1099);
and U2073 (N_2073,N_1907,N_1378);
or U2074 (N_2074,N_1503,N_1997);
xnor U2075 (N_2075,N_1394,N_1133);
nand U2076 (N_2076,N_1506,N_1650);
nor U2077 (N_2077,N_1989,N_1599);
nor U2078 (N_2078,N_1052,N_1462);
and U2079 (N_2079,N_1736,N_1716);
or U2080 (N_2080,N_1967,N_1182);
nor U2081 (N_2081,N_1112,N_1248);
or U2082 (N_2082,N_1320,N_1767);
or U2083 (N_2083,N_1970,N_1927);
nand U2084 (N_2084,N_1890,N_1291);
and U2085 (N_2085,N_1498,N_1196);
xnor U2086 (N_2086,N_1880,N_1138);
xnor U2087 (N_2087,N_1790,N_1110);
nor U2088 (N_2088,N_1738,N_1830);
nand U2089 (N_2089,N_1729,N_1216);
nor U2090 (N_2090,N_1317,N_1246);
xnor U2091 (N_2091,N_1823,N_1935);
nor U2092 (N_2092,N_1040,N_1722);
nand U2093 (N_2093,N_1451,N_1468);
or U2094 (N_2094,N_1264,N_1408);
and U2095 (N_2095,N_1976,N_1331);
nor U2096 (N_2096,N_1377,N_1698);
xor U2097 (N_2097,N_1348,N_1076);
xor U2098 (N_2098,N_1465,N_1297);
or U2099 (N_2099,N_1660,N_1561);
xor U2100 (N_2100,N_1069,N_1481);
xnor U2101 (N_2101,N_1186,N_1527);
xor U2102 (N_2102,N_1852,N_1834);
nor U2103 (N_2103,N_1836,N_1219);
and U2104 (N_2104,N_1058,N_1160);
and U2105 (N_2105,N_1634,N_1427);
xor U2106 (N_2106,N_1089,N_1537);
and U2107 (N_2107,N_1866,N_1543);
xor U2108 (N_2108,N_1701,N_1447);
nand U2109 (N_2109,N_1983,N_1311);
xnor U2110 (N_2110,N_1798,N_1029);
and U2111 (N_2111,N_1461,N_1874);
or U2112 (N_2112,N_1606,N_1280);
nor U2113 (N_2113,N_1888,N_1485);
or U2114 (N_2114,N_1095,N_1309);
xor U2115 (N_2115,N_1185,N_1443);
or U2116 (N_2116,N_1008,N_1452);
and U2117 (N_2117,N_1672,N_1933);
nor U2118 (N_2118,N_1388,N_1104);
xnor U2119 (N_2119,N_1958,N_1153);
and U2120 (N_2120,N_1971,N_1711);
or U2121 (N_2121,N_1034,N_1594);
and U2122 (N_2122,N_1985,N_1018);
nor U2123 (N_2123,N_1600,N_1601);
and U2124 (N_2124,N_1061,N_1275);
xor U2125 (N_2125,N_1082,N_1870);
nand U2126 (N_2126,N_1892,N_1023);
and U2127 (N_2127,N_1307,N_1719);
or U2128 (N_2128,N_1699,N_1885);
xnor U2129 (N_2129,N_1643,N_1355);
xnor U2130 (N_2130,N_1258,N_1369);
xnor U2131 (N_2131,N_1703,N_1632);
and U2132 (N_2132,N_1541,N_1562);
and U2133 (N_2133,N_1635,N_1621);
or U2134 (N_2134,N_1842,N_1811);
xor U2135 (N_2135,N_1163,N_1916);
and U2136 (N_2136,N_1093,N_1864);
or U2137 (N_2137,N_1120,N_1702);
and U2138 (N_2138,N_1205,N_1528);
nand U2139 (N_2139,N_1689,N_1358);
nand U2140 (N_2140,N_1415,N_1912);
nand U2141 (N_2141,N_1324,N_1648);
nor U2142 (N_2142,N_1723,N_1173);
nand U2143 (N_2143,N_1150,N_1257);
xor U2144 (N_2144,N_1457,N_1220);
xnor U2145 (N_2145,N_1117,N_1612);
or U2146 (N_2146,N_1376,N_1563);
or U2147 (N_2147,N_1715,N_1128);
nand U2148 (N_2148,N_1751,N_1484);
nor U2149 (N_2149,N_1202,N_1345);
and U2150 (N_2150,N_1233,N_1166);
and U2151 (N_2151,N_1496,N_1406);
and U2152 (N_2152,N_1809,N_1323);
and U2153 (N_2153,N_1208,N_1303);
xnor U2154 (N_2154,N_1545,N_1550);
xor U2155 (N_2155,N_1906,N_1039);
xnor U2156 (N_2156,N_1760,N_1895);
xnor U2157 (N_2157,N_1992,N_1235);
nor U2158 (N_2158,N_1097,N_1199);
nand U2159 (N_2159,N_1584,N_1360);
nand U2160 (N_2160,N_1222,N_1954);
or U2161 (N_2161,N_1025,N_1181);
nand U2162 (N_2162,N_1618,N_1084);
and U2163 (N_2163,N_1509,N_1158);
xor U2164 (N_2164,N_1241,N_1271);
nand U2165 (N_2165,N_1777,N_1341);
and U2166 (N_2166,N_1318,N_1548);
xor U2167 (N_2167,N_1370,N_1393);
or U2168 (N_2168,N_1062,N_1362);
xor U2169 (N_2169,N_1262,N_1162);
and U2170 (N_2170,N_1841,N_1078);
xor U2171 (N_2171,N_1944,N_1877);
and U2172 (N_2172,N_1032,N_1553);
and U2173 (N_2173,N_1144,N_1934);
xnor U2174 (N_2174,N_1328,N_1686);
and U2175 (N_2175,N_1340,N_1782);
or U2176 (N_2176,N_1668,N_1554);
xnor U2177 (N_2177,N_1367,N_1753);
nor U2178 (N_2178,N_1596,N_1613);
nor U2179 (N_2179,N_1762,N_1131);
or U2180 (N_2180,N_1225,N_1531);
and U2181 (N_2181,N_1558,N_1103);
xnor U2182 (N_2182,N_1856,N_1176);
or U2183 (N_2183,N_1170,N_1015);
nand U2184 (N_2184,N_1828,N_1996);
and U2185 (N_2185,N_1296,N_1590);
xnor U2186 (N_2186,N_1094,N_1420);
xnor U2187 (N_2187,N_1407,N_1449);
xnor U2188 (N_2188,N_1184,N_1681);
xnor U2189 (N_2189,N_1005,N_1342);
xnor U2190 (N_2190,N_1861,N_1141);
and U2191 (N_2191,N_1101,N_1178);
or U2192 (N_2192,N_1765,N_1775);
nor U2193 (N_2193,N_1807,N_1724);
nor U2194 (N_2194,N_1692,N_1766);
nand U2195 (N_2195,N_1445,N_1453);
or U2196 (N_2196,N_1574,N_1801);
and U2197 (N_2197,N_1266,N_1256);
or U2198 (N_2198,N_1893,N_1086);
and U2199 (N_2199,N_1477,N_1243);
nor U2200 (N_2200,N_1577,N_1234);
and U2201 (N_2201,N_1920,N_1608);
or U2202 (N_2202,N_1592,N_1145);
and U2203 (N_2203,N_1924,N_1786);
and U2204 (N_2204,N_1174,N_1146);
nor U2205 (N_2205,N_1418,N_1329);
and U2206 (N_2206,N_1869,N_1544);
or U2207 (N_2207,N_1047,N_1325);
xnor U2208 (N_2208,N_1835,N_1923);
nor U2209 (N_2209,N_1310,N_1665);
and U2210 (N_2210,N_1963,N_1175);
or U2211 (N_2211,N_1791,N_1642);
xor U2212 (N_2212,N_1708,N_1130);
xor U2213 (N_2213,N_1941,N_1147);
xnor U2214 (N_2214,N_1582,N_1441);
nor U2215 (N_2215,N_1994,N_1488);
nor U2216 (N_2216,N_1227,N_1230);
nand U2217 (N_2217,N_1513,N_1404);
nand U2218 (N_2218,N_1579,N_1463);
nand U2219 (N_2219,N_1236,N_1961);
and U2220 (N_2220,N_1087,N_1764);
nand U2221 (N_2221,N_1287,N_1859);
and U2222 (N_2222,N_1867,N_1055);
xnor U2223 (N_2223,N_1609,N_1945);
nor U2224 (N_2224,N_1043,N_1539);
nor U2225 (N_2225,N_1568,N_1625);
xor U2226 (N_2226,N_1051,N_1930);
or U2227 (N_2227,N_1357,N_1494);
nor U2228 (N_2228,N_1007,N_1771);
and U2229 (N_2229,N_1585,N_1414);
nand U2230 (N_2230,N_1213,N_1575);
nor U2231 (N_2231,N_1396,N_1070);
nor U2232 (N_2232,N_1825,N_1981);
nor U2233 (N_2233,N_1067,N_1167);
xnor U2234 (N_2234,N_1359,N_1200);
nand U2235 (N_2235,N_1538,N_1854);
xnor U2236 (N_2236,N_1848,N_1593);
or U2237 (N_2237,N_1884,N_1815);
nor U2238 (N_2238,N_1004,N_1770);
and U2239 (N_2239,N_1464,N_1126);
and U2240 (N_2240,N_1626,N_1334);
nand U2241 (N_2241,N_1743,N_1014);
nand U2242 (N_2242,N_1474,N_1267);
and U2243 (N_2243,N_1428,N_1982);
or U2244 (N_2244,N_1863,N_1470);
nor U2245 (N_2245,N_1832,N_1508);
nand U2246 (N_2246,N_1218,N_1030);
and U2247 (N_2247,N_1068,N_1189);
and U2248 (N_2248,N_1674,N_1567);
and U2249 (N_2249,N_1392,N_1431);
or U2250 (N_2250,N_1459,N_1177);
or U2251 (N_2251,N_1957,N_1768);
nor U2252 (N_2252,N_1604,N_1953);
nor U2253 (N_2253,N_1346,N_1466);
and U2254 (N_2254,N_1605,N_1781);
nor U2255 (N_2255,N_1154,N_1080);
nor U2256 (N_2256,N_1425,N_1614);
xnor U2257 (N_2257,N_1966,N_1458);
and U2258 (N_2258,N_1203,N_1896);
nand U2259 (N_2259,N_1335,N_1519);
and U2260 (N_2260,N_1368,N_1651);
and U2261 (N_2261,N_1207,N_1473);
nand U2262 (N_2262,N_1209,N_1956);
xor U2263 (N_2263,N_1525,N_1135);
nand U2264 (N_2264,N_1808,N_1796);
and U2265 (N_2265,N_1839,N_1695);
and U2266 (N_2266,N_1003,N_1074);
xnor U2267 (N_2267,N_1416,N_1487);
or U2268 (N_2268,N_1529,N_1294);
nand U2269 (N_2269,N_1688,N_1075);
nand U2270 (N_2270,N_1006,N_1444);
and U2271 (N_2271,N_1417,N_1333);
and U2272 (N_2272,N_1217,N_1499);
xnor U2273 (N_2273,N_1083,N_1430);
nand U2274 (N_2274,N_1639,N_1228);
xor U2275 (N_2275,N_1161,N_1833);
or U2276 (N_2276,N_1942,N_1514);
or U2277 (N_2277,N_1497,N_1366);
or U2278 (N_2278,N_1889,N_1033);
nand U2279 (N_2279,N_1017,N_1129);
or U2280 (N_2280,N_1725,N_1330);
nor U2281 (N_2281,N_1125,N_1429);
and U2282 (N_2282,N_1951,N_1769);
or U2283 (N_2283,N_1011,N_1442);
nor U2284 (N_2284,N_1423,N_1857);
or U2285 (N_2285,N_1536,N_1198);
or U2286 (N_2286,N_1255,N_1398);
nor U2287 (N_2287,N_1274,N_1064);
xor U2288 (N_2288,N_1288,N_1785);
nor U2289 (N_2289,N_1685,N_1649);
nor U2290 (N_2290,N_1697,N_1572);
xor U2291 (N_2291,N_1293,N_1565);
nor U2292 (N_2292,N_1027,N_1745);
nor U2293 (N_2293,N_1646,N_1165);
nor U2294 (N_2294,N_1631,N_1111);
nand U2295 (N_2295,N_1873,N_1472);
nor U2296 (N_2296,N_1820,N_1818);
or U2297 (N_2297,N_1270,N_1059);
nor U2298 (N_2298,N_1019,N_1395);
and U2299 (N_2299,N_1837,N_1875);
or U2300 (N_2300,N_1195,N_1540);
or U2301 (N_2301,N_1252,N_1804);
nand U2302 (N_2302,N_1057,N_1986);
nor U2303 (N_2303,N_1844,N_1372);
nor U2304 (N_2304,N_1810,N_1749);
and U2305 (N_2305,N_1399,N_1250);
and U2306 (N_2306,N_1573,N_1779);
and U2307 (N_2307,N_1504,N_1363);
nand U2308 (N_2308,N_1510,N_1433);
or U2309 (N_2309,N_1042,N_1226);
and U2310 (N_2310,N_1321,N_1788);
nand U2311 (N_2311,N_1373,N_1557);
nor U2312 (N_2312,N_1085,N_1286);
xor U2313 (N_2313,N_1113,N_1789);
nor U2314 (N_2314,N_1169,N_1092);
nand U2315 (N_2315,N_1273,N_1386);
nand U2316 (N_2316,N_1846,N_1371);
and U2317 (N_2317,N_1899,N_1010);
or U2318 (N_2318,N_1259,N_1784);
or U2319 (N_2319,N_1589,N_1940);
nand U2320 (N_2320,N_1853,N_1349);
nand U2321 (N_2321,N_1728,N_1720);
and U2322 (N_2322,N_1871,N_1840);
xnor U2323 (N_2323,N_1380,N_1800);
nand U2324 (N_2324,N_1284,N_1903);
or U2325 (N_2325,N_1327,N_1707);
nor U2326 (N_2326,N_1955,N_1677);
xor U2327 (N_2327,N_1615,N_1397);
and U2328 (N_2328,N_1928,N_1633);
xor U2329 (N_2329,N_1718,N_1647);
nor U2330 (N_2330,N_1502,N_1505);
xnor U2331 (N_2331,N_1495,N_1201);
or U2332 (N_2332,N_1090,N_1847);
and U2333 (N_2333,N_1238,N_1192);
or U2334 (N_2334,N_1975,N_1741);
xor U2335 (N_2335,N_1492,N_1036);
nand U2336 (N_2336,N_1115,N_1411);
and U2337 (N_2337,N_1755,N_1949);
nand U2338 (N_2338,N_1242,N_1948);
nor U2339 (N_2339,N_1021,N_1316);
or U2340 (N_2340,N_1232,N_1281);
and U2341 (N_2341,N_1673,N_1754);
and U2342 (N_2342,N_1384,N_1031);
xor U2343 (N_2343,N_1763,N_1727);
or U2344 (N_2344,N_1799,N_1308);
xnor U2345 (N_2345,N_1679,N_1123);
xnor U2346 (N_2346,N_1750,N_1206);
xor U2347 (N_2347,N_1402,N_1434);
and U2348 (N_2348,N_1046,N_1077);
nor U2349 (N_2349,N_1440,N_1439);
xor U2350 (N_2350,N_1298,N_1469);
xnor U2351 (N_2351,N_1410,N_1564);
xor U2352 (N_2352,N_1683,N_1684);
nand U2353 (N_2353,N_1845,N_1587);
and U2354 (N_2354,N_1312,N_1100);
nor U2355 (N_2355,N_1793,N_1352);
and U2356 (N_2356,N_1282,N_1211);
nand U2357 (N_2357,N_1566,N_1424);
xnor U2358 (N_2358,N_1438,N_1116);
or U2359 (N_2359,N_1151,N_1049);
nor U2360 (N_2360,N_1140,N_1619);
nor U2361 (N_2361,N_1486,N_1026);
xor U2362 (N_2362,N_1063,N_1148);
and U2363 (N_2363,N_1965,N_1627);
nand U2364 (N_2364,N_1850,N_1691);
and U2365 (N_2365,N_1805,N_1337);
or U2366 (N_2366,N_1524,N_1803);
nor U2367 (N_2367,N_1879,N_1937);
or U2368 (N_2368,N_1946,N_1114);
or U2369 (N_2369,N_1315,N_1813);
or U2370 (N_2370,N_1156,N_1598);
nand U2371 (N_2371,N_1868,N_1365);
or U2372 (N_2372,N_1670,N_1105);
and U2373 (N_2373,N_1012,N_1515);
or U2374 (N_2374,N_1630,N_1911);
and U2375 (N_2375,N_1422,N_1883);
nor U2376 (N_2376,N_1490,N_1710);
nor U2377 (N_2377,N_1932,N_1471);
nor U2378 (N_2378,N_1822,N_1299);
nand U2379 (N_2379,N_1675,N_1263);
xnor U2380 (N_2380,N_1375,N_1740);
xnor U2381 (N_2381,N_1780,N_1237);
nand U2382 (N_2382,N_1783,N_1595);
nor U2383 (N_2383,N_1164,N_1653);
and U2384 (N_2384,N_1778,N_1733);
or U2385 (N_2385,N_1197,N_1136);
xnor U2386 (N_2386,N_1581,N_1995);
nor U2387 (N_2387,N_1149,N_1343);
nor U2388 (N_2388,N_1645,N_1881);
or U2389 (N_2389,N_1772,N_1187);
nand U2390 (N_2390,N_1221,N_1152);
nand U2391 (N_2391,N_1559,N_1351);
xor U2392 (N_2392,N_1344,N_1050);
xor U2393 (N_2393,N_1454,N_1603);
and U2394 (N_2394,N_1607,N_1391);
nand U2395 (N_2395,N_1663,N_1610);
xor U2396 (N_2396,N_1354,N_1977);
nor U2397 (N_2397,N_1909,N_1338);
and U2398 (N_2398,N_1620,N_1521);
nand U2399 (N_2399,N_1512,N_1053);
and U2400 (N_2400,N_1073,N_1758);
nor U2401 (N_2401,N_1925,N_1523);
or U2402 (N_2402,N_1929,N_1518);
xor U2403 (N_2403,N_1640,N_1364);
and U2404 (N_2404,N_1742,N_1305);
xnor U2405 (N_2405,N_1950,N_1223);
xnor U2406 (N_2406,N_1730,N_1759);
xor U2407 (N_2407,N_1456,N_1214);
nor U2408 (N_2408,N_1931,N_1972);
and U2409 (N_2409,N_1938,N_1143);
and U2410 (N_2410,N_1687,N_1795);
and U2411 (N_2411,N_1882,N_1448);
and U2412 (N_2412,N_1326,N_1578);
xor U2413 (N_2413,N_1066,N_1922);
xor U2414 (N_2414,N_1278,N_1215);
nor U2415 (N_2415,N_1482,N_1522);
or U2416 (N_2416,N_1622,N_1546);
or U2417 (N_2417,N_1959,N_1973);
xnor U2418 (N_2418,N_1731,N_1829);
nand U2419 (N_2419,N_1096,N_1253);
xor U2420 (N_2420,N_1694,N_1926);
and U2421 (N_2421,N_1978,N_1814);
and U2422 (N_2422,N_1666,N_1586);
and U2423 (N_2423,N_1137,N_1060);
or U2424 (N_2424,N_1193,N_1752);
xor U2425 (N_2425,N_1350,N_1726);
and U2426 (N_2426,N_1676,N_1849);
xnor U2427 (N_2427,N_1851,N_1229);
nand U2428 (N_2428,N_1936,N_1106);
xor U2429 (N_2429,N_1044,N_1379);
or U2430 (N_2430,N_1022,N_1098);
nand U2431 (N_2431,N_1898,N_1821);
and U2432 (N_2432,N_1865,N_1412);
nand U2433 (N_2433,N_1797,N_1773);
nor U2434 (N_2434,N_1072,N_1387);
xor U2435 (N_2435,N_1127,N_1212);
and U2436 (N_2436,N_1838,N_1669);
xor U2437 (N_2437,N_1048,N_1637);
nor U2438 (N_2438,N_1001,N_1667);
nor U2439 (N_2439,N_1776,N_1054);
nand U2440 (N_2440,N_1091,N_1552);
nand U2441 (N_2441,N_1993,N_1319);
nand U2442 (N_2442,N_1037,N_1000);
and U2443 (N_2443,N_1897,N_1591);
or U2444 (N_2444,N_1038,N_1757);
nor U2445 (N_2445,N_1188,N_1254);
nand U2446 (N_2446,N_1569,N_1709);
xor U2447 (N_2447,N_1918,N_1435);
nor U2448 (N_2448,N_1964,N_1571);
and U2449 (N_2449,N_1302,N_1616);
nand U2450 (N_2450,N_1507,N_1735);
xor U2451 (N_2451,N_1652,N_1910);
and U2452 (N_2452,N_1132,N_1382);
or U2453 (N_2453,N_1231,N_1385);
or U2454 (N_2454,N_1962,N_1336);
or U2455 (N_2455,N_1381,N_1475);
and U2456 (N_2456,N_1322,N_1081);
or U2457 (N_2457,N_1734,N_1812);
nor U2458 (N_2458,N_1489,N_1292);
nand U2459 (N_2459,N_1479,N_1737);
xnor U2460 (N_2460,N_1450,N_1704);
or U2461 (N_2461,N_1109,N_1313);
nand U2462 (N_2462,N_1744,N_1560);
or U2463 (N_2463,N_1960,N_1261);
and U2464 (N_2464,N_1157,N_1159);
nand U2465 (N_2465,N_1549,N_1139);
xnor U2466 (N_2466,N_1794,N_1712);
nor U2467 (N_2467,N_1204,N_1792);
xor U2468 (N_2468,N_1339,N_1943);
xor U2469 (N_2469,N_1437,N_1747);
and U2470 (N_2470,N_1290,N_1244);
nand U2471 (N_2471,N_1900,N_1016);
nor U2472 (N_2472,N_1872,N_1894);
and U2473 (N_2473,N_1576,N_1706);
nand U2474 (N_2474,N_1824,N_1756);
nor U2475 (N_2475,N_1678,N_1887);
or U2476 (N_2476,N_1919,N_1013);
nor U2477 (N_2477,N_1247,N_1542);
xor U2478 (N_2478,N_1947,N_1361);
nand U2479 (N_2479,N_1056,N_1988);
nor U2480 (N_2480,N_1480,N_1886);
or U2481 (N_2481,N_1774,N_1705);
xnor U2482 (N_2482,N_1939,N_1028);
xor U2483 (N_2483,N_1279,N_1260);
or U2484 (N_2484,N_1356,N_1700);
xnor U2485 (N_2485,N_1405,N_1806);
nand U2486 (N_2486,N_1690,N_1671);
nor U2487 (N_2487,N_1024,N_1347);
xnor U2488 (N_2488,N_1761,N_1002);
xor U2489 (N_2489,N_1180,N_1588);
nand U2490 (N_2490,N_1629,N_1732);
or U2491 (N_2491,N_1065,N_1190);
xor U2492 (N_2492,N_1265,N_1353);
nand U2493 (N_2493,N_1426,N_1662);
or U2494 (N_2494,N_1644,N_1661);
or U2495 (N_2495,N_1389,N_1332);
or U2496 (N_2496,N_1746,N_1251);
nand U2497 (N_2497,N_1045,N_1891);
nand U2498 (N_2498,N_1843,N_1638);
xor U2499 (N_2499,N_1183,N_1240);
xnor U2500 (N_2500,N_1131,N_1782);
nor U2501 (N_2501,N_1447,N_1200);
or U2502 (N_2502,N_1053,N_1944);
and U2503 (N_2503,N_1167,N_1633);
nor U2504 (N_2504,N_1817,N_1223);
and U2505 (N_2505,N_1400,N_1183);
nor U2506 (N_2506,N_1177,N_1654);
nor U2507 (N_2507,N_1592,N_1953);
and U2508 (N_2508,N_1680,N_1253);
xnor U2509 (N_2509,N_1993,N_1317);
nor U2510 (N_2510,N_1239,N_1606);
nand U2511 (N_2511,N_1563,N_1140);
xnor U2512 (N_2512,N_1424,N_1168);
and U2513 (N_2513,N_1855,N_1980);
nand U2514 (N_2514,N_1396,N_1259);
nor U2515 (N_2515,N_1355,N_1505);
nor U2516 (N_2516,N_1425,N_1865);
nor U2517 (N_2517,N_1124,N_1851);
or U2518 (N_2518,N_1004,N_1059);
and U2519 (N_2519,N_1979,N_1805);
nor U2520 (N_2520,N_1668,N_1889);
or U2521 (N_2521,N_1120,N_1682);
nand U2522 (N_2522,N_1237,N_1531);
nor U2523 (N_2523,N_1464,N_1595);
xnor U2524 (N_2524,N_1515,N_1603);
nor U2525 (N_2525,N_1563,N_1440);
xor U2526 (N_2526,N_1642,N_1606);
xnor U2527 (N_2527,N_1704,N_1958);
or U2528 (N_2528,N_1267,N_1909);
and U2529 (N_2529,N_1578,N_1097);
xor U2530 (N_2530,N_1916,N_1228);
or U2531 (N_2531,N_1389,N_1385);
xnor U2532 (N_2532,N_1641,N_1223);
nand U2533 (N_2533,N_1717,N_1826);
or U2534 (N_2534,N_1213,N_1292);
nor U2535 (N_2535,N_1644,N_1819);
xnor U2536 (N_2536,N_1314,N_1945);
or U2537 (N_2537,N_1560,N_1218);
and U2538 (N_2538,N_1418,N_1786);
nor U2539 (N_2539,N_1781,N_1132);
or U2540 (N_2540,N_1100,N_1317);
xnor U2541 (N_2541,N_1832,N_1019);
and U2542 (N_2542,N_1890,N_1985);
and U2543 (N_2543,N_1905,N_1676);
xnor U2544 (N_2544,N_1470,N_1860);
nor U2545 (N_2545,N_1357,N_1410);
nor U2546 (N_2546,N_1543,N_1997);
nand U2547 (N_2547,N_1139,N_1961);
or U2548 (N_2548,N_1145,N_1762);
nor U2549 (N_2549,N_1399,N_1021);
nor U2550 (N_2550,N_1729,N_1021);
nor U2551 (N_2551,N_1912,N_1351);
xor U2552 (N_2552,N_1704,N_1273);
xnor U2553 (N_2553,N_1702,N_1483);
nor U2554 (N_2554,N_1288,N_1647);
and U2555 (N_2555,N_1321,N_1378);
and U2556 (N_2556,N_1938,N_1348);
or U2557 (N_2557,N_1120,N_1487);
nor U2558 (N_2558,N_1748,N_1079);
nor U2559 (N_2559,N_1060,N_1582);
or U2560 (N_2560,N_1121,N_1408);
or U2561 (N_2561,N_1428,N_1766);
nor U2562 (N_2562,N_1671,N_1356);
and U2563 (N_2563,N_1977,N_1386);
nor U2564 (N_2564,N_1767,N_1858);
nand U2565 (N_2565,N_1301,N_1398);
xor U2566 (N_2566,N_1905,N_1242);
nand U2567 (N_2567,N_1754,N_1894);
nor U2568 (N_2568,N_1326,N_1334);
or U2569 (N_2569,N_1118,N_1126);
nor U2570 (N_2570,N_1465,N_1346);
and U2571 (N_2571,N_1983,N_1903);
nand U2572 (N_2572,N_1416,N_1780);
nor U2573 (N_2573,N_1983,N_1289);
xor U2574 (N_2574,N_1659,N_1922);
and U2575 (N_2575,N_1714,N_1437);
nand U2576 (N_2576,N_1437,N_1019);
nor U2577 (N_2577,N_1061,N_1320);
xnor U2578 (N_2578,N_1209,N_1142);
nand U2579 (N_2579,N_1709,N_1975);
nor U2580 (N_2580,N_1370,N_1556);
and U2581 (N_2581,N_1789,N_1414);
nand U2582 (N_2582,N_1391,N_1903);
and U2583 (N_2583,N_1354,N_1686);
nor U2584 (N_2584,N_1325,N_1007);
and U2585 (N_2585,N_1624,N_1550);
nand U2586 (N_2586,N_1065,N_1982);
xor U2587 (N_2587,N_1920,N_1830);
nor U2588 (N_2588,N_1514,N_1611);
nand U2589 (N_2589,N_1727,N_1136);
nor U2590 (N_2590,N_1375,N_1968);
xnor U2591 (N_2591,N_1419,N_1132);
nor U2592 (N_2592,N_1549,N_1401);
nor U2593 (N_2593,N_1151,N_1394);
and U2594 (N_2594,N_1623,N_1857);
or U2595 (N_2595,N_1026,N_1067);
nor U2596 (N_2596,N_1132,N_1043);
nor U2597 (N_2597,N_1151,N_1986);
and U2598 (N_2598,N_1870,N_1150);
xnor U2599 (N_2599,N_1029,N_1354);
nand U2600 (N_2600,N_1557,N_1628);
xor U2601 (N_2601,N_1814,N_1316);
and U2602 (N_2602,N_1918,N_1275);
nor U2603 (N_2603,N_1522,N_1929);
xor U2604 (N_2604,N_1496,N_1230);
and U2605 (N_2605,N_1299,N_1107);
or U2606 (N_2606,N_1376,N_1541);
xnor U2607 (N_2607,N_1612,N_1817);
nand U2608 (N_2608,N_1941,N_1505);
and U2609 (N_2609,N_1398,N_1147);
nand U2610 (N_2610,N_1412,N_1551);
or U2611 (N_2611,N_1963,N_1265);
nand U2612 (N_2612,N_1591,N_1581);
or U2613 (N_2613,N_1966,N_1435);
nor U2614 (N_2614,N_1109,N_1900);
xnor U2615 (N_2615,N_1354,N_1662);
or U2616 (N_2616,N_1127,N_1517);
nand U2617 (N_2617,N_1198,N_1690);
nor U2618 (N_2618,N_1189,N_1399);
nand U2619 (N_2619,N_1558,N_1995);
and U2620 (N_2620,N_1340,N_1698);
xnor U2621 (N_2621,N_1170,N_1273);
nor U2622 (N_2622,N_1110,N_1126);
nor U2623 (N_2623,N_1767,N_1722);
nand U2624 (N_2624,N_1986,N_1414);
xnor U2625 (N_2625,N_1210,N_1329);
and U2626 (N_2626,N_1392,N_1843);
xor U2627 (N_2627,N_1187,N_1126);
or U2628 (N_2628,N_1932,N_1057);
or U2629 (N_2629,N_1601,N_1481);
nand U2630 (N_2630,N_1754,N_1865);
nor U2631 (N_2631,N_1180,N_1894);
and U2632 (N_2632,N_1699,N_1018);
xor U2633 (N_2633,N_1648,N_1117);
nand U2634 (N_2634,N_1560,N_1430);
nor U2635 (N_2635,N_1419,N_1521);
or U2636 (N_2636,N_1347,N_1608);
or U2637 (N_2637,N_1595,N_1800);
or U2638 (N_2638,N_1569,N_1694);
and U2639 (N_2639,N_1164,N_1010);
nand U2640 (N_2640,N_1371,N_1945);
nand U2641 (N_2641,N_1964,N_1978);
nand U2642 (N_2642,N_1117,N_1517);
nand U2643 (N_2643,N_1448,N_1254);
or U2644 (N_2644,N_1629,N_1970);
and U2645 (N_2645,N_1897,N_1974);
nor U2646 (N_2646,N_1152,N_1783);
or U2647 (N_2647,N_1611,N_1674);
and U2648 (N_2648,N_1052,N_1330);
or U2649 (N_2649,N_1372,N_1159);
xor U2650 (N_2650,N_1104,N_1212);
or U2651 (N_2651,N_1673,N_1785);
nand U2652 (N_2652,N_1157,N_1809);
xnor U2653 (N_2653,N_1037,N_1170);
nand U2654 (N_2654,N_1293,N_1499);
xnor U2655 (N_2655,N_1042,N_1965);
xor U2656 (N_2656,N_1642,N_1623);
and U2657 (N_2657,N_1526,N_1834);
nand U2658 (N_2658,N_1184,N_1947);
or U2659 (N_2659,N_1856,N_1356);
nand U2660 (N_2660,N_1443,N_1108);
and U2661 (N_2661,N_1671,N_1777);
or U2662 (N_2662,N_1870,N_1784);
xor U2663 (N_2663,N_1345,N_1530);
nor U2664 (N_2664,N_1895,N_1442);
xor U2665 (N_2665,N_1038,N_1953);
xor U2666 (N_2666,N_1672,N_1004);
and U2667 (N_2667,N_1510,N_1472);
and U2668 (N_2668,N_1236,N_1546);
or U2669 (N_2669,N_1533,N_1374);
xor U2670 (N_2670,N_1856,N_1302);
or U2671 (N_2671,N_1330,N_1655);
nor U2672 (N_2672,N_1782,N_1593);
and U2673 (N_2673,N_1642,N_1150);
nand U2674 (N_2674,N_1686,N_1334);
or U2675 (N_2675,N_1672,N_1278);
nor U2676 (N_2676,N_1336,N_1420);
nor U2677 (N_2677,N_1233,N_1625);
nand U2678 (N_2678,N_1012,N_1771);
or U2679 (N_2679,N_1340,N_1973);
nand U2680 (N_2680,N_1049,N_1404);
xnor U2681 (N_2681,N_1453,N_1597);
or U2682 (N_2682,N_1698,N_1830);
or U2683 (N_2683,N_1834,N_1593);
nand U2684 (N_2684,N_1312,N_1274);
xor U2685 (N_2685,N_1104,N_1381);
nor U2686 (N_2686,N_1213,N_1429);
and U2687 (N_2687,N_1416,N_1833);
and U2688 (N_2688,N_1050,N_1790);
and U2689 (N_2689,N_1913,N_1530);
nor U2690 (N_2690,N_1867,N_1834);
or U2691 (N_2691,N_1664,N_1834);
xnor U2692 (N_2692,N_1036,N_1507);
and U2693 (N_2693,N_1784,N_1438);
or U2694 (N_2694,N_1904,N_1355);
and U2695 (N_2695,N_1547,N_1769);
or U2696 (N_2696,N_1633,N_1512);
nand U2697 (N_2697,N_1043,N_1897);
nor U2698 (N_2698,N_1150,N_1167);
nand U2699 (N_2699,N_1567,N_1457);
nand U2700 (N_2700,N_1805,N_1354);
nand U2701 (N_2701,N_1449,N_1923);
nor U2702 (N_2702,N_1075,N_1237);
and U2703 (N_2703,N_1783,N_1752);
nor U2704 (N_2704,N_1210,N_1604);
xnor U2705 (N_2705,N_1893,N_1635);
xor U2706 (N_2706,N_1518,N_1631);
or U2707 (N_2707,N_1358,N_1412);
or U2708 (N_2708,N_1490,N_1763);
and U2709 (N_2709,N_1804,N_1449);
or U2710 (N_2710,N_1201,N_1002);
nand U2711 (N_2711,N_1272,N_1433);
xnor U2712 (N_2712,N_1520,N_1608);
or U2713 (N_2713,N_1572,N_1248);
xor U2714 (N_2714,N_1289,N_1058);
xor U2715 (N_2715,N_1575,N_1814);
nand U2716 (N_2716,N_1663,N_1519);
xor U2717 (N_2717,N_1101,N_1705);
or U2718 (N_2718,N_1054,N_1518);
or U2719 (N_2719,N_1749,N_1125);
and U2720 (N_2720,N_1616,N_1536);
and U2721 (N_2721,N_1078,N_1060);
nor U2722 (N_2722,N_1862,N_1667);
xnor U2723 (N_2723,N_1099,N_1401);
nand U2724 (N_2724,N_1529,N_1611);
nor U2725 (N_2725,N_1512,N_1934);
and U2726 (N_2726,N_1259,N_1573);
or U2727 (N_2727,N_1129,N_1881);
nand U2728 (N_2728,N_1270,N_1368);
and U2729 (N_2729,N_1746,N_1828);
and U2730 (N_2730,N_1472,N_1816);
and U2731 (N_2731,N_1819,N_1768);
nor U2732 (N_2732,N_1192,N_1374);
nor U2733 (N_2733,N_1569,N_1062);
nand U2734 (N_2734,N_1736,N_1160);
nor U2735 (N_2735,N_1315,N_1631);
and U2736 (N_2736,N_1886,N_1569);
or U2737 (N_2737,N_1377,N_1371);
nand U2738 (N_2738,N_1982,N_1189);
xor U2739 (N_2739,N_1089,N_1394);
and U2740 (N_2740,N_1694,N_1376);
nand U2741 (N_2741,N_1836,N_1455);
nand U2742 (N_2742,N_1546,N_1835);
and U2743 (N_2743,N_1607,N_1331);
and U2744 (N_2744,N_1376,N_1125);
nand U2745 (N_2745,N_1522,N_1484);
xnor U2746 (N_2746,N_1752,N_1498);
and U2747 (N_2747,N_1411,N_1573);
nand U2748 (N_2748,N_1755,N_1406);
or U2749 (N_2749,N_1482,N_1644);
nand U2750 (N_2750,N_1909,N_1221);
nand U2751 (N_2751,N_1582,N_1244);
xor U2752 (N_2752,N_1355,N_1459);
nor U2753 (N_2753,N_1027,N_1870);
and U2754 (N_2754,N_1416,N_1862);
nand U2755 (N_2755,N_1052,N_1405);
and U2756 (N_2756,N_1326,N_1792);
nand U2757 (N_2757,N_1028,N_1822);
nor U2758 (N_2758,N_1029,N_1300);
and U2759 (N_2759,N_1153,N_1457);
nor U2760 (N_2760,N_1475,N_1875);
nand U2761 (N_2761,N_1311,N_1158);
or U2762 (N_2762,N_1699,N_1306);
or U2763 (N_2763,N_1994,N_1154);
nor U2764 (N_2764,N_1092,N_1921);
nor U2765 (N_2765,N_1237,N_1688);
nor U2766 (N_2766,N_1026,N_1248);
nand U2767 (N_2767,N_1622,N_1534);
xor U2768 (N_2768,N_1433,N_1888);
and U2769 (N_2769,N_1315,N_1024);
xor U2770 (N_2770,N_1100,N_1739);
xor U2771 (N_2771,N_1921,N_1980);
nor U2772 (N_2772,N_1823,N_1144);
xor U2773 (N_2773,N_1571,N_1923);
nor U2774 (N_2774,N_1522,N_1449);
nor U2775 (N_2775,N_1128,N_1925);
or U2776 (N_2776,N_1224,N_1035);
and U2777 (N_2777,N_1681,N_1134);
xor U2778 (N_2778,N_1108,N_1095);
nor U2779 (N_2779,N_1264,N_1648);
nor U2780 (N_2780,N_1497,N_1200);
xnor U2781 (N_2781,N_1321,N_1178);
nor U2782 (N_2782,N_1500,N_1656);
nand U2783 (N_2783,N_1407,N_1735);
nor U2784 (N_2784,N_1092,N_1026);
nor U2785 (N_2785,N_1131,N_1237);
xor U2786 (N_2786,N_1754,N_1264);
or U2787 (N_2787,N_1061,N_1130);
nor U2788 (N_2788,N_1112,N_1056);
or U2789 (N_2789,N_1029,N_1979);
nand U2790 (N_2790,N_1567,N_1550);
nor U2791 (N_2791,N_1717,N_1660);
and U2792 (N_2792,N_1407,N_1606);
nor U2793 (N_2793,N_1903,N_1695);
nor U2794 (N_2794,N_1481,N_1340);
nand U2795 (N_2795,N_1454,N_1600);
nor U2796 (N_2796,N_1119,N_1197);
and U2797 (N_2797,N_1941,N_1419);
nand U2798 (N_2798,N_1278,N_1255);
and U2799 (N_2799,N_1107,N_1377);
nand U2800 (N_2800,N_1879,N_1966);
and U2801 (N_2801,N_1505,N_1086);
xnor U2802 (N_2802,N_1950,N_1715);
and U2803 (N_2803,N_1365,N_1058);
nand U2804 (N_2804,N_1520,N_1226);
and U2805 (N_2805,N_1647,N_1907);
nand U2806 (N_2806,N_1031,N_1406);
or U2807 (N_2807,N_1272,N_1606);
or U2808 (N_2808,N_1018,N_1172);
nor U2809 (N_2809,N_1220,N_1617);
nand U2810 (N_2810,N_1521,N_1889);
nor U2811 (N_2811,N_1990,N_1590);
or U2812 (N_2812,N_1117,N_1416);
nor U2813 (N_2813,N_1961,N_1037);
nor U2814 (N_2814,N_1929,N_1927);
nor U2815 (N_2815,N_1147,N_1716);
and U2816 (N_2816,N_1326,N_1194);
nand U2817 (N_2817,N_1714,N_1192);
or U2818 (N_2818,N_1467,N_1200);
xor U2819 (N_2819,N_1807,N_1778);
or U2820 (N_2820,N_1830,N_1204);
nor U2821 (N_2821,N_1155,N_1857);
and U2822 (N_2822,N_1830,N_1245);
or U2823 (N_2823,N_1068,N_1635);
or U2824 (N_2824,N_1972,N_1164);
or U2825 (N_2825,N_1786,N_1561);
and U2826 (N_2826,N_1117,N_1027);
or U2827 (N_2827,N_1375,N_1486);
nor U2828 (N_2828,N_1162,N_1355);
and U2829 (N_2829,N_1280,N_1648);
or U2830 (N_2830,N_1659,N_1973);
and U2831 (N_2831,N_1197,N_1625);
nor U2832 (N_2832,N_1556,N_1889);
nand U2833 (N_2833,N_1718,N_1090);
or U2834 (N_2834,N_1171,N_1328);
nor U2835 (N_2835,N_1622,N_1735);
and U2836 (N_2836,N_1202,N_1676);
nand U2837 (N_2837,N_1900,N_1448);
nor U2838 (N_2838,N_1262,N_1963);
or U2839 (N_2839,N_1831,N_1676);
xnor U2840 (N_2840,N_1279,N_1577);
nand U2841 (N_2841,N_1671,N_1138);
and U2842 (N_2842,N_1056,N_1332);
nor U2843 (N_2843,N_1824,N_1540);
xnor U2844 (N_2844,N_1709,N_1291);
xor U2845 (N_2845,N_1831,N_1239);
or U2846 (N_2846,N_1478,N_1795);
and U2847 (N_2847,N_1869,N_1782);
or U2848 (N_2848,N_1101,N_1661);
nand U2849 (N_2849,N_1158,N_1405);
nor U2850 (N_2850,N_1295,N_1077);
nand U2851 (N_2851,N_1551,N_1432);
and U2852 (N_2852,N_1838,N_1945);
and U2853 (N_2853,N_1417,N_1700);
or U2854 (N_2854,N_1273,N_1598);
nand U2855 (N_2855,N_1597,N_1533);
nand U2856 (N_2856,N_1414,N_1775);
or U2857 (N_2857,N_1220,N_1124);
xor U2858 (N_2858,N_1235,N_1921);
xor U2859 (N_2859,N_1580,N_1227);
or U2860 (N_2860,N_1200,N_1705);
or U2861 (N_2861,N_1780,N_1877);
or U2862 (N_2862,N_1478,N_1407);
or U2863 (N_2863,N_1756,N_1358);
and U2864 (N_2864,N_1777,N_1572);
and U2865 (N_2865,N_1759,N_1475);
or U2866 (N_2866,N_1710,N_1429);
nor U2867 (N_2867,N_1850,N_1860);
nand U2868 (N_2868,N_1488,N_1814);
xor U2869 (N_2869,N_1204,N_1478);
xor U2870 (N_2870,N_1199,N_1000);
nand U2871 (N_2871,N_1659,N_1993);
and U2872 (N_2872,N_1667,N_1131);
xor U2873 (N_2873,N_1768,N_1424);
xor U2874 (N_2874,N_1593,N_1284);
or U2875 (N_2875,N_1304,N_1997);
nor U2876 (N_2876,N_1285,N_1492);
xor U2877 (N_2877,N_1021,N_1691);
and U2878 (N_2878,N_1377,N_1385);
nor U2879 (N_2879,N_1728,N_1037);
xor U2880 (N_2880,N_1761,N_1248);
or U2881 (N_2881,N_1144,N_1164);
nor U2882 (N_2882,N_1081,N_1471);
and U2883 (N_2883,N_1930,N_1293);
nand U2884 (N_2884,N_1308,N_1994);
nor U2885 (N_2885,N_1320,N_1093);
nor U2886 (N_2886,N_1093,N_1058);
nor U2887 (N_2887,N_1588,N_1100);
and U2888 (N_2888,N_1381,N_1641);
nor U2889 (N_2889,N_1513,N_1198);
nand U2890 (N_2890,N_1281,N_1084);
xor U2891 (N_2891,N_1359,N_1809);
or U2892 (N_2892,N_1319,N_1532);
or U2893 (N_2893,N_1436,N_1587);
xnor U2894 (N_2894,N_1497,N_1241);
xnor U2895 (N_2895,N_1186,N_1744);
xor U2896 (N_2896,N_1062,N_1179);
and U2897 (N_2897,N_1960,N_1466);
nor U2898 (N_2898,N_1525,N_1102);
nor U2899 (N_2899,N_1298,N_1562);
or U2900 (N_2900,N_1435,N_1164);
nand U2901 (N_2901,N_1042,N_1013);
or U2902 (N_2902,N_1475,N_1018);
or U2903 (N_2903,N_1629,N_1647);
xnor U2904 (N_2904,N_1153,N_1824);
or U2905 (N_2905,N_1142,N_1784);
nand U2906 (N_2906,N_1074,N_1341);
nand U2907 (N_2907,N_1195,N_1921);
xor U2908 (N_2908,N_1334,N_1299);
and U2909 (N_2909,N_1830,N_1260);
or U2910 (N_2910,N_1535,N_1839);
and U2911 (N_2911,N_1413,N_1046);
or U2912 (N_2912,N_1695,N_1658);
nand U2913 (N_2913,N_1030,N_1241);
nor U2914 (N_2914,N_1646,N_1865);
xnor U2915 (N_2915,N_1087,N_1938);
and U2916 (N_2916,N_1633,N_1905);
or U2917 (N_2917,N_1271,N_1208);
and U2918 (N_2918,N_1074,N_1271);
or U2919 (N_2919,N_1185,N_1458);
and U2920 (N_2920,N_1122,N_1811);
nor U2921 (N_2921,N_1271,N_1152);
nand U2922 (N_2922,N_1930,N_1269);
nor U2923 (N_2923,N_1800,N_1376);
nor U2924 (N_2924,N_1871,N_1670);
nor U2925 (N_2925,N_1813,N_1480);
and U2926 (N_2926,N_1830,N_1501);
and U2927 (N_2927,N_1598,N_1088);
or U2928 (N_2928,N_1501,N_1988);
and U2929 (N_2929,N_1995,N_1263);
and U2930 (N_2930,N_1911,N_1866);
xnor U2931 (N_2931,N_1982,N_1300);
xor U2932 (N_2932,N_1081,N_1314);
nand U2933 (N_2933,N_1644,N_1356);
nor U2934 (N_2934,N_1491,N_1818);
nand U2935 (N_2935,N_1577,N_1557);
xnor U2936 (N_2936,N_1758,N_1173);
and U2937 (N_2937,N_1616,N_1073);
and U2938 (N_2938,N_1122,N_1914);
or U2939 (N_2939,N_1715,N_1909);
or U2940 (N_2940,N_1918,N_1336);
nand U2941 (N_2941,N_1983,N_1740);
or U2942 (N_2942,N_1291,N_1814);
or U2943 (N_2943,N_1476,N_1402);
or U2944 (N_2944,N_1257,N_1288);
and U2945 (N_2945,N_1414,N_1935);
nand U2946 (N_2946,N_1438,N_1816);
nor U2947 (N_2947,N_1005,N_1133);
nand U2948 (N_2948,N_1440,N_1648);
nor U2949 (N_2949,N_1466,N_1385);
xnor U2950 (N_2950,N_1365,N_1718);
and U2951 (N_2951,N_1994,N_1066);
nand U2952 (N_2952,N_1991,N_1941);
nand U2953 (N_2953,N_1299,N_1523);
or U2954 (N_2954,N_1689,N_1026);
nor U2955 (N_2955,N_1643,N_1146);
nor U2956 (N_2956,N_1468,N_1483);
and U2957 (N_2957,N_1418,N_1945);
or U2958 (N_2958,N_1945,N_1094);
xor U2959 (N_2959,N_1437,N_1022);
and U2960 (N_2960,N_1572,N_1841);
or U2961 (N_2961,N_1093,N_1617);
xor U2962 (N_2962,N_1683,N_1812);
nand U2963 (N_2963,N_1408,N_1204);
nor U2964 (N_2964,N_1816,N_1130);
xnor U2965 (N_2965,N_1837,N_1546);
xnor U2966 (N_2966,N_1429,N_1177);
xnor U2967 (N_2967,N_1946,N_1629);
nor U2968 (N_2968,N_1183,N_1051);
and U2969 (N_2969,N_1262,N_1246);
nand U2970 (N_2970,N_1470,N_1400);
nor U2971 (N_2971,N_1715,N_1994);
nand U2972 (N_2972,N_1627,N_1438);
nor U2973 (N_2973,N_1325,N_1074);
or U2974 (N_2974,N_1829,N_1234);
nand U2975 (N_2975,N_1241,N_1128);
xnor U2976 (N_2976,N_1627,N_1964);
or U2977 (N_2977,N_1728,N_1619);
nor U2978 (N_2978,N_1974,N_1125);
or U2979 (N_2979,N_1239,N_1916);
or U2980 (N_2980,N_1240,N_1532);
nor U2981 (N_2981,N_1205,N_1688);
and U2982 (N_2982,N_1139,N_1244);
and U2983 (N_2983,N_1242,N_1779);
or U2984 (N_2984,N_1714,N_1760);
nor U2985 (N_2985,N_1957,N_1573);
or U2986 (N_2986,N_1657,N_1647);
nor U2987 (N_2987,N_1339,N_1768);
and U2988 (N_2988,N_1591,N_1985);
xor U2989 (N_2989,N_1084,N_1658);
nor U2990 (N_2990,N_1518,N_1378);
or U2991 (N_2991,N_1156,N_1513);
nor U2992 (N_2992,N_1533,N_1125);
xnor U2993 (N_2993,N_1441,N_1463);
nand U2994 (N_2994,N_1837,N_1435);
and U2995 (N_2995,N_1724,N_1836);
nand U2996 (N_2996,N_1809,N_1963);
nor U2997 (N_2997,N_1272,N_1826);
or U2998 (N_2998,N_1640,N_1297);
and U2999 (N_2999,N_1655,N_1389);
nor UO_0 (O_0,N_2018,N_2655);
or UO_1 (O_1,N_2036,N_2972);
nor UO_2 (O_2,N_2510,N_2785);
nand UO_3 (O_3,N_2563,N_2906);
or UO_4 (O_4,N_2685,N_2952);
xor UO_5 (O_5,N_2885,N_2632);
xor UO_6 (O_6,N_2545,N_2451);
xnor UO_7 (O_7,N_2198,N_2176);
xor UO_8 (O_8,N_2367,N_2079);
nor UO_9 (O_9,N_2365,N_2267);
or UO_10 (O_10,N_2852,N_2386);
xor UO_11 (O_11,N_2356,N_2435);
or UO_12 (O_12,N_2905,N_2440);
xnor UO_13 (O_13,N_2348,N_2431);
or UO_14 (O_14,N_2195,N_2851);
and UO_15 (O_15,N_2178,N_2713);
and UO_16 (O_16,N_2205,N_2962);
and UO_17 (O_17,N_2899,N_2313);
nand UO_18 (O_18,N_2489,N_2592);
nand UO_19 (O_19,N_2085,N_2555);
nor UO_20 (O_20,N_2997,N_2617);
xor UO_21 (O_21,N_2429,N_2032);
and UO_22 (O_22,N_2849,N_2056);
nand UO_23 (O_23,N_2068,N_2417);
and UO_24 (O_24,N_2770,N_2324);
nor UO_25 (O_25,N_2893,N_2017);
and UO_26 (O_26,N_2715,N_2779);
or UO_27 (O_27,N_2371,N_2477);
nor UO_28 (O_28,N_2109,N_2687);
nor UO_29 (O_29,N_2010,N_2019);
and UO_30 (O_30,N_2066,N_2347);
and UO_31 (O_31,N_2189,N_2642);
nor UO_32 (O_32,N_2524,N_2385);
and UO_33 (O_33,N_2171,N_2706);
nor UO_34 (O_34,N_2294,N_2239);
nand UO_35 (O_35,N_2262,N_2876);
nor UO_36 (O_36,N_2217,N_2160);
nand UO_37 (O_37,N_2305,N_2588);
nor UO_38 (O_38,N_2749,N_2880);
nand UO_39 (O_39,N_2208,N_2117);
or UO_40 (O_40,N_2874,N_2021);
nor UO_41 (O_41,N_2230,N_2135);
xor UO_42 (O_42,N_2025,N_2337);
or UO_43 (O_43,N_2145,N_2657);
xnor UO_44 (O_44,N_2140,N_2264);
nor UO_45 (O_45,N_2295,N_2218);
nor UO_46 (O_46,N_2686,N_2030);
or UO_47 (O_47,N_2043,N_2921);
nand UO_48 (O_48,N_2530,N_2232);
or UO_49 (O_49,N_2448,N_2710);
nand UO_50 (O_50,N_2711,N_2190);
nor UO_51 (O_51,N_2854,N_2001);
and UO_52 (O_52,N_2787,N_2833);
and UO_53 (O_53,N_2860,N_2727);
nor UO_54 (O_54,N_2257,N_2399);
nor UO_55 (O_55,N_2468,N_2151);
nor UO_56 (O_56,N_2863,N_2681);
and UO_57 (O_57,N_2006,N_2162);
nor UO_58 (O_58,N_2502,N_2842);
or UO_59 (O_59,N_2002,N_2163);
or UO_60 (O_60,N_2704,N_2281);
xor UO_61 (O_61,N_2792,N_2603);
and UO_62 (O_62,N_2766,N_2644);
nor UO_63 (O_63,N_2772,N_2283);
or UO_64 (O_64,N_2659,N_2449);
nor UO_65 (O_65,N_2903,N_2654);
nor UO_66 (O_66,N_2321,N_2290);
or UO_67 (O_67,N_2829,N_2971);
or UO_68 (O_68,N_2677,N_2469);
or UO_69 (O_69,N_2045,N_2767);
nor UO_70 (O_70,N_2726,N_2941);
or UO_71 (O_71,N_2862,N_2037);
or UO_72 (O_72,N_2557,N_2776);
or UO_73 (O_73,N_2275,N_2132);
nor UO_74 (O_74,N_2083,N_2302);
xnor UO_75 (O_75,N_2288,N_2457);
nand UO_76 (O_76,N_2932,N_2080);
nor UO_77 (O_77,N_2166,N_2272);
or UO_78 (O_78,N_2547,N_2453);
and UO_79 (O_79,N_2159,N_2988);
or UO_80 (O_80,N_2501,N_2418);
nand UO_81 (O_81,N_2474,N_2495);
nand UO_82 (O_82,N_2948,N_2756);
nor UO_83 (O_83,N_2494,N_2721);
nor UO_84 (O_84,N_2859,N_2268);
xor UO_85 (O_85,N_2165,N_2717);
nand UO_86 (O_86,N_2599,N_2020);
nand UO_87 (O_87,N_2243,N_2044);
nor UO_88 (O_88,N_2558,N_2640);
and UO_89 (O_89,N_2664,N_2630);
and UO_90 (O_90,N_2292,N_2350);
and UO_91 (O_91,N_2662,N_2238);
nor UO_92 (O_92,N_2355,N_2651);
and UO_93 (O_93,N_2693,N_2258);
or UO_94 (O_94,N_2608,N_2291);
nand UO_95 (O_95,N_2134,N_2384);
or UO_96 (O_96,N_2352,N_2936);
and UO_97 (O_97,N_2097,N_2802);
and UO_98 (O_98,N_2696,N_2364);
nand UO_99 (O_99,N_2203,N_2325);
nand UO_100 (O_100,N_2620,N_2867);
nor UO_101 (O_101,N_2795,N_2199);
or UO_102 (O_102,N_2379,N_2894);
nor UO_103 (O_103,N_2922,N_2949);
or UO_104 (O_104,N_2964,N_2411);
nor UO_105 (O_105,N_2222,N_2612);
or UO_106 (O_106,N_2896,N_2820);
or UO_107 (O_107,N_2361,N_2266);
or UO_108 (O_108,N_2855,N_2425);
nand UO_109 (O_109,N_2330,N_2869);
xnor UO_110 (O_110,N_2332,N_2607);
nand UO_111 (O_111,N_2483,N_2844);
nor UO_112 (O_112,N_2298,N_2516);
or UO_113 (O_113,N_2804,N_2720);
and UO_114 (O_114,N_2692,N_2192);
nor UO_115 (O_115,N_2725,N_2938);
and UO_116 (O_116,N_2568,N_2009);
or UO_117 (O_117,N_2096,N_2396);
nand UO_118 (O_118,N_2473,N_2475);
xor UO_119 (O_119,N_2485,N_2590);
nor UO_120 (O_120,N_2926,N_2315);
xor UO_121 (O_121,N_2406,N_2414);
and UO_122 (O_122,N_2426,N_2600);
or UO_123 (O_123,N_2482,N_2575);
nand UO_124 (O_124,N_2335,N_2180);
xnor UO_125 (O_125,N_2175,N_2492);
and UO_126 (O_126,N_2577,N_2416);
nor UO_127 (O_127,N_2280,N_2022);
or UO_128 (O_128,N_2107,N_2616);
nor UO_129 (O_129,N_2168,N_2583);
or UO_130 (O_130,N_2690,N_2004);
and UO_131 (O_131,N_2858,N_2628);
and UO_132 (O_132,N_2979,N_2564);
xnor UO_133 (O_133,N_2441,N_2437);
xnor UO_134 (O_134,N_2119,N_2791);
nand UO_135 (O_135,N_2525,N_2737);
and UO_136 (O_136,N_2256,N_2955);
and UO_137 (O_137,N_2947,N_2843);
nand UO_138 (O_138,N_2318,N_2057);
and UO_139 (O_139,N_2518,N_2063);
or UO_140 (O_140,N_2212,N_2409);
nor UO_141 (O_141,N_2981,N_2177);
nor UO_142 (O_142,N_2179,N_2671);
xnor UO_143 (O_143,N_2888,N_2566);
xnor UO_144 (O_144,N_2382,N_2912);
nor UO_145 (O_145,N_2144,N_2067);
xnor UO_146 (O_146,N_2274,N_2459);
or UO_147 (O_147,N_2788,N_2174);
xor UO_148 (O_148,N_2641,N_2073);
nand UO_149 (O_149,N_2204,N_2108);
nor UO_150 (O_150,N_2974,N_2775);
and UO_151 (O_151,N_2702,N_2937);
or UO_152 (O_152,N_2541,N_2081);
or UO_153 (O_153,N_2241,N_2768);
or UO_154 (O_154,N_2509,N_2086);
or UO_155 (O_155,N_2915,N_2700);
and UO_156 (O_156,N_2570,N_2650);
or UO_157 (O_157,N_2095,N_2764);
xor UO_158 (O_158,N_2075,N_2751);
xor UO_159 (O_159,N_2730,N_2579);
nand UO_160 (O_160,N_2913,N_2456);
xnor UO_161 (O_161,N_2782,N_2211);
xor UO_162 (O_162,N_2158,N_2527);
xnor UO_163 (O_163,N_2622,N_2699);
nand UO_164 (O_164,N_2550,N_2691);
nand UO_165 (O_165,N_2074,N_2580);
nand UO_166 (O_166,N_2419,N_2841);
xor UO_167 (O_167,N_2287,N_2376);
or UO_168 (O_168,N_2918,N_2891);
or UO_169 (O_169,N_2945,N_2601);
nand UO_170 (O_170,N_2434,N_2761);
xnor UO_171 (O_171,N_2346,N_2929);
nand UO_172 (O_172,N_2387,N_2789);
nand UO_173 (O_173,N_2458,N_2040);
and UO_174 (O_174,N_2011,N_2552);
and UO_175 (O_175,N_2811,N_2991);
nor UO_176 (O_176,N_2343,N_2443);
nand UO_177 (O_177,N_2339,N_2391);
xnor UO_178 (O_178,N_2023,N_2289);
or UO_179 (O_179,N_2796,N_2716);
xor UO_180 (O_180,N_2215,N_2856);
xor UO_181 (O_181,N_2410,N_2400);
xnor UO_182 (O_182,N_2742,N_2377);
and UO_183 (O_183,N_2689,N_2614);
or UO_184 (O_184,N_2191,N_2026);
and UO_185 (O_185,N_2923,N_2666);
or UO_186 (O_186,N_2569,N_2070);
nor UO_187 (O_187,N_2278,N_2807);
or UO_188 (O_188,N_2618,N_2263);
nand UO_189 (O_189,N_2142,N_2838);
nand UO_190 (O_190,N_2507,N_2656);
nand UO_191 (O_191,N_2821,N_2977);
or UO_192 (O_192,N_2746,N_2753);
nand UO_193 (O_193,N_2673,N_2794);
nor UO_194 (O_194,N_2672,N_2299);
nand UO_195 (O_195,N_2892,N_2236);
xnor UO_196 (O_196,N_2961,N_2670);
or UO_197 (O_197,N_2832,N_2111);
nand UO_198 (O_198,N_2276,N_2357);
nor UO_199 (O_199,N_2519,N_2279);
nor UO_200 (O_200,N_2878,N_2743);
nand UO_201 (O_201,N_2363,N_2769);
xor UO_202 (O_202,N_2408,N_2994);
nor UO_203 (O_203,N_2549,N_2639);
or UO_204 (O_204,N_2286,N_2015);
nand UO_205 (O_205,N_2529,N_2098);
nor UO_206 (O_206,N_2633,N_2156);
or UO_207 (O_207,N_2837,N_2609);
and UO_208 (O_208,N_2341,N_2900);
xnor UO_209 (O_209,N_2206,N_2989);
or UO_210 (O_210,N_2486,N_2933);
and UO_211 (O_211,N_2593,N_2698);
xnor UO_212 (O_212,N_2835,N_2366);
and UO_213 (O_213,N_2987,N_2029);
xnor UO_214 (O_214,N_2490,N_2170);
or UO_215 (O_215,N_2757,N_2615);
nand UO_216 (O_216,N_2058,N_2805);
nand UO_217 (O_217,N_2983,N_2750);
nand UO_218 (O_218,N_2719,N_2873);
and UO_219 (O_219,N_2871,N_2472);
xor UO_220 (O_220,N_2759,N_2401);
xnor UO_221 (O_221,N_2845,N_2301);
nor UO_222 (O_222,N_2890,N_2164);
or UO_223 (O_223,N_2512,N_2665);
xor UO_224 (O_224,N_2762,N_2797);
nor UO_225 (O_225,N_2173,N_2565);
xor UO_226 (O_226,N_2113,N_2378);
nor UO_227 (O_227,N_2123,N_2819);
nor UO_228 (O_228,N_2423,N_2003);
or UO_229 (O_229,N_2959,N_2567);
nor UO_230 (O_230,N_2760,N_2808);
nand UO_231 (O_231,N_2847,N_2661);
xnor UO_232 (O_232,N_2897,N_2984);
and UO_233 (O_233,N_2216,N_2637);
and UO_234 (O_234,N_2877,N_2823);
xnor UO_235 (O_235,N_2731,N_2147);
or UO_236 (O_236,N_2917,N_2857);
or UO_237 (O_237,N_2993,N_2982);
xnor UO_238 (O_238,N_2210,N_2105);
xnor UO_239 (O_239,N_2733,N_2445);
or UO_240 (O_240,N_2784,N_2901);
nand UO_241 (O_241,N_2319,N_2546);
nor UO_242 (O_242,N_2581,N_2424);
nor UO_243 (O_243,N_2723,N_2528);
nor UO_244 (O_244,N_2783,N_2383);
nor UO_245 (O_245,N_2812,N_2381);
xor UO_246 (O_246,N_2284,N_2604);
xnor UO_247 (O_247,N_2793,N_2621);
and UO_248 (O_248,N_2610,N_2253);
xnor UO_249 (O_249,N_2533,N_2358);
and UO_250 (O_250,N_2428,N_2050);
or UO_251 (O_251,N_2613,N_2504);
nand UO_252 (O_252,N_2985,N_2735);
or UO_253 (O_253,N_2521,N_2157);
xor UO_254 (O_254,N_2016,N_2828);
nand UO_255 (O_255,N_2773,N_2960);
or UO_256 (O_256,N_2186,N_2709);
xnor UO_257 (O_257,N_2311,N_2595);
xnor UO_258 (O_258,N_2722,N_2815);
and UO_259 (O_259,N_2101,N_2513);
nor UO_260 (O_260,N_2831,N_2990);
nor UO_261 (O_261,N_2273,N_2573);
xor UO_262 (O_262,N_2228,N_2996);
nor UO_263 (O_263,N_2125,N_2799);
xnor UO_264 (O_264,N_2488,N_2818);
and UO_265 (O_265,N_2353,N_2141);
or UO_266 (O_266,N_2626,N_2574);
xnor UO_267 (O_267,N_2508,N_2237);
or UO_268 (O_268,N_2118,N_2986);
nor UO_269 (O_269,N_2120,N_2646);
and UO_270 (O_270,N_2219,N_2543);
and UO_271 (O_271,N_2310,N_2139);
and UO_272 (O_272,N_2534,N_2536);
nand UO_273 (O_273,N_2124,N_2957);
nand UO_274 (O_274,N_2094,N_2259);
nor UO_275 (O_275,N_2649,N_2345);
nand UO_276 (O_276,N_2388,N_2827);
nand UO_277 (O_277,N_2196,N_2127);
nand UO_278 (O_278,N_2312,N_2373);
xor UO_279 (O_279,N_2187,N_2925);
and UO_280 (O_280,N_2498,N_2031);
nor UO_281 (O_281,N_2634,N_2479);
and UO_282 (O_282,N_2307,N_2049);
xor UO_283 (O_283,N_2978,N_2729);
or UO_284 (O_284,N_2834,N_2638);
nor UO_285 (O_285,N_2250,N_2830);
and UO_286 (O_286,N_2853,N_2935);
xor UO_287 (O_287,N_2154,N_2559);
and UO_288 (O_288,N_2327,N_2245);
nor UO_289 (O_289,N_2708,N_2576);
nand UO_290 (O_290,N_2668,N_2242);
nand UO_291 (O_291,N_2261,N_2707);
and UO_292 (O_292,N_2244,N_2201);
or UO_293 (O_293,N_2752,N_2875);
nor UO_294 (O_294,N_2653,N_2221);
or UO_295 (O_295,N_2652,N_2738);
xor UO_296 (O_296,N_2801,N_2898);
nor UO_297 (O_297,N_2464,N_2487);
nor UO_298 (O_298,N_2181,N_2155);
nor UO_299 (O_299,N_2397,N_2398);
nor UO_300 (O_300,N_2100,N_2069);
xnor UO_301 (O_301,N_2197,N_2771);
nor UO_302 (O_302,N_2523,N_2596);
xor UO_303 (O_303,N_2229,N_2254);
or UO_304 (O_304,N_2839,N_2447);
and UO_305 (O_305,N_2934,N_2282);
nand UO_306 (O_306,N_2420,N_2334);
and UO_307 (O_307,N_2585,N_2102);
nor UO_308 (O_308,N_2055,N_2910);
and UO_309 (O_309,N_2407,N_2403);
or UO_310 (O_310,N_2390,N_2578);
or UO_311 (O_311,N_2169,N_2824);
and UO_312 (O_312,N_2202,N_2740);
xnor UO_313 (O_313,N_2822,N_2992);
xor UO_314 (O_314,N_2106,N_2556);
nor UO_315 (O_315,N_2598,N_2703);
nor UO_316 (O_316,N_2623,N_2136);
nor UO_317 (O_317,N_2554,N_2968);
nor UO_318 (O_318,N_2514,N_2995);
or UO_319 (O_319,N_2826,N_2039);
or UO_320 (O_320,N_2676,N_2816);
xor UO_321 (O_321,N_2193,N_2980);
nand UO_322 (O_322,N_2911,N_2586);
or UO_323 (O_323,N_2269,N_2946);
nand UO_324 (O_324,N_2354,N_2927);
and UO_325 (O_325,N_2718,N_2452);
nand UO_326 (O_326,N_2744,N_2810);
nor UO_327 (O_327,N_2326,N_2865);
or UO_328 (O_328,N_2053,N_2520);
or UO_329 (O_329,N_2471,N_2806);
xor UO_330 (O_330,N_2088,N_2308);
or UO_331 (O_331,N_2404,N_2780);
nor UO_332 (O_332,N_2303,N_2389);
nor UO_333 (O_333,N_2121,N_2460);
nand UO_334 (O_334,N_2883,N_2248);
or UO_335 (O_335,N_2629,N_2678);
nor UO_336 (O_336,N_2803,N_2825);
xor UO_337 (O_337,N_2270,N_2594);
xnor UO_338 (O_338,N_2701,N_2316);
and UO_339 (O_339,N_2099,N_2958);
nand UO_340 (O_340,N_2148,N_2798);
nor UO_341 (O_341,N_2591,N_2881);
nor UO_342 (O_342,N_2161,N_2882);
and UO_343 (O_343,N_2438,N_2296);
nor UO_344 (O_344,N_2499,N_2684);
nand UO_345 (O_345,N_2370,N_2214);
xor UO_346 (O_346,N_2062,N_2041);
and UO_347 (O_347,N_2129,N_2012);
or UO_348 (O_348,N_2584,N_2333);
and UO_349 (O_349,N_2951,N_2636);
and UO_350 (O_350,N_2736,N_2128);
xnor UO_351 (O_351,N_2679,N_2493);
and UO_352 (O_352,N_2916,N_2694);
xor UO_353 (O_353,N_2943,N_2317);
nor UO_354 (O_354,N_2112,N_2538);
or UO_355 (O_355,N_2647,N_2227);
nor UO_356 (O_356,N_2813,N_2249);
or UO_357 (O_357,N_2252,N_2038);
nand UO_358 (O_358,N_2320,N_2904);
or UO_359 (O_359,N_2745,N_2920);
nor UO_360 (O_360,N_2635,N_2306);
nor UO_361 (O_361,N_2864,N_2589);
or UO_362 (O_362,N_2454,N_2611);
or UO_363 (O_363,N_2660,N_2077);
nor UO_364 (O_364,N_2597,N_2942);
or UO_365 (O_365,N_2571,N_2531);
and UO_366 (O_366,N_2976,N_2602);
nand UO_367 (O_367,N_2505,N_2836);
nand UO_368 (O_368,N_2669,N_2065);
or UO_369 (O_369,N_2146,N_2551);
xor UO_370 (O_370,N_2470,N_2380);
xnor UO_371 (O_371,N_2374,N_2758);
and UO_372 (O_372,N_2809,N_2234);
xor UO_373 (O_373,N_2683,N_2078);
nand UO_374 (O_374,N_2765,N_2969);
nand UO_375 (O_375,N_2393,N_2235);
nand UO_376 (O_376,N_2260,N_2781);
and UO_377 (O_377,N_2465,N_2695);
nand UO_378 (O_378,N_2582,N_2870);
xor UO_379 (O_379,N_2790,N_2532);
and UO_380 (O_380,N_2297,N_2786);
nand UO_381 (O_381,N_2587,N_2480);
nor UO_382 (O_382,N_2246,N_2209);
or UO_383 (O_383,N_2539,N_2497);
nand UO_384 (O_384,N_2506,N_2967);
and UO_385 (O_385,N_2866,N_2028);
and UO_386 (O_386,N_2093,N_2667);
nand UO_387 (O_387,N_2884,N_2104);
nor UO_388 (O_388,N_2402,N_2481);
nor UO_389 (O_389,N_2223,N_2048);
or UO_390 (O_390,N_2331,N_2035);
and UO_391 (O_391,N_2115,N_2777);
nor UO_392 (O_392,N_2553,N_2338);
xnor UO_393 (O_393,N_2143,N_2172);
or UO_394 (O_394,N_2131,N_2110);
and UO_395 (O_395,N_2116,N_2047);
and UO_396 (O_396,N_2375,N_2627);
nor UO_397 (O_397,N_2137,N_2965);
xor UO_398 (O_398,N_2344,N_2271);
nor UO_399 (O_399,N_2183,N_2300);
and UO_400 (O_400,N_2861,N_2625);
nor UO_401 (O_401,N_2940,N_2072);
nor UO_402 (O_402,N_2089,N_2046);
xnor UO_403 (O_403,N_2133,N_2149);
and UO_404 (O_404,N_2998,N_2255);
xnor UO_405 (O_405,N_2277,N_2340);
xor UO_406 (O_406,N_2071,N_2421);
xor UO_407 (O_407,N_2747,N_2150);
xor UO_408 (O_408,N_2060,N_2328);
xnor UO_409 (O_409,N_2846,N_2372);
and UO_410 (O_410,N_2973,N_2362);
or UO_411 (O_411,N_2000,N_2013);
and UO_412 (O_412,N_2741,N_2231);
nor UO_413 (O_413,N_2251,N_2914);
xor UO_414 (O_414,N_2755,N_2442);
or UO_415 (O_415,N_2928,N_2705);
nand UO_416 (O_416,N_2848,N_2034);
nor UO_417 (O_417,N_2999,N_2462);
nand UO_418 (O_418,N_2200,N_2931);
nand UO_419 (O_419,N_2658,N_2194);
and UO_420 (O_420,N_2675,N_2476);
xor UO_421 (O_421,N_2033,N_2122);
xnor UO_422 (O_422,N_2944,N_2349);
nor UO_423 (O_423,N_2526,N_2051);
xnor UO_424 (O_424,N_2966,N_2930);
nand UO_425 (O_425,N_2224,N_2484);
and UO_426 (O_426,N_2413,N_2167);
or UO_427 (O_427,N_2734,N_2535);
and UO_428 (O_428,N_2233,N_2394);
or UO_429 (O_429,N_2908,N_2240);
and UO_430 (O_430,N_2090,N_2084);
xor UO_431 (O_431,N_2293,N_2369);
nand UO_432 (O_432,N_2422,N_2052);
nor UO_433 (O_433,N_2467,N_2027);
or UO_434 (O_434,N_2774,N_2461);
xnor UO_435 (O_435,N_2919,N_2436);
nand UO_436 (O_436,N_2130,N_2061);
xor UO_437 (O_437,N_2950,N_2956);
or UO_438 (O_438,N_2631,N_2213);
xor UO_439 (O_439,N_2184,N_2503);
nand UO_440 (O_440,N_2359,N_2491);
or UO_441 (O_441,N_2909,N_2889);
or UO_442 (O_442,N_2247,N_2103);
xor UO_443 (O_443,N_2225,N_2076);
nand UO_444 (O_444,N_2322,N_2439);
nand UO_445 (O_445,N_2540,N_2091);
xnor UO_446 (O_446,N_2560,N_2392);
and UO_447 (O_447,N_2336,N_2309);
xnor UO_448 (O_448,N_2840,N_2975);
nand UO_449 (O_449,N_2395,N_2415);
or UO_450 (O_450,N_2478,N_2850);
and UO_451 (O_451,N_2561,N_2314);
nand UO_452 (O_452,N_2778,N_2329);
or UO_453 (O_453,N_2872,N_2643);
and UO_454 (O_454,N_2185,N_2496);
xnor UO_455 (O_455,N_2939,N_2024);
nand UO_456 (O_456,N_2511,N_2522);
or UO_457 (O_457,N_2446,N_2342);
xor UO_458 (O_458,N_2542,N_2648);
xor UO_459 (O_459,N_2572,N_2732);
and UO_460 (O_460,N_2087,N_2444);
xor UO_461 (O_461,N_2544,N_2304);
and UO_462 (O_462,N_2887,N_2153);
and UO_463 (O_463,N_2688,N_2970);
nor UO_464 (O_464,N_2152,N_2412);
nand UO_465 (O_465,N_2680,N_2517);
nor UO_466 (O_466,N_2466,N_2817);
nand UO_467 (O_467,N_2005,N_2059);
nand UO_468 (O_468,N_2126,N_2754);
xnor UO_469 (O_469,N_2963,N_2537);
xnor UO_470 (O_470,N_2924,N_2207);
and UO_471 (O_471,N_2285,N_2879);
and UO_472 (O_472,N_2500,N_2220);
or UO_473 (O_473,N_2674,N_2351);
or UO_474 (O_474,N_2728,N_2082);
and UO_475 (O_475,N_2114,N_2954);
or UO_476 (O_476,N_2455,N_2360);
xor UO_477 (O_477,N_2368,N_2663);
nor UO_478 (O_478,N_2606,N_2895);
or UO_479 (O_479,N_2515,N_2007);
and UO_480 (O_480,N_2014,N_2712);
or UO_481 (O_481,N_2562,N_2763);
or UO_482 (O_482,N_2907,N_2748);
nand UO_483 (O_483,N_2008,N_2697);
nand UO_484 (O_484,N_2226,N_2739);
nand UO_485 (O_485,N_2624,N_2548);
xnor UO_486 (O_486,N_2953,N_2800);
or UO_487 (O_487,N_2405,N_2432);
and UO_488 (O_488,N_2902,N_2450);
nand UO_489 (O_489,N_2427,N_2886);
nor UO_490 (O_490,N_2265,N_2064);
xnor UO_491 (O_491,N_2868,N_2814);
or UO_492 (O_492,N_2182,N_2714);
nor UO_493 (O_493,N_2430,N_2619);
nand UO_494 (O_494,N_2645,N_2605);
nand UO_495 (O_495,N_2042,N_2092);
or UO_496 (O_496,N_2433,N_2682);
nand UO_497 (O_497,N_2054,N_2323);
nand UO_498 (O_498,N_2138,N_2463);
xor UO_499 (O_499,N_2724,N_2188);
endmodule