module basic_2500_25000_3000_50_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1383,In_1225);
xnor U1 (N_1,In_151,In_792);
nor U2 (N_2,In_586,In_155);
and U3 (N_3,In_1360,In_641);
nand U4 (N_4,In_1642,In_2063);
xor U5 (N_5,In_2482,In_1773);
nor U6 (N_6,In_725,In_272);
or U7 (N_7,In_2151,In_419);
or U8 (N_8,In_518,In_1960);
nand U9 (N_9,In_1151,In_1638);
and U10 (N_10,In_2322,In_451);
nor U11 (N_11,In_1999,In_2473);
nor U12 (N_12,In_1066,In_1488);
nor U13 (N_13,In_2411,In_2091);
xor U14 (N_14,In_1357,In_143);
or U15 (N_15,In_2280,In_1906);
nor U16 (N_16,In_1430,In_134);
nor U17 (N_17,In_177,In_1484);
xor U18 (N_18,In_2186,In_554);
nor U19 (N_19,In_978,In_539);
xnor U20 (N_20,In_1845,In_1099);
and U21 (N_21,In_604,In_2373);
nand U22 (N_22,In_524,In_1387);
xor U23 (N_23,In_2141,In_2075);
nor U24 (N_24,In_717,In_33);
or U25 (N_25,In_1763,In_1079);
nor U26 (N_26,In_1280,In_1260);
nand U27 (N_27,In_2227,In_653);
or U28 (N_28,In_731,In_907);
nand U29 (N_29,In_1232,In_1180);
nor U30 (N_30,In_2136,In_2226);
nor U31 (N_31,In_1256,In_1457);
and U32 (N_32,In_1563,In_1104);
nand U33 (N_33,In_1121,In_373);
and U34 (N_34,In_395,In_1841);
or U35 (N_35,In_2038,In_443);
xor U36 (N_36,In_1808,In_331);
or U37 (N_37,In_2059,In_489);
nand U38 (N_38,In_1322,In_2429);
or U39 (N_39,In_791,In_1944);
nor U40 (N_40,In_1135,In_1885);
nor U41 (N_41,In_1184,In_469);
nand U42 (N_42,In_313,In_1327);
and U43 (N_43,In_2235,In_1941);
xor U44 (N_44,In_1441,In_1054);
or U45 (N_45,In_316,In_2331);
and U46 (N_46,In_847,In_411);
or U47 (N_47,In_1816,In_242);
nand U48 (N_48,In_32,In_1755);
nand U49 (N_49,In_186,In_96);
or U50 (N_50,In_898,In_2299);
nand U51 (N_51,In_122,In_1794);
nor U52 (N_52,In_1301,In_668);
and U53 (N_53,In_2195,In_1840);
and U54 (N_54,In_71,In_2325);
or U55 (N_55,In_2118,In_1950);
and U56 (N_56,In_2066,In_1905);
and U57 (N_57,In_145,In_528);
nand U58 (N_58,In_1820,In_251);
nor U59 (N_59,In_719,In_977);
nor U60 (N_60,In_1371,In_2272);
or U61 (N_61,In_1230,In_175);
and U62 (N_62,In_1560,In_1014);
or U63 (N_63,In_1183,In_2044);
xnor U64 (N_64,In_2254,In_1328);
xor U65 (N_65,In_2264,In_2407);
and U66 (N_66,In_2001,In_669);
nor U67 (N_67,In_857,In_1416);
nand U68 (N_68,In_1534,In_812);
xnor U69 (N_69,In_249,In_1468);
xnor U70 (N_70,In_1466,In_1966);
or U71 (N_71,In_382,In_1530);
xor U72 (N_72,In_1956,In_658);
nor U73 (N_73,In_809,In_2005);
nor U74 (N_74,In_1163,In_1525);
nand U75 (N_75,In_20,In_1711);
xor U76 (N_76,In_1733,In_91);
nor U77 (N_77,In_2120,In_2218);
and U78 (N_78,In_2403,In_1471);
nor U79 (N_79,In_2347,In_1435);
nand U80 (N_80,In_1164,In_87);
nand U81 (N_81,In_2175,In_499);
or U82 (N_82,In_883,In_1804);
xor U83 (N_83,In_1947,In_1393);
xnor U84 (N_84,In_178,In_1578);
or U85 (N_85,In_2351,In_2165);
nor U86 (N_86,In_1299,In_1681);
nor U87 (N_87,In_2158,In_2378);
nor U88 (N_88,In_775,In_2438);
nand U89 (N_89,In_1427,In_968);
nor U90 (N_90,In_1717,In_612);
and U91 (N_91,In_1548,In_1606);
xor U92 (N_92,In_1541,In_1012);
xor U93 (N_93,In_84,In_1677);
xor U94 (N_94,In_435,In_1922);
nor U95 (N_95,In_227,In_2460);
nor U96 (N_96,In_628,In_463);
nand U97 (N_97,In_187,In_1186);
nor U98 (N_98,In_1772,In_333);
or U99 (N_99,In_222,In_2475);
or U100 (N_100,In_1623,In_1010);
or U101 (N_101,In_467,In_271);
nand U102 (N_102,In_219,In_769);
nand U103 (N_103,In_1146,In_1193);
xor U104 (N_104,In_179,In_329);
nand U105 (N_105,In_2215,In_2340);
nor U106 (N_106,In_825,In_1119);
nand U107 (N_107,In_495,In_594);
xor U108 (N_108,In_2251,In_863);
and U109 (N_109,In_2101,In_1300);
nor U110 (N_110,In_2350,In_1402);
nand U111 (N_111,In_2334,In_292);
and U112 (N_112,In_1660,In_834);
and U113 (N_113,In_2269,In_383);
nor U114 (N_114,In_1353,In_1384);
nor U115 (N_115,In_1628,In_2237);
xnor U116 (N_116,In_1798,In_1889);
and U117 (N_117,In_1108,In_591);
nor U118 (N_118,In_108,In_840);
xor U119 (N_119,In_569,In_284);
or U120 (N_120,In_203,In_264);
xor U121 (N_121,In_1069,In_755);
and U122 (N_122,In_2291,In_1071);
and U123 (N_123,In_889,In_1158);
and U124 (N_124,In_1048,In_1814);
nand U125 (N_125,In_399,In_697);
or U126 (N_126,In_1349,In_2316);
or U127 (N_127,In_148,In_966);
xnor U128 (N_128,In_2238,In_1902);
or U129 (N_129,In_404,In_1639);
xnor U130 (N_130,In_1254,In_2246);
nand U131 (N_131,In_477,In_1378);
nand U132 (N_132,In_959,In_1281);
and U133 (N_133,In_403,In_1728);
xnor U134 (N_134,In_585,In_1882);
or U135 (N_135,In_431,In_502);
nor U136 (N_136,In_1671,In_1325);
xnor U137 (N_137,In_1479,In_2314);
xor U138 (N_138,In_1437,In_957);
or U139 (N_139,In_453,In_273);
nand U140 (N_140,In_1687,In_428);
and U141 (N_141,In_852,In_2140);
nor U142 (N_142,In_1825,In_2479);
nor U143 (N_143,In_380,In_1988);
nor U144 (N_144,In_2148,In_57);
and U145 (N_145,In_1053,In_1451);
xnor U146 (N_146,In_11,In_826);
and U147 (N_147,In_436,In_115);
or U148 (N_148,In_1455,In_2262);
and U149 (N_149,In_1156,In_1134);
and U150 (N_150,In_173,In_929);
or U151 (N_151,In_2400,In_1501);
xor U152 (N_152,In_163,In_39);
and U153 (N_153,In_146,In_745);
xor U154 (N_154,In_1444,In_1702);
nand U155 (N_155,In_818,In_540);
xnor U156 (N_156,In_1324,In_483);
nand U157 (N_157,In_250,In_1990);
and U158 (N_158,In_2494,In_2245);
or U159 (N_159,In_5,In_716);
nand U160 (N_160,In_493,In_2089);
nand U161 (N_161,In_995,In_1921);
and U162 (N_162,In_1699,In_657);
or U163 (N_163,In_80,In_627);
nand U164 (N_164,In_681,In_2448);
and U165 (N_165,In_181,In_2268);
or U166 (N_166,In_1004,In_19);
or U167 (N_167,In_400,In_2150);
nor U168 (N_168,In_934,In_916);
and U169 (N_169,In_1580,In_1105);
or U170 (N_170,In_2297,In_265);
or U171 (N_171,In_507,In_1646);
nor U172 (N_172,In_797,In_202);
nand U173 (N_173,In_1619,In_1552);
xor U174 (N_174,In_83,In_902);
nor U175 (N_175,In_822,In_922);
or U176 (N_176,In_1948,In_293);
nor U177 (N_177,In_261,In_1617);
and U178 (N_178,In_813,In_1070);
nor U179 (N_179,In_2194,In_1751);
and U180 (N_180,In_579,In_777);
xnor U181 (N_181,In_1937,In_76);
xnor U182 (N_182,In_2026,In_1807);
nor U183 (N_183,In_2164,In_1596);
nor U184 (N_184,In_2225,In_319);
nor U185 (N_185,In_1142,In_470);
nand U186 (N_186,In_2058,In_1713);
or U187 (N_187,In_378,In_746);
xor U188 (N_188,In_2317,In_92);
and U189 (N_189,In_2163,In_367);
nand U190 (N_190,In_908,In_109);
and U191 (N_191,In_1945,In_64);
nor U192 (N_192,In_2395,In_666);
or U193 (N_193,In_17,In_672);
xnor U194 (N_194,In_1212,In_2497);
and U195 (N_195,In_113,In_131);
or U196 (N_196,In_1940,In_432);
or U197 (N_197,In_590,In_2304);
nor U198 (N_198,In_1174,In_1269);
xnor U199 (N_199,In_2368,In_1887);
nand U200 (N_200,In_2312,In_938);
xnor U201 (N_201,In_911,In_446);
and U202 (N_202,In_550,In_207);
nor U203 (N_203,In_337,In_2442);
nand U204 (N_204,In_1224,In_307);
or U205 (N_205,In_376,In_674);
and U206 (N_206,In_983,In_1277);
nor U207 (N_207,In_2397,In_675);
xor U208 (N_208,In_632,In_2493);
nor U209 (N_209,In_2160,In_806);
or U210 (N_210,In_1314,In_311);
nor U211 (N_211,In_1631,In_58);
or U212 (N_212,In_936,In_1018);
or U213 (N_213,In_2315,In_1517);
and U214 (N_214,In_671,In_1162);
and U215 (N_215,In_127,In_1460);
nand U216 (N_216,In_1201,In_2109);
and U217 (N_217,In_1476,In_2472);
nor U218 (N_218,In_1866,In_1306);
nand U219 (N_219,In_1914,In_2224);
and U220 (N_220,In_1011,In_1429);
or U221 (N_221,In_947,In_1234);
nor U222 (N_222,In_728,In_593);
xor U223 (N_223,In_101,In_1745);
xnor U224 (N_224,In_858,In_1986);
nor U225 (N_225,In_1392,In_1573);
or U226 (N_226,In_498,In_1729);
and U227 (N_227,In_564,In_2446);
and U228 (N_228,In_37,In_1746);
or U229 (N_229,In_993,In_368);
and U230 (N_230,In_417,In_1629);
nand U231 (N_231,In_758,In_2394);
and U232 (N_232,In_522,In_1523);
and U233 (N_233,In_1493,In_723);
and U234 (N_234,In_991,In_1810);
nand U235 (N_235,In_1795,In_1022);
xor U236 (N_236,In_901,In_2080);
xor U237 (N_237,In_925,In_1089);
xnor U238 (N_238,In_1293,In_1697);
or U239 (N_239,In_1340,In_85);
nor U240 (N_240,In_695,In_690);
or U241 (N_241,In_1673,In_2499);
xnor U242 (N_242,In_111,In_167);
or U243 (N_243,In_1881,In_1620);
and U244 (N_244,In_2426,In_2471);
and U245 (N_245,In_2477,In_2032);
nand U246 (N_246,In_1591,In_1725);
nor U247 (N_247,In_1274,In_1686);
or U248 (N_248,In_615,In_1499);
and U249 (N_249,In_734,In_1526);
nor U250 (N_250,In_1211,In_89);
nor U251 (N_251,In_236,In_2348);
and U252 (N_252,In_866,In_430);
nand U253 (N_253,In_962,In_1284);
xor U254 (N_254,In_9,In_1027);
or U255 (N_255,In_1370,In_183);
and U256 (N_256,In_1038,In_1506);
nand U257 (N_257,In_1756,In_525);
xnor U258 (N_258,In_2391,In_266);
xor U259 (N_259,In_2149,In_2381);
or U260 (N_260,In_1399,In_808);
or U261 (N_261,In_976,In_1282);
and U262 (N_262,In_1992,In_1481);
or U263 (N_263,In_63,In_415);
nand U264 (N_264,In_1528,In_589);
nand U265 (N_265,In_667,In_1006);
xnor U266 (N_266,In_2274,In_280);
and U267 (N_267,In_1157,In_2451);
xnor U268 (N_268,In_1200,In_223);
xor U269 (N_269,In_2084,In_753);
xnor U270 (N_270,In_2388,In_1365);
xnor U271 (N_271,In_2130,In_996);
xnor U272 (N_272,In_82,In_409);
nand U273 (N_273,In_456,In_890);
xor U274 (N_274,In_2017,In_2053);
xnor U275 (N_275,In_783,In_1286);
or U276 (N_276,In_721,In_318);
nor U277 (N_277,In_835,In_379);
xnor U278 (N_278,In_1197,In_2232);
nor U279 (N_279,In_2415,In_239);
nand U280 (N_280,In_1998,In_1559);
nor U281 (N_281,In_2401,In_971);
and U282 (N_282,In_1375,In_1909);
and U283 (N_283,In_2188,In_1590);
xnor U284 (N_284,In_599,In_1233);
nor U285 (N_285,In_751,In_1851);
or U286 (N_286,In_850,In_1716);
or U287 (N_287,In_2319,In_317);
nor U288 (N_288,In_1401,In_1288);
nand U289 (N_289,In_1760,In_1764);
nor U290 (N_290,In_838,In_228);
nor U291 (N_291,In_1724,In_194);
or U292 (N_292,In_478,In_2104);
or U293 (N_293,In_2113,In_2439);
nand U294 (N_294,In_2040,In_182);
and U295 (N_295,In_1228,In_687);
xnor U296 (N_296,In_2092,In_692);
or U297 (N_297,In_747,In_325);
or U298 (N_298,In_192,In_358);
or U299 (N_299,In_2489,In_963);
or U300 (N_300,In_861,In_1955);
xnor U301 (N_301,In_394,In_262);
xor U302 (N_302,In_732,In_268);
or U303 (N_303,In_2128,In_2054);
xnor U304 (N_304,In_1570,In_1969);
and U305 (N_305,In_1267,In_421);
nor U306 (N_306,In_2030,In_1672);
nor U307 (N_307,In_1020,In_831);
xor U308 (N_308,In_128,In_988);
xor U309 (N_309,In_1217,In_263);
nand U310 (N_310,In_1275,In_706);
xnor U311 (N_311,In_1334,In_2288);
nor U312 (N_312,In_1959,In_2321);
and U313 (N_313,In_1210,In_536);
and U314 (N_314,In_1837,In_1458);
nand U315 (N_315,In_1483,In_1019);
nand U316 (N_316,In_1641,In_2060);
or U317 (N_317,In_256,In_2440);
and U318 (N_318,In_789,In_141);
nand U319 (N_319,In_2137,In_2079);
nor U320 (N_320,In_764,In_1077);
or U321 (N_321,In_2057,In_1313);
or U322 (N_322,In_2103,In_166);
and U323 (N_323,In_270,In_452);
and U324 (N_324,In_1005,In_327);
xnor U325 (N_325,In_654,In_2311);
xnor U326 (N_326,In_2432,In_1098);
nor U327 (N_327,In_897,In_644);
xor U328 (N_328,In_1657,In_304);
and U329 (N_329,In_2328,In_2111);
and U330 (N_330,In_2298,In_1783);
or U331 (N_331,In_86,In_575);
nor U332 (N_332,In_660,In_1047);
nand U333 (N_333,In_701,In_881);
xor U334 (N_334,In_759,In_260);
or U335 (N_335,In_696,In_1691);
xnor U336 (N_336,In_2071,In_1985);
nand U337 (N_337,In_2228,In_607);
nor U338 (N_338,In_639,In_827);
nand U339 (N_339,In_1196,In_1597);
nand U340 (N_340,In_1002,In_2016);
nand U341 (N_341,In_2056,In_1386);
and U342 (N_342,In_439,In_1065);
nand U343 (N_343,In_953,In_596);
and U344 (N_344,In_1779,In_1372);
nand U345 (N_345,In_335,In_1718);
nor U346 (N_346,In_56,In_989);
and U347 (N_347,In_506,In_2083);
nand U348 (N_348,In_1490,In_810);
or U349 (N_349,In_1302,In_1522);
and U350 (N_350,In_1759,In_578);
nand U351 (N_351,In_298,In_2453);
nor U352 (N_352,In_1173,In_1787);
nand U353 (N_353,In_2308,In_412);
nor U354 (N_354,In_726,In_1696);
and U355 (N_355,In_1614,In_1358);
or U356 (N_356,In_1305,In_2207);
xnor U357 (N_357,In_1405,In_2413);
and U358 (N_358,In_70,In_1510);
nor U359 (N_359,In_1609,In_2404);
xnor U360 (N_360,In_2003,In_1043);
or U361 (N_361,In_2329,In_209);
xor U362 (N_362,In_1720,In_1740);
nor U363 (N_363,In_1319,In_204);
nand U364 (N_364,In_45,In_150);
and U365 (N_365,In_1754,In_1561);
nand U366 (N_366,In_2229,In_771);
nor U367 (N_367,In_388,In_1218);
nor U368 (N_368,In_22,In_766);
nor U369 (N_369,In_1854,In_299);
nor U370 (N_370,In_225,In_1957);
xor U371 (N_371,In_1843,In_545);
nand U372 (N_372,In_919,In_129);
xor U373 (N_373,In_387,In_1895);
xnor U374 (N_374,In_710,In_1329);
or U375 (N_375,In_975,In_60);
or U376 (N_376,In_1736,In_2356);
xnor U377 (N_377,In_1991,In_1839);
and U378 (N_378,In_1747,In_556);
nor U379 (N_379,In_844,In_1192);
xor U380 (N_380,In_1298,In_548);
nand U381 (N_381,In_40,In_1727);
xor U382 (N_382,In_1930,In_2441);
xnor U383 (N_383,In_2198,In_1678);
or U384 (N_384,In_1369,In_1610);
nand U385 (N_385,In_2015,In_427);
nor U386 (N_386,In_2110,In_1768);
and U387 (N_387,In_1996,In_160);
or U388 (N_388,In_420,In_1209);
nand U389 (N_389,In_987,In_864);
nor U390 (N_390,In_1459,In_75);
nand U391 (N_391,In_1859,In_41);
and U392 (N_392,In_1050,In_2093);
nor U393 (N_393,In_981,In_1583);
or U394 (N_394,In_2098,In_2360);
or U395 (N_395,In_1311,In_762);
and U396 (N_396,In_1635,In_2124);
xnor U397 (N_397,In_1388,In_2041);
and U398 (N_398,In_1704,In_1878);
xnor U399 (N_399,In_2034,In_914);
xor U400 (N_400,In_500,In_1555);
or U401 (N_401,In_676,In_571);
nand U402 (N_402,In_244,In_1502);
nor U403 (N_403,In_398,In_157);
xnor U404 (N_404,In_1901,In_1421);
nand U405 (N_405,In_1817,In_1876);
nor U406 (N_406,In_1422,In_972);
xor U407 (N_407,In_885,In_1867);
nor U408 (N_408,In_459,In_905);
nor U409 (N_409,In_2187,In_1962);
xnor U410 (N_410,In_88,In_680);
nor U411 (N_411,In_69,In_1153);
xnor U412 (N_412,In_1865,In_1860);
nand U413 (N_413,In_1179,In_1425);
xnor U414 (N_414,In_2031,In_1472);
and U415 (N_415,In_26,In_1592);
xor U416 (N_416,In_712,In_2169);
nor U417 (N_417,In_312,In_1929);
nand U418 (N_418,In_42,In_2007);
nand U419 (N_419,In_583,In_872);
and U420 (N_420,In_828,In_752);
or U421 (N_421,In_1424,In_638);
xnor U422 (N_422,In_1191,In_2019);
nand U423 (N_423,In_913,In_900);
nand U424 (N_424,In_274,In_2099);
or U425 (N_425,In_330,In_2168);
and U426 (N_426,In_2081,In_2309);
or U427 (N_427,In_505,In_1214);
xor U428 (N_428,In_1235,In_1853);
nand U429 (N_429,In_1418,In_1781);
nand U430 (N_430,In_1900,In_2156);
nand U431 (N_431,In_1975,In_649);
and U432 (N_432,In_910,In_1447);
and U433 (N_433,In_188,In_2205);
xor U434 (N_434,In_1333,In_1169);
and U435 (N_435,In_156,In_1939);
xor U436 (N_436,In_2202,In_371);
nand U437 (N_437,In_652,In_315);
and U438 (N_438,In_2185,In_1766);
nand U439 (N_439,In_308,In_1055);
nand U440 (N_440,In_1796,In_2339);
and U441 (N_441,In_982,In_1607);
or U442 (N_442,In_133,In_610);
nand U443 (N_443,In_1710,In_501);
xor U444 (N_444,In_1309,In_685);
xnor U445 (N_445,In_2206,In_1464);
and U446 (N_446,In_2418,In_2112);
nor U447 (N_447,In_1809,In_112);
or U448 (N_448,In_2119,In_1240);
xor U449 (N_449,In_1547,In_2219);
nor U450 (N_450,In_275,In_2247);
or U451 (N_451,In_2208,In_365);
and U452 (N_452,In_691,In_72);
xor U453 (N_453,In_413,In_581);
or U454 (N_454,In_1125,In_288);
nand U455 (N_455,In_1084,In_2495);
xor U456 (N_456,In_1793,In_2183);
xnor U457 (N_457,In_1321,In_1128);
nand U458 (N_458,In_1584,In_176);
nand U459 (N_459,In_1812,In_874);
or U460 (N_460,In_2210,In_1974);
and U461 (N_461,In_1245,In_191);
or U462 (N_462,In_43,In_1815);
xnor U463 (N_463,In_803,In_867);
nor U464 (N_464,In_1122,In_942);
and U465 (N_465,In_1127,In_2435);
and U466 (N_466,In_240,In_765);
nor U467 (N_467,In_1175,In_878);
and U468 (N_468,In_281,In_121);
nor U469 (N_469,In_1782,In_1532);
and U470 (N_470,In_2293,In_1533);
and U471 (N_471,In_1222,In_2204);
and U472 (N_472,In_245,In_1542);
nand U473 (N_473,In_1338,In_2182);
or U474 (N_474,In_1467,In_2097);
nand U475 (N_475,In_1161,In_1438);
or U476 (N_476,In_1348,In_455);
or U477 (N_477,In_1935,In_2370);
nand U478 (N_478,In_198,In_1722);
or U479 (N_479,In_1821,In_174);
and U480 (N_480,In_302,In_105);
nor U481 (N_481,In_859,In_730);
and U482 (N_482,In_2458,In_2485);
nand U483 (N_483,In_1304,In_390);
and U484 (N_484,In_515,In_1513);
nor U485 (N_485,In_673,In_933);
or U486 (N_486,In_235,In_2452);
xnor U487 (N_487,In_2303,In_2398);
nor U488 (N_488,In_2197,In_2062);
nor U489 (N_489,In_125,In_782);
nand U490 (N_490,In_1709,In_2402);
or U491 (N_491,In_1739,In_1497);
nand U492 (N_492,In_2474,In_2447);
xor U493 (N_493,In_1040,In_1630);
nand U494 (N_494,In_1732,In_1537);
or U495 (N_495,In_854,In_1827);
or U496 (N_496,In_1096,In_1361);
nand U497 (N_497,In_1095,In_2177);
xor U498 (N_498,In_213,In_1518);
and U499 (N_499,In_119,In_1312);
or U500 (N_500,In_2221,In_2428);
xnor U501 (N_501,N_262,In_18);
or U502 (N_502,In_2082,In_1093);
and U503 (N_503,In_2216,In_29);
xor U504 (N_504,In_2364,In_894);
nand U505 (N_505,In_1317,In_1292);
and U506 (N_506,N_330,In_8);
nand U507 (N_507,N_261,In_2250);
xor U508 (N_508,N_406,In_285);
nand U509 (N_509,N_98,In_1987);
xnor U510 (N_510,N_68,In_2049);
and U511 (N_511,In_1494,In_647);
nor U512 (N_512,In_372,N_90);
nor U513 (N_513,In_1440,N_59);
or U514 (N_514,In_1398,In_1967);
xnor U515 (N_515,In_2295,In_184);
or U516 (N_516,N_316,N_223);
nor U517 (N_517,In_1117,N_19);
nand U518 (N_518,N_88,N_97);
xor U519 (N_519,N_496,In_1953);
or U520 (N_520,In_1916,In_1198);
and U521 (N_521,In_1426,In_1423);
xnor U522 (N_522,In_1356,In_1875);
xor U523 (N_523,In_1166,In_816);
or U524 (N_524,In_2465,In_1017);
nand U525 (N_525,In_1664,In_1056);
nand U526 (N_526,In_1834,N_150);
and U527 (N_527,In_1346,In_2189);
or U528 (N_528,In_761,In_2178);
or U529 (N_529,In_1509,In_1604);
nor U530 (N_530,In_2167,N_39);
xor U531 (N_531,N_289,In_2285);
nand U532 (N_532,In_974,N_385);
xor U533 (N_533,N_38,In_2096);
nand U534 (N_534,In_2013,N_15);
xnor U535 (N_535,In_1403,In_1413);
nand U536 (N_536,In_2199,In_950);
nand U537 (N_537,In_169,In_6);
xnor U538 (N_538,In_1115,In_1241);
or U539 (N_539,In_1981,In_1404);
nor U540 (N_540,N_469,In_336);
xnor U541 (N_541,In_1970,In_1462);
nor U542 (N_542,N_335,In_97);
nor U543 (N_543,In_2072,N_193);
nand U544 (N_544,In_152,In_52);
or U545 (N_545,In_2427,In_278);
nand U546 (N_546,In_1508,In_1636);
xnor U547 (N_547,N_411,In_214);
xor U548 (N_548,In_741,In_2430);
nand U549 (N_549,In_932,N_456);
nand U550 (N_550,N_342,In_619);
nor U551 (N_551,In_253,In_2117);
or U552 (N_552,In_1803,In_682);
xnor U553 (N_553,In_2233,In_899);
or U554 (N_554,In_930,In_1181);
or U555 (N_555,N_485,In_560);
xnor U556 (N_556,N_336,In_1926);
or U557 (N_557,N_177,N_380);
or U558 (N_558,In_1689,N_35);
nor U559 (N_559,In_1652,In_2065);
and U560 (N_560,In_1611,In_1155);
nand U561 (N_561,In_871,In_490);
and U562 (N_562,In_1529,In_1507);
xor U563 (N_563,In_79,In_352);
or U564 (N_564,In_992,In_1296);
and U565 (N_565,In_1454,In_2335);
or U566 (N_566,In_1381,In_126);
nor U567 (N_567,N_477,In_205);
nor U568 (N_568,In_562,In_2336);
and U569 (N_569,In_2457,In_98);
or U570 (N_570,In_1593,In_267);
nand U571 (N_571,N_201,In_714);
or U572 (N_572,In_862,In_1382);
nor U573 (N_573,In_2437,In_664);
xor U574 (N_574,In_891,In_28);
or U575 (N_575,In_1544,In_283);
or U576 (N_576,N_283,N_102);
nand U577 (N_577,N_81,N_155);
xnor U578 (N_578,In_1535,N_26);
nand U579 (N_579,In_970,In_132);
xnor U580 (N_580,N_472,N_435);
or U581 (N_581,In_955,N_136);
and U582 (N_582,In_189,In_832);
nand U583 (N_583,N_227,N_44);
xnor U584 (N_584,In_1589,In_1103);
or U585 (N_585,In_2231,N_263);
or U586 (N_586,N_476,In_2286);
nor U587 (N_587,N_32,N_42);
nor U588 (N_588,In_1107,In_2203);
xor U589 (N_589,In_961,In_801);
or U590 (N_590,In_2282,In_656);
or U591 (N_591,In_147,In_2176);
nor U592 (N_592,In_355,In_778);
nor U593 (N_593,In_2024,N_204);
nand U594 (N_594,In_1489,In_287);
or U595 (N_595,In_1094,In_314);
nand U596 (N_596,In_829,In_2193);
and U597 (N_597,In_798,N_376);
or U598 (N_598,In_2145,N_494);
xor U599 (N_599,In_496,In_2462);
and U600 (N_600,In_918,In_526);
nor U601 (N_601,In_364,In_1046);
or U602 (N_602,In_877,N_224);
and U603 (N_603,In_956,In_1949);
nand U604 (N_604,In_559,In_2357);
and U605 (N_605,In_760,In_1100);
or U606 (N_606,N_270,In_1735);
xnor U607 (N_607,N_251,In_870);
and U608 (N_608,In_2320,In_2095);
and U609 (N_609,In_1081,In_486);
or U610 (N_610,In_1251,In_24);
nand U611 (N_611,In_1654,In_2259);
nand U612 (N_612,In_1194,In_484);
and U613 (N_613,In_2483,N_240);
or U614 (N_614,N_116,In_1202);
nor U615 (N_615,In_1086,In_2008);
xor U616 (N_616,In_138,In_1983);
nand U617 (N_617,In_1354,In_836);
nand U618 (N_618,N_171,In_460);
nand U619 (N_619,N_305,N_301);
and U620 (N_620,In_2278,In_1244);
xnor U621 (N_621,In_2461,In_2217);
or U622 (N_622,In_1666,In_1278);
nor U623 (N_623,N_25,In_2088);
and U624 (N_624,In_2372,In_663);
or U625 (N_625,N_236,N_87);
and U626 (N_626,N_50,In_2252);
nor U627 (N_627,In_1159,N_450);
nor U628 (N_628,In_837,In_2382);
xor U629 (N_629,In_1511,N_37);
xor U630 (N_630,In_1023,In_2078);
xor U631 (N_631,N_388,N_160);
or U632 (N_632,In_1750,In_2018);
nand U633 (N_633,In_1831,In_391);
xnor U634 (N_634,In_1303,In_686);
and U635 (N_635,In_217,In_973);
and U636 (N_636,In_149,N_429);
nand U637 (N_637,In_1973,In_2046);
or U638 (N_638,N_475,N_40);
or U639 (N_639,In_1250,In_2284);
or U640 (N_640,N_448,N_65);
or U641 (N_641,N_445,In_997);
and U642 (N_642,In_2069,In_1670);
xnor U643 (N_643,In_1026,N_51);
xor U644 (N_644,N_460,In_1248);
and U645 (N_645,N_410,In_2342);
nand U646 (N_646,In_2244,In_689);
nor U647 (N_647,In_1343,In_1680);
nand U648 (N_648,N_55,In_1581);
nand U649 (N_649,In_1862,In_165);
or U650 (N_650,In_2425,In_541);
and U651 (N_651,In_865,In_1332);
xor U652 (N_652,In_1075,N_378);
xnor U653 (N_653,In_713,In_1574);
or U654 (N_654,N_11,N_401);
nor U655 (N_655,N_311,In_1886);
nor U656 (N_656,In_124,In_2341);
or U657 (N_657,In_2179,In_2146);
and U658 (N_658,In_2209,In_140);
or U659 (N_659,In_709,In_1540);
and U660 (N_660,In_74,In_1092);
and U661 (N_661,In_842,In_2279);
or U662 (N_662,In_423,In_14);
and U663 (N_663,In_1712,In_1898);
xnor U664 (N_664,In_1456,N_174);
or U665 (N_665,In_1857,In_708);
and U666 (N_666,In_2027,N_161);
and U667 (N_667,In_1565,In_532);
xor U668 (N_668,In_886,In_1035);
nor U669 (N_669,In_153,In_509);
and U670 (N_670,In_1150,In_1595);
xnor U671 (N_671,In_66,In_1872);
nor U672 (N_672,In_363,In_584);
nand U673 (N_673,N_348,N_454);
and U674 (N_674,N_13,In_729);
or U675 (N_675,In_1742,N_396);
nor U676 (N_676,N_156,In_1436);
or U677 (N_677,In_573,In_940);
or U678 (N_678,N_416,In_2490);
xnor U679 (N_679,In_1389,In_2134);
and U680 (N_680,In_416,N_344);
nor U681 (N_681,In_1170,In_237);
nor U682 (N_682,N_182,In_1800);
nand U683 (N_683,In_774,In_449);
or U684 (N_684,In_1041,N_149);
and U685 (N_685,In_356,In_1648);
or U686 (N_686,N_151,In_748);
and U687 (N_687,In_12,In_1824);
nand U688 (N_688,In_1692,N_82);
nand U689 (N_689,In_1283,In_2412);
nand U690 (N_690,In_1613,In_322);
or U691 (N_691,In_2333,N_304);
or U692 (N_692,In_1658,N_5);
nor U693 (N_693,N_284,In_1661);
xor U694 (N_694,N_249,N_77);
nor U695 (N_695,In_2318,N_78);
or U696 (N_696,In_699,In_1083);
and U697 (N_697,In_350,In_1514);
and U698 (N_698,In_1757,In_2061);
nor U699 (N_699,N_157,In_557);
and U700 (N_700,In_1226,In_1861);
and U701 (N_701,In_523,In_2239);
nand U702 (N_702,In_1362,In_1344);
nor U703 (N_703,In_2108,In_2267);
xor U704 (N_704,In_1683,In_1556);
nor U705 (N_705,In_123,In_924);
and U706 (N_706,N_135,In_2480);
or U707 (N_707,N_268,In_616);
nor U708 (N_708,In_2011,In_1688);
and U709 (N_709,In_1879,N_196);
or U710 (N_710,In_1994,In_1058);
and U711 (N_711,In_2042,In_2455);
nand U712 (N_712,In_595,N_427);
nand U713 (N_713,In_1030,In_2289);
nand U714 (N_714,In_551,N_368);
xor U715 (N_715,N_455,In_1243);
and U716 (N_716,N_328,N_257);
and U717 (N_717,In_623,N_95);
and U718 (N_718,In_1470,In_876);
nand U719 (N_719,In_1366,In_2450);
nand U720 (N_720,N_369,In_1706);
and U721 (N_721,In_2366,In_2263);
nand U722 (N_722,In_805,In_221);
or U723 (N_723,In_781,N_382);
xor U724 (N_724,N_395,In_2020);
nor U725 (N_725,In_445,In_195);
and U726 (N_726,In_197,N_239);
nand U727 (N_727,In_2469,In_2463);
or U728 (N_728,N_269,In_520);
or U729 (N_729,In_1715,In_1538);
nand U730 (N_730,N_203,In_892);
xnor U731 (N_731,In_16,N_303);
xor U732 (N_732,In_1262,In_2);
and U733 (N_733,In_2122,In_1685);
nand U734 (N_734,N_139,In_1653);
nand U735 (N_735,N_233,In_2464);
nor U736 (N_736,In_475,In_1374);
xnor U737 (N_737,In_282,In_433);
or U738 (N_738,In_602,N_422);
xor U739 (N_739,In_513,In_1064);
or U740 (N_740,In_2230,In_1237);
nor U741 (N_741,In_31,In_2275);
or U742 (N_742,In_2349,In_441);
nand U743 (N_743,In_1359,In_218);
xnor U744 (N_744,In_1694,In_2073);
nand U745 (N_745,In_1165,In_342);
nand U746 (N_746,In_2258,In_1705);
and U747 (N_747,In_1531,In_1719);
nor U748 (N_748,In_841,In_1714);
or U749 (N_749,In_248,In_770);
xor U750 (N_750,In_2323,In_1287);
nor U751 (N_751,N_295,In_618);
xor U752 (N_752,In_2255,In_1363);
and U753 (N_753,N_22,N_57);
xor U754 (N_754,In_1482,In_1448);
nor U755 (N_755,In_458,In_2090);
or U756 (N_756,N_217,In_485);
and U757 (N_757,In_1612,N_190);
nor U758 (N_758,N_480,In_1698);
or U759 (N_759,In_678,In_1958);
or U760 (N_760,In_1805,In_258);
xnor U761 (N_761,In_1771,In_116);
or U762 (N_762,N_355,N_117);
nand U763 (N_763,N_64,In_819);
nand U764 (N_764,N_384,N_296);
xnor U765 (N_765,In_1176,In_62);
or U766 (N_766,In_1789,In_1024);
or U767 (N_767,In_2371,N_93);
xnor U768 (N_768,In_1871,In_630);
and U769 (N_769,N_219,In_2383);
and U770 (N_770,N_9,In_1154);
nand U771 (N_771,In_2363,In_2243);
nor U772 (N_772,In_2028,N_358);
and U773 (N_773,In_1780,In_497);
nand U774 (N_774,N_158,In_603);
xnor U775 (N_775,In_1776,In_1339);
nor U776 (N_776,In_1778,N_421);
xor U777 (N_777,N_471,In_2260);
and U778 (N_778,In_321,In_1899);
or U779 (N_779,In_357,N_320);
and U780 (N_780,In_1330,In_683);
or U781 (N_781,N_366,In_2487);
nand U782 (N_782,In_464,In_341);
and U783 (N_783,In_1414,In_1933);
xor U784 (N_784,In_1554,In_2343);
xor U785 (N_785,N_465,In_788);
nor U786 (N_786,N_83,In_78);
and U787 (N_787,In_401,N_17);
or U788 (N_788,N_120,In_1391);
nor U789 (N_789,N_488,In_935);
nor U790 (N_790,N_84,In_2115);
or U791 (N_791,In_2352,N_172);
nor U792 (N_792,N_271,In_2393);
nor U793 (N_793,In_2064,In_1074);
nor U794 (N_794,N_275,In_860);
and U795 (N_795,In_10,In_2470);
xor U796 (N_796,In_2374,In_180);
or U797 (N_797,N_423,In_896);
nand U798 (N_798,N_444,N_274);
nand U799 (N_799,N_447,In_2002);
and U800 (N_800,In_450,In_629);
nor U801 (N_801,In_53,In_2443);
and U802 (N_802,In_2296,In_303);
or U803 (N_803,In_1385,In_1982);
or U804 (N_804,N_247,N_357);
nor U805 (N_805,In_510,N_61);
nand U806 (N_806,In_606,In_2408);
nor U807 (N_807,In_21,In_1647);
and U808 (N_808,In_796,In_715);
nand U809 (N_809,In_1883,In_1943);
nor U810 (N_810,In_617,N_212);
or U811 (N_811,In_482,In_102);
or U812 (N_812,In_1474,N_392);
nor U813 (N_813,In_795,N_169);
or U814 (N_814,N_74,In_1297);
or U815 (N_815,In_1236,N_346);
and U816 (N_816,N_487,N_431);
nor U817 (N_817,N_205,In_2488);
nand U818 (N_818,N_122,In_1835);
and U819 (N_819,In_2433,In_1394);
xnor U820 (N_820,N_343,In_1326);
xor U821 (N_821,N_23,N_103);
nor U822 (N_822,N_391,In_2419);
or U823 (N_823,In_1102,N_459);
xor U824 (N_824,N_245,In_802);
and U825 (N_825,In_529,In_1037);
nand U826 (N_826,N_89,In_945);
and U827 (N_827,N_166,In_2144);
or U828 (N_828,N_314,In_1129);
or U829 (N_829,In_1443,In_1428);
and U830 (N_830,In_1039,In_1765);
and U831 (N_831,In_2326,In_817);
nor U832 (N_832,In_1785,In_2172);
xnor U833 (N_833,N_492,In_465);
and U834 (N_834,N_434,In_2010);
or U835 (N_835,In_1221,In_1290);
nand U836 (N_836,N_332,N_92);
xor U837 (N_837,In_2277,In_2087);
nor U838 (N_838,In_1152,In_154);
nand U839 (N_839,In_1106,In_2253);
and U840 (N_840,In_1741,In_2492);
xor U841 (N_841,N_360,In_807);
nor U842 (N_842,In_1477,N_162);
xnor U843 (N_843,In_1553,N_407);
xor U844 (N_844,In_547,In_1503);
nor U845 (N_845,N_367,In_2498);
nor U846 (N_846,N_153,In_2392);
and U847 (N_847,In_1408,In_46);
or U848 (N_848,N_474,In_437);
xnor U849 (N_849,In_2211,In_964);
nand U850 (N_850,In_646,In_1788);
and U851 (N_851,In_1936,In_199);
nand U852 (N_852,N_148,In_276);
nor U853 (N_853,In_2283,In_937);
xnor U854 (N_854,In_1784,In_61);
and U855 (N_855,In_1266,In_824);
nor U856 (N_856,In_1463,In_466);
nor U857 (N_857,In_426,N_114);
xnor U858 (N_858,N_441,N_402);
and U859 (N_859,In_2022,N_417);
xnor U860 (N_860,In_1485,In_1337);
or U861 (N_861,In_565,In_839);
xnor U862 (N_862,In_543,N_21);
or U863 (N_863,In_1364,In_2468);
nor U864 (N_864,In_1830,N_439);
nor U865 (N_865,N_467,N_244);
and U866 (N_866,In_1461,In_369);
xor U867 (N_867,In_620,N_66);
xnor U868 (N_868,In_164,In_568);
or U869 (N_869,In_954,In_1116);
and U870 (N_870,In_15,In_535);
and U871 (N_871,In_454,In_2220);
xnor U872 (N_872,In_1500,In_392);
xor U873 (N_873,In_2107,N_124);
nand U874 (N_874,N_18,In_1893);
xnor U875 (N_875,In_941,In_927);
and U876 (N_876,In_1738,In_665);
or U877 (N_877,In_1,In_1496);
nand U878 (N_878,In_943,In_724);
xnor U879 (N_879,N_106,In_2222);
xnor U880 (N_880,In_648,In_2181);
or U881 (N_881,In_1257,In_855);
xor U882 (N_882,In_1090,In_1434);
xor U883 (N_883,In_1758,In_2367);
or U884 (N_884,In_1568,N_318);
nor U885 (N_885,In_349,In_1307);
or U886 (N_886,N_243,In_224);
or U887 (N_887,In_480,In_2307);
and U888 (N_888,In_1844,N_307);
nor U889 (N_889,In_1880,In_609);
nor U890 (N_890,In_384,N_321);
nor U891 (N_891,In_348,N_256);
xor U892 (N_892,N_420,N_340);
and U893 (N_893,In_487,In_1849);
nor U894 (N_894,In_546,In_2332);
nor U895 (N_895,N_248,N_324);
xor U896 (N_896,N_315,In_434);
nand U897 (N_897,N_277,In_386);
and U898 (N_898,In_2009,In_1924);
and U899 (N_899,In_1925,In_1832);
nand U900 (N_900,In_1918,In_2200);
nor U901 (N_901,In_2417,In_1551);
nor U902 (N_902,In_1519,In_1693);
nor U903 (N_903,In_1761,In_1656);
xor U904 (N_904,In_926,In_106);
and U905 (N_905,In_904,In_514);
nor U906 (N_906,In_2155,In_99);
or U907 (N_907,In_2416,In_793);
nor U908 (N_908,In_533,In_1315);
and U909 (N_909,N_373,In_611);
and U910 (N_910,N_464,In_1059);
xnor U911 (N_911,In_776,N_110);
or U912 (N_912,In_1802,In_2409);
nor U913 (N_913,In_698,In_2422);
nor U914 (N_914,In_1877,In_1062);
nand U915 (N_915,N_10,In_1546);
xor U916 (N_916,In_2138,In_114);
nor U917 (N_917,N_310,N_222);
nand U918 (N_918,N_143,In_915);
xnor U919 (N_919,N_375,In_1615);
and U920 (N_920,In_269,In_662);
or U921 (N_921,In_1701,In_1668);
xnor U922 (N_922,N_176,In_531);
xor U923 (N_923,In_1138,In_856);
nor U924 (N_924,In_2249,In_958);
and U925 (N_925,In_1605,In_1968);
nand U926 (N_926,In_800,In_1318);
nand U927 (N_927,In_1869,In_1978);
nor U928 (N_928,In_743,In_849);
nand U929 (N_929,In_2045,N_430);
or U930 (N_930,In_1752,In_655);
or U931 (N_931,In_1946,In_200);
and U932 (N_932,In_1133,N_491);
or U933 (N_933,N_63,In_1896);
xor U934 (N_934,In_2396,N_409);
xnor U935 (N_935,In_1415,In_81);
nor U936 (N_936,In_1904,In_939);
nor U937 (N_937,In_1730,In_1220);
nand U938 (N_938,In_2266,In_279);
or U939 (N_939,In_2313,N_414);
and U940 (N_940,N_108,N_91);
nand U941 (N_941,In_949,In_1347);
nand U942 (N_942,In_1172,In_1621);
and U943 (N_943,In_77,N_399);
nor U944 (N_944,In_1238,N_178);
nand U945 (N_945,In_2390,In_1249);
nand U946 (N_946,In_1168,N_167);
nand U947 (N_947,In_1675,N_428);
and U948 (N_948,In_1979,In_917);
xor U949 (N_949,N_12,N_134);
and U950 (N_950,In_107,N_379);
and U951 (N_951,In_1025,In_794);
or U952 (N_952,In_504,N_453);
xor U953 (N_953,In_334,In_1618);
or U954 (N_954,In_749,N_131);
or U955 (N_955,In_2174,In_2076);
xor U956 (N_956,In_2306,In_34);
or U957 (N_957,In_521,In_2147);
xnor U958 (N_958,In_252,In_447);
and U959 (N_959,In_986,In_2070);
or U960 (N_960,N_404,In_1097);
xor U961 (N_961,In_226,In_909);
xor U962 (N_962,N_363,In_757);
or U963 (N_963,In_2454,In_1231);
or U964 (N_964,In_1148,In_727);
nor U965 (N_965,N_168,In_2157);
nor U966 (N_966,N_113,N_165);
nor U967 (N_967,In_2449,In_201);
and U968 (N_968,In_1015,In_1345);
nand U969 (N_969,In_171,N_393);
or U970 (N_970,In_2389,N_147);
nor U971 (N_971,In_1190,In_1770);
xor U972 (N_972,In_408,In_985);
nor U973 (N_973,In_2037,In_784);
xnor U974 (N_974,In_2355,In_1579);
xnor U975 (N_975,In_1913,In_2212);
xor U976 (N_976,In_2406,In_1567);
or U977 (N_977,In_1737,In_597);
nand U978 (N_978,In_110,N_229);
nor U979 (N_979,N_192,In_2491);
and U980 (N_980,In_811,In_1446);
nand U981 (N_981,In_1524,In_598);
xor U982 (N_982,N_1,In_2310);
or U983 (N_983,In_1136,In_1625);
nand U984 (N_984,In_104,In_2143);
or U985 (N_985,N_341,In_601);
xnor U986 (N_986,In_2271,In_290);
nand U987 (N_987,In_59,In_2223);
nor U988 (N_988,N_273,In_1253);
and U989 (N_989,N_30,In_1575);
xnor U990 (N_990,N_181,In_1624);
nand U991 (N_991,In_161,In_1667);
nor U992 (N_992,In_694,In_1189);
and U993 (N_993,In_567,In_1662);
or U994 (N_994,In_1976,In_210);
xor U995 (N_995,In_1572,In_1088);
nand U996 (N_996,In_440,In_1131);
and U997 (N_997,In_1308,In_1410);
or U998 (N_998,In_2004,In_2292);
and U999 (N_999,In_1442,N_325);
and U1000 (N_1000,N_706,In_2121);
or U1001 (N_1001,N_532,N_798);
or U1002 (N_1002,N_418,In_1007);
and U1003 (N_1003,In_1919,In_220);
nor U1004 (N_1004,N_911,In_1420);
nor U1005 (N_1005,N_919,In_1826);
and U1006 (N_1006,N_443,N_868);
and U1007 (N_1007,N_645,In_1263);
nor U1008 (N_1008,In_2466,In_1376);
nor U1009 (N_1009,N_468,N_322);
nor U1010 (N_1010,In_1811,N_896);
nor U1011 (N_1011,In_2358,N_505);
nand U1012 (N_1012,In_216,In_1971);
and U1013 (N_1013,N_125,In_2353);
nor U1014 (N_1014,N_976,In_2248);
xnor U1015 (N_1015,N_76,In_1637);
nand U1016 (N_1016,In_1073,In_296);
xnor U1017 (N_1017,N_853,N_512);
and U1018 (N_1018,In_1160,N_554);
xnor U1019 (N_1019,In_737,In_2085);
and U1020 (N_1020,In_1350,In_965);
and U1021 (N_1021,N_821,N_715);
nand U1022 (N_1022,N_990,N_216);
and U1023 (N_1023,In_1598,N_185);
nor U1024 (N_1024,N_985,In_328);
xor U1025 (N_1025,N_962,N_302);
nand U1026 (N_1026,In_2094,N_800);
or U1027 (N_1027,N_2,N_397);
and U1028 (N_1028,In_735,N_637);
nand U1029 (N_1029,N_7,N_924);
nor U1030 (N_1030,N_537,N_795);
nor U1031 (N_1031,N_931,N_56);
xor U1032 (N_1032,In_1295,N_662);
xnor U1033 (N_1033,N_510,N_534);
xnor U1034 (N_1034,N_940,N_914);
or U1035 (N_1035,N_734,N_721);
or U1036 (N_1036,In_1492,N_576);
nand U1037 (N_1037,N_290,N_702);
and U1038 (N_1038,In_1797,N_925);
and U1039 (N_1039,N_617,In_2173);
xnor U1040 (N_1040,In_193,N_438);
nor U1041 (N_1041,N_652,N_632);
nand U1042 (N_1042,N_901,N_85);
or U1043 (N_1043,In_580,N_426);
nand U1044 (N_1044,N_323,In_2257);
nor U1045 (N_1045,In_332,N_685);
or U1046 (N_1046,In_2190,N_881);
nor U1047 (N_1047,N_584,N_980);
nor U1048 (N_1048,In_1395,N_105);
and U1049 (N_1049,N_704,N_829);
xnor U1050 (N_1050,N_299,N_252);
or U1051 (N_1051,N_814,In_1622);
nand U1052 (N_1052,N_761,N_390);
nor U1053 (N_1053,N_747,In_1864);
and U1054 (N_1054,In_1594,In_206);
xor U1055 (N_1055,In_613,N_934);
xor U1056 (N_1056,In_1480,In_1417);
or U1057 (N_1057,In_1989,In_1938);
xor U1058 (N_1058,N_935,In_1052);
and U1059 (N_1059,In_626,N_954);
nor U1060 (N_1060,In_2106,In_326);
nor U1061 (N_1061,N_945,In_241);
or U1062 (N_1062,N_928,In_634);
and U1063 (N_1063,N_361,In_1566);
and U1064 (N_1064,N_973,N_623);
nor U1065 (N_1065,In_882,In_359);
or U1066 (N_1066,In_2486,N_571);
and U1067 (N_1067,N_939,In_255);
or U1068 (N_1068,N_479,N_717);
or U1069 (N_1069,In_234,N_834);
or U1070 (N_1070,In_1608,In_1602);
nor U1071 (N_1071,N_575,N_783);
and U1072 (N_1072,N_29,In_1219);
nor U1073 (N_1073,N_929,In_946);
nor U1074 (N_1074,N_70,In_1208);
nor U1075 (N_1075,N_278,N_350);
and U1076 (N_1076,N_107,N_180);
and U1077 (N_1077,N_878,N_164);
and U1078 (N_1078,N_956,In_739);
nand U1079 (N_1079,N_586,In_172);
xnor U1080 (N_1080,N_827,N_997);
xor U1081 (N_1081,N_432,N_692);
and U1082 (N_1082,In_1078,N_701);
and U1083 (N_1083,N_788,N_874);
or U1084 (N_1084,N_591,In_2369);
xor U1085 (N_1085,In_952,In_1585);
nor U1086 (N_1086,In_1204,N_633);
xor U1087 (N_1087,In_323,In_339);
nand U1088 (N_1088,In_1034,N_313);
xor U1089 (N_1089,N_607,In_1627);
and U1090 (N_1090,In_233,In_377);
or U1091 (N_1091,In_1884,In_1141);
xnor U1092 (N_1092,N_53,In_1268);
nor U1093 (N_1093,N_789,N_808);
nand U1094 (N_1094,N_6,In_47);
and U1095 (N_1095,N_540,In_309);
and U1096 (N_1096,N_944,N_354);
xnor U1097 (N_1097,In_1478,N_62);
or U1098 (N_1098,In_1351,N_173);
nor U1099 (N_1099,In_1915,N_631);
or U1100 (N_1100,N_927,In_305);
or U1101 (N_1101,N_75,N_923);
xor U1102 (N_1102,In_888,In_2126);
or U1103 (N_1103,N_543,N_833);
nand U1104 (N_1104,In_1852,N_894);
xor U1105 (N_1105,In_738,N_280);
nand U1106 (N_1106,In_1178,In_1124);
xor U1107 (N_1107,N_899,In_2431);
nand U1108 (N_1108,In_1515,In_1316);
nor U1109 (N_1109,N_394,In_118);
and U1110 (N_1110,In_1910,N_511);
nor U1111 (N_1111,N_16,In_1995);
nand U1112 (N_1112,N_913,N_41);
xnor U1113 (N_1113,In_2300,In_1744);
or U1114 (N_1114,In_643,In_1060);
and U1115 (N_1115,N_837,N_481);
xor U1116 (N_1116,In_887,N_836);
nand U1117 (N_1117,In_1679,N_958);
or U1118 (N_1118,In_1246,N_895);
nand U1119 (N_1119,In_1650,N_772);
nand U1120 (N_1120,In_117,In_491);
nor U1121 (N_1121,N_96,In_1291);
and U1122 (N_1122,In_542,In_2261);
and U1123 (N_1123,In_1130,In_1726);
and U1124 (N_1124,In_1433,In_948);
xnor U1125 (N_1125,N_977,In_631);
xnor U1126 (N_1126,N_142,In_473);
nand U1127 (N_1127,N_787,N_197);
nor U1128 (N_1128,N_626,In_247);
or U1129 (N_1129,N_767,N_383);
or U1130 (N_1130,N_746,In_1044);
nand U1131 (N_1131,N_792,N_889);
and U1132 (N_1132,N_991,N_200);
nor U1133 (N_1133,In_211,N_806);
and U1134 (N_1134,In_1109,N_415);
or U1135 (N_1135,In_1891,N_345);
nor U1136 (N_1136,N_984,In_1674);
xor U1137 (N_1137,N_649,N_844);
or U1138 (N_1138,N_194,In_651);
and U1139 (N_1139,N_920,In_848);
xnor U1140 (N_1140,In_2100,In_1786);
nor U1141 (N_1141,In_1799,In_301);
nand U1142 (N_1142,N_33,N_877);
or U1143 (N_1143,In_366,In_1273);
nand U1144 (N_1144,In_2287,N_115);
nand U1145 (N_1145,N_989,In_1021);
xor U1146 (N_1146,In_1923,In_2444);
xor U1147 (N_1147,In_229,In_1504);
or U1148 (N_1148,N_625,In_635);
nand U1149 (N_1149,In_2021,N_387);
or U1150 (N_1150,N_687,N_556);
xor U1151 (N_1151,In_2385,N_859);
xor U1152 (N_1152,In_120,N_565);
and U1153 (N_1153,In_633,In_659);
nand U1154 (N_1154,N_14,In_1110);
or U1155 (N_1155,In_306,N_777);
or U1156 (N_1156,In_736,In_2196);
and U1157 (N_1157,In_2241,In_868);
and U1158 (N_1158,N_762,In_1616);
and U1159 (N_1159,N_28,In_2361);
or U1160 (N_1160,In_1001,N_535);
nand U1161 (N_1161,In_1206,N_964);
or U1162 (N_1162,In_1213,In_1649);
or U1163 (N_1163,In_294,N_733);
or U1164 (N_1164,In_2344,N_530);
or U1165 (N_1165,N_862,In_704);
nand U1166 (N_1166,N_739,N_527);
xnor U1167 (N_1167,In_577,In_2276);
or U1168 (N_1168,In_1527,N_582);
nand U1169 (N_1169,In_1259,In_1516);
nor U1170 (N_1170,N_937,In_310);
nor U1171 (N_1171,In_688,In_2302);
nor U1172 (N_1172,In_1373,In_576);
nor U1173 (N_1173,In_1870,In_2476);
or U1174 (N_1174,In_787,N_187);
nor U1175 (N_1175,In_2380,In_879);
nor U1176 (N_1176,N_969,N_965);
and U1177 (N_1177,N_264,In_1847);
and U1178 (N_1178,N_831,N_525);
xor U1179 (N_1179,In_1013,In_815);
and U1180 (N_1180,N_971,N_442);
or U1181 (N_1181,In_1651,N_857);
xor U1182 (N_1182,N_882,N_669);
nand U1183 (N_1183,In_474,In_561);
nand U1184 (N_1184,In_538,N_765);
and U1185 (N_1185,In_1355,In_1265);
and U1186 (N_1186,In_1912,N_774);
nor U1187 (N_1187,In_344,N_559);
nand U1188 (N_1188,N_319,N_646);
nand U1189 (N_1189,In_2006,N_561);
xor U1190 (N_1190,N_842,N_757);
nand U1191 (N_1191,In_1963,In_1846);
or U1192 (N_1192,In_1406,In_530);
and U1193 (N_1193,In_1272,In_1952);
nor U1194 (N_1194,In_1199,N_339);
nor U1195 (N_1195,In_923,N_541);
and U1196 (N_1196,In_471,In_2213);
or U1197 (N_1197,N_672,In_2345);
nand U1198 (N_1198,N_291,N_728);
or U1199 (N_1199,N_654,N_809);
or U1200 (N_1200,N_941,In_1645);
or U1201 (N_1201,In_1111,N_784);
nor U1202 (N_1202,In_2125,N_386);
nor U1203 (N_1203,In_1951,N_546);
nor U1204 (N_1204,In_1412,N_67);
or U1205 (N_1205,N_823,N_689);
and U1206 (N_1206,In_636,In_1261);
nand U1207 (N_1207,N_292,In_1185);
and U1208 (N_1208,N_3,In_410);
or U1209 (N_1209,In_2033,In_1101);
nand U1210 (N_1210,N_916,N_966);
or U1211 (N_1211,In_552,N_604);
nand U1212 (N_1212,In_414,In_2051);
or U1213 (N_1213,In_1144,In_1379);
and U1214 (N_1214,In_999,N_817);
nor U1215 (N_1215,In_786,N_452);
nor U1216 (N_1216,In_2035,N_866);
or U1217 (N_1217,N_647,In_1063);
or U1218 (N_1218,N_111,N_628);
nand U1219 (N_1219,In_1791,In_814);
nand U1220 (N_1220,In_1495,N_907);
nor U1221 (N_1221,In_931,N_946);
nor U1222 (N_1222,N_128,N_666);
and U1223 (N_1223,In_605,N_745);
xnor U1224 (N_1224,In_1690,In_517);
xnor U1225 (N_1225,In_1033,N_752);
nand U1226 (N_1226,N_288,In_2133);
xor U1227 (N_1227,In_1920,In_2036);
or U1228 (N_1228,In_503,N_691);
xor U1229 (N_1229,In_2273,N_329);
xor U1230 (N_1230,N_267,In_1942);
or U1231 (N_1231,N_159,N_812);
xnor U1232 (N_1232,N_684,N_703);
xor U1233 (N_1233,In_1491,In_1965);
or U1234 (N_1234,In_1932,In_1873);
nand U1235 (N_1235,N_499,N_521);
and U1236 (N_1236,In_1858,N_749);
nor U1237 (N_1237,N_635,N_603);
and U1238 (N_1238,N_830,In_2166);
and U1239 (N_1239,In_772,In_884);
nor U1240 (N_1240,In_1432,N_695);
nor U1241 (N_1241,N_562,N_24);
nand U1242 (N_1242,In_340,N_531);
nand U1243 (N_1243,In_2346,In_1143);
nand U1244 (N_1244,N_446,N_548);
nand U1245 (N_1245,In_2290,N_848);
nor U1246 (N_1246,N_519,N_522);
xor U1247 (N_1247,N_760,N_80);
or U1248 (N_1248,N_839,N_594);
nor U1249 (N_1249,In_389,N_675);
nand U1250 (N_1250,N_936,In_375);
nor U1251 (N_1251,N_365,N_726);
xor U1252 (N_1252,N_807,In_429);
and U1253 (N_1253,In_50,N_755);
nor U1254 (N_1254,In_1633,In_1980);
or U1255 (N_1255,In_492,N_636);
or U1256 (N_1256,In_1032,N_599);
or U1257 (N_1257,N_364,In_700);
xnor U1258 (N_1258,In_1061,N_961);
nand U1259 (N_1259,In_49,In_1695);
xnor U1260 (N_1260,In_462,N_130);
and U1261 (N_1261,In_1271,In_1790);
or U1262 (N_1262,N_869,N_890);
xnor U1263 (N_1263,N_298,N_218);
xnor U1264 (N_1264,N_888,In_424);
nor U1265 (N_1265,N_146,In_396);
nor U1266 (N_1266,In_592,N_781);
and U1267 (N_1267,In_1543,In_2421);
nor U1268 (N_1268,N_568,In_2214);
xor U1269 (N_1269,N_744,N_208);
nand U1270 (N_1270,In_1009,N_419);
nor U1271 (N_1271,In_2359,N_738);
or U1272 (N_1272,N_668,N_679);
xor U1273 (N_1273,N_265,N_71);
nand U1274 (N_1274,N_898,In_2424);
nor U1275 (N_1275,N_912,In_1571);
xor U1276 (N_1276,In_2338,In_461);
nor U1277 (N_1277,In_2423,In_1227);
nor U1278 (N_1278,In_1928,In_830);
xor U1279 (N_1279,In_720,In_407);
and U1280 (N_1280,In_1126,In_558);
or U1281 (N_1281,N_211,N_566);
nor U1282 (N_1282,N_644,In_553);
nor U1283 (N_1283,In_508,N_572);
xor U1284 (N_1284,N_905,In_135);
or U1285 (N_1285,N_942,In_346);
or U1286 (N_1286,In_624,In_984);
nand U1287 (N_1287,In_1331,In_846);
xnor U1288 (N_1288,N_871,In_2153);
nand U1289 (N_1289,In_1247,N_611);
and U1290 (N_1290,N_563,N_780);
nor U1291 (N_1291,In_1897,In_1545);
and U1292 (N_1292,N_710,N_850);
nand U1293 (N_1293,N_308,N_595);
and U1294 (N_1294,In_1252,N_921);
and U1295 (N_1295,N_606,N_206);
or U1296 (N_1296,In_1031,In_1767);
xor U1297 (N_1297,In_393,N_520);
or U1298 (N_1298,N_873,In_2478);
xor U1299 (N_1299,In_702,N_822);
and U1300 (N_1300,N_786,In_621);
nand U1301 (N_1301,In_286,In_30);
nor U1302 (N_1302,In_549,N_209);
nand U1303 (N_1303,N_949,In_2399);
xnor U1304 (N_1304,In_1487,N_729);
or U1305 (N_1305,In_130,N_851);
and U1306 (N_1306,N_975,In_1908);
nor U1307 (N_1307,In_2052,N_732);
or U1308 (N_1308,N_605,N_104);
xor U1309 (N_1309,N_588,N_585);
nor U1310 (N_1310,N_838,N_616);
nor U1311 (N_1311,In_136,In_468);
xnor U1312 (N_1312,In_928,In_2171);
nand U1313 (N_1313,In_684,N_903);
and U1314 (N_1314,N_198,N_663);
or U1315 (N_1315,In_1223,In_2362);
and U1316 (N_1316,N_688,In_693);
and U1317 (N_1317,In_1539,N_841);
and U1318 (N_1318,N_673,N_993);
nor U1319 (N_1319,N_943,N_405);
nor U1320 (N_1320,N_722,N_226);
nand U1321 (N_1321,In_1753,N_758);
xnor U1322 (N_1322,In_44,In_1829);
nand U1323 (N_1323,N_819,In_537);
and U1324 (N_1324,In_944,In_1368);
and U1325 (N_1325,N_207,In_2236);
nor U1326 (N_1326,In_1171,In_1341);
nor U1327 (N_1327,In_1137,N_221);
or U1328 (N_1328,In_2132,N_129);
nor U1329 (N_1329,In_481,In_1663);
or U1330 (N_1330,In_215,N_791);
xnor U1331 (N_1331,N_545,In_1439);
nor U1332 (N_1332,N_589,In_25);
or U1333 (N_1333,N_883,N_815);
and U1334 (N_1334,In_1445,In_1964);
nand U1335 (N_1335,In_208,In_2154);
or U1336 (N_1336,In_1396,N_735);
nand U1337 (N_1337,In_773,In_1557);
xor U1338 (N_1338,N_716,N_579);
nor U1339 (N_1339,N_294,N_437);
or U1340 (N_1340,N_489,In_1731);
and U1341 (N_1341,N_658,N_690);
xor U1342 (N_1342,N_775,N_0);
nand U1343 (N_1343,N_119,In_1562);
xor U1344 (N_1344,N_331,N_47);
nand U1345 (N_1345,N_863,In_2191);
or U1346 (N_1346,In_1067,N_141);
nand U1347 (N_1347,In_1588,In_1450);
nand U1348 (N_1348,N_779,In_1700);
and U1349 (N_1349,N_858,N_737);
and U1350 (N_1350,N_707,In_1536);
nor U1351 (N_1351,N_138,N_686);
and U1352 (N_1352,N_213,In_2055);
and U1353 (N_1353,N_970,In_137);
or U1354 (N_1354,N_215,In_231);
xor U1355 (N_1355,N_457,N_253);
nor U1356 (N_1356,In_1828,N_759);
and U1357 (N_1357,In_880,In_1167);
nand U1358 (N_1358,In_1684,In_351);
xor U1359 (N_1359,In_1512,N_337);
or U1360 (N_1360,N_413,N_915);
nor U1361 (N_1361,In_144,N_680);
nor U1362 (N_1362,In_1972,N_816);
or U1363 (N_1363,In_362,N_408);
nand U1364 (N_1364,In_2405,N_979);
and U1365 (N_1365,N_794,In_324);
nor U1366 (N_1366,In_790,N_597);
and U1367 (N_1367,N_766,N_650);
nand U1368 (N_1368,In_479,N_458);
nand U1369 (N_1369,N_897,In_903);
xnor U1370 (N_1370,In_677,In_448);
nor U1371 (N_1371,N_58,In_869);
and U1372 (N_1372,N_598,N_232);
nor U1373 (N_1373,N_643,N_818);
xor U1374 (N_1374,In_1521,In_2159);
nand U1375 (N_1375,N_960,N_371);
nor U1376 (N_1376,In_851,In_642);
and U1377 (N_1377,N_225,In_1669);
nor U1378 (N_1378,In_54,N_656);
nand U1379 (N_1379,In_1118,In_2170);
nand U1380 (N_1380,N_547,N_933);
nand U1381 (N_1381,N_577,N_86);
and U1382 (N_1382,In_1270,N_552);
and U1383 (N_1383,N_720,In_1029);
xnor U1384 (N_1384,In_1558,N_988);
and U1385 (N_1385,N_938,In_1850);
nand U1386 (N_1386,In_1842,N_880);
xor U1387 (N_1387,N_718,N_484);
xor U1388 (N_1388,In_1569,N_214);
xnor U1389 (N_1389,N_667,In_2131);
xor U1390 (N_1390,N_123,N_356);
and U1391 (N_1391,N_891,N_43);
xor U1392 (N_1392,In_2240,In_670);
or U1393 (N_1393,In_1149,N_101);
nand U1394 (N_1394,In_1748,N_580);
nor U1395 (N_1395,In_338,N_152);
and U1396 (N_1396,In_2337,N_524);
nand U1397 (N_1397,N_188,In_27);
nand U1398 (N_1398,N_860,N_449);
nand U1399 (N_1399,In_73,In_744);
and U1400 (N_1400,In_2375,In_622);
nand U1401 (N_1401,N_189,N_992);
and U1402 (N_1402,N_618,N_697);
and U1403 (N_1403,In_162,In_2047);
nand U1404 (N_1404,N_678,In_2068);
or U1405 (N_1405,N_451,In_1264);
or U1406 (N_1406,In_820,In_1655);
xor U1407 (N_1407,In_1049,In_67);
nand U1408 (N_1408,In_1042,In_1961);
xnor U1409 (N_1409,In_425,In_661);
xor U1410 (N_1410,In_1819,In_1626);
xor U1411 (N_1411,N_503,In_1177);
nor U1412 (N_1412,N_237,N_549);
nor U1413 (N_1413,In_1856,N_854);
nor U1414 (N_1414,In_960,In_893);
nor U1415 (N_1415,N_705,N_660);
or U1416 (N_1416,In_979,In_754);
or U1417 (N_1417,N_509,N_309);
nand U1418 (N_1418,In_614,In_2377);
nor U1419 (N_1419,N_875,In_969);
nand U1420 (N_1420,N_998,N_529);
nand U1421 (N_1421,In_343,N_950);
nor U1422 (N_1422,N_242,In_1342);
nor U1423 (N_1423,In_1823,N_910);
nand U1424 (N_1424,N_539,N_900);
xor U1425 (N_1425,N_922,N_978);
or U1426 (N_1426,N_513,In_742);
and U1427 (N_1427,In_259,N_377);
xnor U1428 (N_1428,N_659,In_2039);
or U1429 (N_1429,In_1676,N_184);
nand U1430 (N_1430,In_1072,In_38);
and U1431 (N_1431,N_981,In_895);
or U1432 (N_1432,In_722,In_967);
or U1433 (N_1433,N_250,In_2386);
nor U1434 (N_1434,In_951,In_94);
xnor U1435 (N_1435,N_947,N_601);
nand U1436 (N_1436,N_255,N_764);
nand U1437 (N_1437,In_476,N_849);
nand U1438 (N_1438,N_466,N_374);
xor U1439 (N_1439,In_139,In_1279);
nand U1440 (N_1440,N_648,N_333);
nor U1441 (N_1441,N_664,N_154);
and U1442 (N_1442,In_563,N_968);
and U1443 (N_1443,N_796,In_2459);
nor U1444 (N_1444,In_645,In_246);
nor U1445 (N_1445,N_713,In_1367);
xor U1446 (N_1446,N_79,In_1888);
nor U1447 (N_1447,In_1068,In_1411);
xnor U1448 (N_1448,N_473,N_230);
nand U1449 (N_1449,In_804,In_1903);
nand U1450 (N_1450,In_2376,N_813);
nand U1451 (N_1451,N_754,In_718);
and U1452 (N_1452,In_345,N_653);
nor U1453 (N_1453,In_1486,N_573);
or U1454 (N_1454,In_843,N_258);
nand U1455 (N_1455,N_287,N_145);
nor U1456 (N_1456,N_100,In_1863);
xor U1457 (N_1457,N_996,In_845);
xor U1458 (N_1458,In_1643,N_482);
and U1459 (N_1459,N_655,In_2029);
nand U1460 (N_1460,In_780,In_2481);
or U1461 (N_1461,N_400,In_2445);
and U1462 (N_1462,N_506,N_486);
nor U1463 (N_1463,N_820,N_624);
and U1464 (N_1464,N_54,In_1229);
and U1465 (N_1465,In_1188,In_1498);
xor U1466 (N_1466,In_1549,In_1806);
or U1467 (N_1467,N_619,In_2456);
xor U1468 (N_1468,In_1917,N_478);
nor U1469 (N_1469,N_778,In_1911);
nand U1470 (N_1470,N_297,In_2379);
nand U1471 (N_1471,N_917,N_864);
nand U1472 (N_1472,N_629,In_347);
xor U1473 (N_1473,In_243,In_257);
xnor U1474 (N_1474,N_542,N_671);
xor U1475 (N_1475,In_1890,N_550);
nor U1476 (N_1476,In_381,N_948);
and U1477 (N_1477,N_276,In_1320);
xor U1478 (N_1478,In_1000,N_126);
or U1479 (N_1479,N_627,In_2023);
or U1480 (N_1480,In_1475,In_2043);
nor U1481 (N_1481,N_266,In_1927);
or U1482 (N_1482,N_285,N_564);
nor U1483 (N_1483,In_1016,N_334);
nor U1484 (N_1484,N_551,N_300);
or U1485 (N_1485,In_1195,N_403);
or U1486 (N_1486,N_771,In_833);
and U1487 (N_1487,N_677,N_389);
nor U1488 (N_1488,N_828,N_4);
or U1489 (N_1489,In_2067,N_536);
or U1490 (N_1490,In_1801,In_1600);
nand U1491 (N_1491,N_723,N_872);
and U1492 (N_1492,N_987,In_516);
nor U1493 (N_1493,N_926,In_1140);
and U1494 (N_1494,In_2294,In_1258);
and U1495 (N_1495,In_405,N_381);
nand U1496 (N_1496,In_1576,In_625);
or U1497 (N_1497,In_100,In_1139);
and U1498 (N_1498,N_507,N_740);
and U1499 (N_1499,In_1076,N_112);
or U1500 (N_1500,N_1254,N_1367);
nand U1501 (N_1501,N_699,N_802);
nor U1502 (N_1502,In_570,N_1210);
and U1503 (N_1503,In_2301,N_630);
nand U1504 (N_1504,N_1285,N_1426);
nand U1505 (N_1505,N_1260,N_843);
xor U1506 (N_1506,N_1319,N_1306);
and U1507 (N_1507,N_498,N_1247);
nand U1508 (N_1508,N_1339,N_832);
or U1509 (N_1509,N_1128,N_1373);
xnor U1510 (N_1510,N_338,In_1723);
and U1511 (N_1511,N_570,N_1114);
and U1512 (N_1512,In_587,In_297);
nand U1513 (N_1513,N_1343,N_845);
or U1514 (N_1514,In_444,N_1439);
xor U1515 (N_1515,N_1066,N_1147);
nor U1516 (N_1516,N_202,N_1376);
nand U1517 (N_1517,In_1874,N_1125);
and U1518 (N_1518,N_490,N_1124);
or U1519 (N_1519,In_711,N_500);
and U1520 (N_1520,In_1836,In_422);
nor U1521 (N_1521,N_1051,N_1059);
and U1522 (N_1522,In_51,N_1280);
nand U1523 (N_1523,N_1219,N_175);
xor U1524 (N_1524,N_855,N_1440);
nor U1525 (N_1525,In_1743,In_2105);
nand U1526 (N_1526,In_353,N_1459);
xnor U1527 (N_1527,N_516,N_220);
xor U1528 (N_1528,N_359,N_1305);
and U1529 (N_1529,N_670,N_1121);
and U1530 (N_1530,N_1052,In_1215);
xnor U1531 (N_1531,N_1437,N_1162);
nand U1532 (N_1532,N_1132,N_463);
nand U1533 (N_1533,N_953,N_681);
or U1534 (N_1534,N_1456,N_1360);
and U1535 (N_1535,N_370,N_1103);
or U1536 (N_1536,N_1235,N_1078);
and U1537 (N_1537,N_1488,N_1194);
or U1538 (N_1538,In_488,N_1169);
nor U1539 (N_1539,N_640,In_733);
xor U1540 (N_1540,In_1400,In_1577);
nand U1541 (N_1541,N_1113,N_1203);
and U1542 (N_1542,N_614,In_291);
nand U1543 (N_1543,N_1245,N_567);
nand U1544 (N_1544,N_885,N_1155);
and U1545 (N_1545,N_1045,N_1277);
or U1546 (N_1546,N_1095,N_1183);
or U1547 (N_1547,N_326,N_1093);
nor U1548 (N_1548,N_1393,N_693);
or U1549 (N_1549,In_2414,In_1892);
nand U1550 (N_1550,N_840,N_756);
xnor U1551 (N_1551,N_1071,N_959);
and U1552 (N_1552,N_1171,In_527);
xor U1553 (N_1553,In_1632,In_1123);
xor U1554 (N_1554,In_2234,In_1665);
nor U1555 (N_1555,N_708,N_1275);
nand U1556 (N_1556,N_1218,N_1083);
xnor U1557 (N_1557,N_1036,N_1436);
nor U1558 (N_1558,N_1386,N_1146);
xnor U1559 (N_1559,In_1182,N_1409);
nor U1560 (N_1560,N_1112,N_1214);
nand U1561 (N_1561,In_650,N_1279);
xor U1562 (N_1562,N_1272,In_36);
nor U1563 (N_1563,N_1332,N_1224);
or U1564 (N_1564,In_1028,N_199);
nand U1565 (N_1565,In_300,N_736);
or U1566 (N_1566,N_353,N_1384);
nand U1567 (N_1567,N_621,N_1359);
nand U1568 (N_1568,N_1023,N_1215);
xor U1569 (N_1569,In_159,In_212);
or U1570 (N_1570,N_1312,In_1145);
nand U1571 (N_1571,N_657,N_1079);
nor U1572 (N_1572,N_1227,N_1281);
and U1573 (N_1573,N_1133,In_853);
nor U1574 (N_1574,In_1708,N_1061);
and U1575 (N_1575,In_2135,N_501);
nand U1576 (N_1576,N_751,N_281);
nand U1577 (N_1577,In_1682,In_1838);
and U1578 (N_1578,In_1775,N_1418);
xnor U1579 (N_1579,N_1454,N_1148);
nand U1580 (N_1580,N_1447,N_1410);
or U1581 (N_1581,N_440,N_1388);
nor U1582 (N_1582,In_2116,In_2410);
nor U1583 (N_1583,N_52,N_1389);
nand U1584 (N_1584,N_1434,N_600);
or U1585 (N_1585,N_1407,N_1119);
or U1586 (N_1586,N_1471,N_1463);
or U1587 (N_1587,In_2050,In_906);
or U1588 (N_1588,N_1136,N_1152);
and U1589 (N_1589,N_725,In_1931);
nand U1590 (N_1590,N_1460,N_1018);
and U1591 (N_1591,N_1309,N_955);
xor U1592 (N_1592,In_779,N_1043);
and U1593 (N_1593,N_1381,N_1333);
xnor U1594 (N_1594,N_1302,N_1064);
nand U1595 (N_1595,N_1189,N_1187);
or U1596 (N_1596,N_1355,In_980);
xnor U1597 (N_1597,N_700,N_1361);
or U1598 (N_1598,In_2305,N_1118);
nand U1599 (N_1599,N_893,In_158);
and U1600 (N_1600,N_1056,In_1431);
nor U1601 (N_1601,N_1315,N_694);
and U1602 (N_1602,In_1377,N_665);
or U1603 (N_1603,N_1028,N_1458);
nand U1604 (N_1604,N_260,N_1241);
xor U1605 (N_1605,In_544,N_1427);
nor U1606 (N_1606,In_232,N_495);
or U1607 (N_1607,N_750,In_2180);
nor U1608 (N_1608,In_2270,N_1412);
and U1609 (N_1609,N_1009,N_1135);
nor U1610 (N_1610,N_1089,N_1140);
and U1611 (N_1611,N_1294,N_1259);
and U1612 (N_1612,N_1466,N_1200);
nor U1613 (N_1613,N_1423,N_1229);
nor U1614 (N_1614,N_1372,N_610);
xor U1615 (N_1615,N_1313,In_2077);
and U1616 (N_1616,N_518,N_1337);
nand U1617 (N_1617,N_1138,N_1480);
or U1618 (N_1618,In_1397,N_1461);
xnor U1619 (N_1619,In_534,N_1402);
or U1620 (N_1620,N_231,N_1347);
nand U1621 (N_1621,In_1242,N_1209);
nor U1622 (N_1622,N_1271,N_1230);
or U1623 (N_1623,N_1180,In_1051);
or U1624 (N_1624,In_7,In_1008);
nand U1625 (N_1625,In_1120,N_1398);
nor U1626 (N_1626,N_1211,N_109);
nand U1627 (N_1627,N_1462,N_569);
and U1628 (N_1628,N_696,In_705);
or U1629 (N_1629,N_712,N_1287);
nor U1630 (N_1630,In_1216,N_1340);
and U1631 (N_1631,N_1449,N_1428);
xor U1632 (N_1632,In_1114,In_2434);
or U1633 (N_1633,In_402,In_707);
and U1634 (N_1634,N_259,N_538);
nand U1635 (N_1635,N_1037,N_1293);
nand U1636 (N_1636,N_1493,In_1057);
or U1637 (N_1637,N_560,In_1087);
xor U1638 (N_1638,N_45,N_596);
xnor U1639 (N_1639,N_1476,N_1082);
and U1640 (N_1640,In_990,In_920);
nor U1641 (N_1641,In_1207,N_1295);
or U1642 (N_1642,N_824,In_2467);
nor U1643 (N_1643,N_1481,N_1442);
nand U1644 (N_1644,N_682,N_1318);
nor U1645 (N_1645,N_351,N_241);
nand U1646 (N_1646,N_1243,N_1134);
or U1647 (N_1647,N_1268,In_588);
nor U1648 (N_1648,N_1494,N_797);
xor U1649 (N_1649,In_2123,N_20);
xor U1650 (N_1650,In_1449,N_1199);
nand U1651 (N_1651,N_1429,In_512);
nand U1652 (N_1652,N_1097,In_1634);
xnor U1653 (N_1653,In_1868,N_1239);
nor U1654 (N_1654,N_639,N_362);
nor U1655 (N_1655,N_932,N_1068);
and U1656 (N_1656,N_742,N_312);
and U1657 (N_1657,N_1314,N_1350);
nand U1658 (N_1658,N_1242,In_1113);
nand U1659 (N_1659,N_1202,N_1212);
nand U1660 (N_1660,N_1363,N_1498);
nor U1661 (N_1661,N_69,In_873);
or U1662 (N_1662,In_1813,N_1048);
and U1663 (N_1663,N_553,N_1011);
nor U1664 (N_1664,N_908,N_1098);
and U1665 (N_1665,N_1477,In_821);
xnor U1666 (N_1666,In_823,In_1586);
nand U1667 (N_1667,N_801,N_317);
nand U1668 (N_1668,N_1266,In_2365);
and U1669 (N_1669,N_876,In_2420);
xor U1670 (N_1670,N_612,N_995);
nand U1671 (N_1671,N_1274,N_246);
nand U1672 (N_1672,N_1416,In_168);
and U1673 (N_1673,N_1006,N_1057);
xnor U1674 (N_1674,In_1080,N_1327);
or U1675 (N_1675,N_1117,In_785);
nand U1676 (N_1676,N_1484,In_768);
nor U1677 (N_1677,N_1222,N_1351);
xnor U1678 (N_1678,N_1374,In_555);
and U1679 (N_1679,N_210,N_1468);
and U1680 (N_1680,N_1489,N_1292);
and U1681 (N_1681,In_1419,N_982);
nor U1682 (N_1682,In_566,In_1818);
and U1683 (N_1683,N_578,N_1062);
or U1684 (N_1684,N_1120,N_1096);
xnor U1685 (N_1685,N_1478,In_1855);
nor U1686 (N_1686,N_1019,N_1054);
or U1687 (N_1687,N_1115,N_674);
xor U1688 (N_1688,N_847,N_502);
xnor U1689 (N_1689,N_1004,N_804);
and U1690 (N_1690,N_1411,N_1073);
and U1691 (N_1691,N_951,N_741);
nand U1692 (N_1692,N_1220,In_374);
and U1693 (N_1693,N_1300,In_90);
nand U1694 (N_1694,N_1326,N_835);
and U1695 (N_1695,In_1082,N_1137);
nand U1696 (N_1696,N_986,In_397);
xor U1697 (N_1697,N_1226,N_753);
nand U1698 (N_1698,In_1601,N_293);
or U1699 (N_1699,N_1040,N_1109);
xnor U1700 (N_1700,In_68,N_1485);
nor U1701 (N_1701,N_909,In_1003);
or U1702 (N_1702,N_886,In_1335);
xor U1703 (N_1703,In_998,N_719);
nor U1704 (N_1704,In_921,N_1065);
nor U1705 (N_1705,N_957,N_1086);
xor U1706 (N_1706,In_1762,N_782);
xor U1707 (N_1707,N_557,N_709);
xor U1708 (N_1708,N_1441,N_1238);
and U1709 (N_1709,N_1455,N_1025);
nand U1710 (N_1710,N_974,N_1186);
or U1711 (N_1711,N_228,In_1822);
and U1712 (N_1712,N_1362,N_186);
and U1713 (N_1713,In_103,N_1020);
xor U1714 (N_1714,N_1233,In_2139);
or U1715 (N_1715,N_1320,N_1173);
nor U1716 (N_1716,N_1403,N_555);
and U1717 (N_1717,N_1446,In_1085);
and U1718 (N_1718,N_1445,N_1432);
or U1719 (N_1719,N_526,N_1338);
nand U1720 (N_1720,N_1464,N_1021);
nor U1721 (N_1721,In_2129,In_142);
nor U1722 (N_1722,N_1365,In_1147);
nor U1723 (N_1723,In_1792,N_1284);
xnor U1724 (N_1724,N_1047,In_750);
or U1725 (N_1725,N_642,N_1364);
nand U1726 (N_1726,N_1151,N_1256);
nand U1727 (N_1727,N_514,N_1357);
nor U1728 (N_1728,In_1239,In_1336);
nor U1729 (N_1729,N_1005,N_1430);
xor U1730 (N_1730,N_1431,N_1107);
or U1731 (N_1731,N_1497,In_295);
nor U1732 (N_1732,N_1438,N_1076);
nor U1733 (N_1733,N_1190,N_1371);
xor U1734 (N_1734,N_793,In_2048);
nor U1735 (N_1735,In_1045,N_1131);
nand U1736 (N_1736,N_1049,N_902);
xor U1737 (N_1737,In_1352,N_1033);
nand U1738 (N_1738,N_1164,N_698);
or U1739 (N_1739,N_282,N_412);
and U1740 (N_1740,N_724,In_1833);
xor U1741 (N_1741,In_457,N_1221);
xor U1742 (N_1742,In_1721,N_234);
nor U1743 (N_1743,In_1276,N_1091);
nand U1744 (N_1744,N_811,In_196);
or U1745 (N_1745,N_1225,N_1198);
and U1746 (N_1746,In_3,In_1390);
and U1747 (N_1747,N_1424,N_1165);
and U1748 (N_1748,N_1067,In_1934);
nand U1749 (N_1749,N_856,N_352);
nand U1750 (N_1750,N_1090,N_1369);
and U1751 (N_1751,N_1335,N_558);
or U1752 (N_1752,In_0,N_1077);
nand U1753 (N_1753,N_1304,N_1491);
nand U1754 (N_1754,N_1324,In_230);
or U1755 (N_1755,N_1433,N_286);
nor U1756 (N_1756,In_1091,N_1144);
nand U1757 (N_1757,N_609,N_1094);
or U1758 (N_1758,N_508,N_1311);
or U1759 (N_1759,N_1153,N_805);
xnor U1760 (N_1760,In_640,N_1397);
nor U1761 (N_1761,N_1123,In_2330);
nor U1762 (N_1762,N_347,In_1777);
nor U1763 (N_1763,N_1046,N_622);
xor U1764 (N_1764,N_1316,N_1425);
nor U1765 (N_1765,N_1216,N_1334);
or U1766 (N_1766,N_730,N_1108);
or U1767 (N_1767,In_1977,In_1285);
xor U1768 (N_1768,N_1404,In_406);
nor U1769 (N_1769,N_1201,In_2354);
and U1770 (N_1770,In_608,N_1129);
or U1771 (N_1771,N_27,N_279);
or U1772 (N_1772,N_1443,N_1408);
and U1773 (N_1773,In_1550,N_1297);
nand U1774 (N_1774,N_1392,N_1141);
xnor U1775 (N_1775,N_1116,In_1997);
and U1776 (N_1776,N_1001,N_1263);
nand U1777 (N_1777,N_1378,In_2102);
xnor U1778 (N_1778,N_1007,N_1490);
nor U1779 (N_1779,N_1000,N_1400);
or U1780 (N_1780,N_424,N_651);
nand U1781 (N_1781,N_1396,N_1058);
nand U1782 (N_1782,N_195,N_714);
nand U1783 (N_1783,N_930,In_1848);
or U1784 (N_1784,N_768,N_887);
or U1785 (N_1785,N_590,In_472);
or U1786 (N_1786,N_1331,N_1329);
and U1787 (N_1787,N_1317,N_1237);
xor U1788 (N_1788,N_1496,In_1112);
xnor U1789 (N_1789,N_1448,In_2184);
nand U1790 (N_1790,N_1303,N_602);
xor U1791 (N_1791,N_1188,N_731);
nor U1792 (N_1792,In_2074,In_2152);
nor U1793 (N_1793,N_1008,N_1002);
xnor U1794 (N_1794,N_1253,N_790);
or U1795 (N_1795,N_1413,N_870);
nor U1796 (N_1796,In_48,N_127);
or U1797 (N_1797,N_1422,N_1479);
nor U1798 (N_1798,In_572,N_776);
nor U1799 (N_1799,N_398,In_1310);
nand U1800 (N_1800,N_94,N_1050);
xor U1801 (N_1801,In_2256,N_1204);
nand U1802 (N_1802,N_1264,N_1472);
and U1803 (N_1803,N_46,N_661);
xor U1804 (N_1804,N_1457,N_1348);
nand U1805 (N_1805,N_1358,N_1353);
and U1806 (N_1806,N_1487,N_504);
xor U1807 (N_1807,In_1769,N_770);
nand U1808 (N_1808,In_23,N_179);
or U1809 (N_1809,In_1473,N_1370);
and U1810 (N_1810,In_1205,In_361);
nor U1811 (N_1811,N_683,In_1294);
nor U1812 (N_1812,N_1127,N_1207);
nor U1813 (N_1813,In_385,In_1774);
xnor U1814 (N_1814,In_1599,N_121);
nand U1815 (N_1815,N_31,N_1228);
nand U1816 (N_1816,N_1088,In_1036);
nand U1817 (N_1817,N_1217,N_1349);
or U1818 (N_1818,In_1452,N_1055);
xnor U1819 (N_1819,N_1240,In_190);
nor U1820 (N_1820,N_1177,N_1296);
and U1821 (N_1821,In_1707,N_1232);
and U1822 (N_1822,N_1291,N_1039);
and U1823 (N_1823,N_852,N_1273);
or U1824 (N_1824,N_1383,N_170);
nor U1825 (N_1825,N_1139,N_1453);
nor U1826 (N_1826,N_1244,N_1026);
and U1827 (N_1827,N_349,N_1276);
or U1828 (N_1828,N_634,N_884);
xor U1829 (N_1829,N_1435,N_132);
nand U1830 (N_1830,N_1419,N_773);
nand U1831 (N_1831,In_875,N_1003);
xor U1832 (N_1832,N_1474,In_1407);
nand U1833 (N_1833,N_1181,N_983);
nor U1834 (N_1834,N_1012,N_1366);
nor U1835 (N_1835,N_1150,N_583);
nand U1836 (N_1836,N_1394,N_1070);
xor U1837 (N_1837,In_763,In_1984);
or U1838 (N_1838,In_2281,N_1346);
nand U1839 (N_1839,N_1044,N_879);
and U1840 (N_1840,N_528,N_1444);
or U1841 (N_1841,N_515,N_238);
nand U1842 (N_1842,In_2192,N_1236);
xor U1843 (N_1843,In_1380,N_799);
or U1844 (N_1844,N_436,In_1640);
and U1845 (N_1845,In_93,N_1015);
nand U1846 (N_1846,N_483,In_2127);
nor U1847 (N_1847,N_1197,N_865);
or U1848 (N_1848,N_1014,In_2162);
or U1849 (N_1849,N_1270,In_289);
nor U1850 (N_1850,In_1659,N_1341);
xor U1851 (N_1851,N_183,N_1100);
nor U1852 (N_1852,In_1749,N_1053);
nand U1853 (N_1853,In_2265,N_1246);
and U1854 (N_1854,N_1179,In_442);
xnor U1855 (N_1855,In_2496,In_1323);
nand U1856 (N_1856,N_1145,In_35);
nor U1857 (N_1857,N_1467,N_1031);
and U1858 (N_1858,N_1032,N_1328);
nor U1859 (N_1859,N_272,N_470);
nand U1860 (N_1860,N_517,In_703);
nand U1861 (N_1861,N_1385,In_13);
nand U1862 (N_1862,N_1368,N_1027);
nor U1863 (N_1863,N_1176,N_1074);
xnor U1864 (N_1864,N_1170,N_1105);
nor U1865 (N_1865,In_1203,In_1582);
nand U1866 (N_1866,N_1354,N_1414);
xor U1867 (N_1867,N_1261,In_360);
nand U1868 (N_1868,N_1377,N_620);
or U1869 (N_1869,N_1022,N_1161);
or U1870 (N_1870,In_2086,N_608);
xnor U1871 (N_1871,N_1106,N_1206);
or U1872 (N_1872,N_1182,N_1060);
xor U1873 (N_1873,N_1421,In_320);
xor U1874 (N_1874,In_679,N_1401);
nand U1875 (N_1875,N_163,N_60);
and U1876 (N_1876,In_2012,N_1175);
xnor U1877 (N_1877,In_1453,N_999);
or U1878 (N_1878,N_763,N_1307);
or U1879 (N_1879,N_118,N_1034);
nand U1880 (N_1880,N_861,In_799);
and U1881 (N_1881,N_1192,N_963);
nor U1882 (N_1882,In_2387,In_170);
or U1883 (N_1883,N_711,N_574);
nand U1884 (N_1884,N_846,In_1564);
or U1885 (N_1885,In_1993,N_1142);
nor U1886 (N_1886,N_1080,N_372);
xor U1887 (N_1887,N_1375,N_1234);
or U1888 (N_1888,N_327,N_254);
or U1889 (N_1889,N_73,N_1092);
nor U1890 (N_1890,In_65,In_1644);
xnor U1891 (N_1891,N_1249,In_2384);
and U1892 (N_1892,N_1030,N_1174);
xnor U1893 (N_1893,In_2161,In_1520);
and U1894 (N_1894,N_1063,N_1167);
and U1895 (N_1895,N_1016,N_1356);
xnor U1896 (N_1896,N_1072,N_1017);
nor U1897 (N_1897,In_511,N_1344);
and U1898 (N_1898,N_1085,N_1330);
and U1899 (N_1899,N_1486,N_1231);
nand U1900 (N_1900,In_1469,N_1160);
nor U1901 (N_1901,N_235,N_1417);
nor U1902 (N_1902,N_906,N_1159);
nand U1903 (N_1903,In_582,N_1168);
xor U1904 (N_1904,N_1122,N_1013);
nand U1905 (N_1905,In_1734,N_1166);
or U1906 (N_1906,N_1258,N_1391);
xor U1907 (N_1907,N_1325,N_137);
and U1908 (N_1908,N_904,In_1907);
nand U1909 (N_1909,In_1132,N_1492);
nand U1910 (N_1910,N_1157,In_1255);
and U1911 (N_1911,N_826,N_497);
or U1912 (N_1912,N_1149,N_1267);
or U1913 (N_1913,N_1101,N_1126);
xnor U1914 (N_1914,N_133,N_1390);
xnor U1915 (N_1915,N_638,N_803);
or U1916 (N_1916,In_1894,N_1380);
xnor U1917 (N_1917,In_1703,In_2201);
xor U1918 (N_1918,N_676,N_1099);
xor U1919 (N_1919,N_1255,In_2000);
and U1920 (N_1920,N_748,N_1041);
nor U1921 (N_1921,N_1395,In_2142);
nand U1922 (N_1922,In_2114,N_1475);
or U1923 (N_1923,N_1262,N_967);
and U1924 (N_1924,N_615,N_49);
nand U1925 (N_1925,N_1208,N_1499);
nor U1926 (N_1926,N_1158,N_1075);
or U1927 (N_1927,N_1310,In_740);
nand U1928 (N_1928,N_825,N_727);
nand U1929 (N_1929,N_1298,N_1382);
xnor U1930 (N_1930,N_1178,In_1465);
nor U1931 (N_1931,N_306,N_1248);
or U1932 (N_1932,In_354,N_918);
or U1933 (N_1933,N_1283,N_1290);
and U1934 (N_1934,N_1450,N_48);
and U1935 (N_1935,N_994,N_1193);
nand U1936 (N_1936,N_641,In_600);
and U1937 (N_1937,N_892,In_2484);
xor U1938 (N_1938,N_592,N_1191);
and U1939 (N_1939,N_1278,In_55);
xnor U1940 (N_1940,N_1282,N_1379);
and U1941 (N_1941,N_743,N_1387);
nor U1942 (N_1942,N_1185,N_1087);
nor U1943 (N_1943,N_544,N_1483);
and U1944 (N_1944,N_1196,N_1042);
nor U1945 (N_1945,N_1084,N_1405);
nor U1946 (N_1946,N_1163,In_1187);
and U1947 (N_1947,In_519,N_1289);
or U1948 (N_1948,N_1205,N_1286);
nor U1949 (N_1949,N_1482,In_494);
or U1950 (N_1950,N_8,N_593);
xor U1951 (N_1951,N_1473,N_1081);
and U1952 (N_1952,N_1470,N_533);
and U1953 (N_1953,N_462,In_994);
and U1954 (N_1954,N_1102,N_99);
or U1955 (N_1955,In_238,N_1250);
nor U1956 (N_1956,In_1603,N_144);
and U1957 (N_1957,In_767,N_1451);
and U1958 (N_1958,In_4,N_1038);
nor U1959 (N_1959,N_1399,N_1465);
and U1960 (N_1960,N_140,N_1223);
and U1961 (N_1961,N_587,N_1130);
nand U1962 (N_1962,In_254,In_2324);
or U1963 (N_1963,N_1104,N_461);
nand U1964 (N_1964,N_72,In_277);
nor U1965 (N_1965,N_425,In_185);
or U1966 (N_1966,N_523,N_36);
or U1967 (N_1967,N_1265,In_438);
nand U1968 (N_1968,N_1495,N_810);
nand U1969 (N_1969,In_756,N_1111);
and U1970 (N_1970,N_1469,N_1172);
and U1971 (N_1971,N_867,N_769);
nor U1972 (N_1972,N_1308,In_2327);
and U1973 (N_1973,N_952,N_1301);
or U1974 (N_1974,N_1452,N_1345);
nand U1975 (N_1975,N_1110,N_493);
and U1976 (N_1976,In_1587,N_1195);
or U1977 (N_1977,N_1321,N_785);
and U1978 (N_1978,In_1289,N_972);
nand U1979 (N_1979,N_1257,N_1251);
xnor U1980 (N_1980,N_1252,N_1035);
and U1981 (N_1981,N_1154,In_418);
xor U1982 (N_1982,In_2242,In_1954);
or U1983 (N_1983,N_1213,N_1143);
xor U1984 (N_1984,N_433,N_1323);
and U1985 (N_1985,In_637,N_191);
or U1986 (N_1986,N_1288,N_1299);
or U1987 (N_1987,N_1069,N_581);
nand U1988 (N_1988,In_1409,In_2436);
nor U1989 (N_1989,N_1406,N_1269);
nand U1990 (N_1990,N_1010,N_1184);
xor U1991 (N_1991,In_574,N_1336);
xnor U1992 (N_1992,In_2025,N_34);
nor U1993 (N_1993,In_2014,N_1342);
xnor U1994 (N_1994,In_1505,In_370);
nand U1995 (N_1995,N_1420,N_1322);
xor U1996 (N_1996,N_1156,N_1024);
nand U1997 (N_1997,N_613,N_1415);
nor U1998 (N_1998,In_95,N_1352);
xor U1999 (N_1999,In_912,N_1029);
xor U2000 (N_2000,N_1827,N_1925);
and U2001 (N_2001,N_1942,N_1924);
xor U2002 (N_2002,N_1722,N_1577);
and U2003 (N_2003,N_1703,N_1782);
nand U2004 (N_2004,N_1785,N_1652);
and U2005 (N_2005,N_1920,N_1730);
xor U2006 (N_2006,N_1616,N_1835);
nor U2007 (N_2007,N_1779,N_1916);
or U2008 (N_2008,N_1529,N_1644);
and U2009 (N_2009,N_1811,N_1661);
xnor U2010 (N_2010,N_1553,N_1767);
and U2011 (N_2011,N_1688,N_1950);
nand U2012 (N_2012,N_1989,N_1586);
nor U2013 (N_2013,N_1910,N_1649);
xor U2014 (N_2014,N_1755,N_1512);
xor U2015 (N_2015,N_1580,N_1506);
and U2016 (N_2016,N_1883,N_1682);
nor U2017 (N_2017,N_1640,N_1669);
and U2018 (N_2018,N_1843,N_1588);
nand U2019 (N_2019,N_1839,N_1711);
nand U2020 (N_2020,N_1760,N_1877);
nor U2021 (N_2021,N_1603,N_1706);
nand U2022 (N_2022,N_1845,N_1601);
nor U2023 (N_2023,N_1974,N_1765);
nand U2024 (N_2024,N_1898,N_1926);
or U2025 (N_2025,N_1545,N_1559);
nor U2026 (N_2026,N_1821,N_1912);
xnor U2027 (N_2027,N_1770,N_1733);
or U2028 (N_2028,N_1975,N_1977);
or U2029 (N_2029,N_1532,N_1502);
xor U2030 (N_2030,N_1987,N_1941);
xor U2031 (N_2031,N_1928,N_1995);
xor U2032 (N_2032,N_1943,N_1564);
xor U2033 (N_2033,N_1584,N_1746);
nor U2034 (N_2034,N_1768,N_1732);
or U2035 (N_2035,N_1582,N_1879);
xnor U2036 (N_2036,N_1880,N_1931);
nand U2037 (N_2037,N_1548,N_1633);
nor U2038 (N_2038,N_1922,N_1628);
nor U2039 (N_2039,N_1604,N_1761);
or U2040 (N_2040,N_1713,N_1969);
nand U2041 (N_2041,N_1766,N_1979);
xnor U2042 (N_2042,N_1812,N_1937);
and U2043 (N_2043,N_1986,N_1531);
and U2044 (N_2044,N_1677,N_1623);
or U2045 (N_2045,N_1596,N_1963);
xor U2046 (N_2046,N_1707,N_1508);
and U2047 (N_2047,N_1701,N_1824);
and U2048 (N_2048,N_1595,N_1650);
or U2049 (N_2049,N_1735,N_1891);
xor U2050 (N_2050,N_1547,N_1665);
and U2051 (N_2051,N_1918,N_1863);
nor U2052 (N_2052,N_1887,N_1791);
and U2053 (N_2053,N_1896,N_1878);
xnor U2054 (N_2054,N_1514,N_1959);
nand U2055 (N_2055,N_1727,N_1721);
or U2056 (N_2056,N_1541,N_1752);
and U2057 (N_2057,N_1555,N_1899);
nand U2058 (N_2058,N_1744,N_1729);
or U2059 (N_2059,N_1988,N_1865);
or U2060 (N_2060,N_1813,N_1855);
or U2061 (N_2061,N_1753,N_1662);
xnor U2062 (N_2062,N_1951,N_1698);
and U2063 (N_2063,N_1673,N_1993);
nand U2064 (N_2064,N_1687,N_1645);
and U2065 (N_2065,N_1803,N_1822);
nand U2066 (N_2066,N_1762,N_1915);
nor U2067 (N_2067,N_1589,N_1750);
nand U2068 (N_2068,N_1528,N_1807);
nor U2069 (N_2069,N_1696,N_1914);
and U2070 (N_2070,N_1873,N_1828);
and U2071 (N_2071,N_1534,N_1874);
nor U2072 (N_2072,N_1500,N_1780);
nand U2073 (N_2073,N_1776,N_1758);
xnor U2074 (N_2074,N_1519,N_1570);
or U2075 (N_2075,N_1881,N_1957);
nand U2076 (N_2076,N_1619,N_1647);
nand U2077 (N_2077,N_1850,N_1587);
nor U2078 (N_2078,N_1876,N_1714);
nor U2079 (N_2079,N_1909,N_1686);
xor U2080 (N_2080,N_1870,N_1799);
nor U2081 (N_2081,N_1820,N_1816);
or U2082 (N_2082,N_1819,N_1676);
and U2083 (N_2083,N_1903,N_1535);
nor U2084 (N_2084,N_1517,N_1683);
and U2085 (N_2085,N_1809,N_1970);
xor U2086 (N_2086,N_1771,N_1990);
or U2087 (N_2087,N_1728,N_1847);
and U2088 (N_2088,N_1886,N_1801);
nand U2089 (N_2089,N_1503,N_1756);
nor U2090 (N_2090,N_1818,N_1600);
and U2091 (N_2091,N_1788,N_1948);
xnor U2092 (N_2092,N_1884,N_1826);
xor U2093 (N_2093,N_1862,N_1726);
nand U2094 (N_2094,N_1932,N_1763);
nand U2095 (N_2095,N_1997,N_1590);
nand U2096 (N_2096,N_1594,N_1522);
nor U2097 (N_2097,N_1712,N_1907);
or U2098 (N_2098,N_1634,N_1515);
and U2099 (N_2099,N_1933,N_1944);
and U2100 (N_2100,N_1900,N_1579);
nand U2101 (N_2101,N_1663,N_1784);
or U2102 (N_2102,N_1895,N_1583);
xnor U2103 (N_2103,N_1613,N_1511);
nor U2104 (N_2104,N_1734,N_1953);
and U2105 (N_2105,N_1777,N_1978);
and U2106 (N_2106,N_1680,N_1653);
nor U2107 (N_2107,N_1550,N_1846);
xnor U2108 (N_2108,N_1591,N_1952);
and U2109 (N_2109,N_1982,N_1992);
or U2110 (N_2110,N_1834,N_1871);
xor U2111 (N_2111,N_1888,N_1911);
and U2112 (N_2112,N_1521,N_1804);
nor U2113 (N_2113,N_1983,N_1882);
nor U2114 (N_2114,N_1610,N_1815);
nor U2115 (N_2115,N_1792,N_1842);
xnor U2116 (N_2116,N_1832,N_1708);
or U2117 (N_2117,N_1852,N_1981);
nand U2118 (N_2118,N_1965,N_1674);
nor U2119 (N_2119,N_1923,N_1602);
xor U2120 (N_2120,N_1608,N_1643);
or U2121 (N_2121,N_1611,N_1741);
nand U2122 (N_2122,N_1538,N_1720);
or U2123 (N_2123,N_1985,N_1778);
and U2124 (N_2124,N_1539,N_1636);
nand U2125 (N_2125,N_1802,N_1930);
and U2126 (N_2126,N_1817,N_1738);
nor U2127 (N_2127,N_1569,N_1554);
xnor U2128 (N_2128,N_1516,N_1719);
nand U2129 (N_2129,N_1841,N_1556);
or U2130 (N_2130,N_1654,N_1549);
nand U2131 (N_2131,N_1617,N_1795);
nand U2132 (N_2132,N_1773,N_1858);
nand U2133 (N_2133,N_1501,N_1612);
nor U2134 (N_2134,N_1573,N_1849);
nand U2135 (N_2135,N_1660,N_1523);
xor U2136 (N_2136,N_1793,N_1805);
nand U2137 (N_2137,N_1690,N_1769);
nor U2138 (N_2138,N_1620,N_1798);
and U2139 (N_2139,N_1524,N_1646);
and U2140 (N_2140,N_1540,N_1851);
and U2141 (N_2141,N_1552,N_1685);
and U2142 (N_2142,N_1892,N_1599);
and U2143 (N_2143,N_1837,N_1631);
nor U2144 (N_2144,N_1743,N_1544);
and U2145 (N_2145,N_1679,N_1691);
or U2146 (N_2146,N_1921,N_1621);
nand U2147 (N_2147,N_1867,N_1838);
xor U2148 (N_2148,N_1991,N_1875);
or U2149 (N_2149,N_1563,N_1671);
or U2150 (N_2150,N_1794,N_1740);
nand U2151 (N_2151,N_1964,N_1973);
nand U2152 (N_2152,N_1833,N_1697);
nand U2153 (N_2153,N_1585,N_1861);
xor U2154 (N_2154,N_1605,N_1836);
xor U2155 (N_2155,N_1917,N_1935);
nor U2156 (N_2156,N_1764,N_1542);
xor U2157 (N_2157,N_1783,N_1592);
nor U2158 (N_2158,N_1560,N_1575);
nor U2159 (N_2159,N_1622,N_1715);
and U2160 (N_2160,N_1607,N_1618);
and U2161 (N_2161,N_1772,N_1614);
nand U2162 (N_2162,N_1533,N_1578);
and U2163 (N_2163,N_1906,N_1954);
or U2164 (N_2164,N_1615,N_1658);
nand U2165 (N_2165,N_1936,N_1872);
xor U2166 (N_2166,N_1681,N_1825);
and U2167 (N_2167,N_1551,N_1814);
or U2168 (N_2168,N_1642,N_1929);
xor U2169 (N_2169,N_1704,N_1630);
nand U2170 (N_2170,N_1968,N_1572);
nor U2171 (N_2171,N_1641,N_1913);
nor U2172 (N_2172,N_1561,N_1507);
or U2173 (N_2173,N_1657,N_1829);
nand U2174 (N_2174,N_1518,N_1731);
and U2175 (N_2175,N_1557,N_1939);
and U2176 (N_2176,N_1796,N_1999);
xor U2177 (N_2177,N_1574,N_1629);
or U2178 (N_2178,N_1624,N_1960);
or U2179 (N_2179,N_1510,N_1626);
or U2180 (N_2180,N_1684,N_1857);
nand U2181 (N_2181,N_1659,N_1702);
nand U2182 (N_2182,N_1505,N_1927);
xor U2183 (N_2183,N_1800,N_1971);
xnor U2184 (N_2184,N_1689,N_1759);
and U2185 (N_2185,N_1853,N_1961);
xnor U2186 (N_2186,N_1856,N_1692);
or U2187 (N_2187,N_1955,N_1513);
or U2188 (N_2188,N_1635,N_1894);
and U2189 (N_2189,N_1885,N_1797);
nand U2190 (N_2190,N_1566,N_1754);
or U2191 (N_2191,N_1958,N_1806);
or U2192 (N_2192,N_1725,N_1693);
nor U2193 (N_2193,N_1597,N_1568);
xnor U2194 (N_2194,N_1625,N_1775);
or U2195 (N_2195,N_1637,N_1742);
xnor U2196 (N_2196,N_1901,N_1994);
nor U2197 (N_2197,N_1530,N_1854);
or U2198 (N_2198,N_1748,N_1949);
or U2199 (N_2199,N_1904,N_1581);
and U2200 (N_2200,N_1716,N_1823);
or U2201 (N_2201,N_1695,N_1700);
or U2202 (N_2202,N_1576,N_1739);
nand U2203 (N_2203,N_1667,N_1868);
and U2204 (N_2204,N_1869,N_1786);
nor U2205 (N_2205,N_1908,N_1947);
nand U2206 (N_2206,N_1638,N_1831);
nor U2207 (N_2207,N_1724,N_1723);
xor U2208 (N_2208,N_1527,N_1709);
xnor U2209 (N_2209,N_1787,N_1745);
xor U2210 (N_2210,N_1789,N_1962);
xnor U2211 (N_2211,N_1938,N_1934);
nand U2212 (N_2212,N_1749,N_1537);
or U2213 (N_2213,N_1648,N_1980);
and U2214 (N_2214,N_1526,N_1546);
nand U2215 (N_2215,N_1830,N_1840);
xnor U2216 (N_2216,N_1810,N_1956);
and U2217 (N_2217,N_1897,N_1860);
nor U2218 (N_2218,N_1520,N_1639);
nor U2219 (N_2219,N_1844,N_1672);
and U2220 (N_2220,N_1565,N_1699);
xnor U2221 (N_2221,N_1632,N_1694);
or U2222 (N_2222,N_1774,N_1859);
xor U2223 (N_2223,N_1781,N_1946);
nand U2224 (N_2224,N_1593,N_1670);
and U2225 (N_2225,N_1998,N_1609);
or U2226 (N_2226,N_1790,N_1967);
nand U2227 (N_2227,N_1571,N_1664);
and U2228 (N_2228,N_1678,N_1717);
nor U2229 (N_2229,N_1627,N_1705);
and U2230 (N_2230,N_1558,N_1504);
or U2231 (N_2231,N_1889,N_1675);
nand U2232 (N_2232,N_1606,N_1890);
xnor U2233 (N_2233,N_1864,N_1736);
and U2234 (N_2234,N_1902,N_1718);
and U2235 (N_2235,N_1945,N_1525);
xnor U2236 (N_2236,N_1848,N_1893);
nand U2237 (N_2237,N_1808,N_1972);
nand U2238 (N_2238,N_1567,N_1866);
nor U2239 (N_2239,N_1757,N_1655);
and U2240 (N_2240,N_1940,N_1984);
nor U2241 (N_2241,N_1996,N_1976);
or U2242 (N_2242,N_1966,N_1710);
and U2243 (N_2243,N_1651,N_1656);
or U2244 (N_2244,N_1509,N_1536);
or U2245 (N_2245,N_1751,N_1668);
xor U2246 (N_2246,N_1562,N_1737);
or U2247 (N_2247,N_1543,N_1919);
nor U2248 (N_2248,N_1598,N_1666);
nor U2249 (N_2249,N_1905,N_1747);
and U2250 (N_2250,N_1505,N_1610);
and U2251 (N_2251,N_1992,N_1714);
and U2252 (N_2252,N_1744,N_1625);
or U2253 (N_2253,N_1578,N_1567);
nor U2254 (N_2254,N_1658,N_1536);
nand U2255 (N_2255,N_1764,N_1554);
and U2256 (N_2256,N_1897,N_1701);
xnor U2257 (N_2257,N_1897,N_1726);
nor U2258 (N_2258,N_1824,N_1719);
nor U2259 (N_2259,N_1799,N_1625);
nor U2260 (N_2260,N_1712,N_1519);
nand U2261 (N_2261,N_1938,N_1986);
and U2262 (N_2262,N_1639,N_1991);
nor U2263 (N_2263,N_1995,N_1619);
and U2264 (N_2264,N_1879,N_1659);
and U2265 (N_2265,N_1734,N_1755);
or U2266 (N_2266,N_1984,N_1590);
and U2267 (N_2267,N_1584,N_1698);
nand U2268 (N_2268,N_1787,N_1713);
nor U2269 (N_2269,N_1845,N_1738);
or U2270 (N_2270,N_1925,N_1608);
nor U2271 (N_2271,N_1525,N_1719);
xor U2272 (N_2272,N_1536,N_1635);
and U2273 (N_2273,N_1572,N_1663);
nand U2274 (N_2274,N_1795,N_1905);
nand U2275 (N_2275,N_1809,N_1683);
nor U2276 (N_2276,N_1544,N_1785);
or U2277 (N_2277,N_1996,N_1592);
or U2278 (N_2278,N_1696,N_1728);
and U2279 (N_2279,N_1722,N_1676);
xor U2280 (N_2280,N_1957,N_1931);
nor U2281 (N_2281,N_1851,N_1594);
and U2282 (N_2282,N_1562,N_1869);
nand U2283 (N_2283,N_1558,N_1738);
xnor U2284 (N_2284,N_1886,N_1748);
and U2285 (N_2285,N_1993,N_1800);
nor U2286 (N_2286,N_1530,N_1614);
nor U2287 (N_2287,N_1575,N_1661);
nor U2288 (N_2288,N_1839,N_1546);
nor U2289 (N_2289,N_1667,N_1539);
nor U2290 (N_2290,N_1566,N_1876);
nor U2291 (N_2291,N_1853,N_1557);
and U2292 (N_2292,N_1600,N_1904);
nor U2293 (N_2293,N_1757,N_1661);
nand U2294 (N_2294,N_1995,N_1984);
nor U2295 (N_2295,N_1730,N_1747);
nor U2296 (N_2296,N_1712,N_1759);
nand U2297 (N_2297,N_1693,N_1814);
xnor U2298 (N_2298,N_1524,N_1890);
nand U2299 (N_2299,N_1887,N_1762);
nor U2300 (N_2300,N_1909,N_1985);
xnor U2301 (N_2301,N_1523,N_1879);
xnor U2302 (N_2302,N_1890,N_1649);
or U2303 (N_2303,N_1552,N_1573);
nor U2304 (N_2304,N_1634,N_1848);
xor U2305 (N_2305,N_1896,N_1744);
xnor U2306 (N_2306,N_1833,N_1973);
nand U2307 (N_2307,N_1636,N_1511);
xnor U2308 (N_2308,N_1717,N_1961);
nand U2309 (N_2309,N_1571,N_1972);
or U2310 (N_2310,N_1710,N_1896);
nor U2311 (N_2311,N_1990,N_1531);
xor U2312 (N_2312,N_1914,N_1993);
nand U2313 (N_2313,N_1722,N_1772);
xnor U2314 (N_2314,N_1723,N_1517);
nand U2315 (N_2315,N_1917,N_1648);
nor U2316 (N_2316,N_1648,N_1549);
nor U2317 (N_2317,N_1561,N_1559);
nand U2318 (N_2318,N_1680,N_1789);
nand U2319 (N_2319,N_1890,N_1544);
or U2320 (N_2320,N_1934,N_1866);
and U2321 (N_2321,N_1519,N_1995);
or U2322 (N_2322,N_1726,N_1762);
xor U2323 (N_2323,N_1829,N_1640);
nand U2324 (N_2324,N_1677,N_1723);
or U2325 (N_2325,N_1913,N_1816);
nand U2326 (N_2326,N_1776,N_1640);
nor U2327 (N_2327,N_1952,N_1610);
nand U2328 (N_2328,N_1620,N_1654);
or U2329 (N_2329,N_1782,N_1977);
and U2330 (N_2330,N_1998,N_1650);
or U2331 (N_2331,N_1543,N_1572);
and U2332 (N_2332,N_1969,N_1516);
and U2333 (N_2333,N_1663,N_1692);
and U2334 (N_2334,N_1851,N_1793);
xor U2335 (N_2335,N_1840,N_1786);
or U2336 (N_2336,N_1587,N_1941);
xnor U2337 (N_2337,N_1957,N_1659);
xor U2338 (N_2338,N_1580,N_1668);
or U2339 (N_2339,N_1583,N_1645);
or U2340 (N_2340,N_1746,N_1591);
xor U2341 (N_2341,N_1561,N_1844);
xnor U2342 (N_2342,N_1977,N_1579);
nand U2343 (N_2343,N_1860,N_1854);
or U2344 (N_2344,N_1648,N_1889);
xnor U2345 (N_2345,N_1874,N_1823);
nor U2346 (N_2346,N_1861,N_1532);
and U2347 (N_2347,N_1512,N_1764);
or U2348 (N_2348,N_1809,N_1746);
nor U2349 (N_2349,N_1560,N_1558);
nand U2350 (N_2350,N_1889,N_1639);
or U2351 (N_2351,N_1760,N_1741);
nand U2352 (N_2352,N_1589,N_1724);
xor U2353 (N_2353,N_1637,N_1980);
nor U2354 (N_2354,N_1895,N_1963);
or U2355 (N_2355,N_1734,N_1823);
or U2356 (N_2356,N_1730,N_1974);
or U2357 (N_2357,N_1855,N_1927);
nor U2358 (N_2358,N_1602,N_1920);
xnor U2359 (N_2359,N_1859,N_1788);
nor U2360 (N_2360,N_1511,N_1560);
xor U2361 (N_2361,N_1931,N_1502);
nor U2362 (N_2362,N_1720,N_1952);
xor U2363 (N_2363,N_1938,N_1988);
or U2364 (N_2364,N_1706,N_1683);
or U2365 (N_2365,N_1546,N_1785);
xnor U2366 (N_2366,N_1778,N_1820);
or U2367 (N_2367,N_1723,N_1743);
and U2368 (N_2368,N_1638,N_1510);
and U2369 (N_2369,N_1914,N_1856);
xor U2370 (N_2370,N_1587,N_1702);
xor U2371 (N_2371,N_1598,N_1985);
nand U2372 (N_2372,N_1949,N_1769);
or U2373 (N_2373,N_1897,N_1936);
or U2374 (N_2374,N_1845,N_1684);
nor U2375 (N_2375,N_1965,N_1643);
or U2376 (N_2376,N_1718,N_1669);
xor U2377 (N_2377,N_1912,N_1657);
or U2378 (N_2378,N_1742,N_1739);
nor U2379 (N_2379,N_1595,N_1641);
nand U2380 (N_2380,N_1812,N_1729);
nor U2381 (N_2381,N_1682,N_1748);
nand U2382 (N_2382,N_1501,N_1747);
or U2383 (N_2383,N_1799,N_1982);
xor U2384 (N_2384,N_1859,N_1931);
and U2385 (N_2385,N_1652,N_1774);
nand U2386 (N_2386,N_1801,N_1684);
xor U2387 (N_2387,N_1585,N_1685);
xor U2388 (N_2388,N_1575,N_1797);
and U2389 (N_2389,N_1555,N_1919);
nand U2390 (N_2390,N_1743,N_1855);
nor U2391 (N_2391,N_1566,N_1516);
nor U2392 (N_2392,N_1883,N_1806);
xor U2393 (N_2393,N_1728,N_1573);
nand U2394 (N_2394,N_1803,N_1892);
or U2395 (N_2395,N_1858,N_1559);
nand U2396 (N_2396,N_1512,N_1650);
nand U2397 (N_2397,N_1845,N_1602);
and U2398 (N_2398,N_1765,N_1911);
and U2399 (N_2399,N_1707,N_1721);
and U2400 (N_2400,N_1836,N_1700);
nand U2401 (N_2401,N_1965,N_1683);
nor U2402 (N_2402,N_1602,N_1521);
xor U2403 (N_2403,N_1858,N_1736);
nand U2404 (N_2404,N_1623,N_1506);
xnor U2405 (N_2405,N_1665,N_1863);
or U2406 (N_2406,N_1978,N_1573);
nor U2407 (N_2407,N_1515,N_1541);
nand U2408 (N_2408,N_1834,N_1518);
and U2409 (N_2409,N_1829,N_1553);
or U2410 (N_2410,N_1548,N_1906);
xnor U2411 (N_2411,N_1541,N_1511);
xor U2412 (N_2412,N_1812,N_1916);
nor U2413 (N_2413,N_1849,N_1606);
xnor U2414 (N_2414,N_1701,N_1796);
and U2415 (N_2415,N_1527,N_1855);
nand U2416 (N_2416,N_1611,N_1790);
nand U2417 (N_2417,N_1519,N_1888);
or U2418 (N_2418,N_1766,N_1761);
xnor U2419 (N_2419,N_1570,N_1523);
nand U2420 (N_2420,N_1993,N_1782);
or U2421 (N_2421,N_1968,N_1822);
and U2422 (N_2422,N_1517,N_1666);
or U2423 (N_2423,N_1501,N_1593);
nor U2424 (N_2424,N_1886,N_1639);
nor U2425 (N_2425,N_1712,N_1973);
nor U2426 (N_2426,N_1884,N_1528);
nand U2427 (N_2427,N_1595,N_1981);
nor U2428 (N_2428,N_1788,N_1770);
and U2429 (N_2429,N_1784,N_1823);
and U2430 (N_2430,N_1562,N_1511);
or U2431 (N_2431,N_1681,N_1814);
xor U2432 (N_2432,N_1823,N_1666);
xor U2433 (N_2433,N_1924,N_1688);
or U2434 (N_2434,N_1788,N_1986);
and U2435 (N_2435,N_1655,N_1726);
or U2436 (N_2436,N_1591,N_1709);
nand U2437 (N_2437,N_1805,N_1921);
nor U2438 (N_2438,N_1901,N_1646);
xor U2439 (N_2439,N_1992,N_1770);
or U2440 (N_2440,N_1863,N_1728);
nor U2441 (N_2441,N_1651,N_1559);
nor U2442 (N_2442,N_1996,N_1506);
nor U2443 (N_2443,N_1809,N_1637);
and U2444 (N_2444,N_1510,N_1945);
xnor U2445 (N_2445,N_1801,N_1919);
or U2446 (N_2446,N_1893,N_1960);
nand U2447 (N_2447,N_1871,N_1680);
nand U2448 (N_2448,N_1774,N_1715);
and U2449 (N_2449,N_1737,N_1888);
or U2450 (N_2450,N_1601,N_1897);
or U2451 (N_2451,N_1638,N_1737);
nand U2452 (N_2452,N_1695,N_1967);
or U2453 (N_2453,N_1737,N_1747);
nand U2454 (N_2454,N_1519,N_1719);
or U2455 (N_2455,N_1951,N_1585);
nor U2456 (N_2456,N_1728,N_1987);
and U2457 (N_2457,N_1898,N_1502);
or U2458 (N_2458,N_1643,N_1525);
nor U2459 (N_2459,N_1785,N_1661);
and U2460 (N_2460,N_1945,N_1681);
nand U2461 (N_2461,N_1943,N_1616);
nand U2462 (N_2462,N_1754,N_1611);
nand U2463 (N_2463,N_1667,N_1979);
or U2464 (N_2464,N_1796,N_1976);
nor U2465 (N_2465,N_1817,N_1678);
or U2466 (N_2466,N_1720,N_1540);
nor U2467 (N_2467,N_1543,N_1666);
nand U2468 (N_2468,N_1993,N_1971);
and U2469 (N_2469,N_1729,N_1943);
nor U2470 (N_2470,N_1517,N_1811);
and U2471 (N_2471,N_1724,N_1578);
nor U2472 (N_2472,N_1598,N_1527);
nor U2473 (N_2473,N_1891,N_1699);
nand U2474 (N_2474,N_1739,N_1712);
nor U2475 (N_2475,N_1543,N_1569);
nor U2476 (N_2476,N_1683,N_1872);
nor U2477 (N_2477,N_1566,N_1537);
and U2478 (N_2478,N_1757,N_1734);
or U2479 (N_2479,N_1979,N_1988);
or U2480 (N_2480,N_1938,N_1930);
nand U2481 (N_2481,N_1576,N_1717);
nand U2482 (N_2482,N_1608,N_1548);
or U2483 (N_2483,N_1656,N_1555);
xnor U2484 (N_2484,N_1614,N_1789);
nand U2485 (N_2485,N_1815,N_1934);
xnor U2486 (N_2486,N_1935,N_1711);
xnor U2487 (N_2487,N_1511,N_1976);
nand U2488 (N_2488,N_1604,N_1596);
and U2489 (N_2489,N_1984,N_1584);
nor U2490 (N_2490,N_1735,N_1911);
or U2491 (N_2491,N_1852,N_1688);
nand U2492 (N_2492,N_1802,N_1923);
xor U2493 (N_2493,N_1831,N_1835);
xor U2494 (N_2494,N_1691,N_1730);
nor U2495 (N_2495,N_1910,N_1721);
or U2496 (N_2496,N_1755,N_1673);
and U2497 (N_2497,N_1994,N_1987);
xnor U2498 (N_2498,N_1922,N_1718);
and U2499 (N_2499,N_1596,N_1788);
nor U2500 (N_2500,N_2181,N_2112);
and U2501 (N_2501,N_2089,N_2020);
xor U2502 (N_2502,N_2275,N_2459);
nand U2503 (N_2503,N_2005,N_2482);
and U2504 (N_2504,N_2335,N_2364);
nor U2505 (N_2505,N_2220,N_2159);
or U2506 (N_2506,N_2341,N_2077);
or U2507 (N_2507,N_2237,N_2344);
xor U2508 (N_2508,N_2455,N_2195);
nor U2509 (N_2509,N_2417,N_2423);
xor U2510 (N_2510,N_2067,N_2481);
nand U2511 (N_2511,N_2118,N_2037);
nand U2512 (N_2512,N_2492,N_2257);
xnor U2513 (N_2513,N_2078,N_2437);
xnor U2514 (N_2514,N_2291,N_2164);
nor U2515 (N_2515,N_2125,N_2249);
and U2516 (N_2516,N_2169,N_2352);
nand U2517 (N_2517,N_2387,N_2337);
xor U2518 (N_2518,N_2011,N_2122);
and U2519 (N_2519,N_2339,N_2041);
nor U2520 (N_2520,N_2436,N_2120);
or U2521 (N_2521,N_2449,N_2177);
xnor U2522 (N_2522,N_2151,N_2204);
nand U2523 (N_2523,N_2231,N_2404);
nor U2524 (N_2524,N_2248,N_2408);
and U2525 (N_2525,N_2150,N_2199);
nand U2526 (N_2526,N_2106,N_2167);
nor U2527 (N_2527,N_2245,N_2384);
xnor U2528 (N_2528,N_2431,N_2025);
nor U2529 (N_2529,N_2072,N_2496);
or U2530 (N_2530,N_2043,N_2215);
and U2531 (N_2531,N_2466,N_2317);
and U2532 (N_2532,N_2185,N_2175);
and U2533 (N_2533,N_2391,N_2308);
and U2534 (N_2534,N_2079,N_2233);
and U2535 (N_2535,N_2448,N_2226);
or U2536 (N_2536,N_2196,N_2017);
xor U2537 (N_2537,N_2161,N_2359);
and U2538 (N_2538,N_2109,N_2447);
or U2539 (N_2539,N_2211,N_2365);
and U2540 (N_2540,N_2414,N_2439);
nand U2541 (N_2541,N_2411,N_2480);
and U2542 (N_2542,N_2224,N_2193);
or U2543 (N_2543,N_2280,N_2055);
and U2544 (N_2544,N_2474,N_2093);
xnor U2545 (N_2545,N_2056,N_2381);
xor U2546 (N_2546,N_2018,N_2462);
nand U2547 (N_2547,N_2091,N_2052);
nor U2548 (N_2548,N_2194,N_2172);
xnor U2549 (N_2549,N_2367,N_2271);
nand U2550 (N_2550,N_2269,N_2475);
nor U2551 (N_2551,N_2267,N_2494);
nand U2552 (N_2552,N_2034,N_2350);
and U2553 (N_2553,N_2342,N_2213);
xnor U2554 (N_2554,N_2398,N_2351);
or U2555 (N_2555,N_2382,N_2485);
xor U2556 (N_2556,N_2242,N_2454);
nor U2557 (N_2557,N_2386,N_2318);
nor U2558 (N_2558,N_2276,N_2004);
nand U2559 (N_2559,N_2489,N_2453);
xnor U2560 (N_2560,N_2148,N_2299);
nor U2561 (N_2561,N_2336,N_2095);
nor U2562 (N_2562,N_2380,N_2297);
nor U2563 (N_2563,N_2324,N_2060);
or U2564 (N_2564,N_2035,N_2377);
or U2565 (N_2565,N_2006,N_2426);
and U2566 (N_2566,N_2187,N_2478);
nor U2567 (N_2567,N_2288,N_2270);
nand U2568 (N_2568,N_2107,N_2303);
nor U2569 (N_2569,N_2457,N_2073);
or U2570 (N_2570,N_2312,N_2320);
nand U2571 (N_2571,N_2057,N_2154);
or U2572 (N_2572,N_2407,N_2424);
and U2573 (N_2573,N_2027,N_2302);
and U2574 (N_2574,N_2446,N_2273);
xnor U2575 (N_2575,N_2397,N_2100);
nand U2576 (N_2576,N_2110,N_2098);
nand U2577 (N_2577,N_2022,N_2493);
nor U2578 (N_2578,N_2463,N_2498);
nor U2579 (N_2579,N_2197,N_2347);
or U2580 (N_2580,N_2393,N_2038);
xor U2581 (N_2581,N_2495,N_2266);
or U2582 (N_2582,N_2126,N_2117);
nand U2583 (N_2583,N_2029,N_2223);
or U2584 (N_2584,N_2346,N_2389);
or U2585 (N_2585,N_2392,N_2068);
xor U2586 (N_2586,N_2241,N_2047);
nand U2587 (N_2587,N_2450,N_2321);
xnor U2588 (N_2588,N_2063,N_2418);
and U2589 (N_2589,N_2311,N_2395);
or U2590 (N_2590,N_2435,N_2401);
or U2591 (N_2591,N_2296,N_2440);
xnor U2592 (N_2592,N_2086,N_2180);
xor U2593 (N_2593,N_2028,N_2064);
or U2594 (N_2594,N_2071,N_2059);
xor U2595 (N_2595,N_2490,N_2253);
nand U2596 (N_2596,N_2420,N_2357);
or U2597 (N_2597,N_2258,N_2385);
nand U2598 (N_2598,N_2157,N_2430);
and U2599 (N_2599,N_2042,N_2274);
or U2600 (N_2600,N_2268,N_2353);
and U2601 (N_2601,N_2158,N_2132);
nand U2602 (N_2602,N_2069,N_2304);
or U2603 (N_2603,N_2306,N_2023);
nand U2604 (N_2604,N_2040,N_2484);
nor U2605 (N_2605,N_2432,N_2198);
or U2606 (N_2606,N_2309,N_2356);
nor U2607 (N_2607,N_2143,N_2243);
xnor U2608 (N_2608,N_2121,N_2111);
xor U2609 (N_2609,N_2421,N_2247);
xor U2610 (N_2610,N_2104,N_2039);
nor U2611 (N_2611,N_2166,N_2092);
xnor U2612 (N_2612,N_2360,N_2255);
xor U2613 (N_2613,N_2176,N_2217);
nand U2614 (N_2614,N_2192,N_2183);
nand U2615 (N_2615,N_2066,N_2434);
or U2616 (N_2616,N_2433,N_2361);
nand U2617 (N_2617,N_2378,N_2085);
nor U2618 (N_2618,N_2225,N_2234);
nand U2619 (N_2619,N_2218,N_2451);
nand U2620 (N_2620,N_2103,N_2445);
nand U2621 (N_2621,N_2244,N_2230);
or U2622 (N_2622,N_2141,N_2477);
and U2623 (N_2623,N_2331,N_2413);
or U2624 (N_2624,N_2470,N_2390);
nor U2625 (N_2625,N_2368,N_2362);
nor U2626 (N_2626,N_2314,N_2102);
xnor U2627 (N_2627,N_2239,N_2191);
and U2628 (N_2628,N_2232,N_2240);
xnor U2629 (N_2629,N_2338,N_2115);
nor U2630 (N_2630,N_2214,N_2153);
or U2631 (N_2631,N_2062,N_2082);
and U2632 (N_2632,N_2021,N_2313);
xnor U2633 (N_2633,N_2116,N_2205);
nand U2634 (N_2634,N_2024,N_2476);
and U2635 (N_2635,N_2400,N_2328);
nor U2636 (N_2636,N_2010,N_2325);
or U2637 (N_2637,N_2284,N_2486);
or U2638 (N_2638,N_2155,N_2108);
xor U2639 (N_2639,N_2083,N_2371);
xnor U2640 (N_2640,N_2383,N_2044);
nand U2641 (N_2641,N_2399,N_2084);
nor U2642 (N_2642,N_2265,N_2332);
nand U2643 (N_2643,N_2003,N_2229);
xnor U2644 (N_2644,N_2053,N_2429);
and U2645 (N_2645,N_2279,N_2139);
xnor U2646 (N_2646,N_2261,N_2354);
or U2647 (N_2647,N_2287,N_2412);
and U2648 (N_2648,N_2416,N_2129);
and U2649 (N_2649,N_2286,N_2045);
nor U2650 (N_2650,N_2075,N_2236);
and U2651 (N_2651,N_2008,N_2212);
nor U2652 (N_2652,N_2301,N_2097);
and U2653 (N_2653,N_2326,N_2219);
or U2654 (N_2654,N_2419,N_2246);
nor U2655 (N_2655,N_2144,N_2305);
nor U2656 (N_2656,N_2184,N_2322);
nand U2657 (N_2657,N_2171,N_2259);
xor U2658 (N_2658,N_2165,N_2210);
xor U2659 (N_2659,N_2127,N_2054);
xor U2660 (N_2660,N_2329,N_2289);
and U2661 (N_2661,N_2469,N_2379);
nand U2662 (N_2662,N_2295,N_2315);
nand U2663 (N_2663,N_2394,N_2460);
nand U2664 (N_2664,N_2163,N_2124);
nand U2665 (N_2665,N_2049,N_2088);
xor U2666 (N_2666,N_2499,N_2442);
nor U2667 (N_2667,N_2099,N_2479);
nand U2668 (N_2668,N_2014,N_2061);
or U2669 (N_2669,N_2019,N_2456);
xor U2670 (N_2670,N_2428,N_2000);
nor U2671 (N_2671,N_2156,N_2349);
xor U2672 (N_2672,N_2441,N_2094);
nand U2673 (N_2673,N_2189,N_2202);
or U2674 (N_2674,N_2458,N_2050);
nand U2675 (N_2675,N_2178,N_2396);
and U2676 (N_2676,N_2058,N_2119);
nor U2677 (N_2677,N_2030,N_2201);
nor U2678 (N_2678,N_2190,N_2323);
or U2679 (N_2679,N_2491,N_2046);
nand U2680 (N_2680,N_2101,N_2468);
nor U2681 (N_2681,N_2036,N_2471);
xor U2682 (N_2682,N_2009,N_2294);
or U2683 (N_2683,N_2162,N_2473);
xor U2684 (N_2684,N_2128,N_2300);
nand U2685 (N_2685,N_2130,N_2376);
nor U2686 (N_2686,N_2374,N_2188);
xnor U2687 (N_2687,N_2012,N_2281);
xnor U2688 (N_2688,N_2452,N_2260);
or U2689 (N_2689,N_2209,N_2307);
or U2690 (N_2690,N_2327,N_2403);
or U2691 (N_2691,N_2174,N_2007);
nand U2692 (N_2692,N_2207,N_2142);
xor U2693 (N_2693,N_2074,N_2070);
and U2694 (N_2694,N_2203,N_2206);
xnor U2695 (N_2695,N_2222,N_2032);
and U2696 (N_2696,N_2227,N_2254);
xnor U2697 (N_2697,N_2427,N_2031);
and U2698 (N_2698,N_2136,N_2415);
and U2699 (N_2699,N_2370,N_2298);
xor U2700 (N_2700,N_2497,N_2051);
or U2701 (N_2701,N_2179,N_2355);
nand U2702 (N_2702,N_2147,N_2114);
and U2703 (N_2703,N_2422,N_2334);
or U2704 (N_2704,N_2256,N_2087);
and U2705 (N_2705,N_2221,N_2013);
xor U2706 (N_2706,N_2366,N_2373);
xor U2707 (N_2707,N_2145,N_2293);
nand U2708 (N_2708,N_2002,N_2467);
nor U2709 (N_2709,N_2105,N_2410);
or U2710 (N_2710,N_2251,N_2425);
nand U2711 (N_2711,N_2016,N_2369);
nor U2712 (N_2712,N_2330,N_2443);
nor U2713 (N_2713,N_2090,N_2292);
nor U2714 (N_2714,N_2081,N_2152);
or U2715 (N_2715,N_2080,N_2133);
nor U2716 (N_2716,N_2472,N_2488);
nand U2717 (N_2717,N_2113,N_2208);
nor U2718 (N_2718,N_2388,N_2487);
xnor U2719 (N_2719,N_2228,N_2015);
nand U2720 (N_2720,N_2149,N_2001);
or U2721 (N_2721,N_2343,N_2316);
xor U2722 (N_2722,N_2444,N_2134);
xnor U2723 (N_2723,N_2252,N_2263);
nand U2724 (N_2724,N_2358,N_2235);
and U2725 (N_2725,N_2186,N_2283);
nand U2726 (N_2726,N_2076,N_2402);
xnor U2727 (N_2727,N_2048,N_2406);
xnor U2728 (N_2728,N_2216,N_2135);
and U2729 (N_2729,N_2170,N_2096);
nor U2730 (N_2730,N_2464,N_2465);
xnor U2731 (N_2731,N_2272,N_2173);
and U2732 (N_2732,N_2200,N_2140);
and U2733 (N_2733,N_2123,N_2277);
xnor U2734 (N_2734,N_2138,N_2264);
nor U2735 (N_2735,N_2282,N_2290);
or U2736 (N_2736,N_2319,N_2262);
nor U2737 (N_2737,N_2137,N_2409);
xnor U2738 (N_2738,N_2310,N_2065);
nand U2739 (N_2739,N_2278,N_2285);
and U2740 (N_2740,N_2250,N_2348);
nand U2741 (N_2741,N_2160,N_2372);
and U2742 (N_2742,N_2182,N_2026);
xor U2743 (N_2743,N_2340,N_2438);
or U2744 (N_2744,N_2168,N_2146);
nand U2745 (N_2745,N_2333,N_2461);
xnor U2746 (N_2746,N_2375,N_2405);
or U2747 (N_2747,N_2363,N_2483);
nand U2748 (N_2748,N_2345,N_2238);
nor U2749 (N_2749,N_2131,N_2033);
nor U2750 (N_2750,N_2130,N_2152);
and U2751 (N_2751,N_2478,N_2405);
nand U2752 (N_2752,N_2412,N_2151);
xor U2753 (N_2753,N_2324,N_2264);
nand U2754 (N_2754,N_2221,N_2026);
and U2755 (N_2755,N_2344,N_2149);
and U2756 (N_2756,N_2157,N_2019);
nor U2757 (N_2757,N_2040,N_2394);
nand U2758 (N_2758,N_2035,N_2098);
or U2759 (N_2759,N_2353,N_2281);
and U2760 (N_2760,N_2022,N_2144);
xor U2761 (N_2761,N_2207,N_2196);
and U2762 (N_2762,N_2182,N_2002);
or U2763 (N_2763,N_2274,N_2074);
nand U2764 (N_2764,N_2408,N_2122);
and U2765 (N_2765,N_2131,N_2000);
nor U2766 (N_2766,N_2400,N_2441);
nor U2767 (N_2767,N_2347,N_2402);
nor U2768 (N_2768,N_2071,N_2063);
xnor U2769 (N_2769,N_2329,N_2303);
nand U2770 (N_2770,N_2164,N_2426);
xnor U2771 (N_2771,N_2232,N_2394);
nand U2772 (N_2772,N_2334,N_2042);
nand U2773 (N_2773,N_2241,N_2075);
or U2774 (N_2774,N_2212,N_2241);
or U2775 (N_2775,N_2261,N_2412);
or U2776 (N_2776,N_2499,N_2460);
nor U2777 (N_2777,N_2344,N_2083);
xnor U2778 (N_2778,N_2358,N_2228);
nand U2779 (N_2779,N_2477,N_2013);
nor U2780 (N_2780,N_2067,N_2290);
and U2781 (N_2781,N_2419,N_2302);
nand U2782 (N_2782,N_2153,N_2380);
nand U2783 (N_2783,N_2141,N_2249);
and U2784 (N_2784,N_2469,N_2086);
or U2785 (N_2785,N_2439,N_2278);
nor U2786 (N_2786,N_2418,N_2337);
nor U2787 (N_2787,N_2322,N_2206);
or U2788 (N_2788,N_2478,N_2231);
and U2789 (N_2789,N_2273,N_2150);
and U2790 (N_2790,N_2380,N_2086);
and U2791 (N_2791,N_2347,N_2473);
or U2792 (N_2792,N_2352,N_2219);
nor U2793 (N_2793,N_2095,N_2313);
and U2794 (N_2794,N_2047,N_2418);
and U2795 (N_2795,N_2331,N_2373);
nor U2796 (N_2796,N_2210,N_2356);
xnor U2797 (N_2797,N_2490,N_2155);
nand U2798 (N_2798,N_2125,N_2322);
nand U2799 (N_2799,N_2164,N_2334);
nand U2800 (N_2800,N_2352,N_2093);
nand U2801 (N_2801,N_2389,N_2140);
and U2802 (N_2802,N_2202,N_2055);
or U2803 (N_2803,N_2322,N_2070);
or U2804 (N_2804,N_2182,N_2449);
nor U2805 (N_2805,N_2297,N_2213);
xnor U2806 (N_2806,N_2366,N_2180);
nor U2807 (N_2807,N_2043,N_2076);
and U2808 (N_2808,N_2107,N_2141);
or U2809 (N_2809,N_2182,N_2218);
and U2810 (N_2810,N_2000,N_2254);
nor U2811 (N_2811,N_2077,N_2220);
or U2812 (N_2812,N_2474,N_2380);
xnor U2813 (N_2813,N_2467,N_2093);
or U2814 (N_2814,N_2327,N_2098);
and U2815 (N_2815,N_2254,N_2288);
nor U2816 (N_2816,N_2237,N_2026);
xor U2817 (N_2817,N_2048,N_2231);
or U2818 (N_2818,N_2253,N_2039);
or U2819 (N_2819,N_2364,N_2356);
nand U2820 (N_2820,N_2351,N_2347);
nor U2821 (N_2821,N_2330,N_2046);
or U2822 (N_2822,N_2192,N_2048);
nand U2823 (N_2823,N_2408,N_2339);
nor U2824 (N_2824,N_2238,N_2365);
nor U2825 (N_2825,N_2033,N_2245);
and U2826 (N_2826,N_2236,N_2370);
xnor U2827 (N_2827,N_2281,N_2376);
and U2828 (N_2828,N_2048,N_2252);
xor U2829 (N_2829,N_2266,N_2138);
or U2830 (N_2830,N_2374,N_2171);
xnor U2831 (N_2831,N_2112,N_2213);
and U2832 (N_2832,N_2256,N_2466);
xnor U2833 (N_2833,N_2442,N_2025);
or U2834 (N_2834,N_2390,N_2220);
xor U2835 (N_2835,N_2423,N_2029);
or U2836 (N_2836,N_2248,N_2033);
or U2837 (N_2837,N_2497,N_2016);
or U2838 (N_2838,N_2484,N_2027);
xor U2839 (N_2839,N_2383,N_2425);
xor U2840 (N_2840,N_2100,N_2159);
and U2841 (N_2841,N_2188,N_2275);
nor U2842 (N_2842,N_2050,N_2066);
and U2843 (N_2843,N_2287,N_2365);
and U2844 (N_2844,N_2174,N_2350);
or U2845 (N_2845,N_2268,N_2043);
nor U2846 (N_2846,N_2163,N_2370);
xnor U2847 (N_2847,N_2432,N_2042);
and U2848 (N_2848,N_2342,N_2499);
or U2849 (N_2849,N_2114,N_2001);
and U2850 (N_2850,N_2364,N_2198);
nor U2851 (N_2851,N_2491,N_2187);
and U2852 (N_2852,N_2056,N_2236);
nand U2853 (N_2853,N_2329,N_2030);
xnor U2854 (N_2854,N_2033,N_2351);
or U2855 (N_2855,N_2213,N_2441);
or U2856 (N_2856,N_2363,N_2089);
xnor U2857 (N_2857,N_2193,N_2141);
or U2858 (N_2858,N_2175,N_2447);
nor U2859 (N_2859,N_2398,N_2053);
nand U2860 (N_2860,N_2406,N_2193);
and U2861 (N_2861,N_2231,N_2453);
or U2862 (N_2862,N_2020,N_2166);
nor U2863 (N_2863,N_2415,N_2470);
and U2864 (N_2864,N_2195,N_2468);
and U2865 (N_2865,N_2239,N_2400);
xor U2866 (N_2866,N_2370,N_2157);
and U2867 (N_2867,N_2234,N_2147);
nand U2868 (N_2868,N_2450,N_2136);
and U2869 (N_2869,N_2175,N_2072);
and U2870 (N_2870,N_2272,N_2298);
xnor U2871 (N_2871,N_2464,N_2065);
or U2872 (N_2872,N_2009,N_2494);
and U2873 (N_2873,N_2183,N_2084);
or U2874 (N_2874,N_2366,N_2235);
and U2875 (N_2875,N_2021,N_2245);
xnor U2876 (N_2876,N_2400,N_2247);
and U2877 (N_2877,N_2015,N_2365);
and U2878 (N_2878,N_2012,N_2276);
nand U2879 (N_2879,N_2493,N_2193);
nand U2880 (N_2880,N_2483,N_2028);
nand U2881 (N_2881,N_2143,N_2023);
or U2882 (N_2882,N_2347,N_2439);
or U2883 (N_2883,N_2088,N_2116);
and U2884 (N_2884,N_2232,N_2170);
or U2885 (N_2885,N_2221,N_2178);
nor U2886 (N_2886,N_2316,N_2198);
and U2887 (N_2887,N_2349,N_2330);
or U2888 (N_2888,N_2018,N_2351);
or U2889 (N_2889,N_2441,N_2121);
and U2890 (N_2890,N_2274,N_2180);
and U2891 (N_2891,N_2493,N_2244);
or U2892 (N_2892,N_2324,N_2125);
or U2893 (N_2893,N_2196,N_2012);
nor U2894 (N_2894,N_2350,N_2409);
xnor U2895 (N_2895,N_2491,N_2031);
and U2896 (N_2896,N_2081,N_2079);
xnor U2897 (N_2897,N_2372,N_2335);
xnor U2898 (N_2898,N_2348,N_2370);
and U2899 (N_2899,N_2397,N_2409);
or U2900 (N_2900,N_2264,N_2291);
xor U2901 (N_2901,N_2006,N_2084);
nor U2902 (N_2902,N_2445,N_2444);
nand U2903 (N_2903,N_2430,N_2216);
xor U2904 (N_2904,N_2392,N_2179);
and U2905 (N_2905,N_2105,N_2462);
nand U2906 (N_2906,N_2204,N_2357);
and U2907 (N_2907,N_2265,N_2438);
xnor U2908 (N_2908,N_2064,N_2172);
nor U2909 (N_2909,N_2001,N_2171);
or U2910 (N_2910,N_2437,N_2146);
xnor U2911 (N_2911,N_2101,N_2443);
and U2912 (N_2912,N_2447,N_2171);
and U2913 (N_2913,N_2407,N_2442);
xnor U2914 (N_2914,N_2048,N_2260);
and U2915 (N_2915,N_2495,N_2025);
xnor U2916 (N_2916,N_2059,N_2179);
xnor U2917 (N_2917,N_2153,N_2015);
xnor U2918 (N_2918,N_2201,N_2266);
and U2919 (N_2919,N_2271,N_2108);
and U2920 (N_2920,N_2175,N_2418);
xnor U2921 (N_2921,N_2265,N_2245);
nor U2922 (N_2922,N_2162,N_2309);
and U2923 (N_2923,N_2143,N_2388);
xor U2924 (N_2924,N_2125,N_2151);
and U2925 (N_2925,N_2105,N_2013);
xnor U2926 (N_2926,N_2290,N_2100);
nand U2927 (N_2927,N_2353,N_2246);
nor U2928 (N_2928,N_2112,N_2297);
or U2929 (N_2929,N_2135,N_2226);
or U2930 (N_2930,N_2367,N_2015);
or U2931 (N_2931,N_2293,N_2481);
xnor U2932 (N_2932,N_2099,N_2079);
and U2933 (N_2933,N_2036,N_2358);
or U2934 (N_2934,N_2476,N_2162);
or U2935 (N_2935,N_2462,N_2167);
xor U2936 (N_2936,N_2323,N_2051);
nor U2937 (N_2937,N_2251,N_2389);
or U2938 (N_2938,N_2347,N_2040);
nor U2939 (N_2939,N_2387,N_2281);
xnor U2940 (N_2940,N_2345,N_2472);
xor U2941 (N_2941,N_2126,N_2228);
nor U2942 (N_2942,N_2363,N_2191);
or U2943 (N_2943,N_2308,N_2207);
and U2944 (N_2944,N_2243,N_2149);
nand U2945 (N_2945,N_2300,N_2074);
xnor U2946 (N_2946,N_2328,N_2116);
xnor U2947 (N_2947,N_2426,N_2282);
and U2948 (N_2948,N_2448,N_2177);
nor U2949 (N_2949,N_2341,N_2039);
or U2950 (N_2950,N_2414,N_2308);
and U2951 (N_2951,N_2090,N_2251);
xnor U2952 (N_2952,N_2031,N_2154);
or U2953 (N_2953,N_2136,N_2327);
nor U2954 (N_2954,N_2172,N_2132);
xnor U2955 (N_2955,N_2090,N_2136);
and U2956 (N_2956,N_2330,N_2446);
xnor U2957 (N_2957,N_2364,N_2318);
and U2958 (N_2958,N_2296,N_2390);
and U2959 (N_2959,N_2167,N_2181);
nor U2960 (N_2960,N_2453,N_2405);
and U2961 (N_2961,N_2195,N_2210);
or U2962 (N_2962,N_2401,N_2091);
or U2963 (N_2963,N_2197,N_2377);
and U2964 (N_2964,N_2085,N_2375);
nand U2965 (N_2965,N_2460,N_2176);
nor U2966 (N_2966,N_2255,N_2456);
nor U2967 (N_2967,N_2214,N_2223);
and U2968 (N_2968,N_2069,N_2350);
nand U2969 (N_2969,N_2199,N_2043);
and U2970 (N_2970,N_2339,N_2366);
and U2971 (N_2971,N_2301,N_2137);
nand U2972 (N_2972,N_2154,N_2289);
nand U2973 (N_2973,N_2150,N_2249);
or U2974 (N_2974,N_2400,N_2223);
nor U2975 (N_2975,N_2211,N_2100);
and U2976 (N_2976,N_2460,N_2034);
nor U2977 (N_2977,N_2455,N_2345);
and U2978 (N_2978,N_2395,N_2357);
or U2979 (N_2979,N_2338,N_2283);
nor U2980 (N_2980,N_2064,N_2022);
nor U2981 (N_2981,N_2328,N_2135);
nand U2982 (N_2982,N_2217,N_2265);
or U2983 (N_2983,N_2237,N_2003);
or U2984 (N_2984,N_2014,N_2027);
nor U2985 (N_2985,N_2202,N_2409);
xor U2986 (N_2986,N_2432,N_2396);
or U2987 (N_2987,N_2274,N_2369);
or U2988 (N_2988,N_2304,N_2178);
and U2989 (N_2989,N_2024,N_2278);
xnor U2990 (N_2990,N_2417,N_2433);
xor U2991 (N_2991,N_2104,N_2116);
nor U2992 (N_2992,N_2424,N_2459);
nand U2993 (N_2993,N_2308,N_2197);
xor U2994 (N_2994,N_2427,N_2493);
nor U2995 (N_2995,N_2132,N_2338);
nand U2996 (N_2996,N_2079,N_2304);
xnor U2997 (N_2997,N_2412,N_2331);
xnor U2998 (N_2998,N_2401,N_2399);
and U2999 (N_2999,N_2111,N_2288);
and U3000 (N_3000,N_2690,N_2773);
nor U3001 (N_3001,N_2689,N_2574);
nand U3002 (N_3002,N_2568,N_2671);
nor U3003 (N_3003,N_2927,N_2984);
and U3004 (N_3004,N_2710,N_2623);
xnor U3005 (N_3005,N_2598,N_2964);
and U3006 (N_3006,N_2782,N_2603);
nand U3007 (N_3007,N_2952,N_2570);
nor U3008 (N_3008,N_2756,N_2673);
nor U3009 (N_3009,N_2787,N_2738);
and U3010 (N_3010,N_2641,N_2823);
xor U3011 (N_3011,N_2944,N_2519);
and U3012 (N_3012,N_2726,N_2959);
nor U3013 (N_3013,N_2563,N_2950);
xor U3014 (N_3014,N_2998,N_2708);
xnor U3015 (N_3015,N_2777,N_2810);
and U3016 (N_3016,N_2894,N_2834);
nor U3017 (N_3017,N_2941,N_2926);
or U3018 (N_3018,N_2914,N_2733);
nand U3019 (N_3019,N_2583,N_2801);
nand U3020 (N_3020,N_2813,N_2606);
nand U3021 (N_3021,N_2762,N_2715);
xnor U3022 (N_3022,N_2825,N_2880);
and U3023 (N_3023,N_2901,N_2837);
and U3024 (N_3024,N_2929,N_2989);
nand U3025 (N_3025,N_2879,N_2976);
nor U3026 (N_3026,N_2949,N_2957);
nand U3027 (N_3027,N_2593,N_2676);
xor U3028 (N_3028,N_2804,N_2956);
nand U3029 (N_3029,N_2860,N_2642);
and U3030 (N_3030,N_2900,N_2955);
xnor U3031 (N_3031,N_2831,N_2718);
xnor U3032 (N_3032,N_2930,N_2712);
or U3033 (N_3033,N_2585,N_2584);
xnor U3034 (N_3034,N_2724,N_2592);
xnor U3035 (N_3035,N_2795,N_2702);
nor U3036 (N_3036,N_2717,N_2664);
or U3037 (N_3037,N_2761,N_2903);
xnor U3038 (N_3038,N_2605,N_2505);
xnor U3039 (N_3039,N_2722,N_2776);
xnor U3040 (N_3040,N_2877,N_2991);
nand U3041 (N_3041,N_2672,N_2836);
or U3042 (N_3042,N_2536,N_2802);
nor U3043 (N_3043,N_2772,N_2932);
xor U3044 (N_3044,N_2809,N_2532);
and U3045 (N_3045,N_2633,N_2971);
xnor U3046 (N_3046,N_2943,N_2909);
nor U3047 (N_3047,N_2732,N_2910);
and U3048 (N_3048,N_2750,N_2892);
and U3049 (N_3049,N_2829,N_2681);
nand U3050 (N_3050,N_2812,N_2548);
xnor U3051 (N_3051,N_2752,N_2515);
or U3052 (N_3052,N_2886,N_2791);
or U3053 (N_3053,N_2827,N_2602);
xor U3054 (N_3054,N_2721,N_2890);
or U3055 (N_3055,N_2790,N_2963);
or U3056 (N_3056,N_2631,N_2587);
xnor U3057 (N_3057,N_2815,N_2865);
xor U3058 (N_3058,N_2655,N_2560);
nand U3059 (N_3059,N_2855,N_2609);
nand U3060 (N_3060,N_2685,N_2512);
nor U3061 (N_3061,N_2618,N_2857);
xnor U3062 (N_3062,N_2504,N_2833);
nor U3063 (N_3063,N_2654,N_2818);
nor U3064 (N_3064,N_2911,N_2904);
or U3065 (N_3065,N_2817,N_2597);
and U3066 (N_3066,N_2646,N_2659);
and U3067 (N_3067,N_2805,N_2582);
or U3068 (N_3068,N_2967,N_2948);
and U3069 (N_3069,N_2680,N_2988);
nor U3070 (N_3070,N_2507,N_2799);
and U3071 (N_3071,N_2786,N_2546);
nand U3072 (N_3072,N_2566,N_2628);
nand U3073 (N_3073,N_2595,N_2912);
nor U3074 (N_3074,N_2636,N_2995);
nand U3075 (N_3075,N_2679,N_2906);
or U3076 (N_3076,N_2540,N_2580);
or U3077 (N_3077,N_2530,N_2632);
and U3078 (N_3078,N_2573,N_2543);
xnor U3079 (N_3079,N_2788,N_2538);
and U3080 (N_3080,N_2711,N_2768);
nor U3081 (N_3081,N_2533,N_2703);
nor U3082 (N_3082,N_2862,N_2660);
and U3083 (N_3083,N_2645,N_2819);
nand U3084 (N_3084,N_2841,N_2688);
nand U3085 (N_3085,N_2997,N_2821);
and U3086 (N_3086,N_2590,N_2526);
and U3087 (N_3087,N_2694,N_2897);
nor U3088 (N_3088,N_2621,N_2691);
and U3089 (N_3089,N_2695,N_2946);
nor U3090 (N_3090,N_2518,N_2888);
nor U3091 (N_3091,N_2947,N_2514);
and U3092 (N_3092,N_2578,N_2665);
nor U3093 (N_3093,N_2881,N_2769);
nor U3094 (N_3094,N_2767,N_2760);
xor U3095 (N_3095,N_2610,N_2852);
nor U3096 (N_3096,N_2820,N_2668);
xor U3097 (N_3097,N_2736,N_2936);
or U3098 (N_3098,N_2958,N_2806);
xor U3099 (N_3099,N_2999,N_2960);
nand U3100 (N_3100,N_2569,N_2713);
nand U3101 (N_3101,N_2962,N_2951);
nand U3102 (N_3102,N_2741,N_2678);
xnor U3103 (N_3103,N_2975,N_2896);
or U3104 (N_3104,N_2934,N_2524);
or U3105 (N_3105,N_2567,N_2861);
and U3106 (N_3106,N_2725,N_2581);
or U3107 (N_3107,N_2545,N_2705);
and U3108 (N_3108,N_2516,N_2699);
nor U3109 (N_3109,N_2816,N_2794);
nor U3110 (N_3110,N_2649,N_2882);
or U3111 (N_3111,N_2796,N_2916);
xnor U3112 (N_3112,N_2728,N_2692);
nand U3113 (N_3113,N_2535,N_2828);
xor U3114 (N_3114,N_2883,N_2617);
xnor U3115 (N_3115,N_2990,N_2969);
nand U3116 (N_3116,N_2755,N_2503);
or U3117 (N_3117,N_2928,N_2608);
xnor U3118 (N_3118,N_2634,N_2792);
nand U3119 (N_3119,N_2982,N_2864);
nor U3120 (N_3120,N_2847,N_2553);
nor U3121 (N_3121,N_2870,N_2814);
and U3122 (N_3122,N_2779,N_2965);
and U3123 (N_3123,N_2520,N_2658);
and U3124 (N_3124,N_2968,N_2662);
nor U3125 (N_3125,N_2576,N_2745);
and U3126 (N_3126,N_2562,N_2783);
and U3127 (N_3127,N_2720,N_2933);
or U3128 (N_3128,N_2522,N_2550);
and U3129 (N_3129,N_2838,N_2994);
nor U3130 (N_3130,N_2647,N_2832);
nor U3131 (N_3131,N_2700,N_2523);
xnor U3132 (N_3132,N_2798,N_2940);
or U3133 (N_3133,N_2789,N_2556);
nand U3134 (N_3134,N_2586,N_2552);
or U3135 (N_3135,N_2751,N_2757);
nor U3136 (N_3136,N_2716,N_2867);
or U3137 (N_3137,N_2970,N_2657);
and U3138 (N_3138,N_2542,N_2629);
or U3139 (N_3139,N_2719,N_2701);
xnor U3140 (N_3140,N_2675,N_2992);
nor U3141 (N_3141,N_2978,N_2601);
nor U3142 (N_3142,N_2771,N_2873);
nor U3143 (N_3143,N_2682,N_2754);
or U3144 (N_3144,N_2697,N_2874);
xnor U3145 (N_3145,N_2869,N_2511);
and U3146 (N_3146,N_2571,N_2899);
and U3147 (N_3147,N_2843,N_2961);
nor U3148 (N_3148,N_2666,N_2648);
xor U3149 (N_3149,N_2558,N_2765);
nand U3150 (N_3150,N_2698,N_2669);
nand U3151 (N_3151,N_2902,N_2509);
and U3152 (N_3152,N_2803,N_2594);
nand U3153 (N_3153,N_2945,N_2845);
and U3154 (N_3154,N_2935,N_2624);
and U3155 (N_3155,N_2797,N_2872);
nand U3156 (N_3156,N_2687,N_2577);
or U3157 (N_3157,N_2954,N_2709);
or U3158 (N_3158,N_2541,N_2876);
and U3159 (N_3159,N_2537,N_2600);
xnor U3160 (N_3160,N_2763,N_2746);
nand U3161 (N_3161,N_2527,N_2931);
and U3162 (N_3162,N_2604,N_2878);
and U3163 (N_3163,N_2979,N_2980);
or U3164 (N_3164,N_2729,N_2579);
nand U3165 (N_3165,N_2588,N_2707);
and U3166 (N_3166,N_2517,N_2620);
or U3167 (N_3167,N_2640,N_2793);
nor U3168 (N_3168,N_2921,N_2759);
and U3169 (N_3169,N_2501,N_2974);
or U3170 (N_3170,N_2907,N_2614);
xnor U3171 (N_3171,N_2644,N_2919);
nand U3172 (N_3172,N_2983,N_2652);
nand U3173 (N_3173,N_2774,N_2764);
nand U3174 (N_3174,N_2704,N_2714);
nand U3175 (N_3175,N_2866,N_2639);
nand U3176 (N_3176,N_2730,N_2848);
and U3177 (N_3177,N_2513,N_2723);
and U3178 (N_3178,N_2748,N_2753);
or U3179 (N_3179,N_2740,N_2942);
nor U3180 (N_3180,N_2842,N_2565);
and U3181 (N_3181,N_2973,N_2737);
nand U3182 (N_3182,N_2993,N_2693);
nor U3183 (N_3183,N_2734,N_2706);
nand U3184 (N_3184,N_2742,N_2875);
xnor U3185 (N_3185,N_2844,N_2987);
or U3186 (N_3186,N_2808,N_2525);
xnor U3187 (N_3187,N_2846,N_2922);
or U3188 (N_3188,N_2555,N_2784);
xor U3189 (N_3189,N_2887,N_2822);
or U3190 (N_3190,N_2500,N_2656);
nor U3191 (N_3191,N_2913,N_2529);
nand U3192 (N_3192,N_2607,N_2727);
or U3193 (N_3193,N_2549,N_2811);
nor U3194 (N_3194,N_2667,N_2780);
nand U3195 (N_3195,N_2891,N_2544);
nor U3196 (N_3196,N_2884,N_2651);
or U3197 (N_3197,N_2637,N_2575);
or U3198 (N_3198,N_2981,N_2770);
nand U3199 (N_3199,N_2835,N_2670);
nand U3200 (N_3200,N_2561,N_2889);
nand U3201 (N_3201,N_2938,N_2589);
and U3202 (N_3202,N_2674,N_2826);
xor U3203 (N_3203,N_2622,N_2635);
xnor U3204 (N_3204,N_2638,N_2653);
nand U3205 (N_3205,N_2923,N_2508);
xor U3206 (N_3206,N_2559,N_2905);
xor U3207 (N_3207,N_2807,N_2615);
or U3208 (N_3208,N_2613,N_2591);
or U3209 (N_3209,N_2612,N_2996);
nand U3210 (N_3210,N_2619,N_2856);
and U3211 (N_3211,N_2893,N_2868);
nand U3212 (N_3212,N_2985,N_2557);
and U3213 (N_3213,N_2766,N_2986);
or U3214 (N_3214,N_2800,N_2839);
xnor U3215 (N_3215,N_2551,N_2564);
or U3216 (N_3216,N_2684,N_2966);
nand U3217 (N_3217,N_2677,N_2972);
and U3218 (N_3218,N_2851,N_2824);
nand U3219 (N_3219,N_2686,N_2917);
nand U3220 (N_3220,N_2572,N_2626);
or U3221 (N_3221,N_2506,N_2915);
xnor U3222 (N_3222,N_2663,N_2858);
or U3223 (N_3223,N_2918,N_2683);
or U3224 (N_3224,N_2937,N_2611);
and U3225 (N_3225,N_2739,N_2830);
xor U3226 (N_3226,N_2849,N_2925);
xnor U3227 (N_3227,N_2840,N_2850);
xnor U3228 (N_3228,N_2539,N_2781);
nor U3229 (N_3229,N_2977,N_2953);
nand U3230 (N_3230,N_2920,N_2853);
and U3231 (N_3231,N_2625,N_2885);
nor U3232 (N_3232,N_2528,N_2531);
nor U3233 (N_3233,N_2547,N_2554);
nor U3234 (N_3234,N_2735,N_2924);
nor U3235 (N_3235,N_2627,N_2758);
and U3236 (N_3236,N_2502,N_2599);
and U3237 (N_3237,N_2859,N_2630);
xnor U3238 (N_3238,N_2785,N_2871);
or U3239 (N_3239,N_2616,N_2596);
xnor U3240 (N_3240,N_2898,N_2747);
nor U3241 (N_3241,N_2731,N_2510);
nand U3242 (N_3242,N_2863,N_2521);
or U3243 (N_3243,N_2775,N_2749);
and U3244 (N_3244,N_2778,N_2854);
nand U3245 (N_3245,N_2661,N_2908);
and U3246 (N_3246,N_2743,N_2650);
nand U3247 (N_3247,N_2643,N_2895);
or U3248 (N_3248,N_2744,N_2534);
xor U3249 (N_3249,N_2696,N_2939);
or U3250 (N_3250,N_2822,N_2863);
nor U3251 (N_3251,N_2910,N_2817);
nand U3252 (N_3252,N_2593,N_2673);
nor U3253 (N_3253,N_2509,N_2707);
or U3254 (N_3254,N_2619,N_2511);
xnor U3255 (N_3255,N_2969,N_2535);
xor U3256 (N_3256,N_2773,N_2978);
xnor U3257 (N_3257,N_2845,N_2860);
nor U3258 (N_3258,N_2570,N_2945);
xnor U3259 (N_3259,N_2874,N_2623);
nor U3260 (N_3260,N_2655,N_2969);
and U3261 (N_3261,N_2774,N_2645);
xor U3262 (N_3262,N_2912,N_2529);
nand U3263 (N_3263,N_2586,N_2943);
or U3264 (N_3264,N_2536,N_2735);
and U3265 (N_3265,N_2911,N_2666);
xor U3266 (N_3266,N_2889,N_2510);
nand U3267 (N_3267,N_2955,N_2929);
or U3268 (N_3268,N_2838,N_2921);
nor U3269 (N_3269,N_2511,N_2951);
and U3270 (N_3270,N_2622,N_2689);
nand U3271 (N_3271,N_2909,N_2716);
or U3272 (N_3272,N_2833,N_2806);
and U3273 (N_3273,N_2665,N_2978);
or U3274 (N_3274,N_2693,N_2513);
or U3275 (N_3275,N_2723,N_2881);
nand U3276 (N_3276,N_2513,N_2822);
and U3277 (N_3277,N_2891,N_2600);
or U3278 (N_3278,N_2878,N_2997);
or U3279 (N_3279,N_2589,N_2756);
nand U3280 (N_3280,N_2668,N_2675);
or U3281 (N_3281,N_2578,N_2639);
or U3282 (N_3282,N_2945,N_2980);
and U3283 (N_3283,N_2972,N_2794);
or U3284 (N_3284,N_2764,N_2528);
xor U3285 (N_3285,N_2679,N_2846);
nor U3286 (N_3286,N_2646,N_2892);
nor U3287 (N_3287,N_2747,N_2675);
nand U3288 (N_3288,N_2734,N_2695);
nand U3289 (N_3289,N_2570,N_2887);
xor U3290 (N_3290,N_2898,N_2850);
and U3291 (N_3291,N_2746,N_2743);
and U3292 (N_3292,N_2912,N_2778);
xnor U3293 (N_3293,N_2898,N_2698);
xnor U3294 (N_3294,N_2514,N_2663);
and U3295 (N_3295,N_2918,N_2759);
or U3296 (N_3296,N_2994,N_2956);
or U3297 (N_3297,N_2714,N_2781);
and U3298 (N_3298,N_2698,N_2768);
xor U3299 (N_3299,N_2768,N_2521);
xnor U3300 (N_3300,N_2544,N_2670);
nand U3301 (N_3301,N_2788,N_2934);
and U3302 (N_3302,N_2941,N_2546);
xor U3303 (N_3303,N_2619,N_2707);
or U3304 (N_3304,N_2784,N_2683);
nand U3305 (N_3305,N_2602,N_2959);
and U3306 (N_3306,N_2862,N_2605);
xnor U3307 (N_3307,N_2961,N_2816);
and U3308 (N_3308,N_2860,N_2689);
xor U3309 (N_3309,N_2714,N_2640);
nand U3310 (N_3310,N_2936,N_2523);
or U3311 (N_3311,N_2604,N_2680);
and U3312 (N_3312,N_2850,N_2799);
nor U3313 (N_3313,N_2873,N_2970);
and U3314 (N_3314,N_2803,N_2685);
or U3315 (N_3315,N_2996,N_2784);
or U3316 (N_3316,N_2663,N_2712);
nor U3317 (N_3317,N_2996,N_2888);
nand U3318 (N_3318,N_2516,N_2834);
and U3319 (N_3319,N_2947,N_2507);
nand U3320 (N_3320,N_2922,N_2840);
nor U3321 (N_3321,N_2691,N_2869);
nor U3322 (N_3322,N_2525,N_2694);
or U3323 (N_3323,N_2532,N_2852);
and U3324 (N_3324,N_2616,N_2790);
or U3325 (N_3325,N_2953,N_2786);
and U3326 (N_3326,N_2746,N_2616);
xor U3327 (N_3327,N_2926,N_2697);
nand U3328 (N_3328,N_2552,N_2951);
and U3329 (N_3329,N_2879,N_2809);
nor U3330 (N_3330,N_2775,N_2502);
nand U3331 (N_3331,N_2929,N_2848);
and U3332 (N_3332,N_2922,N_2828);
nand U3333 (N_3333,N_2791,N_2754);
xnor U3334 (N_3334,N_2843,N_2737);
or U3335 (N_3335,N_2516,N_2673);
xnor U3336 (N_3336,N_2942,N_2630);
nand U3337 (N_3337,N_2505,N_2920);
nand U3338 (N_3338,N_2589,N_2621);
nand U3339 (N_3339,N_2828,N_2872);
and U3340 (N_3340,N_2925,N_2801);
nand U3341 (N_3341,N_2521,N_2744);
and U3342 (N_3342,N_2920,N_2870);
or U3343 (N_3343,N_2533,N_2845);
or U3344 (N_3344,N_2641,N_2817);
and U3345 (N_3345,N_2889,N_2973);
nor U3346 (N_3346,N_2567,N_2749);
or U3347 (N_3347,N_2647,N_2689);
and U3348 (N_3348,N_2750,N_2855);
xor U3349 (N_3349,N_2944,N_2679);
nor U3350 (N_3350,N_2584,N_2928);
and U3351 (N_3351,N_2701,N_2557);
and U3352 (N_3352,N_2705,N_2556);
nand U3353 (N_3353,N_2870,N_2567);
or U3354 (N_3354,N_2865,N_2810);
nand U3355 (N_3355,N_2924,N_2645);
nand U3356 (N_3356,N_2714,N_2756);
nand U3357 (N_3357,N_2729,N_2866);
nand U3358 (N_3358,N_2556,N_2963);
nand U3359 (N_3359,N_2602,N_2985);
or U3360 (N_3360,N_2586,N_2874);
nand U3361 (N_3361,N_2936,N_2876);
xnor U3362 (N_3362,N_2717,N_2976);
xnor U3363 (N_3363,N_2628,N_2658);
nand U3364 (N_3364,N_2773,N_2925);
nand U3365 (N_3365,N_2847,N_2953);
nand U3366 (N_3366,N_2907,N_2842);
and U3367 (N_3367,N_2695,N_2983);
nand U3368 (N_3368,N_2917,N_2840);
and U3369 (N_3369,N_2764,N_2890);
and U3370 (N_3370,N_2604,N_2686);
nand U3371 (N_3371,N_2557,N_2586);
xor U3372 (N_3372,N_2772,N_2787);
nor U3373 (N_3373,N_2986,N_2814);
xnor U3374 (N_3374,N_2896,N_2889);
and U3375 (N_3375,N_2828,N_2974);
nor U3376 (N_3376,N_2538,N_2656);
nor U3377 (N_3377,N_2766,N_2590);
nor U3378 (N_3378,N_2649,N_2656);
xor U3379 (N_3379,N_2951,N_2975);
xnor U3380 (N_3380,N_2942,N_2732);
xnor U3381 (N_3381,N_2798,N_2890);
nor U3382 (N_3382,N_2832,N_2516);
xor U3383 (N_3383,N_2634,N_2501);
xor U3384 (N_3384,N_2829,N_2825);
xnor U3385 (N_3385,N_2903,N_2544);
and U3386 (N_3386,N_2878,N_2522);
nand U3387 (N_3387,N_2894,N_2560);
or U3388 (N_3388,N_2924,N_2975);
nand U3389 (N_3389,N_2577,N_2633);
nand U3390 (N_3390,N_2730,N_2761);
and U3391 (N_3391,N_2655,N_2842);
nor U3392 (N_3392,N_2708,N_2767);
and U3393 (N_3393,N_2536,N_2511);
nor U3394 (N_3394,N_2756,N_2659);
and U3395 (N_3395,N_2923,N_2728);
nand U3396 (N_3396,N_2581,N_2628);
xnor U3397 (N_3397,N_2875,N_2815);
or U3398 (N_3398,N_2798,N_2978);
or U3399 (N_3399,N_2662,N_2818);
or U3400 (N_3400,N_2832,N_2730);
and U3401 (N_3401,N_2928,N_2665);
or U3402 (N_3402,N_2636,N_2800);
nand U3403 (N_3403,N_2745,N_2947);
and U3404 (N_3404,N_2832,N_2629);
and U3405 (N_3405,N_2936,N_2555);
xnor U3406 (N_3406,N_2988,N_2947);
nand U3407 (N_3407,N_2874,N_2951);
nand U3408 (N_3408,N_2773,N_2797);
nor U3409 (N_3409,N_2714,N_2514);
nor U3410 (N_3410,N_2776,N_2646);
and U3411 (N_3411,N_2596,N_2847);
xnor U3412 (N_3412,N_2884,N_2788);
and U3413 (N_3413,N_2840,N_2504);
nor U3414 (N_3414,N_2503,N_2887);
and U3415 (N_3415,N_2597,N_2526);
and U3416 (N_3416,N_2609,N_2925);
nand U3417 (N_3417,N_2789,N_2855);
and U3418 (N_3418,N_2706,N_2532);
nor U3419 (N_3419,N_2840,N_2905);
or U3420 (N_3420,N_2597,N_2722);
or U3421 (N_3421,N_2527,N_2537);
xor U3422 (N_3422,N_2711,N_2906);
xnor U3423 (N_3423,N_2732,N_2670);
xor U3424 (N_3424,N_2573,N_2700);
xnor U3425 (N_3425,N_2759,N_2707);
or U3426 (N_3426,N_2658,N_2653);
xor U3427 (N_3427,N_2685,N_2895);
and U3428 (N_3428,N_2589,N_2960);
nor U3429 (N_3429,N_2593,N_2963);
nand U3430 (N_3430,N_2974,N_2977);
nor U3431 (N_3431,N_2809,N_2756);
xnor U3432 (N_3432,N_2959,N_2572);
or U3433 (N_3433,N_2916,N_2638);
xnor U3434 (N_3434,N_2622,N_2973);
nand U3435 (N_3435,N_2730,N_2768);
or U3436 (N_3436,N_2856,N_2964);
or U3437 (N_3437,N_2824,N_2627);
nor U3438 (N_3438,N_2715,N_2592);
nor U3439 (N_3439,N_2533,N_2663);
and U3440 (N_3440,N_2581,N_2847);
xor U3441 (N_3441,N_2712,N_2688);
and U3442 (N_3442,N_2750,N_2547);
or U3443 (N_3443,N_2712,N_2693);
xnor U3444 (N_3444,N_2508,N_2827);
xor U3445 (N_3445,N_2947,N_2815);
nand U3446 (N_3446,N_2868,N_2660);
nor U3447 (N_3447,N_2958,N_2611);
nor U3448 (N_3448,N_2510,N_2723);
and U3449 (N_3449,N_2535,N_2966);
and U3450 (N_3450,N_2845,N_2928);
nand U3451 (N_3451,N_2817,N_2806);
and U3452 (N_3452,N_2510,N_2853);
nor U3453 (N_3453,N_2948,N_2956);
nand U3454 (N_3454,N_2974,N_2522);
and U3455 (N_3455,N_2525,N_2636);
nand U3456 (N_3456,N_2694,N_2839);
nand U3457 (N_3457,N_2928,N_2620);
and U3458 (N_3458,N_2992,N_2821);
nor U3459 (N_3459,N_2884,N_2905);
or U3460 (N_3460,N_2501,N_2554);
xor U3461 (N_3461,N_2950,N_2590);
xnor U3462 (N_3462,N_2984,N_2570);
xor U3463 (N_3463,N_2882,N_2987);
nand U3464 (N_3464,N_2943,N_2963);
and U3465 (N_3465,N_2542,N_2688);
nand U3466 (N_3466,N_2588,N_2582);
xnor U3467 (N_3467,N_2582,N_2553);
nor U3468 (N_3468,N_2708,N_2710);
xnor U3469 (N_3469,N_2618,N_2655);
xnor U3470 (N_3470,N_2688,N_2583);
xor U3471 (N_3471,N_2716,N_2814);
or U3472 (N_3472,N_2620,N_2906);
xor U3473 (N_3473,N_2889,N_2947);
and U3474 (N_3474,N_2949,N_2549);
xnor U3475 (N_3475,N_2588,N_2899);
xnor U3476 (N_3476,N_2646,N_2541);
and U3477 (N_3477,N_2682,N_2983);
and U3478 (N_3478,N_2850,N_2876);
nor U3479 (N_3479,N_2793,N_2897);
nor U3480 (N_3480,N_2514,N_2742);
or U3481 (N_3481,N_2598,N_2660);
nor U3482 (N_3482,N_2821,N_2880);
or U3483 (N_3483,N_2936,N_2687);
and U3484 (N_3484,N_2753,N_2603);
and U3485 (N_3485,N_2805,N_2649);
nor U3486 (N_3486,N_2694,N_2702);
xor U3487 (N_3487,N_2609,N_2705);
and U3488 (N_3488,N_2996,N_2866);
or U3489 (N_3489,N_2793,N_2951);
or U3490 (N_3490,N_2696,N_2631);
xor U3491 (N_3491,N_2675,N_2726);
nand U3492 (N_3492,N_2903,N_2567);
or U3493 (N_3493,N_2783,N_2655);
nand U3494 (N_3494,N_2540,N_2599);
or U3495 (N_3495,N_2545,N_2808);
and U3496 (N_3496,N_2821,N_2709);
and U3497 (N_3497,N_2882,N_2635);
and U3498 (N_3498,N_2933,N_2936);
or U3499 (N_3499,N_2569,N_2704);
nand U3500 (N_3500,N_3404,N_3287);
or U3501 (N_3501,N_3321,N_3037);
xor U3502 (N_3502,N_3405,N_3061);
xor U3503 (N_3503,N_3439,N_3424);
xnor U3504 (N_3504,N_3317,N_3293);
nand U3505 (N_3505,N_3310,N_3279);
xnor U3506 (N_3506,N_3013,N_3094);
nand U3507 (N_3507,N_3022,N_3258);
nand U3508 (N_3508,N_3306,N_3096);
or U3509 (N_3509,N_3472,N_3052);
or U3510 (N_3510,N_3435,N_3031);
or U3511 (N_3511,N_3165,N_3337);
and U3512 (N_3512,N_3179,N_3469);
nor U3513 (N_3513,N_3305,N_3417);
xnor U3514 (N_3514,N_3073,N_3265);
and U3515 (N_3515,N_3480,N_3408);
xnor U3516 (N_3516,N_3401,N_3465);
nor U3517 (N_3517,N_3498,N_3205);
nor U3518 (N_3518,N_3152,N_3479);
nor U3519 (N_3519,N_3230,N_3309);
nand U3520 (N_3520,N_3490,N_3241);
and U3521 (N_3521,N_3026,N_3098);
nand U3522 (N_3522,N_3276,N_3338);
nand U3523 (N_3523,N_3225,N_3206);
nor U3524 (N_3524,N_3430,N_3399);
and U3525 (N_3525,N_3252,N_3455);
xor U3526 (N_3526,N_3215,N_3382);
nor U3527 (N_3527,N_3254,N_3261);
nand U3528 (N_3528,N_3489,N_3175);
nor U3529 (N_3529,N_3053,N_3275);
or U3530 (N_3530,N_3238,N_3048);
xor U3531 (N_3531,N_3441,N_3343);
and U3532 (N_3532,N_3250,N_3297);
and U3533 (N_3533,N_3388,N_3109);
or U3534 (N_3534,N_3466,N_3140);
xor U3535 (N_3535,N_3333,N_3202);
nor U3536 (N_3536,N_3295,N_3302);
nand U3537 (N_3537,N_3386,N_3434);
and U3538 (N_3538,N_3330,N_3186);
nor U3539 (N_3539,N_3045,N_3097);
xor U3540 (N_3540,N_3419,N_3080);
or U3541 (N_3541,N_3390,N_3263);
xnor U3542 (N_3542,N_3444,N_3284);
and U3543 (N_3543,N_3016,N_3128);
xor U3544 (N_3544,N_3020,N_3021);
xnor U3545 (N_3545,N_3339,N_3229);
xor U3546 (N_3546,N_3418,N_3462);
xnor U3547 (N_3547,N_3281,N_3204);
nand U3548 (N_3548,N_3410,N_3454);
xnor U3549 (N_3549,N_3447,N_3428);
xnor U3550 (N_3550,N_3023,N_3234);
and U3551 (N_3551,N_3448,N_3149);
or U3552 (N_3552,N_3180,N_3067);
nand U3553 (N_3553,N_3323,N_3352);
or U3554 (N_3554,N_3446,N_3232);
xor U3555 (N_3555,N_3055,N_3381);
nor U3556 (N_3556,N_3092,N_3062);
nor U3557 (N_3557,N_3001,N_3118);
and U3558 (N_3558,N_3124,N_3197);
nand U3559 (N_3559,N_3355,N_3396);
nand U3560 (N_3560,N_3299,N_3398);
or U3561 (N_3561,N_3086,N_3375);
or U3562 (N_3562,N_3103,N_3363);
xor U3563 (N_3563,N_3283,N_3129);
nor U3564 (N_3564,N_3369,N_3093);
and U3565 (N_3565,N_3360,N_3262);
xor U3566 (N_3566,N_3237,N_3416);
and U3567 (N_3567,N_3458,N_3029);
nand U3568 (N_3568,N_3332,N_3312);
nand U3569 (N_3569,N_3028,N_3070);
xor U3570 (N_3570,N_3464,N_3395);
or U3571 (N_3571,N_3366,N_3420);
nand U3572 (N_3572,N_3264,N_3210);
nor U3573 (N_3573,N_3119,N_3136);
or U3574 (N_3574,N_3426,N_3325);
and U3575 (N_3575,N_3496,N_3292);
nor U3576 (N_3576,N_3101,N_3046);
nor U3577 (N_3577,N_3174,N_3161);
nand U3578 (N_3578,N_3437,N_3207);
xnor U3579 (N_3579,N_3088,N_3245);
xor U3580 (N_3580,N_3056,N_3269);
xor U3581 (N_3581,N_3125,N_3078);
and U3582 (N_3582,N_3414,N_3361);
xor U3583 (N_3583,N_3342,N_3195);
nor U3584 (N_3584,N_3365,N_3138);
nand U3585 (N_3585,N_3126,N_3249);
xnor U3586 (N_3586,N_3148,N_3137);
nand U3587 (N_3587,N_3108,N_3139);
or U3588 (N_3588,N_3383,N_3286);
xnor U3589 (N_3589,N_3300,N_3164);
nand U3590 (N_3590,N_3378,N_3329);
or U3591 (N_3591,N_3142,N_3107);
and U3592 (N_3592,N_3289,N_3389);
nor U3593 (N_3593,N_3181,N_3331);
nor U3594 (N_3594,N_3074,N_3173);
xnor U3595 (N_3595,N_3423,N_3167);
xor U3596 (N_3596,N_3168,N_3120);
nand U3597 (N_3597,N_3006,N_3208);
xnor U3598 (N_3598,N_3453,N_3268);
nand U3599 (N_3599,N_3411,N_3193);
nor U3600 (N_3600,N_3248,N_3456);
nor U3601 (N_3601,N_3433,N_3451);
nor U3602 (N_3602,N_3224,N_3171);
nor U3603 (N_3603,N_3066,N_3012);
nand U3604 (N_3604,N_3047,N_3150);
or U3605 (N_3605,N_3247,N_3327);
nor U3606 (N_3606,N_3182,N_3384);
nand U3607 (N_3607,N_3198,N_3117);
xor U3608 (N_3608,N_3328,N_3387);
xnor U3609 (N_3609,N_3253,N_3304);
and U3610 (N_3610,N_3183,N_3421);
xnor U3611 (N_3611,N_3482,N_3019);
nor U3612 (N_3612,N_3461,N_3445);
or U3613 (N_3613,N_3320,N_3166);
and U3614 (N_3614,N_3176,N_3135);
nor U3615 (N_3615,N_3222,N_3002);
and U3616 (N_3616,N_3372,N_3064);
xor U3617 (N_3617,N_3223,N_3110);
nand U3618 (N_3618,N_3014,N_3259);
and U3619 (N_3619,N_3051,N_3474);
or U3620 (N_3620,N_3005,N_3218);
xor U3621 (N_3621,N_3009,N_3228);
nand U3622 (N_3622,N_3425,N_3475);
and U3623 (N_3623,N_3121,N_3442);
or U3624 (N_3624,N_3484,N_3082);
xnor U3625 (N_3625,N_3463,N_3000);
nand U3626 (N_3626,N_3111,N_3069);
nand U3627 (N_3627,N_3298,N_3102);
nor U3628 (N_3628,N_3402,N_3314);
or U3629 (N_3629,N_3038,N_3294);
or U3630 (N_3630,N_3359,N_3227);
or U3631 (N_3631,N_3169,N_3160);
xnor U3632 (N_3632,N_3374,N_3406);
xnor U3633 (N_3633,N_3468,N_3364);
nand U3634 (N_3634,N_3192,N_3316);
xor U3635 (N_3635,N_3219,N_3071);
xnor U3636 (N_3636,N_3041,N_3345);
or U3637 (N_3637,N_3178,N_3170);
nor U3638 (N_3638,N_3353,N_3007);
or U3639 (N_3639,N_3471,N_3003);
nand U3640 (N_3640,N_3290,N_3172);
and U3641 (N_3641,N_3100,N_3141);
xor U3642 (N_3642,N_3032,N_3033);
nor U3643 (N_3643,N_3089,N_3270);
nand U3644 (N_3644,N_3058,N_3087);
nor U3645 (N_3645,N_3004,N_3060);
nand U3646 (N_3646,N_3081,N_3079);
nor U3647 (N_3647,N_3274,N_3499);
xor U3648 (N_3648,N_3334,N_3194);
and U3649 (N_3649,N_3385,N_3185);
or U3650 (N_3650,N_3256,N_3188);
xor U3651 (N_3651,N_3449,N_3257);
xor U3652 (N_3652,N_3477,N_3481);
xor U3653 (N_3653,N_3341,N_3362);
nand U3654 (N_3654,N_3367,N_3350);
nor U3655 (N_3655,N_3349,N_3260);
and U3656 (N_3656,N_3478,N_3091);
xor U3657 (N_3657,N_3162,N_3266);
and U3658 (N_3658,N_3151,N_3476);
nor U3659 (N_3659,N_3049,N_3340);
xnor U3660 (N_3660,N_3123,N_3470);
and U3661 (N_3661,N_3054,N_3407);
and U3662 (N_3662,N_3273,N_3042);
and U3663 (N_3663,N_3243,N_3035);
or U3664 (N_3664,N_3459,N_3090);
nor U3665 (N_3665,N_3377,N_3409);
nand U3666 (N_3666,N_3158,N_3467);
xnor U3667 (N_3667,N_3072,N_3116);
xor U3668 (N_3668,N_3301,N_3282);
and U3669 (N_3669,N_3065,N_3485);
xor U3670 (N_3670,N_3356,N_3285);
and U3671 (N_3671,N_3212,N_3131);
nor U3672 (N_3672,N_3491,N_3348);
xnor U3673 (N_3673,N_3422,N_3379);
nand U3674 (N_3674,N_3015,N_3075);
and U3675 (N_3675,N_3104,N_3400);
nand U3676 (N_3676,N_3190,N_3068);
or U3677 (N_3677,N_3017,N_3039);
or U3678 (N_3678,N_3153,N_3085);
and U3679 (N_3679,N_3412,N_3358);
or U3680 (N_3680,N_3246,N_3144);
or U3681 (N_3681,N_3099,N_3267);
nor U3682 (N_3682,N_3373,N_3115);
nand U3683 (N_3683,N_3209,N_3440);
and U3684 (N_3684,N_3050,N_3191);
xor U3685 (N_3685,N_3313,N_3059);
and U3686 (N_3686,N_3127,N_3211);
xnor U3687 (N_3687,N_3213,N_3403);
nor U3688 (N_3688,N_3226,N_3011);
xnor U3689 (N_3689,N_3235,N_3319);
nor U3690 (N_3690,N_3380,N_3030);
and U3691 (N_3691,N_3322,N_3106);
nor U3692 (N_3692,N_3105,N_3145);
nor U3693 (N_3693,N_3271,N_3495);
and U3694 (N_3694,N_3397,N_3436);
nor U3695 (N_3695,N_3196,N_3077);
nand U3696 (N_3696,N_3163,N_3351);
and U3697 (N_3697,N_3457,N_3443);
nand U3698 (N_3698,N_3326,N_3429);
or U3699 (N_3699,N_3307,N_3024);
or U3700 (N_3700,N_3233,N_3156);
and U3701 (N_3701,N_3244,N_3239);
and U3702 (N_3702,N_3147,N_3483);
and U3703 (N_3703,N_3114,N_3392);
nor U3704 (N_3704,N_3280,N_3057);
nand U3705 (N_3705,N_3157,N_3272);
nand U3706 (N_3706,N_3251,N_3113);
nand U3707 (N_3707,N_3393,N_3354);
and U3708 (N_3708,N_3084,N_3189);
or U3709 (N_3709,N_3036,N_3217);
xnor U3710 (N_3710,N_3154,N_3347);
and U3711 (N_3711,N_3199,N_3460);
and U3712 (N_3712,N_3200,N_3308);
and U3713 (N_3713,N_3303,N_3155);
nand U3714 (N_3714,N_3291,N_3255);
nor U3715 (N_3715,N_3083,N_3143);
nand U3716 (N_3716,N_3277,N_3452);
xnor U3717 (N_3717,N_3018,N_3368);
nand U3718 (N_3718,N_3335,N_3438);
xor U3719 (N_3719,N_3376,N_3315);
and U3720 (N_3720,N_3432,N_3415);
or U3721 (N_3721,N_3493,N_3242);
nor U3722 (N_3722,N_3450,N_3159);
nand U3723 (N_3723,N_3371,N_3214);
xor U3724 (N_3724,N_3220,N_3132);
xor U3725 (N_3725,N_3203,N_3043);
nor U3726 (N_3726,N_3044,N_3201);
nor U3727 (N_3727,N_3177,N_3431);
xnor U3728 (N_3728,N_3278,N_3008);
and U3729 (N_3729,N_3010,N_3318);
nor U3730 (N_3730,N_3497,N_3311);
nand U3731 (N_3731,N_3288,N_3240);
and U3732 (N_3732,N_3346,N_3324);
nand U3733 (N_3733,N_3063,N_3025);
or U3734 (N_3734,N_3357,N_3095);
or U3735 (N_3735,N_3027,N_3187);
or U3736 (N_3736,N_3122,N_3487);
nor U3737 (N_3737,N_3112,N_3336);
nor U3738 (N_3738,N_3216,N_3486);
xor U3739 (N_3739,N_3492,N_3130);
nand U3740 (N_3740,N_3040,N_3231);
and U3741 (N_3741,N_3391,N_3370);
and U3742 (N_3742,N_3394,N_3134);
xnor U3743 (N_3743,N_3221,N_3184);
and U3744 (N_3744,N_3427,N_3146);
and U3745 (N_3745,N_3076,N_3236);
xor U3746 (N_3746,N_3488,N_3494);
xnor U3747 (N_3747,N_3133,N_3413);
nor U3748 (N_3748,N_3034,N_3344);
or U3749 (N_3749,N_3473,N_3296);
xnor U3750 (N_3750,N_3077,N_3472);
or U3751 (N_3751,N_3349,N_3224);
nor U3752 (N_3752,N_3092,N_3486);
and U3753 (N_3753,N_3278,N_3137);
nor U3754 (N_3754,N_3410,N_3014);
nor U3755 (N_3755,N_3491,N_3377);
or U3756 (N_3756,N_3258,N_3041);
nand U3757 (N_3757,N_3077,N_3262);
nor U3758 (N_3758,N_3450,N_3249);
xnor U3759 (N_3759,N_3157,N_3232);
xnor U3760 (N_3760,N_3216,N_3367);
or U3761 (N_3761,N_3024,N_3245);
xnor U3762 (N_3762,N_3277,N_3329);
and U3763 (N_3763,N_3484,N_3359);
and U3764 (N_3764,N_3411,N_3114);
nand U3765 (N_3765,N_3246,N_3423);
or U3766 (N_3766,N_3477,N_3372);
nor U3767 (N_3767,N_3303,N_3265);
nor U3768 (N_3768,N_3075,N_3202);
and U3769 (N_3769,N_3467,N_3045);
nor U3770 (N_3770,N_3438,N_3496);
and U3771 (N_3771,N_3452,N_3176);
and U3772 (N_3772,N_3370,N_3138);
xor U3773 (N_3773,N_3074,N_3157);
xnor U3774 (N_3774,N_3287,N_3327);
xnor U3775 (N_3775,N_3379,N_3270);
and U3776 (N_3776,N_3037,N_3068);
nand U3777 (N_3777,N_3399,N_3249);
and U3778 (N_3778,N_3320,N_3465);
and U3779 (N_3779,N_3466,N_3267);
nor U3780 (N_3780,N_3348,N_3262);
xor U3781 (N_3781,N_3370,N_3277);
or U3782 (N_3782,N_3398,N_3049);
nand U3783 (N_3783,N_3488,N_3127);
xor U3784 (N_3784,N_3406,N_3306);
nor U3785 (N_3785,N_3480,N_3154);
nor U3786 (N_3786,N_3164,N_3080);
nand U3787 (N_3787,N_3313,N_3216);
nand U3788 (N_3788,N_3311,N_3344);
and U3789 (N_3789,N_3322,N_3388);
or U3790 (N_3790,N_3006,N_3482);
and U3791 (N_3791,N_3487,N_3416);
and U3792 (N_3792,N_3480,N_3015);
or U3793 (N_3793,N_3074,N_3387);
or U3794 (N_3794,N_3429,N_3440);
nor U3795 (N_3795,N_3295,N_3476);
or U3796 (N_3796,N_3169,N_3484);
nor U3797 (N_3797,N_3229,N_3098);
nand U3798 (N_3798,N_3266,N_3052);
xor U3799 (N_3799,N_3327,N_3189);
nand U3800 (N_3800,N_3065,N_3307);
xor U3801 (N_3801,N_3359,N_3427);
nor U3802 (N_3802,N_3421,N_3226);
and U3803 (N_3803,N_3024,N_3487);
and U3804 (N_3804,N_3448,N_3496);
nand U3805 (N_3805,N_3201,N_3401);
nand U3806 (N_3806,N_3311,N_3447);
nand U3807 (N_3807,N_3170,N_3391);
xor U3808 (N_3808,N_3031,N_3307);
xnor U3809 (N_3809,N_3264,N_3166);
and U3810 (N_3810,N_3345,N_3394);
nor U3811 (N_3811,N_3066,N_3456);
nor U3812 (N_3812,N_3045,N_3431);
or U3813 (N_3813,N_3279,N_3269);
and U3814 (N_3814,N_3346,N_3066);
nor U3815 (N_3815,N_3168,N_3004);
and U3816 (N_3816,N_3073,N_3461);
and U3817 (N_3817,N_3357,N_3034);
xor U3818 (N_3818,N_3304,N_3299);
and U3819 (N_3819,N_3314,N_3023);
xor U3820 (N_3820,N_3380,N_3492);
nor U3821 (N_3821,N_3069,N_3464);
xnor U3822 (N_3822,N_3209,N_3012);
or U3823 (N_3823,N_3302,N_3086);
and U3824 (N_3824,N_3467,N_3328);
or U3825 (N_3825,N_3342,N_3259);
xor U3826 (N_3826,N_3158,N_3051);
or U3827 (N_3827,N_3430,N_3028);
or U3828 (N_3828,N_3105,N_3284);
or U3829 (N_3829,N_3437,N_3329);
or U3830 (N_3830,N_3232,N_3126);
nand U3831 (N_3831,N_3200,N_3305);
nand U3832 (N_3832,N_3341,N_3193);
nand U3833 (N_3833,N_3455,N_3459);
xnor U3834 (N_3834,N_3329,N_3311);
xnor U3835 (N_3835,N_3461,N_3254);
nor U3836 (N_3836,N_3023,N_3238);
nand U3837 (N_3837,N_3260,N_3415);
xnor U3838 (N_3838,N_3004,N_3150);
and U3839 (N_3839,N_3122,N_3390);
nor U3840 (N_3840,N_3360,N_3343);
and U3841 (N_3841,N_3193,N_3207);
nand U3842 (N_3842,N_3402,N_3197);
xor U3843 (N_3843,N_3148,N_3380);
and U3844 (N_3844,N_3330,N_3320);
xnor U3845 (N_3845,N_3418,N_3048);
nor U3846 (N_3846,N_3064,N_3328);
nor U3847 (N_3847,N_3073,N_3239);
and U3848 (N_3848,N_3185,N_3180);
nor U3849 (N_3849,N_3332,N_3498);
nand U3850 (N_3850,N_3394,N_3422);
xnor U3851 (N_3851,N_3134,N_3430);
or U3852 (N_3852,N_3138,N_3176);
nand U3853 (N_3853,N_3173,N_3276);
or U3854 (N_3854,N_3220,N_3007);
or U3855 (N_3855,N_3272,N_3242);
nor U3856 (N_3856,N_3314,N_3122);
and U3857 (N_3857,N_3285,N_3277);
or U3858 (N_3858,N_3146,N_3319);
and U3859 (N_3859,N_3027,N_3163);
nor U3860 (N_3860,N_3189,N_3002);
and U3861 (N_3861,N_3036,N_3285);
nor U3862 (N_3862,N_3057,N_3114);
and U3863 (N_3863,N_3494,N_3421);
xor U3864 (N_3864,N_3148,N_3129);
and U3865 (N_3865,N_3014,N_3443);
nor U3866 (N_3866,N_3040,N_3463);
and U3867 (N_3867,N_3391,N_3115);
nand U3868 (N_3868,N_3051,N_3072);
nor U3869 (N_3869,N_3454,N_3303);
nor U3870 (N_3870,N_3392,N_3477);
and U3871 (N_3871,N_3139,N_3494);
nand U3872 (N_3872,N_3466,N_3068);
and U3873 (N_3873,N_3242,N_3471);
xnor U3874 (N_3874,N_3210,N_3153);
or U3875 (N_3875,N_3159,N_3400);
xor U3876 (N_3876,N_3475,N_3378);
xnor U3877 (N_3877,N_3234,N_3254);
and U3878 (N_3878,N_3457,N_3039);
xor U3879 (N_3879,N_3318,N_3228);
xor U3880 (N_3880,N_3384,N_3134);
and U3881 (N_3881,N_3458,N_3379);
or U3882 (N_3882,N_3440,N_3156);
xnor U3883 (N_3883,N_3490,N_3311);
xnor U3884 (N_3884,N_3163,N_3046);
nand U3885 (N_3885,N_3467,N_3072);
nand U3886 (N_3886,N_3282,N_3443);
and U3887 (N_3887,N_3305,N_3496);
nor U3888 (N_3888,N_3384,N_3063);
and U3889 (N_3889,N_3251,N_3453);
or U3890 (N_3890,N_3007,N_3278);
nor U3891 (N_3891,N_3337,N_3032);
nor U3892 (N_3892,N_3477,N_3359);
xor U3893 (N_3893,N_3195,N_3174);
and U3894 (N_3894,N_3081,N_3109);
or U3895 (N_3895,N_3424,N_3212);
or U3896 (N_3896,N_3209,N_3322);
xnor U3897 (N_3897,N_3330,N_3054);
nor U3898 (N_3898,N_3061,N_3370);
xnor U3899 (N_3899,N_3359,N_3263);
nor U3900 (N_3900,N_3090,N_3114);
nor U3901 (N_3901,N_3360,N_3489);
nor U3902 (N_3902,N_3003,N_3361);
xor U3903 (N_3903,N_3217,N_3225);
nand U3904 (N_3904,N_3478,N_3125);
and U3905 (N_3905,N_3308,N_3140);
or U3906 (N_3906,N_3248,N_3084);
nor U3907 (N_3907,N_3314,N_3084);
xor U3908 (N_3908,N_3210,N_3416);
nand U3909 (N_3909,N_3348,N_3481);
and U3910 (N_3910,N_3402,N_3199);
nand U3911 (N_3911,N_3239,N_3339);
nand U3912 (N_3912,N_3083,N_3121);
nand U3913 (N_3913,N_3335,N_3047);
xnor U3914 (N_3914,N_3127,N_3335);
and U3915 (N_3915,N_3443,N_3487);
xnor U3916 (N_3916,N_3366,N_3276);
and U3917 (N_3917,N_3120,N_3094);
xnor U3918 (N_3918,N_3046,N_3263);
and U3919 (N_3919,N_3427,N_3351);
and U3920 (N_3920,N_3473,N_3101);
nor U3921 (N_3921,N_3460,N_3418);
nor U3922 (N_3922,N_3300,N_3296);
xor U3923 (N_3923,N_3269,N_3433);
nand U3924 (N_3924,N_3020,N_3385);
or U3925 (N_3925,N_3319,N_3276);
nand U3926 (N_3926,N_3143,N_3299);
or U3927 (N_3927,N_3133,N_3232);
nor U3928 (N_3928,N_3263,N_3318);
nor U3929 (N_3929,N_3071,N_3115);
or U3930 (N_3930,N_3128,N_3007);
nand U3931 (N_3931,N_3302,N_3004);
and U3932 (N_3932,N_3165,N_3361);
or U3933 (N_3933,N_3327,N_3332);
or U3934 (N_3934,N_3086,N_3061);
and U3935 (N_3935,N_3458,N_3044);
nand U3936 (N_3936,N_3441,N_3317);
xnor U3937 (N_3937,N_3182,N_3325);
nand U3938 (N_3938,N_3409,N_3303);
nand U3939 (N_3939,N_3017,N_3035);
nor U3940 (N_3940,N_3356,N_3291);
and U3941 (N_3941,N_3316,N_3208);
nor U3942 (N_3942,N_3031,N_3458);
or U3943 (N_3943,N_3135,N_3491);
nand U3944 (N_3944,N_3266,N_3302);
or U3945 (N_3945,N_3497,N_3035);
nor U3946 (N_3946,N_3032,N_3039);
xnor U3947 (N_3947,N_3494,N_3195);
nand U3948 (N_3948,N_3199,N_3453);
or U3949 (N_3949,N_3345,N_3463);
and U3950 (N_3950,N_3284,N_3062);
and U3951 (N_3951,N_3244,N_3252);
and U3952 (N_3952,N_3107,N_3387);
xnor U3953 (N_3953,N_3174,N_3443);
and U3954 (N_3954,N_3245,N_3362);
and U3955 (N_3955,N_3198,N_3258);
or U3956 (N_3956,N_3380,N_3067);
nand U3957 (N_3957,N_3154,N_3469);
xor U3958 (N_3958,N_3073,N_3045);
xor U3959 (N_3959,N_3068,N_3283);
nand U3960 (N_3960,N_3487,N_3073);
and U3961 (N_3961,N_3455,N_3492);
and U3962 (N_3962,N_3187,N_3435);
nand U3963 (N_3963,N_3257,N_3042);
xor U3964 (N_3964,N_3302,N_3332);
xor U3965 (N_3965,N_3379,N_3091);
xnor U3966 (N_3966,N_3390,N_3417);
and U3967 (N_3967,N_3402,N_3253);
and U3968 (N_3968,N_3239,N_3355);
nor U3969 (N_3969,N_3074,N_3168);
and U3970 (N_3970,N_3075,N_3082);
xnor U3971 (N_3971,N_3430,N_3299);
and U3972 (N_3972,N_3369,N_3110);
and U3973 (N_3973,N_3333,N_3322);
nand U3974 (N_3974,N_3493,N_3465);
xor U3975 (N_3975,N_3041,N_3147);
nor U3976 (N_3976,N_3481,N_3359);
nand U3977 (N_3977,N_3176,N_3254);
nor U3978 (N_3978,N_3325,N_3419);
xnor U3979 (N_3979,N_3414,N_3370);
xnor U3980 (N_3980,N_3418,N_3080);
or U3981 (N_3981,N_3103,N_3220);
nand U3982 (N_3982,N_3384,N_3111);
and U3983 (N_3983,N_3334,N_3394);
and U3984 (N_3984,N_3281,N_3286);
or U3985 (N_3985,N_3214,N_3109);
and U3986 (N_3986,N_3115,N_3479);
or U3987 (N_3987,N_3229,N_3189);
and U3988 (N_3988,N_3416,N_3100);
nand U3989 (N_3989,N_3357,N_3425);
xor U3990 (N_3990,N_3115,N_3392);
nor U3991 (N_3991,N_3437,N_3308);
nand U3992 (N_3992,N_3168,N_3137);
or U3993 (N_3993,N_3483,N_3181);
or U3994 (N_3994,N_3352,N_3444);
xor U3995 (N_3995,N_3396,N_3016);
and U3996 (N_3996,N_3129,N_3302);
xor U3997 (N_3997,N_3113,N_3429);
xnor U3998 (N_3998,N_3120,N_3289);
xor U3999 (N_3999,N_3448,N_3025);
nor U4000 (N_4000,N_3880,N_3999);
xnor U4001 (N_4001,N_3682,N_3833);
nand U4002 (N_4002,N_3524,N_3981);
or U4003 (N_4003,N_3852,N_3867);
xor U4004 (N_4004,N_3707,N_3713);
nor U4005 (N_4005,N_3757,N_3684);
or U4006 (N_4006,N_3797,N_3886);
nand U4007 (N_4007,N_3868,N_3950);
or U4008 (N_4008,N_3882,N_3862);
and U4009 (N_4009,N_3541,N_3975);
nor U4010 (N_4010,N_3946,N_3941);
nand U4011 (N_4011,N_3835,N_3515);
and U4012 (N_4012,N_3751,N_3562);
nand U4013 (N_4013,N_3896,N_3702);
and U4014 (N_4014,N_3724,N_3501);
nor U4015 (N_4015,N_3934,N_3727);
and U4016 (N_4016,N_3508,N_3506);
nor U4017 (N_4017,N_3874,N_3722);
nand U4018 (N_4018,N_3526,N_3692);
or U4019 (N_4019,N_3641,N_3669);
nand U4020 (N_4020,N_3772,N_3790);
nand U4021 (N_4021,N_3788,N_3634);
and U4022 (N_4022,N_3918,N_3924);
nand U4023 (N_4023,N_3601,N_3770);
xor U4024 (N_4024,N_3542,N_3813);
xnor U4025 (N_4025,N_3728,N_3741);
and U4026 (N_4026,N_3588,N_3858);
or U4027 (N_4027,N_3709,N_3939);
nand U4028 (N_4028,N_3746,N_3584);
xnor U4029 (N_4029,N_3533,N_3875);
or U4030 (N_4030,N_3881,N_3899);
nor U4031 (N_4031,N_3587,N_3949);
xor U4032 (N_4032,N_3830,N_3642);
and U4033 (N_4033,N_3943,N_3839);
or U4034 (N_4034,N_3814,N_3937);
xnor U4035 (N_4035,N_3805,N_3905);
xor U4036 (N_4036,N_3894,N_3661);
nor U4037 (N_4037,N_3982,N_3958);
xnor U4038 (N_4038,N_3804,N_3631);
and U4039 (N_4039,N_3556,N_3566);
nand U4040 (N_4040,N_3753,N_3603);
or U4041 (N_4041,N_3683,N_3764);
xor U4042 (N_4042,N_3820,N_3983);
and U4043 (N_4043,N_3885,N_3694);
xnor U4044 (N_4044,N_3523,N_3745);
or U4045 (N_4045,N_3717,N_3645);
and U4046 (N_4046,N_3915,N_3596);
nor U4047 (N_4047,N_3824,N_3942);
xor U4048 (N_4048,N_3961,N_3914);
xor U4049 (N_4049,N_3926,N_3655);
xor U4050 (N_4050,N_3838,N_3505);
nand U4051 (N_4051,N_3701,N_3929);
xnor U4052 (N_4052,N_3966,N_3906);
nor U4053 (N_4053,N_3628,N_3768);
xnor U4054 (N_4054,N_3968,N_3917);
nor U4055 (N_4055,N_3734,N_3627);
nand U4056 (N_4056,N_3602,N_3763);
nand U4057 (N_4057,N_3554,N_3795);
xnor U4058 (N_4058,N_3671,N_3612);
nor U4059 (N_4059,N_3643,N_3743);
nand U4060 (N_4060,N_3887,N_3986);
nor U4061 (N_4061,N_3545,N_3831);
xor U4062 (N_4062,N_3715,N_3582);
nor U4063 (N_4063,N_3985,N_3590);
nand U4064 (N_4064,N_3555,N_3619);
xor U4065 (N_4065,N_3606,N_3739);
xnor U4066 (N_4066,N_3599,N_3513);
nor U4067 (N_4067,N_3687,N_3546);
and U4068 (N_4068,N_3898,N_3577);
xnor U4069 (N_4069,N_3570,N_3615);
or U4070 (N_4070,N_3581,N_3654);
and U4071 (N_4071,N_3879,N_3931);
or U4072 (N_4072,N_3689,N_3826);
xnor U4073 (N_4073,N_3793,N_3580);
nor U4074 (N_4074,N_3696,N_3605);
nor U4075 (N_4075,N_3691,N_3752);
nand U4076 (N_4076,N_3668,N_3823);
and U4077 (N_4077,N_3667,N_3877);
nand U4078 (N_4078,N_3940,N_3973);
nor U4079 (N_4079,N_3796,N_3552);
and U4080 (N_4080,N_3547,N_3571);
nor U4081 (N_4081,N_3510,N_3742);
nor U4082 (N_4082,N_3923,N_3889);
and U4083 (N_4083,N_3652,N_3507);
or U4084 (N_4084,N_3632,N_3543);
xor U4085 (N_4085,N_3732,N_3700);
or U4086 (N_4086,N_3676,N_3851);
xnor U4087 (N_4087,N_3716,N_3800);
xor U4088 (N_4088,N_3675,N_3551);
or U4089 (N_4089,N_3609,N_3569);
xnor U4090 (N_4090,N_3616,N_3540);
or U4091 (N_4091,N_3792,N_3598);
nor U4092 (N_4092,N_3686,N_3829);
xor U4093 (N_4093,N_3884,N_3677);
nor U4094 (N_4094,N_3821,N_3782);
nand U4095 (N_4095,N_3725,N_3892);
or U4096 (N_4096,N_3840,N_3553);
xnor U4097 (N_4097,N_3807,N_3780);
and U4098 (N_4098,N_3964,N_3936);
and U4099 (N_4099,N_3878,N_3784);
nand U4100 (N_4100,N_3567,N_3902);
xnor U4101 (N_4101,N_3980,N_3626);
or U4102 (N_4102,N_3591,N_3955);
nand U4103 (N_4103,N_3754,N_3673);
and U4104 (N_4104,N_3954,N_3729);
xnor U4105 (N_4105,N_3514,N_3520);
xor U4106 (N_4106,N_3697,N_3565);
xnor U4107 (N_4107,N_3624,N_3842);
or U4108 (N_4108,N_3965,N_3883);
nor U4109 (N_4109,N_3978,N_3657);
nor U4110 (N_4110,N_3895,N_3748);
nand U4111 (N_4111,N_3910,N_3756);
nand U4112 (N_4112,N_3731,N_3576);
nor U4113 (N_4113,N_3620,N_3815);
or U4114 (N_4114,N_3755,N_3922);
nand U4115 (N_4115,N_3783,N_3802);
and U4116 (N_4116,N_3798,N_3903);
nor U4117 (N_4117,N_3575,N_3749);
xor U4118 (N_4118,N_3776,N_3803);
or U4119 (N_4119,N_3809,N_3561);
nor U4120 (N_4120,N_3549,N_3614);
or U4121 (N_4121,N_3993,N_3572);
and U4122 (N_4122,N_3819,N_3679);
nand U4123 (N_4123,N_3818,N_3633);
or U4124 (N_4124,N_3738,N_3623);
nand U4125 (N_4125,N_3859,N_3557);
or U4126 (N_4126,N_3618,N_3998);
and U4127 (N_4127,N_3947,N_3512);
nand U4128 (N_4128,N_3647,N_3503);
and U4129 (N_4129,N_3951,N_3919);
and U4130 (N_4130,N_3997,N_3927);
and U4131 (N_4131,N_3876,N_3908);
and U4132 (N_4132,N_3733,N_3854);
nor U4133 (N_4133,N_3989,N_3573);
and U4134 (N_4134,N_3737,N_3629);
nor U4135 (N_4135,N_3843,N_3608);
xor U4136 (N_4136,N_3900,N_3970);
and U4137 (N_4137,N_3856,N_3688);
xnor U4138 (N_4138,N_3786,N_3967);
nand U4139 (N_4139,N_3944,N_3904);
nand U4140 (N_4140,N_3893,N_3718);
xor U4141 (N_4141,N_3644,N_3777);
or U4142 (N_4142,N_3962,N_3848);
nand U4143 (N_4143,N_3959,N_3604);
or U4144 (N_4144,N_3550,N_3538);
and U4145 (N_4145,N_3656,N_3670);
nor U4146 (N_4146,N_3680,N_3617);
xnor U4147 (N_4147,N_3622,N_3744);
and U4148 (N_4148,N_3646,N_3897);
nand U4149 (N_4149,N_3866,N_3945);
and U4150 (N_4150,N_3834,N_3960);
nor U4151 (N_4151,N_3522,N_3971);
nand U4152 (N_4152,N_3853,N_3963);
xor U4153 (N_4153,N_3518,N_3630);
nor U4154 (N_4154,N_3594,N_3911);
nand U4155 (N_4155,N_3850,N_3695);
nor U4156 (N_4156,N_3789,N_3771);
or U4157 (N_4157,N_3791,N_3828);
nor U4158 (N_4158,N_3996,N_3901);
and U4159 (N_4159,N_3909,N_3787);
and U4160 (N_4160,N_3698,N_3650);
and U4161 (N_4161,N_3593,N_3560);
or U4162 (N_4162,N_3952,N_3761);
nor U4163 (N_4163,N_3595,N_3703);
nor U4164 (N_4164,N_3600,N_3665);
and U4165 (N_4165,N_3990,N_3736);
nand U4166 (N_4166,N_3636,N_3544);
nand U4167 (N_4167,N_3504,N_3649);
nand U4168 (N_4168,N_3871,N_3855);
xor U4169 (N_4169,N_3660,N_3706);
and U4170 (N_4170,N_3579,N_3583);
and U4171 (N_4171,N_3810,N_3648);
nand U4172 (N_4172,N_3653,N_3511);
nand U4173 (N_4173,N_3827,N_3864);
or U4174 (N_4174,N_3953,N_3863);
nand U4175 (N_4175,N_3747,N_3708);
xor U4176 (N_4176,N_3585,N_3726);
or U4177 (N_4177,N_3625,N_3563);
xor U4178 (N_4178,N_3516,N_3502);
xor U4179 (N_4179,N_3638,N_3607);
nor U4180 (N_4180,N_3740,N_3735);
nand U4181 (N_4181,N_3832,N_3872);
and U4182 (N_4182,N_3844,N_3811);
and U4183 (N_4183,N_3509,N_3532);
nand U4184 (N_4184,N_3935,N_3586);
and U4185 (N_4185,N_3711,N_3956);
nand U4186 (N_4186,N_3597,N_3710);
and U4187 (N_4187,N_3765,N_3837);
nor U4188 (N_4188,N_3678,N_3979);
or U4189 (N_4189,N_3521,N_3925);
and U4190 (N_4190,N_3912,N_3558);
nand U4191 (N_4191,N_3822,N_3773);
nor U4192 (N_4192,N_3760,N_3801);
and U4193 (N_4193,N_3666,N_3992);
or U4194 (N_4194,N_3613,N_3991);
xor U4195 (N_4195,N_3775,N_3530);
xnor U4196 (N_4196,N_3988,N_3564);
and U4197 (N_4197,N_3534,N_3976);
nand U4198 (N_4198,N_3995,N_3723);
nor U4199 (N_4199,N_3778,N_3681);
nand U4200 (N_4200,N_3559,N_3704);
and U4201 (N_4201,N_3930,N_3948);
and U4202 (N_4202,N_3860,N_3535);
nand U4203 (N_4203,N_3719,N_3674);
xnor U4204 (N_4204,N_3525,N_3519);
xnor U4205 (N_4205,N_3799,N_3816);
and U4206 (N_4206,N_3621,N_3640);
and U4207 (N_4207,N_3994,N_3610);
and U4208 (N_4208,N_3658,N_3846);
or U4209 (N_4209,N_3869,N_3500);
nor U4210 (N_4210,N_3536,N_3664);
xor U4211 (N_4211,N_3779,N_3766);
or U4212 (N_4212,N_3517,N_3977);
nand U4213 (N_4213,N_3712,N_3806);
nand U4214 (N_4214,N_3750,N_3891);
nor U4215 (N_4215,N_3865,N_3984);
nand U4216 (N_4216,N_3699,N_3527);
or U4217 (N_4217,N_3920,N_3888);
and U4218 (N_4218,N_3913,N_3662);
nand U4219 (N_4219,N_3932,N_3651);
xnor U4220 (N_4220,N_3589,N_3714);
nand U4221 (N_4221,N_3825,N_3721);
nor U4222 (N_4222,N_3812,N_3857);
nand U4223 (N_4223,N_3663,N_3672);
or U4224 (N_4224,N_3592,N_3916);
xnor U4225 (N_4225,N_3759,N_3568);
nand U4226 (N_4226,N_3861,N_3528);
xnor U4227 (N_4227,N_3957,N_3873);
xnor U4228 (N_4228,N_3836,N_3921);
nand U4229 (N_4229,N_3987,N_3529);
xnor U4230 (N_4230,N_3659,N_3890);
or U4231 (N_4231,N_3774,N_3767);
nand U4232 (N_4232,N_3972,N_3637);
nor U4233 (N_4233,N_3578,N_3537);
nor U4234 (N_4234,N_3611,N_3685);
nor U4235 (N_4235,N_3730,N_3781);
and U4236 (N_4236,N_3847,N_3928);
nor U4237 (N_4237,N_3762,N_3974);
or U4238 (N_4238,N_3548,N_3639);
or U4239 (N_4239,N_3794,N_3969);
xor U4240 (N_4240,N_3635,N_3817);
or U4241 (N_4241,N_3841,N_3531);
nand U4242 (N_4242,N_3539,N_3870);
nand U4243 (N_4243,N_3938,N_3690);
nand U4244 (N_4244,N_3808,N_3785);
and U4245 (N_4245,N_3769,N_3845);
and U4246 (N_4246,N_3720,N_3705);
nand U4247 (N_4247,N_3907,N_3758);
or U4248 (N_4248,N_3933,N_3693);
or U4249 (N_4249,N_3849,N_3574);
or U4250 (N_4250,N_3510,N_3889);
xor U4251 (N_4251,N_3827,N_3662);
and U4252 (N_4252,N_3888,N_3795);
and U4253 (N_4253,N_3905,N_3932);
or U4254 (N_4254,N_3983,N_3919);
and U4255 (N_4255,N_3969,N_3653);
nor U4256 (N_4256,N_3544,N_3845);
nand U4257 (N_4257,N_3617,N_3791);
and U4258 (N_4258,N_3661,N_3891);
or U4259 (N_4259,N_3542,N_3854);
or U4260 (N_4260,N_3685,N_3937);
or U4261 (N_4261,N_3713,N_3855);
xor U4262 (N_4262,N_3913,N_3858);
or U4263 (N_4263,N_3756,N_3688);
nand U4264 (N_4264,N_3665,N_3814);
nor U4265 (N_4265,N_3533,N_3628);
nand U4266 (N_4266,N_3927,N_3756);
nand U4267 (N_4267,N_3763,N_3867);
nand U4268 (N_4268,N_3940,N_3513);
nand U4269 (N_4269,N_3635,N_3673);
nand U4270 (N_4270,N_3905,N_3506);
nor U4271 (N_4271,N_3577,N_3546);
xnor U4272 (N_4272,N_3724,N_3809);
nor U4273 (N_4273,N_3842,N_3808);
nand U4274 (N_4274,N_3916,N_3887);
and U4275 (N_4275,N_3734,N_3635);
or U4276 (N_4276,N_3720,N_3728);
and U4277 (N_4277,N_3918,N_3732);
nor U4278 (N_4278,N_3740,N_3596);
or U4279 (N_4279,N_3812,N_3526);
and U4280 (N_4280,N_3944,N_3892);
nand U4281 (N_4281,N_3754,N_3669);
and U4282 (N_4282,N_3937,N_3890);
or U4283 (N_4283,N_3655,N_3703);
or U4284 (N_4284,N_3929,N_3623);
or U4285 (N_4285,N_3636,N_3852);
and U4286 (N_4286,N_3800,N_3586);
or U4287 (N_4287,N_3577,N_3523);
or U4288 (N_4288,N_3967,N_3690);
nand U4289 (N_4289,N_3941,N_3640);
xnor U4290 (N_4290,N_3627,N_3836);
nor U4291 (N_4291,N_3550,N_3688);
or U4292 (N_4292,N_3523,N_3512);
nor U4293 (N_4293,N_3600,N_3664);
and U4294 (N_4294,N_3646,N_3825);
or U4295 (N_4295,N_3652,N_3842);
nor U4296 (N_4296,N_3519,N_3915);
or U4297 (N_4297,N_3801,N_3750);
nor U4298 (N_4298,N_3724,N_3731);
nand U4299 (N_4299,N_3617,N_3926);
and U4300 (N_4300,N_3955,N_3825);
nor U4301 (N_4301,N_3936,N_3624);
nor U4302 (N_4302,N_3971,N_3891);
nand U4303 (N_4303,N_3872,N_3729);
or U4304 (N_4304,N_3570,N_3894);
and U4305 (N_4305,N_3632,N_3607);
or U4306 (N_4306,N_3934,N_3604);
xnor U4307 (N_4307,N_3531,N_3661);
or U4308 (N_4308,N_3702,N_3784);
xnor U4309 (N_4309,N_3935,N_3795);
and U4310 (N_4310,N_3553,N_3946);
and U4311 (N_4311,N_3530,N_3503);
nor U4312 (N_4312,N_3893,N_3625);
nand U4313 (N_4313,N_3944,N_3529);
and U4314 (N_4314,N_3632,N_3949);
xnor U4315 (N_4315,N_3588,N_3637);
xnor U4316 (N_4316,N_3652,N_3581);
or U4317 (N_4317,N_3797,N_3707);
and U4318 (N_4318,N_3577,N_3760);
or U4319 (N_4319,N_3525,N_3845);
or U4320 (N_4320,N_3571,N_3917);
xor U4321 (N_4321,N_3908,N_3965);
and U4322 (N_4322,N_3639,N_3913);
xor U4323 (N_4323,N_3522,N_3548);
nand U4324 (N_4324,N_3729,N_3558);
nand U4325 (N_4325,N_3927,N_3773);
xnor U4326 (N_4326,N_3981,N_3850);
nand U4327 (N_4327,N_3888,N_3897);
nor U4328 (N_4328,N_3824,N_3655);
xnor U4329 (N_4329,N_3540,N_3615);
nor U4330 (N_4330,N_3521,N_3866);
and U4331 (N_4331,N_3998,N_3944);
nor U4332 (N_4332,N_3768,N_3734);
xor U4333 (N_4333,N_3501,N_3883);
and U4334 (N_4334,N_3891,N_3716);
and U4335 (N_4335,N_3753,N_3882);
and U4336 (N_4336,N_3518,N_3613);
nand U4337 (N_4337,N_3991,N_3521);
xor U4338 (N_4338,N_3808,N_3876);
nand U4339 (N_4339,N_3718,N_3596);
nand U4340 (N_4340,N_3626,N_3889);
xor U4341 (N_4341,N_3961,N_3660);
and U4342 (N_4342,N_3792,N_3846);
and U4343 (N_4343,N_3909,N_3548);
nor U4344 (N_4344,N_3542,N_3601);
nand U4345 (N_4345,N_3871,N_3712);
nor U4346 (N_4346,N_3855,N_3612);
nand U4347 (N_4347,N_3992,N_3789);
nand U4348 (N_4348,N_3602,N_3719);
nand U4349 (N_4349,N_3885,N_3818);
or U4350 (N_4350,N_3909,N_3862);
and U4351 (N_4351,N_3552,N_3845);
nand U4352 (N_4352,N_3760,N_3579);
nand U4353 (N_4353,N_3522,N_3992);
xnor U4354 (N_4354,N_3918,N_3851);
nand U4355 (N_4355,N_3996,N_3719);
nand U4356 (N_4356,N_3980,N_3659);
and U4357 (N_4357,N_3505,N_3631);
and U4358 (N_4358,N_3657,N_3909);
or U4359 (N_4359,N_3656,N_3778);
nor U4360 (N_4360,N_3915,N_3965);
nor U4361 (N_4361,N_3883,N_3897);
and U4362 (N_4362,N_3934,N_3628);
or U4363 (N_4363,N_3807,N_3573);
nand U4364 (N_4364,N_3646,N_3925);
or U4365 (N_4365,N_3514,N_3657);
or U4366 (N_4366,N_3936,N_3687);
and U4367 (N_4367,N_3905,N_3672);
nand U4368 (N_4368,N_3687,N_3859);
or U4369 (N_4369,N_3904,N_3848);
and U4370 (N_4370,N_3970,N_3799);
or U4371 (N_4371,N_3610,N_3667);
nor U4372 (N_4372,N_3742,N_3814);
nand U4373 (N_4373,N_3990,N_3652);
or U4374 (N_4374,N_3903,N_3632);
xnor U4375 (N_4375,N_3534,N_3999);
xnor U4376 (N_4376,N_3622,N_3662);
xor U4377 (N_4377,N_3791,N_3940);
nand U4378 (N_4378,N_3759,N_3528);
xor U4379 (N_4379,N_3570,N_3790);
xor U4380 (N_4380,N_3962,N_3500);
xnor U4381 (N_4381,N_3948,N_3718);
xnor U4382 (N_4382,N_3684,N_3953);
or U4383 (N_4383,N_3962,N_3616);
nand U4384 (N_4384,N_3601,N_3781);
and U4385 (N_4385,N_3703,N_3542);
and U4386 (N_4386,N_3624,N_3650);
xnor U4387 (N_4387,N_3959,N_3887);
or U4388 (N_4388,N_3968,N_3647);
and U4389 (N_4389,N_3929,N_3520);
xnor U4390 (N_4390,N_3821,N_3904);
nor U4391 (N_4391,N_3572,N_3746);
nor U4392 (N_4392,N_3890,N_3566);
and U4393 (N_4393,N_3831,N_3747);
xor U4394 (N_4394,N_3984,N_3540);
nor U4395 (N_4395,N_3506,N_3538);
nor U4396 (N_4396,N_3676,N_3945);
and U4397 (N_4397,N_3550,N_3677);
xnor U4398 (N_4398,N_3642,N_3560);
nand U4399 (N_4399,N_3796,N_3531);
nor U4400 (N_4400,N_3929,N_3928);
and U4401 (N_4401,N_3788,N_3949);
nand U4402 (N_4402,N_3767,N_3899);
xnor U4403 (N_4403,N_3521,N_3667);
nor U4404 (N_4404,N_3977,N_3661);
or U4405 (N_4405,N_3771,N_3629);
xor U4406 (N_4406,N_3966,N_3753);
or U4407 (N_4407,N_3701,N_3656);
xnor U4408 (N_4408,N_3928,N_3672);
nand U4409 (N_4409,N_3994,N_3560);
and U4410 (N_4410,N_3701,N_3930);
nand U4411 (N_4411,N_3526,N_3677);
nand U4412 (N_4412,N_3545,N_3760);
nand U4413 (N_4413,N_3599,N_3801);
nand U4414 (N_4414,N_3898,N_3695);
and U4415 (N_4415,N_3604,N_3750);
or U4416 (N_4416,N_3532,N_3643);
or U4417 (N_4417,N_3922,N_3911);
or U4418 (N_4418,N_3968,N_3726);
and U4419 (N_4419,N_3786,N_3918);
or U4420 (N_4420,N_3833,N_3673);
or U4421 (N_4421,N_3655,N_3865);
nand U4422 (N_4422,N_3645,N_3562);
and U4423 (N_4423,N_3657,N_3925);
nand U4424 (N_4424,N_3648,N_3511);
or U4425 (N_4425,N_3627,N_3992);
xnor U4426 (N_4426,N_3525,N_3685);
xor U4427 (N_4427,N_3900,N_3593);
or U4428 (N_4428,N_3523,N_3655);
nor U4429 (N_4429,N_3698,N_3882);
or U4430 (N_4430,N_3742,N_3993);
nor U4431 (N_4431,N_3700,N_3886);
nand U4432 (N_4432,N_3537,N_3544);
xnor U4433 (N_4433,N_3710,N_3888);
nor U4434 (N_4434,N_3853,N_3882);
nor U4435 (N_4435,N_3635,N_3718);
and U4436 (N_4436,N_3733,N_3932);
nor U4437 (N_4437,N_3627,N_3804);
or U4438 (N_4438,N_3631,N_3838);
and U4439 (N_4439,N_3956,N_3519);
nand U4440 (N_4440,N_3506,N_3938);
nor U4441 (N_4441,N_3817,N_3908);
nor U4442 (N_4442,N_3962,N_3889);
and U4443 (N_4443,N_3857,N_3643);
nand U4444 (N_4444,N_3622,N_3532);
xnor U4445 (N_4445,N_3625,N_3780);
or U4446 (N_4446,N_3891,N_3824);
xnor U4447 (N_4447,N_3688,N_3968);
and U4448 (N_4448,N_3927,N_3763);
nand U4449 (N_4449,N_3905,N_3615);
or U4450 (N_4450,N_3915,N_3806);
nor U4451 (N_4451,N_3896,N_3961);
nor U4452 (N_4452,N_3563,N_3983);
nor U4453 (N_4453,N_3941,N_3676);
xor U4454 (N_4454,N_3919,N_3599);
and U4455 (N_4455,N_3884,N_3776);
nand U4456 (N_4456,N_3796,N_3919);
and U4457 (N_4457,N_3806,N_3616);
nor U4458 (N_4458,N_3685,N_3631);
and U4459 (N_4459,N_3802,N_3923);
nand U4460 (N_4460,N_3687,N_3560);
or U4461 (N_4461,N_3738,N_3823);
and U4462 (N_4462,N_3552,N_3968);
or U4463 (N_4463,N_3661,N_3611);
xor U4464 (N_4464,N_3549,N_3851);
or U4465 (N_4465,N_3598,N_3760);
nor U4466 (N_4466,N_3654,N_3897);
xor U4467 (N_4467,N_3854,N_3992);
and U4468 (N_4468,N_3526,N_3724);
nor U4469 (N_4469,N_3649,N_3617);
and U4470 (N_4470,N_3857,N_3879);
and U4471 (N_4471,N_3679,N_3793);
nor U4472 (N_4472,N_3807,N_3525);
nand U4473 (N_4473,N_3994,N_3792);
and U4474 (N_4474,N_3897,N_3934);
xor U4475 (N_4475,N_3685,N_3647);
or U4476 (N_4476,N_3541,N_3634);
nor U4477 (N_4477,N_3677,N_3820);
xor U4478 (N_4478,N_3737,N_3537);
nand U4479 (N_4479,N_3709,N_3820);
nor U4480 (N_4480,N_3693,N_3805);
or U4481 (N_4481,N_3799,N_3710);
and U4482 (N_4482,N_3848,N_3718);
xnor U4483 (N_4483,N_3826,N_3662);
nor U4484 (N_4484,N_3651,N_3947);
and U4485 (N_4485,N_3760,N_3999);
nand U4486 (N_4486,N_3517,N_3926);
nor U4487 (N_4487,N_3564,N_3573);
or U4488 (N_4488,N_3662,N_3512);
xor U4489 (N_4489,N_3627,N_3806);
or U4490 (N_4490,N_3738,N_3504);
nor U4491 (N_4491,N_3576,N_3645);
nand U4492 (N_4492,N_3545,N_3598);
or U4493 (N_4493,N_3936,N_3562);
or U4494 (N_4494,N_3887,N_3828);
nor U4495 (N_4495,N_3677,N_3993);
nand U4496 (N_4496,N_3972,N_3505);
nand U4497 (N_4497,N_3607,N_3652);
and U4498 (N_4498,N_3995,N_3759);
or U4499 (N_4499,N_3962,N_3766);
nand U4500 (N_4500,N_4275,N_4453);
nor U4501 (N_4501,N_4331,N_4293);
xnor U4502 (N_4502,N_4068,N_4299);
xor U4503 (N_4503,N_4088,N_4037);
nand U4504 (N_4504,N_4337,N_4350);
xnor U4505 (N_4505,N_4481,N_4261);
nand U4506 (N_4506,N_4228,N_4124);
and U4507 (N_4507,N_4263,N_4060);
or U4508 (N_4508,N_4038,N_4149);
or U4509 (N_4509,N_4262,N_4449);
nand U4510 (N_4510,N_4399,N_4456);
nand U4511 (N_4511,N_4126,N_4433);
and U4512 (N_4512,N_4265,N_4097);
nor U4513 (N_4513,N_4345,N_4113);
nand U4514 (N_4514,N_4001,N_4008);
nand U4515 (N_4515,N_4317,N_4315);
and U4516 (N_4516,N_4328,N_4286);
or U4517 (N_4517,N_4282,N_4365);
and U4518 (N_4518,N_4170,N_4191);
xnor U4519 (N_4519,N_4464,N_4268);
or U4520 (N_4520,N_4138,N_4305);
or U4521 (N_4521,N_4306,N_4118);
nand U4522 (N_4522,N_4376,N_4098);
and U4523 (N_4523,N_4329,N_4128);
or U4524 (N_4524,N_4388,N_4135);
nand U4525 (N_4525,N_4493,N_4393);
nor U4526 (N_4526,N_4253,N_4358);
nand U4527 (N_4527,N_4221,N_4071);
nand U4528 (N_4528,N_4308,N_4499);
nand U4529 (N_4529,N_4448,N_4183);
or U4530 (N_4530,N_4014,N_4136);
nand U4531 (N_4531,N_4385,N_4454);
nand U4532 (N_4532,N_4168,N_4485);
xnor U4533 (N_4533,N_4112,N_4394);
nor U4534 (N_4534,N_4109,N_4470);
nor U4535 (N_4535,N_4383,N_4378);
and U4536 (N_4536,N_4058,N_4141);
nand U4537 (N_4537,N_4259,N_4336);
nand U4538 (N_4538,N_4437,N_4023);
nand U4539 (N_4539,N_4266,N_4412);
xor U4540 (N_4540,N_4207,N_4372);
nand U4541 (N_4541,N_4373,N_4167);
or U4542 (N_4542,N_4420,N_4443);
xnor U4543 (N_4543,N_4432,N_4404);
xor U4544 (N_4544,N_4173,N_4201);
nand U4545 (N_4545,N_4411,N_4226);
and U4546 (N_4546,N_4356,N_4123);
and U4547 (N_4547,N_4015,N_4447);
xor U4548 (N_4548,N_4450,N_4018);
nor U4549 (N_4549,N_4452,N_4127);
and U4550 (N_4550,N_4289,N_4083);
and U4551 (N_4551,N_4190,N_4327);
and U4552 (N_4552,N_4232,N_4090);
nand U4553 (N_4553,N_4162,N_4415);
and U4554 (N_4554,N_4197,N_4475);
nand U4555 (N_4555,N_4072,N_4219);
nor U4556 (N_4556,N_4033,N_4290);
xor U4557 (N_4557,N_4302,N_4175);
or U4558 (N_4558,N_4333,N_4359);
xor U4559 (N_4559,N_4177,N_4076);
nand U4560 (N_4560,N_4227,N_4387);
nand U4561 (N_4561,N_4321,N_4067);
nand U4562 (N_4562,N_4439,N_4081);
xnor U4563 (N_4563,N_4156,N_4044);
or U4564 (N_4564,N_4422,N_4478);
nor U4565 (N_4565,N_4442,N_4052);
nand U4566 (N_4566,N_4248,N_4476);
and U4567 (N_4567,N_4380,N_4445);
and U4568 (N_4568,N_4313,N_4419);
nand U4569 (N_4569,N_4487,N_4099);
xnor U4570 (N_4570,N_4210,N_4055);
or U4571 (N_4571,N_4473,N_4355);
and U4572 (N_4572,N_4320,N_4225);
nand U4573 (N_4573,N_4129,N_4349);
nor U4574 (N_4574,N_4322,N_4028);
nor U4575 (N_4575,N_4264,N_4494);
nand U4576 (N_4576,N_4012,N_4427);
xnor U4577 (N_4577,N_4272,N_4389);
nand U4578 (N_4578,N_4184,N_4298);
xnor U4579 (N_4579,N_4395,N_4063);
nor U4580 (N_4580,N_4276,N_4239);
and U4581 (N_4581,N_4495,N_4243);
and U4582 (N_4582,N_4054,N_4034);
and U4583 (N_4583,N_4451,N_4117);
or U4584 (N_4584,N_4270,N_4474);
or U4585 (N_4585,N_4338,N_4105);
xor U4586 (N_4586,N_4413,N_4229);
nand U4587 (N_4587,N_4017,N_4379);
or U4588 (N_4588,N_4429,N_4431);
xnor U4589 (N_4589,N_4403,N_4424);
or U4590 (N_4590,N_4150,N_4391);
and U4591 (N_4591,N_4472,N_4161);
xor U4592 (N_4592,N_4005,N_4425);
nand U4593 (N_4593,N_4347,N_4163);
nor U4594 (N_4594,N_4213,N_4301);
xnor U4595 (N_4595,N_4295,N_4222);
nor U4596 (N_4596,N_4371,N_4004);
or U4597 (N_4597,N_4486,N_4155);
nor U4598 (N_4598,N_4164,N_4457);
and U4599 (N_4599,N_4152,N_4077);
or U4600 (N_4600,N_4196,N_4455);
nor U4601 (N_4601,N_4362,N_4288);
xnor U4602 (N_4602,N_4115,N_4143);
nor U4603 (N_4603,N_4468,N_4323);
nor U4604 (N_4604,N_4461,N_4212);
and U4605 (N_4605,N_4217,N_4325);
nor U4606 (N_4606,N_4215,N_4179);
and U4607 (N_4607,N_4006,N_4198);
or U4608 (N_4608,N_4381,N_4285);
and U4609 (N_4609,N_4312,N_4384);
nand U4610 (N_4610,N_4087,N_4193);
nand U4611 (N_4611,N_4480,N_4459);
or U4612 (N_4612,N_4497,N_4339);
xnor U4613 (N_4613,N_4482,N_4353);
or U4614 (N_4614,N_4182,N_4280);
nor U4615 (N_4615,N_4319,N_4430);
or U4616 (N_4616,N_4334,N_4057);
and U4617 (N_4617,N_4107,N_4340);
xnor U4618 (N_4618,N_4114,N_4223);
and U4619 (N_4619,N_4477,N_4185);
xnor U4620 (N_4620,N_4418,N_4354);
nor U4621 (N_4621,N_4199,N_4296);
or U4622 (N_4622,N_4051,N_4428);
xor U4623 (N_4623,N_4142,N_4498);
or U4624 (N_4624,N_4157,N_4133);
nor U4625 (N_4625,N_4016,N_4463);
or U4626 (N_4626,N_4318,N_4056);
nor U4627 (N_4627,N_4026,N_4483);
xnor U4628 (N_4628,N_4096,N_4370);
or U4629 (N_4629,N_4174,N_4255);
and U4630 (N_4630,N_4279,N_4120);
nor U4631 (N_4631,N_4277,N_4409);
nand U4632 (N_4632,N_4211,N_4209);
nand U4633 (N_4633,N_4351,N_4400);
nor U4634 (N_4634,N_4416,N_4111);
or U4635 (N_4635,N_4310,N_4045);
and U4636 (N_4636,N_4307,N_4132);
nor U4637 (N_4637,N_4440,N_4086);
nor U4638 (N_4638,N_4267,N_4390);
or U4639 (N_4639,N_4119,N_4062);
or U4640 (N_4640,N_4042,N_4047);
nor U4641 (N_4641,N_4151,N_4160);
or U4642 (N_4642,N_4417,N_4241);
or U4643 (N_4643,N_4093,N_4031);
nand U4644 (N_4644,N_4147,N_4316);
nand U4645 (N_4645,N_4176,N_4407);
or U4646 (N_4646,N_4116,N_4467);
or U4647 (N_4647,N_4080,N_4234);
xnor U4648 (N_4648,N_4091,N_4311);
nand U4649 (N_4649,N_4094,N_4125);
nor U4650 (N_4650,N_4027,N_4029);
and U4651 (N_4651,N_4396,N_4484);
nand U4652 (N_4652,N_4144,N_4491);
nand U4653 (N_4653,N_4187,N_4224);
and U4654 (N_4654,N_4146,N_4220);
and U4655 (N_4655,N_4375,N_4025);
or U4656 (N_4656,N_4260,N_4466);
xnor U4657 (N_4657,N_4079,N_4330);
xnor U4658 (N_4658,N_4247,N_4292);
nor U4659 (N_4659,N_4022,N_4165);
or U4660 (N_4660,N_4332,N_4352);
nand U4661 (N_4661,N_4324,N_4172);
xnor U4662 (N_4662,N_4139,N_4314);
xnor U4663 (N_4663,N_4019,N_4050);
nor U4664 (N_4664,N_4496,N_4195);
xor U4665 (N_4665,N_4368,N_4131);
nand U4666 (N_4666,N_4078,N_4249);
or U4667 (N_4667,N_4471,N_4250);
or U4668 (N_4668,N_4344,N_4284);
xnor U4669 (N_4669,N_4148,N_4095);
xnor U4670 (N_4670,N_4252,N_4106);
or U4671 (N_4671,N_4009,N_4397);
and U4672 (N_4672,N_4122,N_4188);
or U4673 (N_4673,N_4341,N_4204);
or U4674 (N_4674,N_4434,N_4271);
and U4675 (N_4675,N_4377,N_4200);
nor U4676 (N_4676,N_4216,N_4066);
and U4677 (N_4677,N_4154,N_4238);
xnor U4678 (N_4678,N_4303,N_4102);
nand U4679 (N_4679,N_4065,N_4092);
nor U4680 (N_4680,N_4242,N_4049);
nor U4681 (N_4681,N_4040,N_4069);
and U4682 (N_4682,N_4140,N_4064);
and U4683 (N_4683,N_4010,N_4231);
or U4684 (N_4684,N_4030,N_4269);
or U4685 (N_4685,N_4089,N_4438);
xor U4686 (N_4686,N_4364,N_4405);
nand U4687 (N_4687,N_4061,N_4460);
nand U4688 (N_4688,N_4203,N_4110);
and U4689 (N_4689,N_4246,N_4257);
and U4690 (N_4690,N_4085,N_4205);
nand U4691 (N_4691,N_4348,N_4300);
xor U4692 (N_4692,N_4366,N_4367);
or U4693 (N_4693,N_4342,N_4178);
xnor U4694 (N_4694,N_4007,N_4240);
or U4695 (N_4695,N_4360,N_4297);
xor U4696 (N_4696,N_4043,N_4256);
and U4697 (N_4697,N_4281,N_4488);
nand U4698 (N_4698,N_4479,N_4011);
nand U4699 (N_4699,N_4075,N_4003);
and U4700 (N_4700,N_4166,N_4233);
nor U4701 (N_4701,N_4465,N_4032);
xor U4702 (N_4702,N_4024,N_4335);
or U4703 (N_4703,N_4103,N_4489);
nand U4704 (N_4704,N_4206,N_4082);
and U4705 (N_4705,N_4251,N_4421);
xnor U4706 (N_4706,N_4283,N_4053);
or U4707 (N_4707,N_4194,N_4244);
xnor U4708 (N_4708,N_4100,N_4258);
or U4709 (N_4709,N_4492,N_4369);
and U4710 (N_4710,N_4214,N_4073);
and U4711 (N_4711,N_4374,N_4153);
nor U4712 (N_4712,N_4361,N_4108);
nand U4713 (N_4713,N_4294,N_4408);
or U4714 (N_4714,N_4462,N_4230);
nand U4715 (N_4715,N_4181,N_4189);
nand U4716 (N_4716,N_4208,N_4423);
and U4717 (N_4717,N_4130,N_4134);
nor U4718 (N_4718,N_4039,N_4382);
and U4719 (N_4719,N_4402,N_4309);
nor U4720 (N_4720,N_4444,N_4346);
or U4721 (N_4721,N_4273,N_4158);
nand U4722 (N_4722,N_4104,N_4202);
xor U4723 (N_4723,N_4036,N_4070);
or U4724 (N_4724,N_4287,N_4159);
nor U4725 (N_4725,N_4013,N_4121);
xor U4726 (N_4726,N_4020,N_4235);
or U4727 (N_4727,N_4021,N_4469);
nand U4728 (N_4728,N_4357,N_4101);
and U4729 (N_4729,N_4046,N_4304);
nor U4730 (N_4730,N_4436,N_4410);
and U4731 (N_4731,N_4145,N_4278);
or U4732 (N_4732,N_4274,N_4169);
nor U4733 (N_4733,N_4035,N_4041);
nor U4734 (N_4734,N_4002,N_4435);
or U4735 (N_4735,N_4291,N_4084);
xor U4736 (N_4736,N_4245,N_4392);
nand U4737 (N_4737,N_4406,N_4398);
xor U4738 (N_4738,N_4137,N_4074);
xnor U4739 (N_4739,N_4363,N_4186);
and U4740 (N_4740,N_4000,N_4254);
xnor U4741 (N_4741,N_4386,N_4180);
nor U4742 (N_4742,N_4490,N_4441);
xnor U4743 (N_4743,N_4326,N_4236);
nor U4744 (N_4744,N_4171,N_4059);
xor U4745 (N_4745,N_4048,N_4237);
xor U4746 (N_4746,N_4458,N_4343);
or U4747 (N_4747,N_4446,N_4218);
nand U4748 (N_4748,N_4192,N_4414);
nor U4749 (N_4749,N_4401,N_4426);
xnor U4750 (N_4750,N_4115,N_4443);
xor U4751 (N_4751,N_4228,N_4353);
nor U4752 (N_4752,N_4260,N_4393);
nor U4753 (N_4753,N_4436,N_4121);
nor U4754 (N_4754,N_4319,N_4174);
xnor U4755 (N_4755,N_4316,N_4096);
or U4756 (N_4756,N_4011,N_4483);
and U4757 (N_4757,N_4245,N_4406);
xor U4758 (N_4758,N_4003,N_4139);
or U4759 (N_4759,N_4294,N_4239);
and U4760 (N_4760,N_4173,N_4039);
nand U4761 (N_4761,N_4141,N_4188);
and U4762 (N_4762,N_4101,N_4108);
and U4763 (N_4763,N_4154,N_4301);
nand U4764 (N_4764,N_4127,N_4165);
and U4765 (N_4765,N_4386,N_4254);
or U4766 (N_4766,N_4202,N_4195);
nand U4767 (N_4767,N_4106,N_4423);
and U4768 (N_4768,N_4392,N_4074);
and U4769 (N_4769,N_4368,N_4083);
nand U4770 (N_4770,N_4490,N_4095);
nor U4771 (N_4771,N_4426,N_4304);
or U4772 (N_4772,N_4048,N_4384);
and U4773 (N_4773,N_4343,N_4001);
nand U4774 (N_4774,N_4491,N_4225);
nor U4775 (N_4775,N_4340,N_4465);
or U4776 (N_4776,N_4412,N_4243);
nor U4777 (N_4777,N_4176,N_4413);
and U4778 (N_4778,N_4210,N_4383);
xnor U4779 (N_4779,N_4486,N_4313);
or U4780 (N_4780,N_4473,N_4429);
xor U4781 (N_4781,N_4294,N_4079);
nor U4782 (N_4782,N_4477,N_4261);
or U4783 (N_4783,N_4247,N_4044);
xor U4784 (N_4784,N_4231,N_4108);
xnor U4785 (N_4785,N_4211,N_4001);
nand U4786 (N_4786,N_4031,N_4066);
nand U4787 (N_4787,N_4188,N_4330);
or U4788 (N_4788,N_4232,N_4225);
nand U4789 (N_4789,N_4141,N_4447);
and U4790 (N_4790,N_4449,N_4494);
and U4791 (N_4791,N_4480,N_4347);
or U4792 (N_4792,N_4390,N_4453);
nor U4793 (N_4793,N_4263,N_4190);
nand U4794 (N_4794,N_4483,N_4194);
nand U4795 (N_4795,N_4140,N_4356);
and U4796 (N_4796,N_4051,N_4379);
or U4797 (N_4797,N_4128,N_4487);
nor U4798 (N_4798,N_4464,N_4389);
nor U4799 (N_4799,N_4333,N_4311);
and U4800 (N_4800,N_4410,N_4005);
xor U4801 (N_4801,N_4148,N_4311);
nand U4802 (N_4802,N_4319,N_4457);
xnor U4803 (N_4803,N_4134,N_4354);
nor U4804 (N_4804,N_4134,N_4294);
nor U4805 (N_4805,N_4116,N_4447);
and U4806 (N_4806,N_4080,N_4394);
nor U4807 (N_4807,N_4175,N_4405);
nor U4808 (N_4808,N_4020,N_4219);
xor U4809 (N_4809,N_4364,N_4177);
nand U4810 (N_4810,N_4216,N_4319);
and U4811 (N_4811,N_4237,N_4221);
nor U4812 (N_4812,N_4164,N_4393);
nor U4813 (N_4813,N_4413,N_4262);
or U4814 (N_4814,N_4308,N_4060);
xnor U4815 (N_4815,N_4110,N_4271);
or U4816 (N_4816,N_4212,N_4136);
or U4817 (N_4817,N_4469,N_4037);
nand U4818 (N_4818,N_4442,N_4430);
and U4819 (N_4819,N_4377,N_4314);
nand U4820 (N_4820,N_4101,N_4295);
and U4821 (N_4821,N_4105,N_4154);
or U4822 (N_4822,N_4413,N_4044);
xor U4823 (N_4823,N_4171,N_4316);
nand U4824 (N_4824,N_4275,N_4049);
nand U4825 (N_4825,N_4220,N_4193);
or U4826 (N_4826,N_4360,N_4356);
xnor U4827 (N_4827,N_4286,N_4240);
and U4828 (N_4828,N_4313,N_4073);
nand U4829 (N_4829,N_4196,N_4134);
nand U4830 (N_4830,N_4365,N_4091);
and U4831 (N_4831,N_4002,N_4497);
and U4832 (N_4832,N_4386,N_4027);
and U4833 (N_4833,N_4210,N_4381);
nor U4834 (N_4834,N_4076,N_4469);
nand U4835 (N_4835,N_4253,N_4366);
nor U4836 (N_4836,N_4321,N_4045);
nand U4837 (N_4837,N_4072,N_4154);
or U4838 (N_4838,N_4179,N_4092);
and U4839 (N_4839,N_4236,N_4130);
and U4840 (N_4840,N_4499,N_4429);
and U4841 (N_4841,N_4499,N_4419);
or U4842 (N_4842,N_4398,N_4338);
and U4843 (N_4843,N_4177,N_4320);
nand U4844 (N_4844,N_4058,N_4443);
xor U4845 (N_4845,N_4130,N_4259);
nand U4846 (N_4846,N_4257,N_4351);
nor U4847 (N_4847,N_4234,N_4398);
nor U4848 (N_4848,N_4379,N_4006);
and U4849 (N_4849,N_4413,N_4199);
or U4850 (N_4850,N_4399,N_4271);
nor U4851 (N_4851,N_4047,N_4378);
or U4852 (N_4852,N_4374,N_4019);
xor U4853 (N_4853,N_4268,N_4468);
and U4854 (N_4854,N_4284,N_4443);
and U4855 (N_4855,N_4484,N_4467);
nand U4856 (N_4856,N_4311,N_4220);
nand U4857 (N_4857,N_4153,N_4343);
nand U4858 (N_4858,N_4228,N_4024);
xnor U4859 (N_4859,N_4390,N_4221);
nor U4860 (N_4860,N_4192,N_4363);
or U4861 (N_4861,N_4027,N_4423);
or U4862 (N_4862,N_4029,N_4049);
xnor U4863 (N_4863,N_4040,N_4452);
or U4864 (N_4864,N_4385,N_4432);
nand U4865 (N_4865,N_4133,N_4493);
or U4866 (N_4866,N_4447,N_4024);
or U4867 (N_4867,N_4216,N_4444);
and U4868 (N_4868,N_4325,N_4379);
nand U4869 (N_4869,N_4383,N_4215);
nor U4870 (N_4870,N_4470,N_4008);
and U4871 (N_4871,N_4223,N_4428);
nand U4872 (N_4872,N_4052,N_4425);
or U4873 (N_4873,N_4432,N_4071);
nor U4874 (N_4874,N_4498,N_4140);
or U4875 (N_4875,N_4498,N_4460);
xor U4876 (N_4876,N_4248,N_4219);
nand U4877 (N_4877,N_4369,N_4402);
or U4878 (N_4878,N_4233,N_4244);
xor U4879 (N_4879,N_4209,N_4451);
nand U4880 (N_4880,N_4484,N_4247);
xnor U4881 (N_4881,N_4246,N_4082);
nand U4882 (N_4882,N_4171,N_4195);
nor U4883 (N_4883,N_4261,N_4341);
or U4884 (N_4884,N_4395,N_4456);
xor U4885 (N_4885,N_4182,N_4225);
or U4886 (N_4886,N_4459,N_4136);
and U4887 (N_4887,N_4193,N_4381);
or U4888 (N_4888,N_4064,N_4455);
or U4889 (N_4889,N_4246,N_4210);
xnor U4890 (N_4890,N_4133,N_4411);
or U4891 (N_4891,N_4069,N_4343);
xnor U4892 (N_4892,N_4351,N_4206);
nor U4893 (N_4893,N_4270,N_4194);
and U4894 (N_4894,N_4278,N_4077);
nor U4895 (N_4895,N_4184,N_4061);
xnor U4896 (N_4896,N_4065,N_4362);
nor U4897 (N_4897,N_4178,N_4121);
nand U4898 (N_4898,N_4357,N_4064);
nand U4899 (N_4899,N_4070,N_4389);
xnor U4900 (N_4900,N_4128,N_4042);
and U4901 (N_4901,N_4411,N_4020);
nor U4902 (N_4902,N_4347,N_4321);
or U4903 (N_4903,N_4303,N_4402);
or U4904 (N_4904,N_4091,N_4150);
nand U4905 (N_4905,N_4202,N_4055);
and U4906 (N_4906,N_4364,N_4483);
nor U4907 (N_4907,N_4408,N_4000);
or U4908 (N_4908,N_4418,N_4151);
and U4909 (N_4909,N_4384,N_4058);
nor U4910 (N_4910,N_4280,N_4187);
nand U4911 (N_4911,N_4228,N_4113);
or U4912 (N_4912,N_4347,N_4406);
nand U4913 (N_4913,N_4285,N_4460);
xnor U4914 (N_4914,N_4276,N_4367);
nand U4915 (N_4915,N_4326,N_4183);
or U4916 (N_4916,N_4374,N_4388);
and U4917 (N_4917,N_4187,N_4441);
nand U4918 (N_4918,N_4271,N_4338);
nand U4919 (N_4919,N_4030,N_4165);
nand U4920 (N_4920,N_4221,N_4172);
or U4921 (N_4921,N_4261,N_4253);
xnor U4922 (N_4922,N_4487,N_4138);
nand U4923 (N_4923,N_4457,N_4259);
nor U4924 (N_4924,N_4179,N_4195);
nor U4925 (N_4925,N_4307,N_4486);
xnor U4926 (N_4926,N_4497,N_4120);
nand U4927 (N_4927,N_4213,N_4110);
and U4928 (N_4928,N_4210,N_4245);
and U4929 (N_4929,N_4432,N_4214);
xor U4930 (N_4930,N_4340,N_4304);
and U4931 (N_4931,N_4075,N_4044);
nor U4932 (N_4932,N_4080,N_4067);
xor U4933 (N_4933,N_4497,N_4082);
and U4934 (N_4934,N_4495,N_4071);
nand U4935 (N_4935,N_4441,N_4437);
nor U4936 (N_4936,N_4384,N_4314);
nand U4937 (N_4937,N_4423,N_4300);
nand U4938 (N_4938,N_4100,N_4039);
nand U4939 (N_4939,N_4156,N_4098);
or U4940 (N_4940,N_4369,N_4496);
nor U4941 (N_4941,N_4307,N_4204);
nand U4942 (N_4942,N_4302,N_4278);
xor U4943 (N_4943,N_4097,N_4430);
nor U4944 (N_4944,N_4239,N_4347);
and U4945 (N_4945,N_4319,N_4193);
or U4946 (N_4946,N_4243,N_4444);
nand U4947 (N_4947,N_4419,N_4126);
xor U4948 (N_4948,N_4099,N_4307);
nor U4949 (N_4949,N_4381,N_4331);
xnor U4950 (N_4950,N_4020,N_4327);
nor U4951 (N_4951,N_4106,N_4094);
nand U4952 (N_4952,N_4393,N_4444);
or U4953 (N_4953,N_4477,N_4058);
or U4954 (N_4954,N_4080,N_4165);
or U4955 (N_4955,N_4157,N_4460);
or U4956 (N_4956,N_4258,N_4445);
and U4957 (N_4957,N_4403,N_4494);
xor U4958 (N_4958,N_4228,N_4217);
and U4959 (N_4959,N_4475,N_4233);
nor U4960 (N_4960,N_4230,N_4263);
xor U4961 (N_4961,N_4444,N_4423);
or U4962 (N_4962,N_4048,N_4087);
nand U4963 (N_4963,N_4276,N_4238);
or U4964 (N_4964,N_4316,N_4342);
nor U4965 (N_4965,N_4301,N_4060);
and U4966 (N_4966,N_4135,N_4474);
and U4967 (N_4967,N_4108,N_4391);
nor U4968 (N_4968,N_4378,N_4063);
nand U4969 (N_4969,N_4396,N_4115);
xor U4970 (N_4970,N_4181,N_4362);
and U4971 (N_4971,N_4288,N_4129);
and U4972 (N_4972,N_4427,N_4486);
nor U4973 (N_4973,N_4288,N_4297);
and U4974 (N_4974,N_4043,N_4006);
nand U4975 (N_4975,N_4411,N_4074);
nor U4976 (N_4976,N_4411,N_4044);
nand U4977 (N_4977,N_4161,N_4405);
and U4978 (N_4978,N_4473,N_4340);
nor U4979 (N_4979,N_4268,N_4344);
and U4980 (N_4980,N_4197,N_4210);
xor U4981 (N_4981,N_4191,N_4346);
or U4982 (N_4982,N_4128,N_4318);
and U4983 (N_4983,N_4086,N_4310);
or U4984 (N_4984,N_4186,N_4102);
or U4985 (N_4985,N_4395,N_4094);
xor U4986 (N_4986,N_4018,N_4179);
xor U4987 (N_4987,N_4055,N_4325);
nand U4988 (N_4988,N_4319,N_4370);
xor U4989 (N_4989,N_4434,N_4353);
nor U4990 (N_4990,N_4460,N_4310);
nor U4991 (N_4991,N_4304,N_4176);
nand U4992 (N_4992,N_4184,N_4407);
xor U4993 (N_4993,N_4407,N_4403);
nor U4994 (N_4994,N_4404,N_4241);
xnor U4995 (N_4995,N_4189,N_4163);
or U4996 (N_4996,N_4225,N_4423);
xnor U4997 (N_4997,N_4372,N_4125);
xnor U4998 (N_4998,N_4434,N_4232);
nor U4999 (N_4999,N_4155,N_4477);
or U5000 (N_5000,N_4566,N_4617);
nor U5001 (N_5001,N_4679,N_4711);
and U5002 (N_5002,N_4789,N_4696);
xnor U5003 (N_5003,N_4864,N_4845);
and U5004 (N_5004,N_4992,N_4808);
or U5005 (N_5005,N_4543,N_4717);
nor U5006 (N_5006,N_4535,N_4561);
or U5007 (N_5007,N_4893,N_4903);
or U5008 (N_5008,N_4769,N_4874);
nand U5009 (N_5009,N_4965,N_4879);
and U5010 (N_5010,N_4590,N_4862);
nand U5011 (N_5011,N_4866,N_4658);
nand U5012 (N_5012,N_4757,N_4923);
xor U5013 (N_5013,N_4783,N_4790);
xnor U5014 (N_5014,N_4603,N_4883);
and U5015 (N_5015,N_4718,N_4576);
nor U5016 (N_5016,N_4506,N_4601);
nand U5017 (N_5017,N_4564,N_4650);
or U5018 (N_5018,N_4557,N_4641);
nand U5019 (N_5019,N_4987,N_4526);
nor U5020 (N_5020,N_4985,N_4675);
and U5021 (N_5021,N_4512,N_4528);
nand U5022 (N_5022,N_4639,N_4976);
xor U5023 (N_5023,N_4645,N_4916);
and U5024 (N_5024,N_4915,N_4761);
nor U5025 (N_5025,N_4887,N_4755);
xor U5026 (N_5026,N_4742,N_4597);
nor U5027 (N_5027,N_4867,N_4969);
and U5028 (N_5028,N_4981,N_4787);
and U5029 (N_5029,N_4998,N_4710);
and U5030 (N_5030,N_4766,N_4937);
or U5031 (N_5031,N_4542,N_4517);
nand U5032 (N_5032,N_4765,N_4530);
xor U5033 (N_5033,N_4740,N_4665);
nor U5034 (N_5034,N_4609,N_4667);
nand U5035 (N_5035,N_4607,N_4505);
nor U5036 (N_5036,N_4792,N_4890);
and U5037 (N_5037,N_4759,N_4818);
nand U5038 (N_5038,N_4620,N_4660);
and U5039 (N_5039,N_4515,N_4882);
and U5040 (N_5040,N_4863,N_4572);
nand U5041 (N_5041,N_4956,N_4853);
and U5042 (N_5042,N_4736,N_4584);
or U5043 (N_5043,N_4606,N_4955);
or U5044 (N_5044,N_4995,N_4944);
and U5045 (N_5045,N_4756,N_4546);
xor U5046 (N_5046,N_4527,N_4712);
xnor U5047 (N_5047,N_4720,N_4832);
or U5048 (N_5048,N_4647,N_4691);
or U5049 (N_5049,N_4860,N_4669);
xor U5050 (N_5050,N_4913,N_4846);
xor U5051 (N_5051,N_4516,N_4685);
nand U5052 (N_5052,N_4681,N_4537);
nand U5053 (N_5053,N_4621,N_4966);
or U5054 (N_5054,N_4994,N_4906);
xnor U5055 (N_5055,N_4582,N_4744);
xnor U5056 (N_5056,N_4773,N_4522);
or U5057 (N_5057,N_4697,N_4855);
nand U5058 (N_5058,N_4507,N_4677);
nor U5059 (N_5059,N_4967,N_4805);
nor U5060 (N_5060,N_4531,N_4539);
and U5061 (N_5061,N_4676,N_4555);
nor U5062 (N_5062,N_4749,N_4559);
nand U5063 (N_5063,N_4803,N_4794);
and U5064 (N_5064,N_4727,N_4917);
or U5065 (N_5065,N_4936,N_4648);
xnor U5066 (N_5066,N_4703,N_4578);
and U5067 (N_5067,N_4837,N_4904);
or U5068 (N_5068,N_4826,N_4802);
and U5069 (N_5069,N_4975,N_4991);
xor U5070 (N_5070,N_4571,N_4778);
or U5071 (N_5071,N_4637,N_4532);
and U5072 (N_5072,N_4586,N_4960);
or U5073 (N_5073,N_4624,N_4980);
xor U5074 (N_5074,N_4941,N_4735);
and U5075 (N_5075,N_4630,N_4569);
xnor U5076 (N_5076,N_4666,N_4694);
nor U5077 (N_5077,N_4693,N_4961);
or U5078 (N_5078,N_4947,N_4661);
xnor U5079 (N_5079,N_4841,N_4653);
xnor U5080 (N_5080,N_4610,N_4689);
nor U5081 (N_5081,N_4682,N_4804);
or U5082 (N_5082,N_4593,N_4678);
or U5083 (N_5083,N_4743,N_4951);
nand U5084 (N_5084,N_4894,N_4733);
nor U5085 (N_5085,N_4737,N_4554);
and U5086 (N_5086,N_4798,N_4950);
nor U5087 (N_5087,N_4556,N_4716);
xor U5088 (N_5088,N_4702,N_4823);
and U5089 (N_5089,N_4908,N_4668);
nand U5090 (N_5090,N_4806,N_4519);
or U5091 (N_5091,N_4780,N_4785);
and U5092 (N_5092,N_4560,N_4786);
or U5093 (N_5093,N_4581,N_4671);
nor U5094 (N_5094,N_4589,N_4840);
xnor U5095 (N_5095,N_4723,N_4945);
and U5096 (N_5096,N_4988,N_4738);
and U5097 (N_5097,N_4629,N_4767);
nand U5098 (N_5098,N_4705,N_4799);
and U5099 (N_5099,N_4807,N_4549);
nand U5100 (N_5100,N_4508,N_4633);
xor U5101 (N_5101,N_4814,N_4538);
and U5102 (N_5102,N_4847,N_4898);
or U5103 (N_5103,N_4844,N_4541);
or U5104 (N_5104,N_4587,N_4871);
nor U5105 (N_5105,N_4970,N_4760);
nor U5106 (N_5106,N_4605,N_4642);
xnor U5107 (N_5107,N_4984,N_4521);
or U5108 (N_5108,N_4745,N_4927);
or U5109 (N_5109,N_4509,N_4873);
nand U5110 (N_5110,N_4649,N_4911);
or U5111 (N_5111,N_4553,N_4878);
and U5112 (N_5112,N_4880,N_4858);
or U5113 (N_5113,N_4910,N_4895);
nand U5114 (N_5114,N_4623,N_4851);
nor U5115 (N_5115,N_4654,N_4524);
and U5116 (N_5116,N_4848,N_4585);
xnor U5117 (N_5117,N_4713,N_4729);
and U5118 (N_5118,N_4815,N_4771);
or U5119 (N_5119,N_4817,N_4791);
and U5120 (N_5120,N_4615,N_4510);
and U5121 (N_5121,N_4536,N_4636);
xor U5122 (N_5122,N_4869,N_4575);
or U5123 (N_5123,N_4626,N_4739);
or U5124 (N_5124,N_4776,N_4954);
nand U5125 (N_5125,N_4835,N_4881);
and U5126 (N_5126,N_4672,N_4953);
xnor U5127 (N_5127,N_4925,N_4670);
xor U5128 (N_5128,N_4540,N_4920);
and U5129 (N_5129,N_4747,N_4750);
xnor U5130 (N_5130,N_4831,N_4709);
xor U5131 (N_5131,N_4959,N_4978);
or U5132 (N_5132,N_4859,N_4940);
nor U5133 (N_5133,N_4812,N_4690);
xor U5134 (N_5134,N_4754,N_4914);
nand U5135 (N_5135,N_4828,N_4868);
nand U5136 (N_5136,N_4502,N_4811);
nor U5137 (N_5137,N_4876,N_4656);
nand U5138 (N_5138,N_4958,N_4591);
nand U5139 (N_5139,N_4550,N_4779);
nor U5140 (N_5140,N_4640,N_4608);
nand U5141 (N_5141,N_4973,N_4875);
xnor U5142 (N_5142,N_4632,N_4905);
xnor U5143 (N_5143,N_4619,N_4938);
nand U5144 (N_5144,N_4926,N_4957);
xor U5145 (N_5145,N_4731,N_4545);
xnor U5146 (N_5146,N_4918,N_4664);
xnor U5147 (N_5147,N_4644,N_4652);
and U5148 (N_5148,N_4824,N_4999);
or U5149 (N_5149,N_4795,N_4662);
and U5150 (N_5150,N_4796,N_4594);
nand U5151 (N_5151,N_4612,N_4722);
nor U5152 (N_5152,N_4663,N_4673);
nand U5153 (N_5153,N_4686,N_4870);
nor U5154 (N_5154,N_4513,N_4809);
xnor U5155 (N_5155,N_4793,N_4854);
xnor U5156 (N_5156,N_4892,N_4884);
or U5157 (N_5157,N_4565,N_4627);
nor U5158 (N_5158,N_4930,N_4674);
nand U5159 (N_5159,N_4820,N_4701);
or U5160 (N_5160,N_4503,N_4708);
nand U5161 (N_5161,N_4500,N_4752);
xnor U5162 (N_5162,N_4788,N_4889);
and U5163 (N_5163,N_4872,N_4628);
nand U5164 (N_5164,N_4625,N_4520);
xnor U5165 (N_5165,N_4996,N_4816);
xnor U5166 (N_5166,N_4849,N_4562);
xnor U5167 (N_5167,N_4935,N_4891);
xnor U5168 (N_5168,N_4852,N_4643);
and U5169 (N_5169,N_4730,N_4775);
nor U5170 (N_5170,N_4877,N_4638);
and U5171 (N_5171,N_4774,N_4827);
xnor U5172 (N_5172,N_4688,N_4635);
and U5173 (N_5173,N_4772,N_4968);
xor U5174 (N_5174,N_4762,N_4583);
nor U5175 (N_5175,N_4912,N_4631);
nand U5176 (N_5176,N_4983,N_4657);
nand U5177 (N_5177,N_4568,N_4746);
nand U5178 (N_5178,N_4551,N_4948);
or U5179 (N_5179,N_4886,N_4721);
nand U5180 (N_5180,N_4700,N_4782);
nand U5181 (N_5181,N_4659,N_4932);
xnor U5182 (N_5182,N_4800,N_4924);
nand U5183 (N_5183,N_4901,N_4714);
and U5184 (N_5184,N_4829,N_4896);
or U5185 (N_5185,N_4986,N_4579);
nand U5186 (N_5186,N_4602,N_4810);
and U5187 (N_5187,N_4850,N_4834);
nor U5188 (N_5188,N_4725,N_4616);
nor U5189 (N_5189,N_4753,N_4900);
nor U5190 (N_5190,N_4595,N_4573);
nor U5191 (N_5191,N_4529,N_4687);
and U5192 (N_5192,N_4533,N_4833);
xnor U5193 (N_5193,N_4952,N_4504);
or U5194 (N_5194,N_4843,N_4614);
nor U5195 (N_5195,N_4784,N_4839);
or U5196 (N_5196,N_4801,N_4706);
xor U5197 (N_5197,N_4990,N_4797);
nand U5198 (N_5198,N_4919,N_4715);
xnor U5199 (N_5199,N_4604,N_4857);
nor U5200 (N_5200,N_4993,N_4768);
nand U5201 (N_5201,N_4558,N_4523);
and U5202 (N_5202,N_4764,N_4949);
nor U5203 (N_5203,N_4865,N_4751);
or U5204 (N_5204,N_4634,N_4683);
nor U5205 (N_5205,N_4518,N_4726);
and U5206 (N_5206,N_4974,N_4741);
and U5207 (N_5207,N_4698,N_4728);
or U5208 (N_5208,N_4813,N_4548);
xnor U5209 (N_5209,N_4724,N_4838);
xor U5210 (N_5210,N_4963,N_4971);
and U5211 (N_5211,N_4707,N_4611);
nand U5212 (N_5212,N_4931,N_4622);
nor U5213 (N_5213,N_4934,N_4692);
and U5214 (N_5214,N_4680,N_4939);
xor U5215 (N_5215,N_4942,N_4684);
xor U5216 (N_5216,N_4972,N_4929);
nor U5217 (N_5217,N_4836,N_4655);
or U5218 (N_5218,N_4501,N_4699);
nor U5219 (N_5219,N_4618,N_4598);
nor U5220 (N_5220,N_4781,N_4646);
nand U5221 (N_5221,N_4748,N_4830);
and U5222 (N_5222,N_4819,N_4909);
and U5223 (N_5223,N_4822,N_4982);
nor U5224 (N_5224,N_4962,N_4577);
and U5225 (N_5225,N_4651,N_4599);
nor U5226 (N_5226,N_4928,N_4964);
xor U5227 (N_5227,N_4885,N_4600);
nand U5228 (N_5228,N_4592,N_4534);
and U5229 (N_5229,N_4899,N_4770);
nand U5230 (N_5230,N_4588,N_4946);
and U5231 (N_5231,N_4902,N_4704);
and U5232 (N_5232,N_4719,N_4547);
nor U5233 (N_5233,N_4821,N_4574);
xor U5234 (N_5234,N_4544,N_4570);
or U5235 (N_5235,N_4856,N_4888);
xor U5236 (N_5236,N_4732,N_4580);
nor U5237 (N_5237,N_4933,N_4511);
nand U5238 (N_5238,N_4695,N_4563);
or U5239 (N_5239,N_4596,N_4734);
nand U5240 (N_5240,N_4763,N_4567);
nor U5241 (N_5241,N_4907,N_4921);
or U5242 (N_5242,N_4989,N_4552);
or U5243 (N_5243,N_4979,N_4525);
nor U5244 (N_5244,N_4825,N_4613);
nand U5245 (N_5245,N_4943,N_4922);
xor U5246 (N_5246,N_4861,N_4897);
nor U5247 (N_5247,N_4758,N_4997);
nor U5248 (N_5248,N_4842,N_4514);
xnor U5249 (N_5249,N_4977,N_4777);
or U5250 (N_5250,N_4702,N_4572);
nor U5251 (N_5251,N_4723,N_4592);
and U5252 (N_5252,N_4994,N_4817);
or U5253 (N_5253,N_4835,N_4721);
or U5254 (N_5254,N_4600,N_4976);
xor U5255 (N_5255,N_4603,N_4668);
or U5256 (N_5256,N_4530,N_4583);
nor U5257 (N_5257,N_4672,N_4807);
xor U5258 (N_5258,N_4975,N_4532);
xor U5259 (N_5259,N_4509,N_4850);
or U5260 (N_5260,N_4738,N_4756);
or U5261 (N_5261,N_4779,N_4621);
or U5262 (N_5262,N_4645,N_4723);
or U5263 (N_5263,N_4870,N_4967);
or U5264 (N_5264,N_4835,N_4600);
or U5265 (N_5265,N_4690,N_4862);
or U5266 (N_5266,N_4618,N_4749);
nor U5267 (N_5267,N_4856,N_4568);
or U5268 (N_5268,N_4954,N_4877);
nor U5269 (N_5269,N_4577,N_4739);
or U5270 (N_5270,N_4701,N_4669);
or U5271 (N_5271,N_4787,N_4824);
nor U5272 (N_5272,N_4579,N_4984);
nand U5273 (N_5273,N_4673,N_4579);
nand U5274 (N_5274,N_4562,N_4636);
and U5275 (N_5275,N_4771,N_4575);
and U5276 (N_5276,N_4753,N_4698);
and U5277 (N_5277,N_4998,N_4538);
nand U5278 (N_5278,N_4810,N_4752);
and U5279 (N_5279,N_4636,N_4996);
nor U5280 (N_5280,N_4808,N_4776);
xor U5281 (N_5281,N_4836,N_4961);
and U5282 (N_5282,N_4932,N_4577);
xnor U5283 (N_5283,N_4683,N_4509);
and U5284 (N_5284,N_4548,N_4509);
or U5285 (N_5285,N_4570,N_4897);
nand U5286 (N_5286,N_4870,N_4685);
nor U5287 (N_5287,N_4626,N_4558);
and U5288 (N_5288,N_4549,N_4754);
nand U5289 (N_5289,N_4578,N_4783);
nand U5290 (N_5290,N_4924,N_4703);
nor U5291 (N_5291,N_4659,N_4595);
nor U5292 (N_5292,N_4597,N_4664);
and U5293 (N_5293,N_4987,N_4742);
nand U5294 (N_5294,N_4790,N_4505);
and U5295 (N_5295,N_4857,N_4990);
nand U5296 (N_5296,N_4588,N_4997);
xor U5297 (N_5297,N_4585,N_4831);
xor U5298 (N_5298,N_4570,N_4817);
nor U5299 (N_5299,N_4572,N_4583);
and U5300 (N_5300,N_4622,N_4913);
and U5301 (N_5301,N_4739,N_4865);
xor U5302 (N_5302,N_4588,N_4751);
xnor U5303 (N_5303,N_4772,N_4934);
or U5304 (N_5304,N_4561,N_4750);
nor U5305 (N_5305,N_4951,N_4642);
nor U5306 (N_5306,N_4965,N_4872);
or U5307 (N_5307,N_4617,N_4993);
nand U5308 (N_5308,N_4536,N_4970);
nand U5309 (N_5309,N_4544,N_4902);
or U5310 (N_5310,N_4831,N_4562);
and U5311 (N_5311,N_4604,N_4541);
nor U5312 (N_5312,N_4670,N_4603);
nor U5313 (N_5313,N_4691,N_4597);
nor U5314 (N_5314,N_4580,N_4941);
nand U5315 (N_5315,N_4898,N_4842);
nand U5316 (N_5316,N_4965,N_4816);
nor U5317 (N_5317,N_4575,N_4824);
and U5318 (N_5318,N_4983,N_4866);
xnor U5319 (N_5319,N_4965,N_4746);
xnor U5320 (N_5320,N_4736,N_4530);
or U5321 (N_5321,N_4532,N_4586);
nand U5322 (N_5322,N_4709,N_4793);
xnor U5323 (N_5323,N_4581,N_4707);
xnor U5324 (N_5324,N_4897,N_4628);
nand U5325 (N_5325,N_4515,N_4834);
nand U5326 (N_5326,N_4676,N_4873);
nand U5327 (N_5327,N_4997,N_4698);
nor U5328 (N_5328,N_4856,N_4757);
or U5329 (N_5329,N_4993,N_4573);
xnor U5330 (N_5330,N_4613,N_4923);
and U5331 (N_5331,N_4656,N_4650);
nor U5332 (N_5332,N_4772,N_4886);
xor U5333 (N_5333,N_4775,N_4892);
xnor U5334 (N_5334,N_4686,N_4674);
and U5335 (N_5335,N_4692,N_4674);
nor U5336 (N_5336,N_4764,N_4532);
nor U5337 (N_5337,N_4988,N_4800);
nand U5338 (N_5338,N_4790,N_4778);
nand U5339 (N_5339,N_4856,N_4734);
or U5340 (N_5340,N_4811,N_4534);
nor U5341 (N_5341,N_4965,N_4947);
nor U5342 (N_5342,N_4579,N_4603);
or U5343 (N_5343,N_4635,N_4734);
nand U5344 (N_5344,N_4950,N_4901);
or U5345 (N_5345,N_4638,N_4799);
xor U5346 (N_5346,N_4639,N_4732);
or U5347 (N_5347,N_4865,N_4958);
nand U5348 (N_5348,N_4859,N_4794);
nand U5349 (N_5349,N_4989,N_4520);
or U5350 (N_5350,N_4851,N_4893);
nor U5351 (N_5351,N_4541,N_4623);
xor U5352 (N_5352,N_4796,N_4819);
nor U5353 (N_5353,N_4801,N_4639);
xor U5354 (N_5354,N_4700,N_4734);
and U5355 (N_5355,N_4506,N_4697);
xnor U5356 (N_5356,N_4898,N_4669);
nand U5357 (N_5357,N_4594,N_4693);
xnor U5358 (N_5358,N_4617,N_4768);
or U5359 (N_5359,N_4920,N_4702);
nor U5360 (N_5360,N_4777,N_4513);
nor U5361 (N_5361,N_4844,N_4907);
or U5362 (N_5362,N_4699,N_4832);
and U5363 (N_5363,N_4500,N_4994);
and U5364 (N_5364,N_4618,N_4608);
nor U5365 (N_5365,N_4849,N_4628);
or U5366 (N_5366,N_4691,N_4888);
nand U5367 (N_5367,N_4527,N_4874);
xnor U5368 (N_5368,N_4854,N_4564);
nand U5369 (N_5369,N_4998,N_4907);
xnor U5370 (N_5370,N_4644,N_4955);
and U5371 (N_5371,N_4555,N_4631);
nand U5372 (N_5372,N_4673,N_4585);
nand U5373 (N_5373,N_4982,N_4995);
and U5374 (N_5374,N_4753,N_4565);
nand U5375 (N_5375,N_4805,N_4524);
nand U5376 (N_5376,N_4978,N_4560);
or U5377 (N_5377,N_4917,N_4517);
xnor U5378 (N_5378,N_4748,N_4755);
nor U5379 (N_5379,N_4772,N_4741);
xnor U5380 (N_5380,N_4697,N_4717);
and U5381 (N_5381,N_4779,N_4647);
and U5382 (N_5382,N_4810,N_4623);
and U5383 (N_5383,N_4816,N_4999);
nor U5384 (N_5384,N_4975,N_4994);
nand U5385 (N_5385,N_4705,N_4663);
and U5386 (N_5386,N_4622,N_4783);
and U5387 (N_5387,N_4535,N_4747);
or U5388 (N_5388,N_4721,N_4744);
and U5389 (N_5389,N_4993,N_4968);
and U5390 (N_5390,N_4793,N_4827);
xnor U5391 (N_5391,N_4626,N_4754);
xor U5392 (N_5392,N_4948,N_4777);
and U5393 (N_5393,N_4579,N_4599);
and U5394 (N_5394,N_4556,N_4696);
nand U5395 (N_5395,N_4741,N_4553);
or U5396 (N_5396,N_4709,N_4547);
nor U5397 (N_5397,N_4932,N_4554);
xor U5398 (N_5398,N_4504,N_4827);
and U5399 (N_5399,N_4584,N_4999);
and U5400 (N_5400,N_4626,N_4764);
and U5401 (N_5401,N_4748,N_4730);
and U5402 (N_5402,N_4665,N_4710);
or U5403 (N_5403,N_4830,N_4553);
nor U5404 (N_5404,N_4586,N_4542);
nand U5405 (N_5405,N_4884,N_4606);
or U5406 (N_5406,N_4555,N_4603);
nand U5407 (N_5407,N_4602,N_4717);
nor U5408 (N_5408,N_4532,N_4548);
xnor U5409 (N_5409,N_4661,N_4951);
or U5410 (N_5410,N_4812,N_4935);
and U5411 (N_5411,N_4720,N_4742);
nand U5412 (N_5412,N_4934,N_4529);
and U5413 (N_5413,N_4716,N_4561);
nor U5414 (N_5414,N_4540,N_4843);
nand U5415 (N_5415,N_4908,N_4640);
xnor U5416 (N_5416,N_4595,N_4710);
and U5417 (N_5417,N_4809,N_4654);
nand U5418 (N_5418,N_4554,N_4866);
and U5419 (N_5419,N_4804,N_4903);
or U5420 (N_5420,N_4771,N_4854);
and U5421 (N_5421,N_4777,N_4786);
xor U5422 (N_5422,N_4810,N_4946);
or U5423 (N_5423,N_4714,N_4947);
or U5424 (N_5424,N_4915,N_4844);
nand U5425 (N_5425,N_4574,N_4665);
and U5426 (N_5426,N_4779,N_4834);
xor U5427 (N_5427,N_4848,N_4689);
or U5428 (N_5428,N_4886,N_4972);
nor U5429 (N_5429,N_4905,N_4643);
xor U5430 (N_5430,N_4849,N_4954);
xnor U5431 (N_5431,N_4893,N_4593);
nand U5432 (N_5432,N_4647,N_4523);
nor U5433 (N_5433,N_4963,N_4547);
nand U5434 (N_5434,N_4689,N_4681);
or U5435 (N_5435,N_4783,N_4949);
xnor U5436 (N_5436,N_4657,N_4940);
xor U5437 (N_5437,N_4613,N_4704);
xor U5438 (N_5438,N_4996,N_4707);
xor U5439 (N_5439,N_4928,N_4929);
nor U5440 (N_5440,N_4872,N_4956);
nand U5441 (N_5441,N_4584,N_4793);
nor U5442 (N_5442,N_4877,N_4650);
nor U5443 (N_5443,N_4975,N_4850);
and U5444 (N_5444,N_4930,N_4722);
nand U5445 (N_5445,N_4908,N_4957);
or U5446 (N_5446,N_4678,N_4643);
and U5447 (N_5447,N_4865,N_4660);
nand U5448 (N_5448,N_4773,N_4897);
and U5449 (N_5449,N_4529,N_4856);
xor U5450 (N_5450,N_4556,N_4515);
nand U5451 (N_5451,N_4968,N_4623);
xor U5452 (N_5452,N_4539,N_4942);
and U5453 (N_5453,N_4997,N_4935);
nand U5454 (N_5454,N_4819,N_4959);
or U5455 (N_5455,N_4629,N_4641);
xor U5456 (N_5456,N_4717,N_4650);
xnor U5457 (N_5457,N_4853,N_4616);
nor U5458 (N_5458,N_4940,N_4767);
or U5459 (N_5459,N_4755,N_4904);
xor U5460 (N_5460,N_4727,N_4603);
xor U5461 (N_5461,N_4692,N_4568);
or U5462 (N_5462,N_4966,N_4978);
nand U5463 (N_5463,N_4514,N_4857);
or U5464 (N_5464,N_4858,N_4763);
nand U5465 (N_5465,N_4689,N_4698);
or U5466 (N_5466,N_4797,N_4732);
and U5467 (N_5467,N_4500,N_4896);
or U5468 (N_5468,N_4746,N_4896);
or U5469 (N_5469,N_4924,N_4994);
nor U5470 (N_5470,N_4953,N_4761);
and U5471 (N_5471,N_4710,N_4536);
nand U5472 (N_5472,N_4931,N_4988);
nand U5473 (N_5473,N_4596,N_4810);
nand U5474 (N_5474,N_4693,N_4919);
nor U5475 (N_5475,N_4555,N_4640);
or U5476 (N_5476,N_4607,N_4982);
nand U5477 (N_5477,N_4840,N_4798);
nand U5478 (N_5478,N_4515,N_4682);
nor U5479 (N_5479,N_4692,N_4857);
nand U5480 (N_5480,N_4748,N_4547);
xnor U5481 (N_5481,N_4972,N_4995);
or U5482 (N_5482,N_4619,N_4670);
nor U5483 (N_5483,N_4782,N_4913);
nor U5484 (N_5484,N_4532,N_4559);
nor U5485 (N_5485,N_4820,N_4587);
nand U5486 (N_5486,N_4567,N_4938);
xor U5487 (N_5487,N_4875,N_4619);
xor U5488 (N_5488,N_4813,N_4848);
nand U5489 (N_5489,N_4963,N_4858);
nand U5490 (N_5490,N_4679,N_4898);
or U5491 (N_5491,N_4959,N_4893);
or U5492 (N_5492,N_4792,N_4530);
and U5493 (N_5493,N_4962,N_4842);
nand U5494 (N_5494,N_4951,N_4702);
and U5495 (N_5495,N_4755,N_4954);
nand U5496 (N_5496,N_4640,N_4528);
nor U5497 (N_5497,N_4921,N_4538);
nand U5498 (N_5498,N_4779,N_4934);
nor U5499 (N_5499,N_4799,N_4601);
nand U5500 (N_5500,N_5100,N_5211);
and U5501 (N_5501,N_5095,N_5156);
xnor U5502 (N_5502,N_5213,N_5007);
or U5503 (N_5503,N_5191,N_5099);
nand U5504 (N_5504,N_5217,N_5404);
or U5505 (N_5505,N_5143,N_5473);
or U5506 (N_5506,N_5197,N_5267);
or U5507 (N_5507,N_5270,N_5113);
and U5508 (N_5508,N_5277,N_5078);
or U5509 (N_5509,N_5260,N_5126);
or U5510 (N_5510,N_5476,N_5196);
and U5511 (N_5511,N_5447,N_5451);
and U5512 (N_5512,N_5210,N_5180);
and U5513 (N_5513,N_5269,N_5232);
nor U5514 (N_5514,N_5075,N_5487);
nand U5515 (N_5515,N_5496,N_5157);
xnor U5516 (N_5516,N_5306,N_5389);
or U5517 (N_5517,N_5429,N_5309);
or U5518 (N_5518,N_5322,N_5106);
nor U5519 (N_5519,N_5062,N_5367);
and U5520 (N_5520,N_5227,N_5424);
nor U5521 (N_5521,N_5441,N_5365);
nor U5522 (N_5522,N_5033,N_5202);
nand U5523 (N_5523,N_5460,N_5030);
nor U5524 (N_5524,N_5163,N_5419);
or U5525 (N_5525,N_5125,N_5042);
and U5526 (N_5526,N_5304,N_5248);
nor U5527 (N_5527,N_5082,N_5250);
nand U5528 (N_5528,N_5205,N_5034);
and U5529 (N_5529,N_5194,N_5142);
xnor U5530 (N_5530,N_5313,N_5076);
and U5531 (N_5531,N_5357,N_5264);
nand U5532 (N_5532,N_5006,N_5107);
and U5533 (N_5533,N_5225,N_5065);
or U5534 (N_5534,N_5430,N_5437);
nor U5535 (N_5535,N_5017,N_5321);
or U5536 (N_5536,N_5491,N_5284);
and U5537 (N_5537,N_5040,N_5302);
or U5538 (N_5538,N_5330,N_5218);
nor U5539 (N_5539,N_5031,N_5358);
and U5540 (N_5540,N_5059,N_5381);
and U5541 (N_5541,N_5041,N_5026);
nand U5542 (N_5542,N_5010,N_5458);
nor U5543 (N_5543,N_5454,N_5391);
or U5544 (N_5544,N_5016,N_5360);
and U5545 (N_5545,N_5161,N_5150);
or U5546 (N_5546,N_5370,N_5188);
or U5547 (N_5547,N_5448,N_5146);
and U5548 (N_5548,N_5052,N_5477);
xnor U5549 (N_5549,N_5485,N_5344);
nor U5550 (N_5550,N_5400,N_5054);
xnor U5551 (N_5551,N_5296,N_5254);
xor U5552 (N_5552,N_5499,N_5081);
nor U5553 (N_5553,N_5114,N_5317);
and U5554 (N_5554,N_5453,N_5275);
nand U5555 (N_5555,N_5085,N_5325);
nand U5556 (N_5556,N_5350,N_5061);
xor U5557 (N_5557,N_5044,N_5170);
nand U5558 (N_5558,N_5333,N_5292);
or U5559 (N_5559,N_5395,N_5092);
or U5560 (N_5560,N_5377,N_5077);
nand U5561 (N_5561,N_5204,N_5220);
and U5562 (N_5562,N_5393,N_5459);
and U5563 (N_5563,N_5425,N_5167);
xor U5564 (N_5564,N_5049,N_5481);
or U5565 (N_5565,N_5411,N_5449);
or U5566 (N_5566,N_5489,N_5402);
and U5567 (N_5567,N_5199,N_5039);
or U5568 (N_5568,N_5435,N_5467);
nand U5569 (N_5569,N_5127,N_5004);
and U5570 (N_5570,N_5000,N_5193);
nand U5571 (N_5571,N_5410,N_5490);
and U5572 (N_5572,N_5261,N_5186);
or U5573 (N_5573,N_5116,N_5238);
nand U5574 (N_5574,N_5450,N_5427);
nand U5575 (N_5575,N_5074,N_5329);
nand U5576 (N_5576,N_5339,N_5366);
and U5577 (N_5577,N_5298,N_5242);
nor U5578 (N_5578,N_5070,N_5035);
nor U5579 (N_5579,N_5145,N_5421);
nand U5580 (N_5580,N_5086,N_5417);
nand U5581 (N_5581,N_5474,N_5209);
xnor U5582 (N_5582,N_5368,N_5198);
nand U5583 (N_5583,N_5356,N_5120);
nand U5584 (N_5584,N_5256,N_5064);
and U5585 (N_5585,N_5324,N_5266);
and U5586 (N_5586,N_5274,N_5349);
nor U5587 (N_5587,N_5137,N_5201);
or U5588 (N_5588,N_5183,N_5245);
xnor U5589 (N_5589,N_5109,N_5436);
nor U5590 (N_5590,N_5463,N_5177);
nand U5591 (N_5591,N_5282,N_5397);
or U5592 (N_5592,N_5222,N_5392);
xnor U5593 (N_5593,N_5223,N_5015);
nand U5594 (N_5594,N_5090,N_5305);
and U5595 (N_5595,N_5228,N_5221);
nor U5596 (N_5596,N_5008,N_5179);
and U5597 (N_5597,N_5363,N_5399);
or U5598 (N_5598,N_5159,N_5431);
nor U5599 (N_5599,N_5046,N_5405);
and U5600 (N_5600,N_5002,N_5452);
nor U5601 (N_5601,N_5158,N_5129);
nor U5602 (N_5602,N_5401,N_5243);
or U5603 (N_5603,N_5257,N_5140);
xor U5604 (N_5604,N_5434,N_5083);
or U5605 (N_5605,N_5244,N_5051);
xnor U5606 (N_5606,N_5440,N_5318);
and U5607 (N_5607,N_5475,N_5268);
or U5608 (N_5608,N_5406,N_5048);
or U5609 (N_5609,N_5111,N_5214);
nand U5610 (N_5610,N_5272,N_5438);
or U5611 (N_5611,N_5375,N_5479);
or U5612 (N_5612,N_5276,N_5340);
or U5613 (N_5613,N_5373,N_5239);
and U5614 (N_5614,N_5294,N_5301);
or U5615 (N_5615,N_5480,N_5029);
xor U5616 (N_5616,N_5484,N_5383);
and U5617 (N_5617,N_5005,N_5045);
or U5618 (N_5618,N_5172,N_5018);
and U5619 (N_5619,N_5295,N_5439);
nor U5620 (N_5620,N_5493,N_5098);
nor U5621 (N_5621,N_5422,N_5025);
or U5622 (N_5622,N_5128,N_5303);
or U5623 (N_5623,N_5396,N_5009);
xnor U5624 (N_5624,N_5038,N_5148);
and U5625 (N_5625,N_5206,N_5465);
xnor U5626 (N_5626,N_5273,N_5027);
nand U5627 (N_5627,N_5043,N_5162);
nor U5628 (N_5628,N_5182,N_5253);
or U5629 (N_5629,N_5153,N_5003);
or U5630 (N_5630,N_5249,N_5192);
and U5631 (N_5631,N_5262,N_5311);
nand U5632 (N_5632,N_5320,N_5297);
and U5633 (N_5633,N_5293,N_5247);
and U5634 (N_5634,N_5011,N_5104);
nor U5635 (N_5635,N_5445,N_5428);
nand U5636 (N_5636,N_5118,N_5079);
xor U5637 (N_5637,N_5184,N_5251);
xnor U5638 (N_5638,N_5073,N_5139);
nand U5639 (N_5639,N_5337,N_5335);
or U5640 (N_5640,N_5338,N_5168);
or U5641 (N_5641,N_5382,N_5415);
or U5642 (N_5642,N_5271,N_5135);
nand U5643 (N_5643,N_5147,N_5088);
and U5644 (N_5644,N_5123,N_5133);
and U5645 (N_5645,N_5319,N_5328);
nand U5646 (N_5646,N_5130,N_5498);
nor U5647 (N_5647,N_5331,N_5461);
nor U5648 (N_5648,N_5121,N_5110);
or U5649 (N_5649,N_5200,N_5160);
or U5650 (N_5650,N_5495,N_5355);
or U5651 (N_5651,N_5105,N_5470);
nor U5652 (N_5652,N_5001,N_5281);
nand U5653 (N_5653,N_5134,N_5055);
and U5654 (N_5654,N_5229,N_5108);
and U5655 (N_5655,N_5021,N_5394);
nand U5656 (N_5656,N_5345,N_5359);
and U5657 (N_5657,N_5386,N_5068);
nor U5658 (N_5658,N_5216,N_5326);
and U5659 (N_5659,N_5144,N_5056);
and U5660 (N_5660,N_5084,N_5066);
nor U5661 (N_5661,N_5283,N_5036);
nand U5662 (N_5662,N_5483,N_5327);
xor U5663 (N_5663,N_5285,N_5478);
xnor U5664 (N_5664,N_5444,N_5057);
and U5665 (N_5665,N_5291,N_5390);
nand U5666 (N_5666,N_5175,N_5224);
nand U5667 (N_5667,N_5014,N_5050);
xor U5668 (N_5668,N_5181,N_5091);
or U5669 (N_5669,N_5067,N_5376);
and U5670 (N_5670,N_5259,N_5246);
and U5671 (N_5671,N_5351,N_5418);
or U5672 (N_5672,N_5323,N_5426);
nand U5673 (N_5673,N_5455,N_5252);
nand U5674 (N_5674,N_5403,N_5132);
nor U5675 (N_5675,N_5456,N_5233);
xor U5676 (N_5676,N_5019,N_5255);
nand U5677 (N_5677,N_5115,N_5384);
nor U5678 (N_5678,N_5346,N_5412);
xor U5679 (N_5679,N_5165,N_5013);
or U5680 (N_5680,N_5122,N_5028);
or U5681 (N_5681,N_5315,N_5492);
xnor U5682 (N_5682,N_5457,N_5387);
or U5683 (N_5683,N_5385,N_5316);
nor U5684 (N_5684,N_5169,N_5408);
nand U5685 (N_5685,N_5190,N_5388);
nand U5686 (N_5686,N_5258,N_5471);
nand U5687 (N_5687,N_5300,N_5378);
and U5688 (N_5688,N_5189,N_5203);
xor U5689 (N_5689,N_5497,N_5053);
nor U5690 (N_5690,N_5468,N_5069);
nor U5691 (N_5691,N_5174,N_5494);
or U5692 (N_5692,N_5080,N_5173);
nor U5693 (N_5693,N_5012,N_5290);
nand U5694 (N_5694,N_5187,N_5094);
or U5695 (N_5695,N_5280,N_5101);
or U5696 (N_5696,N_5379,N_5195);
and U5697 (N_5697,N_5486,N_5409);
nand U5698 (N_5698,N_5097,N_5185);
nor U5699 (N_5699,N_5208,N_5149);
nand U5700 (N_5700,N_5372,N_5307);
or U5701 (N_5701,N_5347,N_5265);
nand U5702 (N_5702,N_5093,N_5263);
or U5703 (N_5703,N_5234,N_5063);
and U5704 (N_5704,N_5374,N_5420);
nor U5705 (N_5705,N_5332,N_5362);
nand U5706 (N_5706,N_5155,N_5141);
or U5707 (N_5707,N_5171,N_5136);
nand U5708 (N_5708,N_5380,N_5124);
xnor U5709 (N_5709,N_5354,N_5288);
xor U5710 (N_5710,N_5341,N_5071);
and U5711 (N_5711,N_5348,N_5154);
nand U5712 (N_5712,N_5219,N_5237);
and U5713 (N_5713,N_5022,N_5231);
nand U5714 (N_5714,N_5353,N_5020);
nor U5715 (N_5715,N_5310,N_5215);
nor U5716 (N_5716,N_5235,N_5464);
and U5717 (N_5717,N_5230,N_5442);
and U5718 (N_5718,N_5112,N_5037);
nand U5719 (N_5719,N_5087,N_5236);
nand U5720 (N_5720,N_5212,N_5369);
nor U5721 (N_5721,N_5072,N_5089);
and U5722 (N_5722,N_5024,N_5466);
nor U5723 (N_5723,N_5023,N_5096);
and U5724 (N_5724,N_5102,N_5416);
xor U5725 (N_5725,N_5278,N_5407);
and U5726 (N_5726,N_5166,N_5414);
or U5727 (N_5727,N_5289,N_5240);
nand U5728 (N_5728,N_5151,N_5178);
and U5729 (N_5729,N_5432,N_5152);
and U5730 (N_5730,N_5446,N_5287);
or U5731 (N_5731,N_5308,N_5103);
xor U5732 (N_5732,N_5342,N_5286);
and U5733 (N_5733,N_5164,N_5058);
nand U5734 (N_5734,N_5482,N_5241);
nand U5735 (N_5735,N_5032,N_5207);
nor U5736 (N_5736,N_5226,N_5314);
and U5737 (N_5737,N_5352,N_5488);
nor U5738 (N_5738,N_5462,N_5364);
nor U5739 (N_5739,N_5131,N_5423);
and U5740 (N_5740,N_5138,N_5472);
nand U5741 (N_5741,N_5398,N_5433);
xnor U5742 (N_5742,N_5443,N_5279);
xnor U5743 (N_5743,N_5334,N_5336);
nand U5744 (N_5744,N_5117,N_5176);
and U5745 (N_5745,N_5343,N_5119);
xor U5746 (N_5746,N_5047,N_5361);
or U5747 (N_5747,N_5299,N_5312);
and U5748 (N_5748,N_5060,N_5413);
and U5749 (N_5749,N_5469,N_5371);
xor U5750 (N_5750,N_5240,N_5246);
or U5751 (N_5751,N_5405,N_5266);
nand U5752 (N_5752,N_5397,N_5338);
nand U5753 (N_5753,N_5401,N_5484);
and U5754 (N_5754,N_5205,N_5158);
or U5755 (N_5755,N_5300,N_5295);
nor U5756 (N_5756,N_5299,N_5180);
or U5757 (N_5757,N_5148,N_5447);
nand U5758 (N_5758,N_5395,N_5447);
xnor U5759 (N_5759,N_5174,N_5270);
and U5760 (N_5760,N_5349,N_5169);
or U5761 (N_5761,N_5243,N_5193);
and U5762 (N_5762,N_5396,N_5018);
nand U5763 (N_5763,N_5496,N_5056);
xnor U5764 (N_5764,N_5492,N_5149);
and U5765 (N_5765,N_5352,N_5306);
xnor U5766 (N_5766,N_5440,N_5419);
and U5767 (N_5767,N_5352,N_5097);
xor U5768 (N_5768,N_5249,N_5183);
and U5769 (N_5769,N_5223,N_5447);
nor U5770 (N_5770,N_5025,N_5230);
nand U5771 (N_5771,N_5065,N_5319);
nand U5772 (N_5772,N_5310,N_5294);
xor U5773 (N_5773,N_5321,N_5344);
xor U5774 (N_5774,N_5298,N_5048);
or U5775 (N_5775,N_5136,N_5341);
nand U5776 (N_5776,N_5377,N_5148);
xnor U5777 (N_5777,N_5157,N_5373);
xnor U5778 (N_5778,N_5351,N_5195);
nand U5779 (N_5779,N_5323,N_5387);
nor U5780 (N_5780,N_5378,N_5336);
xor U5781 (N_5781,N_5106,N_5244);
nor U5782 (N_5782,N_5432,N_5471);
nand U5783 (N_5783,N_5063,N_5327);
or U5784 (N_5784,N_5235,N_5207);
or U5785 (N_5785,N_5341,N_5295);
nand U5786 (N_5786,N_5289,N_5044);
nor U5787 (N_5787,N_5120,N_5019);
nor U5788 (N_5788,N_5176,N_5210);
nand U5789 (N_5789,N_5001,N_5123);
nand U5790 (N_5790,N_5235,N_5272);
nand U5791 (N_5791,N_5046,N_5489);
nand U5792 (N_5792,N_5213,N_5032);
nand U5793 (N_5793,N_5287,N_5451);
and U5794 (N_5794,N_5324,N_5395);
xor U5795 (N_5795,N_5274,N_5493);
nand U5796 (N_5796,N_5175,N_5242);
nor U5797 (N_5797,N_5115,N_5049);
xor U5798 (N_5798,N_5239,N_5304);
and U5799 (N_5799,N_5094,N_5166);
and U5800 (N_5800,N_5085,N_5433);
or U5801 (N_5801,N_5161,N_5354);
or U5802 (N_5802,N_5295,N_5051);
xnor U5803 (N_5803,N_5314,N_5255);
nor U5804 (N_5804,N_5392,N_5421);
nor U5805 (N_5805,N_5026,N_5104);
or U5806 (N_5806,N_5126,N_5390);
or U5807 (N_5807,N_5322,N_5155);
nor U5808 (N_5808,N_5347,N_5411);
nor U5809 (N_5809,N_5113,N_5167);
nand U5810 (N_5810,N_5289,N_5290);
nor U5811 (N_5811,N_5496,N_5401);
nor U5812 (N_5812,N_5171,N_5404);
nor U5813 (N_5813,N_5376,N_5198);
xnor U5814 (N_5814,N_5427,N_5324);
xor U5815 (N_5815,N_5433,N_5099);
nor U5816 (N_5816,N_5148,N_5285);
and U5817 (N_5817,N_5134,N_5261);
nand U5818 (N_5818,N_5414,N_5031);
or U5819 (N_5819,N_5419,N_5019);
and U5820 (N_5820,N_5149,N_5448);
and U5821 (N_5821,N_5145,N_5047);
nand U5822 (N_5822,N_5229,N_5422);
or U5823 (N_5823,N_5114,N_5018);
nor U5824 (N_5824,N_5488,N_5199);
nor U5825 (N_5825,N_5204,N_5054);
and U5826 (N_5826,N_5382,N_5413);
and U5827 (N_5827,N_5258,N_5095);
nand U5828 (N_5828,N_5205,N_5177);
or U5829 (N_5829,N_5476,N_5437);
nand U5830 (N_5830,N_5119,N_5099);
xor U5831 (N_5831,N_5416,N_5348);
or U5832 (N_5832,N_5383,N_5175);
nor U5833 (N_5833,N_5365,N_5118);
or U5834 (N_5834,N_5081,N_5195);
nand U5835 (N_5835,N_5489,N_5311);
nor U5836 (N_5836,N_5277,N_5086);
nand U5837 (N_5837,N_5412,N_5207);
and U5838 (N_5838,N_5340,N_5105);
nand U5839 (N_5839,N_5073,N_5051);
or U5840 (N_5840,N_5323,N_5101);
nor U5841 (N_5841,N_5001,N_5426);
nand U5842 (N_5842,N_5290,N_5175);
nor U5843 (N_5843,N_5483,N_5066);
nor U5844 (N_5844,N_5293,N_5497);
or U5845 (N_5845,N_5304,N_5173);
or U5846 (N_5846,N_5401,N_5134);
xnor U5847 (N_5847,N_5261,N_5105);
or U5848 (N_5848,N_5228,N_5425);
xnor U5849 (N_5849,N_5359,N_5475);
xor U5850 (N_5850,N_5486,N_5224);
nand U5851 (N_5851,N_5380,N_5311);
nor U5852 (N_5852,N_5240,N_5428);
nand U5853 (N_5853,N_5427,N_5124);
and U5854 (N_5854,N_5380,N_5049);
nand U5855 (N_5855,N_5492,N_5043);
nor U5856 (N_5856,N_5078,N_5126);
nor U5857 (N_5857,N_5241,N_5456);
nor U5858 (N_5858,N_5495,N_5175);
and U5859 (N_5859,N_5001,N_5056);
nor U5860 (N_5860,N_5048,N_5111);
or U5861 (N_5861,N_5210,N_5356);
nor U5862 (N_5862,N_5092,N_5259);
nand U5863 (N_5863,N_5497,N_5443);
nand U5864 (N_5864,N_5424,N_5144);
and U5865 (N_5865,N_5124,N_5144);
nor U5866 (N_5866,N_5395,N_5394);
nand U5867 (N_5867,N_5120,N_5346);
or U5868 (N_5868,N_5070,N_5421);
and U5869 (N_5869,N_5488,N_5082);
and U5870 (N_5870,N_5379,N_5025);
and U5871 (N_5871,N_5042,N_5372);
nor U5872 (N_5872,N_5389,N_5246);
or U5873 (N_5873,N_5430,N_5369);
or U5874 (N_5874,N_5417,N_5065);
nor U5875 (N_5875,N_5362,N_5479);
or U5876 (N_5876,N_5326,N_5358);
nand U5877 (N_5877,N_5345,N_5023);
and U5878 (N_5878,N_5441,N_5115);
nand U5879 (N_5879,N_5422,N_5041);
or U5880 (N_5880,N_5306,N_5173);
and U5881 (N_5881,N_5405,N_5356);
nor U5882 (N_5882,N_5184,N_5356);
nand U5883 (N_5883,N_5369,N_5330);
or U5884 (N_5884,N_5350,N_5288);
and U5885 (N_5885,N_5416,N_5460);
and U5886 (N_5886,N_5059,N_5368);
nand U5887 (N_5887,N_5229,N_5222);
nor U5888 (N_5888,N_5459,N_5045);
or U5889 (N_5889,N_5056,N_5464);
nor U5890 (N_5890,N_5014,N_5081);
xor U5891 (N_5891,N_5170,N_5194);
and U5892 (N_5892,N_5125,N_5008);
nand U5893 (N_5893,N_5211,N_5150);
or U5894 (N_5894,N_5227,N_5238);
nand U5895 (N_5895,N_5426,N_5470);
or U5896 (N_5896,N_5362,N_5307);
xor U5897 (N_5897,N_5220,N_5020);
xor U5898 (N_5898,N_5449,N_5048);
xnor U5899 (N_5899,N_5067,N_5495);
and U5900 (N_5900,N_5408,N_5352);
nand U5901 (N_5901,N_5094,N_5047);
or U5902 (N_5902,N_5331,N_5000);
xor U5903 (N_5903,N_5066,N_5057);
or U5904 (N_5904,N_5382,N_5008);
nand U5905 (N_5905,N_5146,N_5453);
and U5906 (N_5906,N_5143,N_5101);
xor U5907 (N_5907,N_5336,N_5189);
xnor U5908 (N_5908,N_5094,N_5300);
or U5909 (N_5909,N_5245,N_5067);
nand U5910 (N_5910,N_5274,N_5271);
or U5911 (N_5911,N_5144,N_5160);
nor U5912 (N_5912,N_5196,N_5104);
nand U5913 (N_5913,N_5322,N_5247);
xor U5914 (N_5914,N_5089,N_5145);
or U5915 (N_5915,N_5211,N_5480);
nor U5916 (N_5916,N_5322,N_5440);
xor U5917 (N_5917,N_5107,N_5099);
xnor U5918 (N_5918,N_5024,N_5179);
nand U5919 (N_5919,N_5250,N_5296);
and U5920 (N_5920,N_5050,N_5299);
xnor U5921 (N_5921,N_5394,N_5026);
or U5922 (N_5922,N_5032,N_5191);
or U5923 (N_5923,N_5283,N_5433);
and U5924 (N_5924,N_5432,N_5151);
and U5925 (N_5925,N_5339,N_5181);
and U5926 (N_5926,N_5277,N_5484);
or U5927 (N_5927,N_5083,N_5103);
or U5928 (N_5928,N_5206,N_5103);
and U5929 (N_5929,N_5070,N_5009);
xor U5930 (N_5930,N_5293,N_5470);
nand U5931 (N_5931,N_5290,N_5314);
nand U5932 (N_5932,N_5208,N_5494);
nor U5933 (N_5933,N_5333,N_5438);
nor U5934 (N_5934,N_5159,N_5201);
nor U5935 (N_5935,N_5070,N_5116);
xnor U5936 (N_5936,N_5375,N_5040);
nor U5937 (N_5937,N_5324,N_5020);
and U5938 (N_5938,N_5036,N_5285);
and U5939 (N_5939,N_5444,N_5428);
nand U5940 (N_5940,N_5402,N_5371);
nand U5941 (N_5941,N_5329,N_5430);
and U5942 (N_5942,N_5477,N_5329);
xor U5943 (N_5943,N_5171,N_5060);
nor U5944 (N_5944,N_5215,N_5254);
xnor U5945 (N_5945,N_5218,N_5243);
xnor U5946 (N_5946,N_5498,N_5315);
nor U5947 (N_5947,N_5489,N_5193);
nand U5948 (N_5948,N_5087,N_5010);
nand U5949 (N_5949,N_5245,N_5158);
xnor U5950 (N_5950,N_5266,N_5294);
nand U5951 (N_5951,N_5171,N_5453);
xnor U5952 (N_5952,N_5487,N_5441);
and U5953 (N_5953,N_5102,N_5321);
and U5954 (N_5954,N_5297,N_5003);
xnor U5955 (N_5955,N_5072,N_5204);
xor U5956 (N_5956,N_5342,N_5003);
nand U5957 (N_5957,N_5290,N_5264);
or U5958 (N_5958,N_5416,N_5219);
and U5959 (N_5959,N_5225,N_5250);
xor U5960 (N_5960,N_5482,N_5065);
or U5961 (N_5961,N_5092,N_5052);
nor U5962 (N_5962,N_5015,N_5056);
nor U5963 (N_5963,N_5432,N_5308);
nand U5964 (N_5964,N_5027,N_5138);
xor U5965 (N_5965,N_5427,N_5033);
and U5966 (N_5966,N_5179,N_5111);
nand U5967 (N_5967,N_5008,N_5085);
or U5968 (N_5968,N_5186,N_5238);
nand U5969 (N_5969,N_5478,N_5197);
nand U5970 (N_5970,N_5030,N_5405);
or U5971 (N_5971,N_5420,N_5328);
or U5972 (N_5972,N_5289,N_5308);
or U5973 (N_5973,N_5027,N_5194);
or U5974 (N_5974,N_5487,N_5227);
and U5975 (N_5975,N_5264,N_5482);
xnor U5976 (N_5976,N_5134,N_5410);
and U5977 (N_5977,N_5432,N_5256);
nand U5978 (N_5978,N_5187,N_5487);
nor U5979 (N_5979,N_5385,N_5382);
xnor U5980 (N_5980,N_5307,N_5305);
or U5981 (N_5981,N_5479,N_5452);
nor U5982 (N_5982,N_5488,N_5329);
nor U5983 (N_5983,N_5259,N_5158);
or U5984 (N_5984,N_5105,N_5095);
and U5985 (N_5985,N_5114,N_5423);
or U5986 (N_5986,N_5240,N_5498);
xor U5987 (N_5987,N_5296,N_5284);
nor U5988 (N_5988,N_5193,N_5452);
and U5989 (N_5989,N_5351,N_5114);
nand U5990 (N_5990,N_5434,N_5046);
nor U5991 (N_5991,N_5227,N_5486);
xor U5992 (N_5992,N_5387,N_5402);
xor U5993 (N_5993,N_5016,N_5408);
or U5994 (N_5994,N_5057,N_5171);
and U5995 (N_5995,N_5263,N_5203);
and U5996 (N_5996,N_5010,N_5309);
nor U5997 (N_5997,N_5456,N_5361);
nor U5998 (N_5998,N_5421,N_5062);
and U5999 (N_5999,N_5363,N_5174);
nand U6000 (N_6000,N_5746,N_5723);
nand U6001 (N_6001,N_5636,N_5698);
nand U6002 (N_6002,N_5719,N_5946);
or U6003 (N_6003,N_5691,N_5917);
and U6004 (N_6004,N_5867,N_5998);
nand U6005 (N_6005,N_5891,N_5561);
nor U6006 (N_6006,N_5855,N_5679);
and U6007 (N_6007,N_5965,N_5780);
nor U6008 (N_6008,N_5995,N_5713);
nor U6009 (N_6009,N_5554,N_5774);
xnor U6010 (N_6010,N_5744,N_5624);
and U6011 (N_6011,N_5957,N_5770);
xnor U6012 (N_6012,N_5631,N_5926);
or U6013 (N_6013,N_5531,N_5503);
nand U6014 (N_6014,N_5593,N_5854);
xnor U6015 (N_6015,N_5889,N_5704);
and U6016 (N_6016,N_5528,N_5865);
xnor U6017 (N_6017,N_5737,N_5586);
or U6018 (N_6018,N_5573,N_5844);
xor U6019 (N_6019,N_5654,N_5875);
and U6020 (N_6020,N_5981,N_5763);
nor U6021 (N_6021,N_5600,N_5539);
xor U6022 (N_6022,N_5546,N_5640);
nor U6023 (N_6023,N_5784,N_5976);
xnor U6024 (N_6024,N_5726,N_5545);
nand U6025 (N_6025,N_5595,N_5899);
xor U6026 (N_6026,N_5734,N_5563);
or U6027 (N_6027,N_5846,N_5836);
and U6028 (N_6028,N_5582,N_5896);
and U6029 (N_6029,N_5900,N_5847);
and U6030 (N_6030,N_5789,N_5630);
nand U6031 (N_6031,N_5575,N_5699);
or U6032 (N_6032,N_5978,N_5923);
or U6033 (N_6033,N_5859,N_5681);
nor U6034 (N_6034,N_5868,N_5930);
nor U6035 (N_6035,N_5626,N_5556);
or U6036 (N_6036,N_5783,N_5937);
xnor U6037 (N_6037,N_5715,N_5623);
or U6038 (N_6038,N_5757,N_5851);
nand U6039 (N_6039,N_5835,N_5838);
and U6040 (N_6040,N_5710,N_5524);
and U6041 (N_6041,N_5878,N_5898);
nor U6042 (N_6042,N_5842,N_5897);
or U6043 (N_6043,N_5864,N_5509);
or U6044 (N_6044,N_5741,N_5906);
xnor U6045 (N_6045,N_5729,N_5559);
xnor U6046 (N_6046,N_5692,N_5728);
nand U6047 (N_6047,N_5607,N_5647);
and U6048 (N_6048,N_5638,N_5544);
nor U6049 (N_6049,N_5912,N_5580);
and U6050 (N_6050,N_5622,N_5797);
xnor U6051 (N_6051,N_5931,N_5673);
xnor U6052 (N_6052,N_5814,N_5806);
xnor U6053 (N_6053,N_5819,N_5525);
nor U6054 (N_6054,N_5656,N_5961);
and U6055 (N_6055,N_5667,N_5547);
and U6056 (N_6056,N_5823,N_5648);
and U6057 (N_6057,N_5802,N_5657);
or U6058 (N_6058,N_5615,N_5787);
and U6059 (N_6059,N_5739,N_5581);
xor U6060 (N_6060,N_5845,N_5954);
and U6061 (N_6061,N_5807,N_5996);
and U6062 (N_6062,N_5584,N_5949);
nor U6063 (N_6063,N_5672,N_5821);
nand U6064 (N_6064,N_5888,N_5629);
xor U6065 (N_6065,N_5651,N_5948);
xor U6066 (N_6066,N_5754,N_5810);
or U6067 (N_6067,N_5986,N_5568);
and U6068 (N_6068,N_5570,N_5676);
or U6069 (N_6069,N_5796,N_5975);
xnor U6070 (N_6070,N_5853,N_5811);
or U6071 (N_6071,N_5705,N_5655);
or U6072 (N_6072,N_5639,N_5934);
and U6073 (N_6073,N_5773,N_5759);
nand U6074 (N_6074,N_5733,N_5992);
or U6075 (N_6075,N_5738,N_5566);
nand U6076 (N_6076,N_5702,N_5960);
or U6077 (N_6077,N_5767,N_5512);
and U6078 (N_6078,N_5979,N_5879);
nand U6079 (N_6079,N_5680,N_5689);
and U6080 (N_6080,N_5997,N_5579);
xor U6081 (N_6081,N_5985,N_5781);
nor U6082 (N_6082,N_5971,N_5943);
nand U6083 (N_6083,N_5758,N_5771);
xor U6084 (N_6084,N_5808,N_5688);
or U6085 (N_6085,N_5766,N_5952);
nor U6086 (N_6086,N_5536,N_5519);
or U6087 (N_6087,N_5837,N_5678);
nor U6088 (N_6088,N_5550,N_5721);
or U6089 (N_6089,N_5760,N_5685);
nor U6090 (N_6090,N_5518,N_5974);
and U6091 (N_6091,N_5942,N_5703);
xnor U6092 (N_6092,N_5701,N_5765);
nor U6093 (N_6093,N_5990,N_5786);
or U6094 (N_6094,N_5884,N_5552);
and U6095 (N_6095,N_5506,N_5714);
xor U6096 (N_6096,N_5972,N_5696);
nor U6097 (N_6097,N_5973,N_5583);
and U6098 (N_6098,N_5747,N_5591);
nand U6099 (N_6099,N_5502,N_5542);
and U6100 (N_6100,N_5801,N_5970);
and U6101 (N_6101,N_5893,N_5769);
nand U6102 (N_6102,N_5813,N_5516);
xor U6103 (N_6103,N_5826,N_5827);
xor U6104 (N_6104,N_5824,N_5597);
and U6105 (N_6105,N_5939,N_5871);
nor U6106 (N_6106,N_5791,N_5849);
xnor U6107 (N_6107,N_5523,N_5700);
nand U6108 (N_6108,N_5543,N_5508);
xnor U6109 (N_6109,N_5812,N_5989);
nor U6110 (N_6110,N_5850,N_5727);
and U6111 (N_6111,N_5904,N_5594);
and U6112 (N_6112,N_5905,N_5914);
xor U6113 (N_6113,N_5510,N_5890);
xnor U6114 (N_6114,N_5565,N_5541);
nor U6115 (N_6115,N_5576,N_5772);
nand U6116 (N_6116,N_5664,N_5799);
or U6117 (N_6117,N_5574,N_5686);
nor U6118 (N_6118,N_5944,N_5947);
nor U6119 (N_6119,N_5732,N_5907);
xor U6120 (N_6120,N_5620,N_5562);
xor U6121 (N_6121,N_5841,N_5751);
and U6122 (N_6122,N_5936,N_5611);
and U6123 (N_6123,N_5677,N_5590);
nand U6124 (N_6124,N_5832,N_5668);
nor U6125 (N_6125,N_5618,N_5921);
nand U6126 (N_6126,N_5538,N_5553);
or U6127 (N_6127,N_5895,N_5885);
xnor U6128 (N_6128,N_5963,N_5848);
xnor U6129 (N_6129,N_5643,N_5745);
xnor U6130 (N_6130,N_5980,N_5507);
and U6131 (N_6131,N_5804,N_5782);
xor U6132 (N_6132,N_5609,N_5652);
or U6133 (N_6133,N_5788,N_5964);
nand U6134 (N_6134,N_5669,N_5852);
nor U6135 (N_6135,N_5828,N_5614);
nand U6136 (N_6136,N_5722,N_5604);
nor U6137 (N_6137,N_5716,N_5522);
or U6138 (N_6138,N_5924,N_5792);
or U6139 (N_6139,N_5682,N_5549);
or U6140 (N_6140,N_5641,N_5857);
nand U6141 (N_6141,N_5916,N_5551);
nor U6142 (N_6142,N_5925,N_5709);
nand U6143 (N_6143,N_5589,N_5775);
or U6144 (N_6144,N_5613,N_5564);
or U6145 (N_6145,N_5794,N_5612);
and U6146 (N_6146,N_5929,N_5927);
nor U6147 (N_6147,N_5752,N_5743);
nor U6148 (N_6148,N_5778,N_5911);
nor U6149 (N_6149,N_5762,N_5987);
and U6150 (N_6150,N_5953,N_5817);
or U6151 (N_6151,N_5874,N_5683);
nand U6152 (N_6152,N_5515,N_5616);
xnor U6153 (N_6153,N_5511,N_5560);
nor U6154 (N_6154,N_5894,N_5798);
or U6155 (N_6155,N_5818,N_5596);
nand U6156 (N_6156,N_5910,N_5717);
xor U6157 (N_6157,N_5659,N_5687);
or U6158 (N_6158,N_5736,N_5605);
nand U6159 (N_6159,N_5977,N_5650);
and U6160 (N_6160,N_5578,N_5517);
nor U6161 (N_6161,N_5843,N_5860);
and U6162 (N_6162,N_5708,N_5598);
nor U6163 (N_6163,N_5585,N_5628);
nor U6164 (N_6164,N_5940,N_5532);
nand U6165 (N_6165,N_5902,N_5634);
or U6166 (N_6166,N_5645,N_5764);
xnor U6167 (N_6167,N_5920,N_5742);
xor U6168 (N_6168,N_5839,N_5740);
or U6169 (N_6169,N_5666,N_5922);
xnor U6170 (N_6170,N_5505,N_5919);
nand U6171 (N_6171,N_5617,N_5822);
nor U6172 (N_6172,N_5969,N_5880);
and U6173 (N_6173,N_5557,N_5815);
and U6174 (N_6174,N_5540,N_5635);
or U6175 (N_6175,N_5803,N_5913);
and U6176 (N_6176,N_5671,N_5637);
and U6177 (N_6177,N_5886,N_5707);
nor U6178 (N_6178,N_5606,N_5500);
nand U6179 (N_6179,N_5950,N_5777);
and U6180 (N_6180,N_5514,N_5994);
nor U6181 (N_6181,N_5756,N_5935);
nand U6182 (N_6182,N_5951,N_5809);
and U6183 (N_6183,N_5873,N_5697);
nor U6184 (N_6184,N_5833,N_5627);
or U6185 (N_6185,N_5501,N_5881);
or U6186 (N_6186,N_5735,N_5993);
xor U6187 (N_6187,N_5670,N_5632);
nand U6188 (N_6188,N_5805,N_5928);
nor U6189 (N_6189,N_5675,N_5693);
nand U6190 (N_6190,N_5530,N_5856);
or U6191 (N_6191,N_5959,N_5753);
or U6192 (N_6192,N_5933,N_5755);
nand U6193 (N_6193,N_5903,N_5908);
or U6194 (N_6194,N_5711,N_5588);
xnor U6195 (N_6195,N_5958,N_5862);
and U6196 (N_6196,N_5674,N_5649);
nand U6197 (N_6197,N_5730,N_5748);
and U6198 (N_6198,N_5684,N_5941);
or U6199 (N_6199,N_5555,N_5779);
xnor U6200 (N_6200,N_5520,N_5962);
and U6201 (N_6201,N_5869,N_5840);
and U6202 (N_6202,N_5537,N_5776);
nor U6203 (N_6203,N_5535,N_5870);
xnor U6204 (N_6204,N_5863,N_5548);
nor U6205 (N_6205,N_5877,N_5527);
xnor U6206 (N_6206,N_5861,N_5619);
nor U6207 (N_6207,N_5829,N_5621);
and U6208 (N_6208,N_5724,N_5866);
nand U6209 (N_6209,N_5558,N_5984);
xnor U6210 (N_6210,N_5572,N_5909);
or U6211 (N_6211,N_5882,N_5642);
nand U6212 (N_6212,N_5800,N_5661);
nand U6213 (N_6213,N_5533,N_5915);
xnor U6214 (N_6214,N_5695,N_5599);
nor U6215 (N_6215,N_5610,N_5571);
nor U6216 (N_6216,N_5785,N_5749);
nor U6217 (N_6217,N_5956,N_5831);
xor U6218 (N_6218,N_5725,N_5901);
nor U6219 (N_6219,N_5662,N_5587);
nor U6220 (N_6220,N_5938,N_5663);
nor U6221 (N_6221,N_5968,N_5602);
nor U6222 (N_6222,N_5718,N_5768);
xnor U6223 (N_6223,N_5665,N_5750);
nand U6224 (N_6224,N_5694,N_5633);
nand U6225 (N_6225,N_5982,N_5534);
nor U6226 (N_6226,N_5816,N_5592);
nor U6227 (N_6227,N_5706,N_5999);
xor U6228 (N_6228,N_5988,N_5690);
and U6229 (N_6229,N_5513,N_5529);
and U6230 (N_6230,N_5601,N_5983);
nand U6231 (N_6231,N_5761,N_5646);
nor U6232 (N_6232,N_5653,N_5567);
xnor U6233 (N_6233,N_5955,N_5603);
nand U6234 (N_6234,N_5712,N_5504);
nand U6235 (N_6235,N_5918,N_5577);
nand U6236 (N_6236,N_5883,N_5872);
nor U6237 (N_6237,N_5731,N_5887);
and U6238 (N_6238,N_5876,N_5569);
xor U6239 (N_6239,N_5790,N_5991);
or U6240 (N_6240,N_5521,N_5825);
and U6241 (N_6241,N_5795,N_5660);
and U6242 (N_6242,N_5625,N_5820);
xor U6243 (N_6243,N_5644,N_5793);
nand U6244 (N_6244,N_5658,N_5967);
nand U6245 (N_6245,N_5834,N_5526);
or U6246 (N_6246,N_5892,N_5945);
or U6247 (N_6247,N_5608,N_5932);
xor U6248 (N_6248,N_5966,N_5830);
or U6249 (N_6249,N_5858,N_5720);
xnor U6250 (N_6250,N_5565,N_5854);
nor U6251 (N_6251,N_5622,N_5911);
nand U6252 (N_6252,N_5535,N_5590);
nor U6253 (N_6253,N_5825,N_5665);
xor U6254 (N_6254,N_5738,N_5746);
xnor U6255 (N_6255,N_5590,N_5760);
nand U6256 (N_6256,N_5947,N_5555);
nor U6257 (N_6257,N_5510,N_5976);
or U6258 (N_6258,N_5903,N_5764);
and U6259 (N_6259,N_5891,N_5873);
and U6260 (N_6260,N_5761,N_5848);
nor U6261 (N_6261,N_5981,N_5650);
or U6262 (N_6262,N_5968,N_5892);
nand U6263 (N_6263,N_5912,N_5835);
or U6264 (N_6264,N_5641,N_5967);
or U6265 (N_6265,N_5527,N_5930);
and U6266 (N_6266,N_5937,N_5975);
nor U6267 (N_6267,N_5547,N_5983);
nand U6268 (N_6268,N_5871,N_5655);
and U6269 (N_6269,N_5618,N_5567);
xnor U6270 (N_6270,N_5860,N_5585);
and U6271 (N_6271,N_5530,N_5614);
and U6272 (N_6272,N_5989,N_5863);
or U6273 (N_6273,N_5596,N_5968);
xnor U6274 (N_6274,N_5902,N_5910);
nor U6275 (N_6275,N_5873,N_5941);
nor U6276 (N_6276,N_5783,N_5749);
and U6277 (N_6277,N_5992,N_5669);
or U6278 (N_6278,N_5699,N_5577);
and U6279 (N_6279,N_5834,N_5853);
nor U6280 (N_6280,N_5783,N_5869);
xnor U6281 (N_6281,N_5602,N_5514);
or U6282 (N_6282,N_5782,N_5676);
or U6283 (N_6283,N_5759,N_5877);
or U6284 (N_6284,N_5902,N_5755);
and U6285 (N_6285,N_5633,N_5634);
xor U6286 (N_6286,N_5829,N_5766);
xnor U6287 (N_6287,N_5570,N_5663);
and U6288 (N_6288,N_5802,N_5728);
and U6289 (N_6289,N_5722,N_5959);
xnor U6290 (N_6290,N_5682,N_5899);
or U6291 (N_6291,N_5711,N_5855);
and U6292 (N_6292,N_5618,N_5823);
nor U6293 (N_6293,N_5770,N_5827);
nand U6294 (N_6294,N_5720,N_5812);
nand U6295 (N_6295,N_5538,N_5906);
nand U6296 (N_6296,N_5861,N_5683);
nand U6297 (N_6297,N_5602,N_5876);
xor U6298 (N_6298,N_5512,N_5630);
and U6299 (N_6299,N_5949,N_5937);
nand U6300 (N_6300,N_5695,N_5758);
and U6301 (N_6301,N_5809,N_5662);
and U6302 (N_6302,N_5687,N_5825);
or U6303 (N_6303,N_5965,N_5525);
and U6304 (N_6304,N_5573,N_5805);
nor U6305 (N_6305,N_5542,N_5629);
xor U6306 (N_6306,N_5825,N_5612);
xnor U6307 (N_6307,N_5717,N_5659);
nor U6308 (N_6308,N_5930,N_5788);
xor U6309 (N_6309,N_5673,N_5622);
xnor U6310 (N_6310,N_5699,N_5880);
or U6311 (N_6311,N_5561,N_5817);
and U6312 (N_6312,N_5731,N_5831);
or U6313 (N_6313,N_5988,N_5963);
or U6314 (N_6314,N_5882,N_5720);
nor U6315 (N_6315,N_5944,N_5801);
or U6316 (N_6316,N_5640,N_5777);
and U6317 (N_6317,N_5939,N_5840);
or U6318 (N_6318,N_5778,N_5676);
nor U6319 (N_6319,N_5578,N_5914);
or U6320 (N_6320,N_5970,N_5600);
xor U6321 (N_6321,N_5559,N_5553);
nand U6322 (N_6322,N_5767,N_5976);
or U6323 (N_6323,N_5709,N_5656);
nand U6324 (N_6324,N_5599,N_5821);
or U6325 (N_6325,N_5549,N_5711);
or U6326 (N_6326,N_5831,N_5760);
or U6327 (N_6327,N_5980,N_5721);
xor U6328 (N_6328,N_5942,N_5965);
nand U6329 (N_6329,N_5991,N_5740);
xnor U6330 (N_6330,N_5736,N_5745);
or U6331 (N_6331,N_5793,N_5831);
xor U6332 (N_6332,N_5628,N_5697);
or U6333 (N_6333,N_5874,N_5509);
nor U6334 (N_6334,N_5718,N_5970);
nor U6335 (N_6335,N_5930,N_5643);
nor U6336 (N_6336,N_5861,N_5584);
and U6337 (N_6337,N_5983,N_5539);
nor U6338 (N_6338,N_5760,N_5833);
xnor U6339 (N_6339,N_5993,N_5798);
or U6340 (N_6340,N_5870,N_5818);
or U6341 (N_6341,N_5753,N_5675);
nand U6342 (N_6342,N_5897,N_5778);
and U6343 (N_6343,N_5617,N_5866);
xnor U6344 (N_6344,N_5788,N_5870);
and U6345 (N_6345,N_5598,N_5887);
or U6346 (N_6346,N_5660,N_5877);
nor U6347 (N_6347,N_5961,N_5521);
xor U6348 (N_6348,N_5720,N_5908);
nor U6349 (N_6349,N_5890,N_5948);
nor U6350 (N_6350,N_5528,N_5999);
xnor U6351 (N_6351,N_5575,N_5551);
and U6352 (N_6352,N_5998,N_5644);
or U6353 (N_6353,N_5892,N_5673);
and U6354 (N_6354,N_5890,N_5965);
and U6355 (N_6355,N_5877,N_5796);
xor U6356 (N_6356,N_5881,N_5722);
nand U6357 (N_6357,N_5601,N_5617);
nor U6358 (N_6358,N_5972,N_5835);
xor U6359 (N_6359,N_5975,N_5914);
xor U6360 (N_6360,N_5568,N_5730);
and U6361 (N_6361,N_5605,N_5715);
xor U6362 (N_6362,N_5571,N_5764);
nor U6363 (N_6363,N_5823,N_5767);
or U6364 (N_6364,N_5604,N_5814);
and U6365 (N_6365,N_5758,N_5554);
xnor U6366 (N_6366,N_5720,N_5893);
and U6367 (N_6367,N_5759,N_5745);
and U6368 (N_6368,N_5822,N_5887);
xnor U6369 (N_6369,N_5615,N_5517);
and U6370 (N_6370,N_5626,N_5918);
nand U6371 (N_6371,N_5821,N_5899);
or U6372 (N_6372,N_5672,N_5910);
xnor U6373 (N_6373,N_5703,N_5817);
nor U6374 (N_6374,N_5995,N_5695);
or U6375 (N_6375,N_5731,N_5752);
nor U6376 (N_6376,N_5983,N_5815);
or U6377 (N_6377,N_5704,N_5807);
nand U6378 (N_6378,N_5958,N_5628);
xor U6379 (N_6379,N_5936,N_5709);
xnor U6380 (N_6380,N_5607,N_5969);
xor U6381 (N_6381,N_5670,N_5862);
nor U6382 (N_6382,N_5755,N_5825);
nand U6383 (N_6383,N_5864,N_5733);
nand U6384 (N_6384,N_5509,N_5881);
xnor U6385 (N_6385,N_5950,N_5871);
or U6386 (N_6386,N_5651,N_5807);
or U6387 (N_6387,N_5752,N_5833);
nand U6388 (N_6388,N_5593,N_5650);
and U6389 (N_6389,N_5924,N_5872);
or U6390 (N_6390,N_5556,N_5962);
or U6391 (N_6391,N_5942,N_5991);
or U6392 (N_6392,N_5912,N_5751);
nand U6393 (N_6393,N_5585,N_5974);
nand U6394 (N_6394,N_5780,N_5679);
nand U6395 (N_6395,N_5538,N_5618);
nor U6396 (N_6396,N_5625,N_5931);
or U6397 (N_6397,N_5952,N_5543);
xor U6398 (N_6398,N_5870,N_5531);
nor U6399 (N_6399,N_5705,N_5687);
xnor U6400 (N_6400,N_5677,N_5989);
nand U6401 (N_6401,N_5694,N_5604);
xor U6402 (N_6402,N_5672,N_5922);
nor U6403 (N_6403,N_5653,N_5710);
and U6404 (N_6404,N_5510,N_5708);
and U6405 (N_6405,N_5733,N_5604);
and U6406 (N_6406,N_5960,N_5784);
and U6407 (N_6407,N_5846,N_5924);
or U6408 (N_6408,N_5545,N_5608);
or U6409 (N_6409,N_5643,N_5973);
nand U6410 (N_6410,N_5754,N_5570);
and U6411 (N_6411,N_5618,N_5531);
nand U6412 (N_6412,N_5506,N_5541);
xor U6413 (N_6413,N_5923,N_5864);
nand U6414 (N_6414,N_5578,N_5827);
nand U6415 (N_6415,N_5935,N_5950);
or U6416 (N_6416,N_5803,N_5775);
or U6417 (N_6417,N_5537,N_5690);
nor U6418 (N_6418,N_5963,N_5697);
or U6419 (N_6419,N_5504,N_5843);
and U6420 (N_6420,N_5540,N_5868);
nand U6421 (N_6421,N_5769,N_5700);
nand U6422 (N_6422,N_5573,N_5643);
and U6423 (N_6423,N_5516,N_5922);
nor U6424 (N_6424,N_5990,N_5683);
nand U6425 (N_6425,N_5509,N_5773);
nand U6426 (N_6426,N_5884,N_5844);
or U6427 (N_6427,N_5541,N_5803);
nor U6428 (N_6428,N_5850,N_5535);
nand U6429 (N_6429,N_5652,N_5514);
and U6430 (N_6430,N_5907,N_5722);
nor U6431 (N_6431,N_5991,N_5792);
nand U6432 (N_6432,N_5973,N_5741);
xnor U6433 (N_6433,N_5626,N_5971);
or U6434 (N_6434,N_5661,N_5956);
nor U6435 (N_6435,N_5793,N_5525);
nor U6436 (N_6436,N_5892,N_5664);
and U6437 (N_6437,N_5611,N_5625);
and U6438 (N_6438,N_5730,N_5673);
xor U6439 (N_6439,N_5817,N_5795);
or U6440 (N_6440,N_5962,N_5739);
or U6441 (N_6441,N_5828,N_5894);
and U6442 (N_6442,N_5910,N_5519);
nand U6443 (N_6443,N_5557,N_5519);
or U6444 (N_6444,N_5632,N_5773);
or U6445 (N_6445,N_5893,N_5984);
or U6446 (N_6446,N_5904,N_5994);
nand U6447 (N_6447,N_5773,N_5820);
or U6448 (N_6448,N_5740,N_5651);
nand U6449 (N_6449,N_5504,N_5745);
xnor U6450 (N_6450,N_5904,N_5753);
nand U6451 (N_6451,N_5803,N_5745);
and U6452 (N_6452,N_5888,N_5942);
or U6453 (N_6453,N_5877,N_5999);
xor U6454 (N_6454,N_5579,N_5699);
or U6455 (N_6455,N_5699,N_5515);
nor U6456 (N_6456,N_5788,N_5850);
nand U6457 (N_6457,N_5569,N_5856);
or U6458 (N_6458,N_5945,N_5888);
or U6459 (N_6459,N_5942,N_5850);
nand U6460 (N_6460,N_5816,N_5609);
and U6461 (N_6461,N_5535,N_5941);
nand U6462 (N_6462,N_5860,N_5976);
nor U6463 (N_6463,N_5587,N_5715);
xor U6464 (N_6464,N_5684,N_5910);
xor U6465 (N_6465,N_5503,N_5601);
nor U6466 (N_6466,N_5740,N_5605);
or U6467 (N_6467,N_5621,N_5791);
or U6468 (N_6468,N_5868,N_5815);
or U6469 (N_6469,N_5822,N_5982);
xor U6470 (N_6470,N_5768,N_5563);
xor U6471 (N_6471,N_5574,N_5666);
nor U6472 (N_6472,N_5827,N_5866);
xor U6473 (N_6473,N_5576,N_5544);
xnor U6474 (N_6474,N_5845,N_5658);
or U6475 (N_6475,N_5726,N_5947);
nand U6476 (N_6476,N_5573,N_5519);
xor U6477 (N_6477,N_5703,N_5739);
and U6478 (N_6478,N_5776,N_5977);
xor U6479 (N_6479,N_5713,N_5512);
or U6480 (N_6480,N_5973,N_5977);
nand U6481 (N_6481,N_5878,N_5988);
nor U6482 (N_6482,N_5966,N_5539);
and U6483 (N_6483,N_5821,N_5866);
xnor U6484 (N_6484,N_5853,N_5753);
nand U6485 (N_6485,N_5647,N_5826);
nor U6486 (N_6486,N_5664,N_5631);
or U6487 (N_6487,N_5653,N_5717);
nand U6488 (N_6488,N_5567,N_5614);
or U6489 (N_6489,N_5556,N_5754);
nor U6490 (N_6490,N_5918,N_5563);
and U6491 (N_6491,N_5983,N_5624);
nand U6492 (N_6492,N_5642,N_5525);
xor U6493 (N_6493,N_5870,N_5762);
xnor U6494 (N_6494,N_5761,N_5894);
or U6495 (N_6495,N_5573,N_5616);
nor U6496 (N_6496,N_5509,N_5941);
xnor U6497 (N_6497,N_5538,N_5989);
xnor U6498 (N_6498,N_5725,N_5721);
nor U6499 (N_6499,N_5617,N_5997);
or U6500 (N_6500,N_6385,N_6044);
xor U6501 (N_6501,N_6437,N_6239);
or U6502 (N_6502,N_6312,N_6011);
nand U6503 (N_6503,N_6473,N_6001);
and U6504 (N_6504,N_6339,N_6463);
and U6505 (N_6505,N_6207,N_6096);
and U6506 (N_6506,N_6337,N_6230);
nor U6507 (N_6507,N_6277,N_6025);
and U6508 (N_6508,N_6480,N_6326);
nor U6509 (N_6509,N_6389,N_6004);
nor U6510 (N_6510,N_6432,N_6322);
xnor U6511 (N_6511,N_6137,N_6447);
or U6512 (N_6512,N_6106,N_6219);
nand U6513 (N_6513,N_6059,N_6186);
nand U6514 (N_6514,N_6058,N_6206);
or U6515 (N_6515,N_6095,N_6193);
and U6516 (N_6516,N_6279,N_6017);
and U6517 (N_6517,N_6350,N_6080);
or U6518 (N_6518,N_6470,N_6183);
nand U6519 (N_6519,N_6005,N_6194);
xnor U6520 (N_6520,N_6321,N_6085);
and U6521 (N_6521,N_6115,N_6391);
nor U6522 (N_6522,N_6212,N_6367);
or U6523 (N_6523,N_6126,N_6411);
and U6524 (N_6524,N_6346,N_6377);
nor U6525 (N_6525,N_6063,N_6236);
xor U6526 (N_6526,N_6185,N_6233);
nor U6527 (N_6527,N_6290,N_6468);
or U6528 (N_6528,N_6021,N_6332);
or U6529 (N_6529,N_6049,N_6048);
nand U6530 (N_6530,N_6408,N_6160);
nor U6531 (N_6531,N_6423,N_6174);
nand U6532 (N_6532,N_6338,N_6288);
nor U6533 (N_6533,N_6162,N_6157);
and U6534 (N_6534,N_6073,N_6429);
and U6535 (N_6535,N_6268,N_6336);
nor U6536 (N_6536,N_6150,N_6294);
or U6537 (N_6537,N_6135,N_6184);
nor U6538 (N_6538,N_6110,N_6242);
or U6539 (N_6539,N_6146,N_6291);
xor U6540 (N_6540,N_6421,N_6000);
nor U6541 (N_6541,N_6484,N_6287);
or U6542 (N_6542,N_6167,N_6091);
xor U6543 (N_6543,N_6072,N_6472);
and U6544 (N_6544,N_6077,N_6070);
xnor U6545 (N_6545,N_6410,N_6306);
xor U6546 (N_6546,N_6122,N_6226);
and U6547 (N_6547,N_6192,N_6246);
or U6548 (N_6548,N_6003,N_6462);
nor U6549 (N_6549,N_6248,N_6204);
nand U6550 (N_6550,N_6127,N_6170);
and U6551 (N_6551,N_6498,N_6442);
nor U6552 (N_6552,N_6453,N_6075);
nand U6553 (N_6553,N_6347,N_6330);
or U6554 (N_6554,N_6151,N_6022);
nor U6555 (N_6555,N_6384,N_6360);
nor U6556 (N_6556,N_6344,N_6315);
xor U6557 (N_6557,N_6222,N_6349);
nand U6558 (N_6558,N_6187,N_6314);
nor U6559 (N_6559,N_6008,N_6300);
nand U6560 (N_6560,N_6060,N_6234);
nor U6561 (N_6561,N_6262,N_6489);
xor U6562 (N_6562,N_6431,N_6313);
nor U6563 (N_6563,N_6179,N_6396);
nand U6564 (N_6564,N_6030,N_6199);
nor U6565 (N_6565,N_6276,N_6419);
or U6566 (N_6566,N_6253,N_6018);
xor U6567 (N_6567,N_6490,N_6220);
xnor U6568 (N_6568,N_6256,N_6166);
xnor U6569 (N_6569,N_6380,N_6323);
or U6570 (N_6570,N_6412,N_6494);
xnor U6571 (N_6571,N_6343,N_6238);
nand U6572 (N_6572,N_6175,N_6153);
nor U6573 (N_6573,N_6272,N_6040);
and U6574 (N_6574,N_6409,N_6295);
nand U6575 (N_6575,N_6352,N_6356);
nor U6576 (N_6576,N_6196,N_6200);
xor U6577 (N_6577,N_6086,N_6348);
and U6578 (N_6578,N_6034,N_6416);
nor U6579 (N_6579,N_6228,N_6145);
nand U6580 (N_6580,N_6168,N_6031);
and U6581 (N_6581,N_6016,N_6460);
or U6582 (N_6582,N_6052,N_6247);
nor U6583 (N_6583,N_6152,N_6090);
and U6584 (N_6584,N_6020,N_6491);
xnor U6585 (N_6585,N_6231,N_6033);
nor U6586 (N_6586,N_6123,N_6041);
and U6587 (N_6587,N_6109,N_6210);
or U6588 (N_6588,N_6088,N_6013);
xor U6589 (N_6589,N_6101,N_6173);
xor U6590 (N_6590,N_6138,N_6099);
or U6591 (N_6591,N_6042,N_6303);
xor U6592 (N_6592,N_6370,N_6397);
and U6593 (N_6593,N_6083,N_6198);
xnor U6594 (N_6594,N_6263,N_6057);
nor U6595 (N_6595,N_6172,N_6188);
nor U6596 (N_6596,N_6414,N_6171);
and U6597 (N_6597,N_6444,N_6324);
nand U6598 (N_6598,N_6482,N_6074);
and U6599 (N_6599,N_6136,N_6359);
and U6600 (N_6600,N_6098,N_6217);
xor U6601 (N_6601,N_6467,N_6364);
nor U6602 (N_6602,N_6366,N_6358);
or U6603 (N_6603,N_6297,N_6430);
nor U6604 (N_6604,N_6285,N_6250);
or U6605 (N_6605,N_6235,N_6158);
nor U6606 (N_6606,N_6014,N_6395);
nand U6607 (N_6607,N_6144,N_6037);
xnor U6608 (N_6608,N_6108,N_6402);
and U6609 (N_6609,N_6307,N_6069);
or U6610 (N_6610,N_6165,N_6425);
and U6611 (N_6611,N_6215,N_6213);
or U6612 (N_6612,N_6134,N_6131);
or U6613 (N_6613,N_6325,N_6032);
and U6614 (N_6614,N_6148,N_6441);
and U6615 (N_6615,N_6113,N_6399);
xnor U6616 (N_6616,N_6181,N_6007);
xnor U6617 (N_6617,N_6273,N_6012);
xnor U6618 (N_6618,N_6319,N_6378);
nand U6619 (N_6619,N_6093,N_6459);
or U6620 (N_6620,N_6120,N_6245);
xor U6621 (N_6621,N_6404,N_6465);
nand U6622 (N_6622,N_6082,N_6129);
nand U6623 (N_6623,N_6114,N_6401);
nor U6624 (N_6624,N_6026,N_6061);
nand U6625 (N_6625,N_6365,N_6054);
nor U6626 (N_6626,N_6392,N_6289);
nor U6627 (N_6627,N_6164,N_6045);
nand U6628 (N_6628,N_6433,N_6269);
nand U6629 (N_6629,N_6182,N_6439);
and U6630 (N_6630,N_6050,N_6438);
or U6631 (N_6631,N_6499,N_6147);
and U6632 (N_6632,N_6039,N_6124);
nand U6633 (N_6633,N_6311,N_6284);
xnor U6634 (N_6634,N_6149,N_6400);
and U6635 (N_6635,N_6418,N_6161);
xnor U6636 (N_6636,N_6481,N_6112);
nor U6637 (N_6637,N_6225,N_6002);
and U6638 (N_6638,N_6374,N_6451);
or U6639 (N_6639,N_6260,N_6329);
nand U6640 (N_6640,N_6201,N_6267);
nand U6641 (N_6641,N_6125,N_6156);
and U6642 (N_6642,N_6483,N_6195);
or U6643 (N_6643,N_6117,N_6116);
nand U6644 (N_6644,N_6296,N_6105);
nand U6645 (N_6645,N_6232,N_6251);
or U6646 (N_6646,N_6216,N_6051);
and U6647 (N_6647,N_6353,N_6477);
nand U6648 (N_6648,N_6141,N_6218);
xor U6649 (N_6649,N_6104,N_6316);
and U6650 (N_6650,N_6068,N_6208);
nor U6651 (N_6651,N_6487,N_6413);
xnor U6652 (N_6652,N_6205,N_6372);
xnor U6653 (N_6653,N_6055,N_6202);
nand U6654 (N_6654,N_6209,N_6043);
nor U6655 (N_6655,N_6363,N_6027);
and U6656 (N_6656,N_6286,N_6440);
nand U6657 (N_6657,N_6293,N_6244);
xor U6658 (N_6658,N_6282,N_6373);
nor U6659 (N_6659,N_6422,N_6426);
or U6660 (N_6660,N_6169,N_6275);
nand U6661 (N_6661,N_6143,N_6038);
nor U6662 (N_6662,N_6456,N_6065);
nor U6663 (N_6663,N_6434,N_6028);
xnor U6664 (N_6664,N_6351,N_6254);
xnor U6665 (N_6665,N_6229,N_6062);
and U6666 (N_6666,N_6006,N_6066);
nand U6667 (N_6667,N_6318,N_6428);
or U6668 (N_6668,N_6457,N_6203);
and U6669 (N_6669,N_6130,N_6274);
and U6670 (N_6670,N_6092,N_6492);
xnor U6671 (N_6671,N_6355,N_6403);
and U6672 (N_6672,N_6495,N_6299);
nand U6673 (N_6673,N_6255,N_6094);
nor U6674 (N_6674,N_6476,N_6118);
xnor U6675 (N_6675,N_6335,N_6393);
nand U6676 (N_6676,N_6067,N_6461);
nand U6677 (N_6677,N_6308,N_6159);
nor U6678 (N_6678,N_6446,N_6280);
nand U6679 (N_6679,N_6420,N_6121);
xor U6680 (N_6680,N_6331,N_6455);
and U6681 (N_6681,N_6310,N_6452);
xor U6682 (N_6682,N_6024,N_6278);
and U6683 (N_6683,N_6304,N_6496);
nor U6684 (N_6684,N_6298,N_6478);
xnor U6685 (N_6685,N_6394,N_6227);
xor U6686 (N_6686,N_6089,N_6435);
xnor U6687 (N_6687,N_6271,N_6261);
and U6688 (N_6688,N_6076,N_6493);
nand U6689 (N_6689,N_6197,N_6371);
or U6690 (N_6690,N_6047,N_6265);
xor U6691 (N_6691,N_6485,N_6317);
xor U6692 (N_6692,N_6163,N_6281);
nand U6693 (N_6693,N_6376,N_6375);
and U6694 (N_6694,N_6379,N_6191);
or U6695 (N_6695,N_6368,N_6270);
nor U6696 (N_6696,N_6214,N_6252);
nand U6697 (N_6697,N_6301,N_6383);
and U6698 (N_6698,N_6128,N_6388);
nor U6699 (N_6699,N_6327,N_6223);
or U6700 (N_6700,N_6398,N_6340);
nor U6701 (N_6701,N_6139,N_6479);
or U6702 (N_6702,N_6464,N_6454);
xnor U6703 (N_6703,N_6333,N_6320);
nand U6704 (N_6704,N_6176,N_6241);
nor U6705 (N_6705,N_6087,N_6053);
nor U6706 (N_6706,N_6341,N_6056);
nor U6707 (N_6707,N_6180,N_6458);
and U6708 (N_6708,N_6382,N_6436);
and U6709 (N_6709,N_6450,N_6036);
nor U6710 (N_6710,N_6097,N_6107);
and U6711 (N_6711,N_6249,N_6142);
or U6712 (N_6712,N_6334,N_6009);
nor U6713 (N_6713,N_6100,N_6305);
nand U6714 (N_6714,N_6427,N_6081);
nand U6715 (N_6715,N_6445,N_6140);
nand U6716 (N_6716,N_6119,N_6357);
and U6717 (N_6717,N_6240,N_6309);
and U6718 (N_6718,N_6010,N_6448);
and U6719 (N_6719,N_6475,N_6471);
nor U6720 (N_6720,N_6497,N_6019);
nand U6721 (N_6721,N_6466,N_6342);
nor U6722 (N_6722,N_6362,N_6474);
or U6723 (N_6723,N_6102,N_6103);
nor U6724 (N_6724,N_6415,N_6133);
or U6725 (N_6725,N_6071,N_6029);
or U6726 (N_6726,N_6211,N_6023);
nand U6727 (N_6727,N_6224,N_6190);
nand U6728 (N_6728,N_6424,N_6486);
or U6729 (N_6729,N_6243,N_6406);
nor U6730 (N_6730,N_6257,N_6035);
and U6731 (N_6731,N_6258,N_6407);
or U6732 (N_6732,N_6488,N_6266);
or U6733 (N_6733,N_6302,N_6015);
xnor U6734 (N_6734,N_6155,N_6443);
xnor U6735 (N_6735,N_6417,N_6328);
and U6736 (N_6736,N_6189,N_6111);
nor U6737 (N_6737,N_6387,N_6078);
or U6738 (N_6738,N_6079,N_6369);
nor U6739 (N_6739,N_6154,N_6177);
nor U6740 (N_6740,N_6064,N_6361);
nor U6741 (N_6741,N_6292,N_6449);
or U6742 (N_6742,N_6354,N_6381);
xnor U6743 (N_6743,N_6405,N_6084);
or U6744 (N_6744,N_6221,N_6132);
or U6745 (N_6745,N_6386,N_6046);
nor U6746 (N_6746,N_6283,N_6345);
nor U6747 (N_6747,N_6259,N_6237);
nand U6748 (N_6748,N_6264,N_6390);
xnor U6749 (N_6749,N_6178,N_6469);
and U6750 (N_6750,N_6289,N_6400);
nor U6751 (N_6751,N_6420,N_6353);
nand U6752 (N_6752,N_6090,N_6289);
and U6753 (N_6753,N_6163,N_6219);
nor U6754 (N_6754,N_6286,N_6053);
or U6755 (N_6755,N_6045,N_6027);
or U6756 (N_6756,N_6282,N_6070);
xor U6757 (N_6757,N_6452,N_6164);
or U6758 (N_6758,N_6025,N_6028);
xor U6759 (N_6759,N_6372,N_6127);
nor U6760 (N_6760,N_6470,N_6404);
xor U6761 (N_6761,N_6390,N_6051);
xnor U6762 (N_6762,N_6363,N_6434);
and U6763 (N_6763,N_6146,N_6413);
nor U6764 (N_6764,N_6086,N_6464);
and U6765 (N_6765,N_6115,N_6206);
nand U6766 (N_6766,N_6220,N_6256);
xnor U6767 (N_6767,N_6097,N_6420);
or U6768 (N_6768,N_6223,N_6386);
and U6769 (N_6769,N_6170,N_6293);
nand U6770 (N_6770,N_6150,N_6438);
and U6771 (N_6771,N_6128,N_6332);
or U6772 (N_6772,N_6095,N_6393);
xnor U6773 (N_6773,N_6382,N_6050);
nor U6774 (N_6774,N_6216,N_6168);
nand U6775 (N_6775,N_6217,N_6079);
nand U6776 (N_6776,N_6380,N_6208);
nor U6777 (N_6777,N_6466,N_6306);
or U6778 (N_6778,N_6067,N_6255);
nand U6779 (N_6779,N_6240,N_6270);
nand U6780 (N_6780,N_6429,N_6149);
xor U6781 (N_6781,N_6036,N_6247);
or U6782 (N_6782,N_6097,N_6185);
or U6783 (N_6783,N_6115,N_6014);
or U6784 (N_6784,N_6038,N_6464);
and U6785 (N_6785,N_6152,N_6322);
xor U6786 (N_6786,N_6464,N_6415);
xnor U6787 (N_6787,N_6378,N_6063);
xor U6788 (N_6788,N_6141,N_6442);
or U6789 (N_6789,N_6449,N_6252);
nor U6790 (N_6790,N_6000,N_6061);
or U6791 (N_6791,N_6471,N_6117);
nand U6792 (N_6792,N_6257,N_6080);
nor U6793 (N_6793,N_6087,N_6097);
and U6794 (N_6794,N_6377,N_6221);
xnor U6795 (N_6795,N_6144,N_6447);
nor U6796 (N_6796,N_6060,N_6052);
xor U6797 (N_6797,N_6147,N_6217);
nor U6798 (N_6798,N_6002,N_6052);
nor U6799 (N_6799,N_6035,N_6354);
and U6800 (N_6800,N_6254,N_6423);
xnor U6801 (N_6801,N_6287,N_6483);
nand U6802 (N_6802,N_6253,N_6114);
nor U6803 (N_6803,N_6391,N_6370);
and U6804 (N_6804,N_6244,N_6312);
nor U6805 (N_6805,N_6307,N_6030);
and U6806 (N_6806,N_6181,N_6227);
and U6807 (N_6807,N_6374,N_6454);
and U6808 (N_6808,N_6443,N_6207);
and U6809 (N_6809,N_6427,N_6375);
nor U6810 (N_6810,N_6029,N_6056);
nand U6811 (N_6811,N_6274,N_6067);
and U6812 (N_6812,N_6468,N_6000);
nand U6813 (N_6813,N_6410,N_6281);
or U6814 (N_6814,N_6337,N_6133);
and U6815 (N_6815,N_6136,N_6120);
and U6816 (N_6816,N_6207,N_6277);
nor U6817 (N_6817,N_6139,N_6036);
or U6818 (N_6818,N_6180,N_6148);
nor U6819 (N_6819,N_6489,N_6154);
xnor U6820 (N_6820,N_6328,N_6431);
nand U6821 (N_6821,N_6061,N_6178);
or U6822 (N_6822,N_6198,N_6252);
nand U6823 (N_6823,N_6146,N_6141);
nor U6824 (N_6824,N_6476,N_6238);
and U6825 (N_6825,N_6294,N_6399);
nand U6826 (N_6826,N_6146,N_6462);
xor U6827 (N_6827,N_6135,N_6487);
or U6828 (N_6828,N_6196,N_6189);
and U6829 (N_6829,N_6409,N_6088);
and U6830 (N_6830,N_6039,N_6123);
nor U6831 (N_6831,N_6176,N_6455);
xor U6832 (N_6832,N_6318,N_6433);
and U6833 (N_6833,N_6112,N_6160);
and U6834 (N_6834,N_6332,N_6197);
nor U6835 (N_6835,N_6449,N_6262);
and U6836 (N_6836,N_6230,N_6346);
xnor U6837 (N_6837,N_6369,N_6113);
nor U6838 (N_6838,N_6424,N_6260);
xor U6839 (N_6839,N_6164,N_6459);
nor U6840 (N_6840,N_6223,N_6034);
nor U6841 (N_6841,N_6351,N_6156);
and U6842 (N_6842,N_6087,N_6058);
or U6843 (N_6843,N_6344,N_6431);
nand U6844 (N_6844,N_6198,N_6055);
xor U6845 (N_6845,N_6077,N_6412);
and U6846 (N_6846,N_6339,N_6037);
or U6847 (N_6847,N_6316,N_6139);
nor U6848 (N_6848,N_6426,N_6067);
and U6849 (N_6849,N_6290,N_6325);
and U6850 (N_6850,N_6436,N_6052);
xor U6851 (N_6851,N_6338,N_6263);
nor U6852 (N_6852,N_6112,N_6113);
nor U6853 (N_6853,N_6149,N_6093);
nor U6854 (N_6854,N_6477,N_6278);
nor U6855 (N_6855,N_6363,N_6340);
or U6856 (N_6856,N_6224,N_6237);
nand U6857 (N_6857,N_6433,N_6228);
xnor U6858 (N_6858,N_6459,N_6336);
xor U6859 (N_6859,N_6388,N_6099);
and U6860 (N_6860,N_6421,N_6039);
or U6861 (N_6861,N_6484,N_6493);
xnor U6862 (N_6862,N_6371,N_6069);
xor U6863 (N_6863,N_6061,N_6170);
xor U6864 (N_6864,N_6147,N_6212);
nor U6865 (N_6865,N_6002,N_6384);
xnor U6866 (N_6866,N_6161,N_6176);
and U6867 (N_6867,N_6329,N_6328);
xor U6868 (N_6868,N_6373,N_6034);
xor U6869 (N_6869,N_6209,N_6040);
nand U6870 (N_6870,N_6057,N_6236);
nand U6871 (N_6871,N_6154,N_6171);
nor U6872 (N_6872,N_6179,N_6350);
nand U6873 (N_6873,N_6116,N_6382);
xor U6874 (N_6874,N_6010,N_6311);
and U6875 (N_6875,N_6056,N_6274);
and U6876 (N_6876,N_6009,N_6189);
nand U6877 (N_6877,N_6228,N_6182);
xnor U6878 (N_6878,N_6212,N_6459);
nor U6879 (N_6879,N_6486,N_6351);
and U6880 (N_6880,N_6204,N_6383);
nand U6881 (N_6881,N_6030,N_6365);
xor U6882 (N_6882,N_6469,N_6120);
nor U6883 (N_6883,N_6359,N_6374);
nor U6884 (N_6884,N_6484,N_6199);
xnor U6885 (N_6885,N_6155,N_6052);
nand U6886 (N_6886,N_6170,N_6217);
nand U6887 (N_6887,N_6324,N_6425);
nand U6888 (N_6888,N_6251,N_6443);
nor U6889 (N_6889,N_6101,N_6497);
xor U6890 (N_6890,N_6325,N_6334);
and U6891 (N_6891,N_6185,N_6407);
or U6892 (N_6892,N_6455,N_6188);
or U6893 (N_6893,N_6118,N_6097);
or U6894 (N_6894,N_6148,N_6095);
or U6895 (N_6895,N_6363,N_6180);
nor U6896 (N_6896,N_6380,N_6367);
nand U6897 (N_6897,N_6236,N_6099);
and U6898 (N_6898,N_6244,N_6207);
xnor U6899 (N_6899,N_6331,N_6456);
xnor U6900 (N_6900,N_6255,N_6301);
nand U6901 (N_6901,N_6217,N_6230);
nand U6902 (N_6902,N_6188,N_6034);
or U6903 (N_6903,N_6330,N_6061);
and U6904 (N_6904,N_6424,N_6144);
nor U6905 (N_6905,N_6095,N_6490);
and U6906 (N_6906,N_6010,N_6181);
xnor U6907 (N_6907,N_6167,N_6123);
or U6908 (N_6908,N_6146,N_6089);
nor U6909 (N_6909,N_6359,N_6232);
or U6910 (N_6910,N_6360,N_6369);
and U6911 (N_6911,N_6432,N_6337);
nand U6912 (N_6912,N_6069,N_6402);
nand U6913 (N_6913,N_6474,N_6318);
and U6914 (N_6914,N_6055,N_6480);
xnor U6915 (N_6915,N_6157,N_6327);
and U6916 (N_6916,N_6023,N_6158);
or U6917 (N_6917,N_6449,N_6228);
nand U6918 (N_6918,N_6266,N_6213);
or U6919 (N_6919,N_6365,N_6420);
xor U6920 (N_6920,N_6241,N_6185);
and U6921 (N_6921,N_6338,N_6282);
nand U6922 (N_6922,N_6346,N_6232);
and U6923 (N_6923,N_6254,N_6466);
and U6924 (N_6924,N_6006,N_6201);
nand U6925 (N_6925,N_6088,N_6460);
nor U6926 (N_6926,N_6212,N_6456);
xnor U6927 (N_6927,N_6164,N_6096);
and U6928 (N_6928,N_6070,N_6081);
nor U6929 (N_6929,N_6101,N_6251);
or U6930 (N_6930,N_6313,N_6450);
xnor U6931 (N_6931,N_6281,N_6136);
xor U6932 (N_6932,N_6098,N_6030);
nand U6933 (N_6933,N_6352,N_6214);
and U6934 (N_6934,N_6062,N_6064);
nand U6935 (N_6935,N_6468,N_6084);
nand U6936 (N_6936,N_6417,N_6311);
and U6937 (N_6937,N_6174,N_6047);
nor U6938 (N_6938,N_6308,N_6219);
nand U6939 (N_6939,N_6383,N_6117);
or U6940 (N_6940,N_6345,N_6323);
nand U6941 (N_6941,N_6375,N_6279);
or U6942 (N_6942,N_6197,N_6375);
nor U6943 (N_6943,N_6463,N_6171);
nand U6944 (N_6944,N_6481,N_6424);
xnor U6945 (N_6945,N_6434,N_6242);
nand U6946 (N_6946,N_6314,N_6265);
xnor U6947 (N_6947,N_6239,N_6006);
and U6948 (N_6948,N_6329,N_6088);
nand U6949 (N_6949,N_6170,N_6228);
and U6950 (N_6950,N_6350,N_6445);
nand U6951 (N_6951,N_6282,N_6224);
or U6952 (N_6952,N_6305,N_6332);
and U6953 (N_6953,N_6043,N_6195);
nand U6954 (N_6954,N_6412,N_6460);
and U6955 (N_6955,N_6291,N_6029);
or U6956 (N_6956,N_6020,N_6390);
nor U6957 (N_6957,N_6232,N_6440);
nor U6958 (N_6958,N_6332,N_6139);
or U6959 (N_6959,N_6083,N_6185);
nor U6960 (N_6960,N_6116,N_6350);
xnor U6961 (N_6961,N_6110,N_6468);
nand U6962 (N_6962,N_6151,N_6021);
xor U6963 (N_6963,N_6398,N_6141);
nor U6964 (N_6964,N_6090,N_6164);
nand U6965 (N_6965,N_6161,N_6423);
xor U6966 (N_6966,N_6165,N_6367);
or U6967 (N_6967,N_6135,N_6275);
nor U6968 (N_6968,N_6051,N_6145);
xor U6969 (N_6969,N_6454,N_6045);
xnor U6970 (N_6970,N_6002,N_6051);
nor U6971 (N_6971,N_6446,N_6030);
nand U6972 (N_6972,N_6203,N_6005);
nand U6973 (N_6973,N_6326,N_6428);
or U6974 (N_6974,N_6416,N_6279);
xor U6975 (N_6975,N_6356,N_6428);
or U6976 (N_6976,N_6330,N_6316);
nor U6977 (N_6977,N_6355,N_6333);
nor U6978 (N_6978,N_6030,N_6326);
nor U6979 (N_6979,N_6298,N_6083);
nand U6980 (N_6980,N_6426,N_6469);
and U6981 (N_6981,N_6202,N_6249);
nand U6982 (N_6982,N_6188,N_6383);
or U6983 (N_6983,N_6326,N_6444);
nor U6984 (N_6984,N_6368,N_6186);
nand U6985 (N_6985,N_6427,N_6046);
xnor U6986 (N_6986,N_6132,N_6309);
nor U6987 (N_6987,N_6406,N_6109);
and U6988 (N_6988,N_6249,N_6476);
and U6989 (N_6989,N_6247,N_6277);
nor U6990 (N_6990,N_6321,N_6488);
and U6991 (N_6991,N_6084,N_6032);
nor U6992 (N_6992,N_6122,N_6374);
xnor U6993 (N_6993,N_6236,N_6148);
or U6994 (N_6994,N_6363,N_6318);
nor U6995 (N_6995,N_6258,N_6066);
and U6996 (N_6996,N_6288,N_6208);
or U6997 (N_6997,N_6062,N_6284);
nor U6998 (N_6998,N_6317,N_6050);
nor U6999 (N_6999,N_6315,N_6061);
nand U7000 (N_7000,N_6590,N_6752);
or U7001 (N_7001,N_6797,N_6878);
or U7002 (N_7002,N_6984,N_6769);
nand U7003 (N_7003,N_6598,N_6925);
nor U7004 (N_7004,N_6945,N_6975);
xor U7005 (N_7005,N_6504,N_6754);
or U7006 (N_7006,N_6978,N_6856);
nand U7007 (N_7007,N_6882,N_6720);
xnor U7008 (N_7008,N_6500,N_6879);
nor U7009 (N_7009,N_6520,N_6521);
nor U7010 (N_7010,N_6583,N_6656);
nand U7011 (N_7011,N_6963,N_6663);
and U7012 (N_7012,N_6540,N_6643);
xor U7013 (N_7013,N_6632,N_6671);
nand U7014 (N_7014,N_6582,N_6693);
and U7015 (N_7015,N_6696,N_6745);
or U7016 (N_7016,N_6743,N_6898);
or U7017 (N_7017,N_6639,N_6547);
nand U7018 (N_7018,N_6753,N_6832);
and U7019 (N_7019,N_6997,N_6516);
or U7020 (N_7020,N_6911,N_6537);
or U7021 (N_7021,N_6750,N_6608);
nor U7022 (N_7022,N_6541,N_6721);
or U7023 (N_7023,N_6679,N_6680);
xor U7024 (N_7024,N_6550,N_6712);
nand U7025 (N_7025,N_6788,N_6654);
and U7026 (N_7026,N_6615,N_6999);
or U7027 (N_7027,N_6606,N_6989);
nor U7028 (N_7028,N_6969,N_6722);
nand U7029 (N_7029,N_6888,N_6740);
nand U7030 (N_7030,N_6692,N_6585);
xnor U7031 (N_7031,N_6939,N_6518);
xnor U7032 (N_7032,N_6938,N_6528);
or U7033 (N_7033,N_6777,N_6869);
xor U7034 (N_7034,N_6770,N_6662);
nand U7035 (N_7035,N_6886,N_6688);
nor U7036 (N_7036,N_6717,N_6725);
and U7037 (N_7037,N_6954,N_6936);
or U7038 (N_7038,N_6628,N_6804);
and U7039 (N_7039,N_6714,N_6655);
xnor U7040 (N_7040,N_6806,N_6915);
and U7041 (N_7041,N_6588,N_6556);
and U7042 (N_7042,N_6928,N_6567);
nand U7043 (N_7043,N_6814,N_6649);
nand U7044 (N_7044,N_6600,N_6668);
nor U7045 (N_7045,N_6953,N_6546);
nand U7046 (N_7046,N_6914,N_6811);
xor U7047 (N_7047,N_6695,N_6626);
nor U7048 (N_7048,N_6799,N_6738);
xnor U7049 (N_7049,N_6858,N_6774);
xor U7050 (N_7050,N_6545,N_6605);
xor U7051 (N_7051,N_6783,N_6706);
and U7052 (N_7052,N_6872,N_6973);
xor U7053 (N_7053,N_6621,N_6789);
xnor U7054 (N_7054,N_6943,N_6507);
nor U7055 (N_7055,N_6813,N_6843);
xnor U7056 (N_7056,N_6702,N_6673);
and U7057 (N_7057,N_6609,N_6839);
xor U7058 (N_7058,N_6847,N_6990);
nand U7059 (N_7059,N_6617,N_6559);
and U7060 (N_7060,N_6798,N_6986);
xor U7061 (N_7061,N_6652,N_6513);
or U7062 (N_7062,N_6890,N_6514);
or U7063 (N_7063,N_6708,N_6509);
nor U7064 (N_7064,N_6996,N_6601);
nor U7065 (N_7065,N_6909,N_6863);
or U7066 (N_7066,N_6751,N_6635);
xor U7067 (N_7067,N_6711,N_6565);
or U7068 (N_7068,N_6530,N_6836);
and U7069 (N_7069,N_6912,N_6658);
nor U7070 (N_7070,N_6759,N_6553);
xnor U7071 (N_7071,N_6794,N_6737);
or U7072 (N_7072,N_6848,N_6744);
nor U7073 (N_7073,N_6616,N_6803);
or U7074 (N_7074,N_6614,N_6694);
and U7075 (N_7075,N_6849,N_6758);
and U7076 (N_7076,N_6795,N_6913);
xnor U7077 (N_7077,N_6883,N_6991);
nor U7078 (N_7078,N_6979,N_6646);
or U7079 (N_7079,N_6723,N_6503);
or U7080 (N_7080,N_6589,N_6968);
and U7081 (N_7081,N_6768,N_6526);
xnor U7082 (N_7082,N_6833,N_6860);
nand U7083 (N_7083,N_6709,N_6866);
nand U7084 (N_7084,N_6665,N_6531);
nand U7085 (N_7085,N_6841,N_6964);
or U7086 (N_7086,N_6884,N_6596);
xnor U7087 (N_7087,N_6876,N_6602);
or U7088 (N_7088,N_6701,N_6767);
xor U7089 (N_7089,N_6527,N_6718);
or U7090 (N_7090,N_6785,N_6577);
nand U7091 (N_7091,N_6987,N_6641);
nor U7092 (N_7092,N_6746,N_6942);
xnor U7093 (N_7093,N_6930,N_6686);
or U7094 (N_7094,N_6620,N_6874);
or U7095 (N_7095,N_6733,N_6892);
and U7096 (N_7096,N_6624,N_6690);
nand U7097 (N_7097,N_6682,N_6881);
nor U7098 (N_7098,N_6897,N_6908);
or U7099 (N_7099,N_6985,N_6837);
and U7100 (N_7100,N_6724,N_6793);
and U7101 (N_7101,N_6956,N_6960);
nor U7102 (N_7102,N_6887,N_6916);
nand U7103 (N_7103,N_6926,N_6967);
nand U7104 (N_7104,N_6691,N_6749);
and U7105 (N_7105,N_6716,N_6631);
nand U7106 (N_7106,N_6684,N_6747);
or U7107 (N_7107,N_6861,N_6851);
or U7108 (N_7108,N_6757,N_6659);
or U7109 (N_7109,N_6773,N_6675);
xor U7110 (N_7110,N_6742,N_6780);
xnor U7111 (N_7111,N_6625,N_6638);
nor U7112 (N_7112,N_6604,N_6670);
or U7113 (N_7113,N_6927,N_6959);
or U7114 (N_7114,N_6561,N_6707);
nand U7115 (N_7115,N_6900,N_6756);
nor U7116 (N_7116,N_6735,N_6533);
and U7117 (N_7117,N_6816,N_6891);
xnor U7118 (N_7118,N_6579,N_6636);
nand U7119 (N_7119,N_6937,N_6760);
nor U7120 (N_7120,N_6957,N_6506);
nor U7121 (N_7121,N_6958,N_6918);
xor U7122 (N_7122,N_6845,N_6512);
nand U7123 (N_7123,N_6554,N_6895);
nand U7124 (N_7124,N_6787,N_6569);
nand U7125 (N_7125,N_6681,N_6705);
nand U7126 (N_7126,N_6764,N_6988);
and U7127 (N_7127,N_6940,N_6840);
nor U7128 (N_7128,N_6505,N_6970);
nor U7129 (N_7129,N_6877,N_6657);
xnor U7130 (N_7130,N_6563,N_6552);
and U7131 (N_7131,N_6854,N_6575);
nand U7132 (N_7132,N_6834,N_6573);
nand U7133 (N_7133,N_6919,N_6697);
or U7134 (N_7134,N_6801,N_6594);
xnor U7135 (N_7135,N_6951,N_6805);
or U7136 (N_7136,N_6782,N_6525);
or U7137 (N_7137,N_6995,N_6826);
nor U7138 (N_7138,N_6762,N_6634);
nand U7139 (N_7139,N_6775,N_6972);
and U7140 (N_7140,N_6593,N_6700);
and U7141 (N_7141,N_6535,N_6522);
and U7142 (N_7142,N_6824,N_6835);
nand U7143 (N_7143,N_6727,N_6906);
or U7144 (N_7144,N_6728,N_6946);
nor U7145 (N_7145,N_6935,N_6555);
nand U7146 (N_7146,N_6574,N_6544);
nor U7147 (N_7147,N_6532,N_6651);
or U7148 (N_7148,N_6704,N_6664);
nor U7149 (N_7149,N_6580,N_6611);
nor U7150 (N_7150,N_6977,N_6821);
and U7151 (N_7151,N_6903,N_6548);
xnor U7152 (N_7152,N_6570,N_6812);
nor U7153 (N_7153,N_6944,N_6729);
xor U7154 (N_7154,N_6618,N_6992);
nor U7155 (N_7155,N_6901,N_6599);
and U7156 (N_7156,N_6807,N_6699);
nor U7157 (N_7157,N_6976,N_6962);
and U7158 (N_7158,N_6543,N_6713);
and U7159 (N_7159,N_6850,N_6980);
or U7160 (N_7160,N_6633,N_6873);
nand U7161 (N_7161,N_6560,N_6647);
and U7162 (N_7162,N_6676,N_6660);
or U7163 (N_7163,N_6581,N_6859);
nor U7164 (N_7164,N_6678,N_6784);
or U7165 (N_7165,N_6934,N_6831);
nand U7166 (N_7166,N_6862,N_6549);
nand U7167 (N_7167,N_6644,N_6519);
nor U7168 (N_7168,N_6674,N_6542);
or U7169 (N_7169,N_6687,N_6571);
xnor U7170 (N_7170,N_6640,N_6653);
and U7171 (N_7171,N_6515,N_6523);
and U7172 (N_7172,N_6661,N_6949);
xnor U7173 (N_7173,N_6994,N_6648);
nand U7174 (N_7174,N_6855,N_6904);
and U7175 (N_7175,N_6689,N_6623);
xnor U7176 (N_7176,N_6981,N_6965);
xor U7177 (N_7177,N_6779,N_6572);
or U7178 (N_7178,N_6867,N_6677);
or U7179 (N_7179,N_6823,N_6667);
nand U7180 (N_7180,N_6741,N_6922);
xor U7181 (N_7181,N_6776,N_6950);
and U7182 (N_7182,N_6905,N_6539);
nor U7183 (N_7183,N_6961,N_6810);
xor U7184 (N_7184,N_6966,N_6932);
nand U7185 (N_7185,N_6917,N_6853);
xor U7186 (N_7186,N_6685,N_6819);
nor U7187 (N_7187,N_6672,N_6838);
xor U7188 (N_7188,N_6993,N_6586);
xor U7189 (N_7189,N_6587,N_6698);
nor U7190 (N_7190,N_6578,N_6766);
xnor U7191 (N_7191,N_6731,N_6511);
or U7192 (N_7192,N_6846,N_6557);
xor U7193 (N_7193,N_6790,N_6924);
or U7194 (N_7194,N_6558,N_6896);
and U7195 (N_7195,N_6645,N_6510);
nand U7196 (N_7196,N_6844,N_6865);
or U7197 (N_7197,N_6864,N_6899);
and U7198 (N_7198,N_6564,N_6734);
nor U7199 (N_7199,N_6827,N_6683);
nor U7200 (N_7200,N_6726,N_6818);
nor U7201 (N_7201,N_6591,N_6948);
or U7202 (N_7202,N_6982,N_6893);
nor U7203 (N_7203,N_6830,N_6719);
nor U7204 (N_7204,N_6894,N_6748);
and U7205 (N_7205,N_6947,N_6730);
or U7206 (N_7206,N_6820,N_6931);
or U7207 (N_7207,N_6971,N_6871);
nor U7208 (N_7208,N_6815,N_6627);
and U7209 (N_7209,N_6666,N_6595);
or U7210 (N_7210,N_6923,N_6796);
nor U7211 (N_7211,N_6902,N_6629);
or U7212 (N_7212,N_6929,N_6584);
xor U7213 (N_7213,N_6857,N_6619);
and U7214 (N_7214,N_6603,N_6524);
and U7215 (N_7215,N_6755,N_6610);
or U7216 (N_7216,N_6808,N_6817);
nand U7217 (N_7217,N_6889,N_6669);
and U7218 (N_7218,N_6763,N_6568);
or U7219 (N_7219,N_6800,N_6612);
and U7220 (N_7220,N_6566,N_6974);
xnor U7221 (N_7221,N_6809,N_6842);
nand U7222 (N_7222,N_6642,N_6715);
xnor U7223 (N_7223,N_6517,N_6870);
or U7224 (N_7224,N_6822,N_6761);
xor U7225 (N_7225,N_6739,N_6952);
or U7226 (N_7226,N_6825,N_6732);
xor U7227 (N_7227,N_6921,N_6534);
nor U7228 (N_7228,N_6786,N_6650);
nor U7229 (N_7229,N_6529,N_6792);
or U7230 (N_7230,N_6910,N_6765);
nor U7231 (N_7231,N_6562,N_6868);
nor U7232 (N_7232,N_6933,N_6983);
or U7233 (N_7233,N_6791,N_6501);
nor U7234 (N_7234,N_6781,N_6630);
and U7235 (N_7235,N_6955,N_6736);
nor U7236 (N_7236,N_6885,N_6597);
or U7237 (N_7237,N_6907,N_6613);
xnor U7238 (N_7238,N_6508,N_6875);
nor U7239 (N_7239,N_6880,N_6941);
nand U7240 (N_7240,N_6551,N_6778);
xnor U7241 (N_7241,N_6772,N_6852);
xnor U7242 (N_7242,N_6920,N_6536);
nor U7243 (N_7243,N_6622,N_6802);
xnor U7244 (N_7244,N_6998,N_6538);
and U7245 (N_7245,N_6828,N_6502);
nor U7246 (N_7246,N_6771,N_6607);
xnor U7247 (N_7247,N_6829,N_6703);
nand U7248 (N_7248,N_6576,N_6592);
and U7249 (N_7249,N_6637,N_6710);
xnor U7250 (N_7250,N_6703,N_6579);
nor U7251 (N_7251,N_6858,N_6660);
nor U7252 (N_7252,N_6629,N_6630);
or U7253 (N_7253,N_6527,N_6940);
or U7254 (N_7254,N_6887,N_6520);
xnor U7255 (N_7255,N_6615,N_6873);
nor U7256 (N_7256,N_6524,N_6501);
nor U7257 (N_7257,N_6520,N_6519);
and U7258 (N_7258,N_6500,N_6786);
nor U7259 (N_7259,N_6729,N_6994);
nand U7260 (N_7260,N_6702,N_6854);
and U7261 (N_7261,N_6954,N_6719);
nor U7262 (N_7262,N_6811,N_6745);
xor U7263 (N_7263,N_6860,N_6609);
xnor U7264 (N_7264,N_6513,N_6603);
xnor U7265 (N_7265,N_6912,N_6852);
nor U7266 (N_7266,N_6857,N_6607);
xor U7267 (N_7267,N_6923,N_6843);
xor U7268 (N_7268,N_6888,N_6787);
nand U7269 (N_7269,N_6503,N_6527);
and U7270 (N_7270,N_6506,N_6657);
nor U7271 (N_7271,N_6919,N_6807);
and U7272 (N_7272,N_6962,N_6605);
nor U7273 (N_7273,N_6851,N_6680);
nor U7274 (N_7274,N_6811,N_6754);
nor U7275 (N_7275,N_6845,N_6791);
nor U7276 (N_7276,N_6657,N_6704);
nand U7277 (N_7277,N_6635,N_6726);
and U7278 (N_7278,N_6565,N_6615);
nand U7279 (N_7279,N_6575,N_6568);
or U7280 (N_7280,N_6827,N_6925);
nor U7281 (N_7281,N_6649,N_6907);
xor U7282 (N_7282,N_6863,N_6752);
nand U7283 (N_7283,N_6634,N_6722);
xor U7284 (N_7284,N_6995,N_6980);
nand U7285 (N_7285,N_6963,N_6919);
xnor U7286 (N_7286,N_6778,N_6598);
nor U7287 (N_7287,N_6999,N_6806);
nand U7288 (N_7288,N_6931,N_6610);
xnor U7289 (N_7289,N_6772,N_6888);
xnor U7290 (N_7290,N_6737,N_6988);
and U7291 (N_7291,N_6937,N_6790);
nor U7292 (N_7292,N_6540,N_6661);
and U7293 (N_7293,N_6707,N_6510);
or U7294 (N_7294,N_6806,N_6538);
xor U7295 (N_7295,N_6735,N_6929);
xnor U7296 (N_7296,N_6522,N_6926);
and U7297 (N_7297,N_6801,N_6699);
nor U7298 (N_7298,N_6778,N_6668);
xor U7299 (N_7299,N_6862,N_6900);
nand U7300 (N_7300,N_6508,N_6822);
nor U7301 (N_7301,N_6752,N_6882);
xor U7302 (N_7302,N_6920,N_6986);
and U7303 (N_7303,N_6827,N_6679);
and U7304 (N_7304,N_6670,N_6852);
xor U7305 (N_7305,N_6974,N_6587);
nor U7306 (N_7306,N_6731,N_6778);
or U7307 (N_7307,N_6866,N_6947);
nand U7308 (N_7308,N_6599,N_6820);
nor U7309 (N_7309,N_6669,N_6928);
and U7310 (N_7310,N_6652,N_6731);
xnor U7311 (N_7311,N_6889,N_6534);
or U7312 (N_7312,N_6587,N_6731);
or U7313 (N_7313,N_6677,N_6563);
xnor U7314 (N_7314,N_6548,N_6858);
or U7315 (N_7315,N_6709,N_6892);
and U7316 (N_7316,N_6685,N_6666);
nor U7317 (N_7317,N_6567,N_6626);
and U7318 (N_7318,N_6635,N_6844);
and U7319 (N_7319,N_6826,N_6978);
or U7320 (N_7320,N_6964,N_6756);
and U7321 (N_7321,N_6617,N_6744);
xnor U7322 (N_7322,N_6822,N_6631);
nor U7323 (N_7323,N_6817,N_6527);
xnor U7324 (N_7324,N_6641,N_6928);
nor U7325 (N_7325,N_6961,N_6787);
nand U7326 (N_7326,N_6755,N_6740);
nor U7327 (N_7327,N_6641,N_6855);
nor U7328 (N_7328,N_6744,N_6904);
and U7329 (N_7329,N_6982,N_6634);
and U7330 (N_7330,N_6927,N_6706);
nand U7331 (N_7331,N_6949,N_6887);
nor U7332 (N_7332,N_6903,N_6940);
nand U7333 (N_7333,N_6926,N_6700);
xor U7334 (N_7334,N_6661,N_6807);
or U7335 (N_7335,N_6674,N_6706);
and U7336 (N_7336,N_6521,N_6817);
xnor U7337 (N_7337,N_6799,N_6923);
xor U7338 (N_7338,N_6906,N_6776);
nand U7339 (N_7339,N_6922,N_6944);
nor U7340 (N_7340,N_6976,N_6959);
xor U7341 (N_7341,N_6989,N_6880);
nor U7342 (N_7342,N_6835,N_6686);
nor U7343 (N_7343,N_6889,N_6576);
and U7344 (N_7344,N_6999,N_6586);
xnor U7345 (N_7345,N_6664,N_6641);
and U7346 (N_7346,N_6520,N_6547);
or U7347 (N_7347,N_6544,N_6529);
nor U7348 (N_7348,N_6778,N_6511);
nor U7349 (N_7349,N_6541,N_6636);
or U7350 (N_7350,N_6643,N_6982);
and U7351 (N_7351,N_6514,N_6581);
xor U7352 (N_7352,N_6804,N_6884);
or U7353 (N_7353,N_6740,N_6973);
nand U7354 (N_7354,N_6635,N_6578);
nand U7355 (N_7355,N_6802,N_6862);
and U7356 (N_7356,N_6636,N_6892);
nand U7357 (N_7357,N_6517,N_6502);
and U7358 (N_7358,N_6583,N_6965);
or U7359 (N_7359,N_6881,N_6546);
xor U7360 (N_7360,N_6720,N_6561);
nor U7361 (N_7361,N_6938,N_6592);
or U7362 (N_7362,N_6963,N_6774);
and U7363 (N_7363,N_6510,N_6970);
and U7364 (N_7364,N_6766,N_6538);
xnor U7365 (N_7365,N_6697,N_6849);
nor U7366 (N_7366,N_6505,N_6691);
xnor U7367 (N_7367,N_6722,N_6845);
and U7368 (N_7368,N_6800,N_6758);
nor U7369 (N_7369,N_6506,N_6940);
and U7370 (N_7370,N_6521,N_6778);
nor U7371 (N_7371,N_6883,N_6652);
xor U7372 (N_7372,N_6509,N_6535);
or U7373 (N_7373,N_6623,N_6654);
nor U7374 (N_7374,N_6950,N_6676);
and U7375 (N_7375,N_6559,N_6882);
nor U7376 (N_7376,N_6935,N_6506);
or U7377 (N_7377,N_6615,N_6715);
or U7378 (N_7378,N_6609,N_6660);
nor U7379 (N_7379,N_6692,N_6516);
nand U7380 (N_7380,N_6780,N_6675);
or U7381 (N_7381,N_6855,N_6871);
or U7382 (N_7382,N_6665,N_6999);
xnor U7383 (N_7383,N_6980,N_6506);
and U7384 (N_7384,N_6695,N_6936);
or U7385 (N_7385,N_6645,N_6891);
xor U7386 (N_7386,N_6915,N_6770);
nand U7387 (N_7387,N_6649,N_6981);
and U7388 (N_7388,N_6661,N_6795);
xnor U7389 (N_7389,N_6770,N_6842);
nor U7390 (N_7390,N_6814,N_6607);
nor U7391 (N_7391,N_6803,N_6916);
nand U7392 (N_7392,N_6585,N_6529);
xor U7393 (N_7393,N_6961,N_6698);
nand U7394 (N_7394,N_6545,N_6767);
nand U7395 (N_7395,N_6653,N_6625);
or U7396 (N_7396,N_6718,N_6557);
and U7397 (N_7397,N_6956,N_6647);
nor U7398 (N_7398,N_6538,N_6713);
nand U7399 (N_7399,N_6720,N_6687);
nand U7400 (N_7400,N_6716,N_6950);
and U7401 (N_7401,N_6737,N_6609);
and U7402 (N_7402,N_6835,N_6831);
nand U7403 (N_7403,N_6885,N_6930);
and U7404 (N_7404,N_6986,N_6801);
nand U7405 (N_7405,N_6881,N_6551);
or U7406 (N_7406,N_6592,N_6522);
and U7407 (N_7407,N_6695,N_6840);
nor U7408 (N_7408,N_6958,N_6536);
nor U7409 (N_7409,N_6926,N_6643);
and U7410 (N_7410,N_6935,N_6676);
xnor U7411 (N_7411,N_6743,N_6833);
nor U7412 (N_7412,N_6625,N_6529);
nor U7413 (N_7413,N_6763,N_6944);
nor U7414 (N_7414,N_6842,N_6704);
nand U7415 (N_7415,N_6625,N_6612);
xor U7416 (N_7416,N_6743,N_6716);
and U7417 (N_7417,N_6674,N_6991);
or U7418 (N_7418,N_6881,N_6951);
or U7419 (N_7419,N_6539,N_6915);
xnor U7420 (N_7420,N_6849,N_6824);
nand U7421 (N_7421,N_6851,N_6528);
or U7422 (N_7422,N_6784,N_6916);
nor U7423 (N_7423,N_6748,N_6684);
or U7424 (N_7424,N_6652,N_6643);
nor U7425 (N_7425,N_6930,N_6692);
xor U7426 (N_7426,N_6501,N_6590);
or U7427 (N_7427,N_6607,N_6533);
nand U7428 (N_7428,N_6873,N_6789);
xor U7429 (N_7429,N_6751,N_6603);
xor U7430 (N_7430,N_6625,N_6814);
or U7431 (N_7431,N_6709,N_6795);
nor U7432 (N_7432,N_6861,N_6784);
nand U7433 (N_7433,N_6867,N_6726);
or U7434 (N_7434,N_6734,N_6589);
xor U7435 (N_7435,N_6678,N_6555);
nand U7436 (N_7436,N_6634,N_6847);
and U7437 (N_7437,N_6754,N_6501);
nand U7438 (N_7438,N_6868,N_6818);
nor U7439 (N_7439,N_6929,N_6586);
or U7440 (N_7440,N_6619,N_6801);
nor U7441 (N_7441,N_6633,N_6884);
xnor U7442 (N_7442,N_6962,N_6506);
and U7443 (N_7443,N_6616,N_6744);
xnor U7444 (N_7444,N_6540,N_6610);
nor U7445 (N_7445,N_6706,N_6617);
nand U7446 (N_7446,N_6872,N_6592);
or U7447 (N_7447,N_6528,N_6767);
nand U7448 (N_7448,N_6927,N_6685);
nand U7449 (N_7449,N_6723,N_6677);
nand U7450 (N_7450,N_6704,N_6917);
xnor U7451 (N_7451,N_6743,N_6792);
or U7452 (N_7452,N_6757,N_6992);
nand U7453 (N_7453,N_6833,N_6694);
nor U7454 (N_7454,N_6661,N_6658);
xor U7455 (N_7455,N_6522,N_6814);
and U7456 (N_7456,N_6775,N_6922);
and U7457 (N_7457,N_6721,N_6997);
and U7458 (N_7458,N_6574,N_6834);
xor U7459 (N_7459,N_6941,N_6804);
xor U7460 (N_7460,N_6549,N_6787);
nor U7461 (N_7461,N_6539,N_6947);
or U7462 (N_7462,N_6567,N_6801);
nand U7463 (N_7463,N_6882,N_6543);
and U7464 (N_7464,N_6853,N_6957);
nor U7465 (N_7465,N_6535,N_6900);
or U7466 (N_7466,N_6612,N_6596);
xnor U7467 (N_7467,N_6986,N_6961);
or U7468 (N_7468,N_6875,N_6978);
nand U7469 (N_7469,N_6654,N_6926);
xor U7470 (N_7470,N_6698,N_6518);
nor U7471 (N_7471,N_6973,N_6999);
nand U7472 (N_7472,N_6847,N_6583);
or U7473 (N_7473,N_6879,N_6555);
nand U7474 (N_7474,N_6584,N_6821);
nor U7475 (N_7475,N_6651,N_6503);
or U7476 (N_7476,N_6797,N_6580);
or U7477 (N_7477,N_6747,N_6965);
or U7478 (N_7478,N_6547,N_6665);
and U7479 (N_7479,N_6933,N_6988);
nor U7480 (N_7480,N_6537,N_6966);
xnor U7481 (N_7481,N_6929,N_6731);
and U7482 (N_7482,N_6744,N_6725);
nand U7483 (N_7483,N_6890,N_6545);
nand U7484 (N_7484,N_6634,N_6975);
nor U7485 (N_7485,N_6958,N_6966);
nor U7486 (N_7486,N_6713,N_6525);
and U7487 (N_7487,N_6823,N_6822);
xor U7488 (N_7488,N_6575,N_6526);
xor U7489 (N_7489,N_6922,N_6744);
and U7490 (N_7490,N_6742,N_6681);
or U7491 (N_7491,N_6691,N_6989);
or U7492 (N_7492,N_6741,N_6718);
nand U7493 (N_7493,N_6840,N_6982);
xnor U7494 (N_7494,N_6617,N_6511);
nor U7495 (N_7495,N_6845,N_6837);
or U7496 (N_7496,N_6898,N_6870);
nand U7497 (N_7497,N_6507,N_6531);
nand U7498 (N_7498,N_6704,N_6695);
xnor U7499 (N_7499,N_6806,N_6642);
or U7500 (N_7500,N_7241,N_7191);
nor U7501 (N_7501,N_7473,N_7278);
nor U7502 (N_7502,N_7470,N_7378);
or U7503 (N_7503,N_7367,N_7067);
or U7504 (N_7504,N_7076,N_7031);
nand U7505 (N_7505,N_7298,N_7214);
xnor U7506 (N_7506,N_7426,N_7442);
nand U7507 (N_7507,N_7102,N_7326);
and U7508 (N_7508,N_7487,N_7145);
and U7509 (N_7509,N_7055,N_7292);
nor U7510 (N_7510,N_7228,N_7119);
xor U7511 (N_7511,N_7484,N_7064);
nand U7512 (N_7512,N_7182,N_7094);
nor U7513 (N_7513,N_7331,N_7411);
nor U7514 (N_7514,N_7423,N_7417);
or U7515 (N_7515,N_7015,N_7133);
nor U7516 (N_7516,N_7143,N_7202);
and U7517 (N_7517,N_7343,N_7208);
or U7518 (N_7518,N_7234,N_7203);
xnor U7519 (N_7519,N_7497,N_7270);
xnor U7520 (N_7520,N_7020,N_7335);
and U7521 (N_7521,N_7181,N_7400);
nand U7522 (N_7522,N_7163,N_7036);
or U7523 (N_7523,N_7482,N_7025);
and U7524 (N_7524,N_7238,N_7457);
and U7525 (N_7525,N_7110,N_7434);
and U7526 (N_7526,N_7200,N_7466);
or U7527 (N_7527,N_7138,N_7256);
nor U7528 (N_7528,N_7439,N_7491);
nor U7529 (N_7529,N_7149,N_7364);
nor U7530 (N_7530,N_7391,N_7167);
nor U7531 (N_7531,N_7140,N_7130);
or U7532 (N_7532,N_7296,N_7082);
nor U7533 (N_7533,N_7425,N_7356);
xnor U7534 (N_7534,N_7271,N_7369);
nor U7535 (N_7535,N_7481,N_7247);
and U7536 (N_7536,N_7339,N_7101);
nor U7537 (N_7537,N_7150,N_7061);
nand U7538 (N_7538,N_7360,N_7069);
xnor U7539 (N_7539,N_7489,N_7363);
xor U7540 (N_7540,N_7332,N_7000);
xnor U7541 (N_7541,N_7173,N_7037);
xnor U7542 (N_7542,N_7250,N_7257);
nand U7543 (N_7543,N_7154,N_7348);
or U7544 (N_7544,N_7449,N_7035);
and U7545 (N_7545,N_7223,N_7351);
or U7546 (N_7546,N_7224,N_7258);
nand U7547 (N_7547,N_7229,N_7019);
nor U7548 (N_7548,N_7324,N_7353);
or U7549 (N_7549,N_7317,N_7003);
xor U7550 (N_7550,N_7006,N_7329);
or U7551 (N_7551,N_7413,N_7265);
and U7552 (N_7552,N_7105,N_7476);
and U7553 (N_7553,N_7153,N_7245);
and U7554 (N_7554,N_7085,N_7034);
nand U7555 (N_7555,N_7168,N_7472);
xnor U7556 (N_7556,N_7027,N_7050);
nor U7557 (N_7557,N_7295,N_7211);
xor U7558 (N_7558,N_7029,N_7284);
or U7559 (N_7559,N_7416,N_7079);
and U7560 (N_7560,N_7393,N_7325);
nand U7561 (N_7561,N_7017,N_7040);
nor U7562 (N_7562,N_7045,N_7291);
or U7563 (N_7563,N_7398,N_7249);
nand U7564 (N_7564,N_7465,N_7243);
nor U7565 (N_7565,N_7454,N_7212);
nor U7566 (N_7566,N_7300,N_7078);
or U7567 (N_7567,N_7347,N_7240);
nor U7568 (N_7568,N_7118,N_7207);
nor U7569 (N_7569,N_7009,N_7396);
nand U7570 (N_7570,N_7023,N_7408);
and U7571 (N_7571,N_7113,N_7178);
nor U7572 (N_7572,N_7436,N_7221);
nand U7573 (N_7573,N_7308,N_7059);
nor U7574 (N_7574,N_7225,N_7390);
nand U7575 (N_7575,N_7022,N_7362);
xor U7576 (N_7576,N_7453,N_7340);
xnor U7577 (N_7577,N_7299,N_7451);
xnor U7578 (N_7578,N_7410,N_7230);
and U7579 (N_7579,N_7456,N_7267);
nand U7580 (N_7580,N_7441,N_7498);
nand U7581 (N_7581,N_7169,N_7345);
nand U7582 (N_7582,N_7137,N_7049);
nor U7583 (N_7583,N_7205,N_7021);
nand U7584 (N_7584,N_7060,N_7054);
xor U7585 (N_7585,N_7183,N_7158);
xnor U7586 (N_7586,N_7496,N_7337);
and U7587 (N_7587,N_7114,N_7260);
nand U7588 (N_7588,N_7159,N_7316);
or U7589 (N_7589,N_7122,N_7013);
nand U7590 (N_7590,N_7033,N_7002);
and U7591 (N_7591,N_7379,N_7170);
nor U7592 (N_7592,N_7071,N_7446);
xor U7593 (N_7593,N_7327,N_7084);
and U7594 (N_7594,N_7272,N_7172);
xnor U7595 (N_7595,N_7231,N_7438);
xnor U7596 (N_7596,N_7310,N_7262);
nand U7597 (N_7597,N_7192,N_7461);
nor U7598 (N_7598,N_7160,N_7415);
nand U7599 (N_7599,N_7458,N_7232);
or U7600 (N_7600,N_7171,N_7459);
nand U7601 (N_7601,N_7155,N_7039);
nand U7602 (N_7602,N_7279,N_7198);
xor U7603 (N_7603,N_7239,N_7407);
and U7604 (N_7604,N_7406,N_7385);
xor U7605 (N_7605,N_7199,N_7201);
xor U7606 (N_7606,N_7273,N_7443);
nor U7607 (N_7607,N_7156,N_7072);
nand U7608 (N_7608,N_7188,N_7342);
nor U7609 (N_7609,N_7103,N_7264);
or U7610 (N_7610,N_7433,N_7414);
or U7611 (N_7611,N_7179,N_7285);
and U7612 (N_7612,N_7321,N_7405);
nor U7613 (N_7613,N_7399,N_7334);
or U7614 (N_7614,N_7125,N_7161);
and U7615 (N_7615,N_7280,N_7185);
or U7616 (N_7616,N_7366,N_7128);
nand U7617 (N_7617,N_7246,N_7121);
nand U7618 (N_7618,N_7124,N_7100);
nand U7619 (N_7619,N_7237,N_7336);
nand U7620 (N_7620,N_7311,N_7215);
xnor U7621 (N_7621,N_7194,N_7307);
nand U7622 (N_7622,N_7255,N_7152);
xor U7623 (N_7623,N_7297,N_7089);
or U7624 (N_7624,N_7139,N_7395);
nor U7625 (N_7625,N_7252,N_7314);
and U7626 (N_7626,N_7112,N_7402);
xnor U7627 (N_7627,N_7312,N_7359);
nand U7628 (N_7628,N_7219,N_7431);
nor U7629 (N_7629,N_7404,N_7287);
nor U7630 (N_7630,N_7403,N_7065);
nor U7631 (N_7631,N_7261,N_7432);
or U7632 (N_7632,N_7127,N_7204);
or U7633 (N_7633,N_7350,N_7422);
or U7634 (N_7634,N_7490,N_7471);
or U7635 (N_7635,N_7095,N_7355);
xor U7636 (N_7636,N_7032,N_7141);
nand U7637 (N_7637,N_7077,N_7098);
xnor U7638 (N_7638,N_7075,N_7104);
or U7639 (N_7639,N_7135,N_7445);
and U7640 (N_7640,N_7401,N_7372);
xor U7641 (N_7641,N_7387,N_7376);
or U7642 (N_7642,N_7444,N_7389);
or U7643 (N_7643,N_7242,N_7365);
nand U7644 (N_7644,N_7233,N_7305);
nand U7645 (N_7645,N_7475,N_7357);
or U7646 (N_7646,N_7375,N_7217);
or U7647 (N_7647,N_7001,N_7437);
and U7648 (N_7648,N_7056,N_7419);
and U7649 (N_7649,N_7197,N_7288);
nor U7650 (N_7650,N_7485,N_7302);
xnor U7651 (N_7651,N_7136,N_7048);
xnor U7652 (N_7652,N_7097,N_7480);
nor U7653 (N_7653,N_7107,N_7106);
nor U7654 (N_7654,N_7165,N_7176);
and U7655 (N_7655,N_7309,N_7189);
xnor U7656 (N_7656,N_7010,N_7290);
xnor U7657 (N_7657,N_7266,N_7397);
nand U7658 (N_7658,N_7477,N_7174);
nor U7659 (N_7659,N_7304,N_7109);
nand U7660 (N_7660,N_7129,N_7184);
and U7661 (N_7661,N_7455,N_7384);
and U7662 (N_7662,N_7358,N_7062);
or U7663 (N_7663,N_7263,N_7248);
xor U7664 (N_7664,N_7051,N_7142);
and U7665 (N_7665,N_7004,N_7134);
xnor U7666 (N_7666,N_7320,N_7361);
nand U7667 (N_7667,N_7282,N_7474);
nand U7668 (N_7668,N_7117,N_7464);
xor U7669 (N_7669,N_7467,N_7042);
and U7670 (N_7670,N_7463,N_7452);
or U7671 (N_7671,N_7486,N_7063);
xnor U7672 (N_7672,N_7052,N_7175);
nor U7673 (N_7673,N_7016,N_7053);
nor U7674 (N_7674,N_7083,N_7014);
nand U7675 (N_7675,N_7421,N_7483);
xnor U7676 (N_7676,N_7303,N_7274);
nand U7677 (N_7677,N_7058,N_7008);
nor U7678 (N_7678,N_7381,N_7333);
nor U7679 (N_7679,N_7044,N_7494);
nand U7680 (N_7680,N_7392,N_7218);
or U7681 (N_7681,N_7478,N_7253);
nand U7682 (N_7682,N_7328,N_7126);
nand U7683 (N_7683,N_7057,N_7306);
or U7684 (N_7684,N_7047,N_7386);
and U7685 (N_7685,N_7227,N_7440);
or U7686 (N_7686,N_7499,N_7388);
and U7687 (N_7687,N_7024,N_7157);
and U7688 (N_7688,N_7373,N_7216);
nand U7689 (N_7689,N_7070,N_7206);
nor U7690 (N_7690,N_7090,N_7382);
xor U7691 (N_7691,N_7315,N_7092);
xor U7692 (N_7692,N_7294,N_7151);
and U7693 (N_7693,N_7074,N_7226);
and U7694 (N_7694,N_7322,N_7283);
xnor U7695 (N_7695,N_7111,N_7220);
nand U7696 (N_7696,N_7268,N_7383);
and U7697 (N_7697,N_7093,N_7429);
or U7698 (N_7698,N_7495,N_7447);
nand U7699 (N_7699,N_7277,N_7468);
nand U7700 (N_7700,N_7374,N_7177);
and U7701 (N_7701,N_7099,N_7349);
nand U7702 (N_7702,N_7193,N_7043);
nand U7703 (N_7703,N_7275,N_7435);
and U7704 (N_7704,N_7005,N_7346);
nor U7705 (N_7705,N_7195,N_7115);
nand U7706 (N_7706,N_7028,N_7018);
or U7707 (N_7707,N_7038,N_7412);
nor U7708 (N_7708,N_7254,N_7338);
nor U7709 (N_7709,N_7080,N_7148);
nor U7710 (N_7710,N_7081,N_7144);
or U7711 (N_7711,N_7088,N_7026);
nor U7712 (N_7712,N_7493,N_7318);
nor U7713 (N_7713,N_7424,N_7488);
nand U7714 (N_7714,N_7091,N_7132);
xnor U7715 (N_7715,N_7073,N_7492);
or U7716 (N_7716,N_7086,N_7190);
nand U7717 (N_7717,N_7187,N_7213);
nand U7718 (N_7718,N_7409,N_7068);
and U7719 (N_7719,N_7380,N_7269);
nor U7720 (N_7720,N_7281,N_7196);
nor U7721 (N_7721,N_7236,N_7344);
nand U7722 (N_7722,N_7131,N_7319);
xor U7723 (N_7723,N_7354,N_7259);
or U7724 (N_7724,N_7146,N_7377);
or U7725 (N_7725,N_7450,N_7222);
nor U7726 (N_7726,N_7276,N_7286);
nand U7727 (N_7727,N_7479,N_7186);
nor U7728 (N_7728,N_7244,N_7066);
xnor U7729 (N_7729,N_7120,N_7030);
or U7730 (N_7730,N_7323,N_7427);
or U7731 (N_7731,N_7108,N_7209);
xnor U7732 (N_7732,N_7046,N_7394);
or U7733 (N_7733,N_7352,N_7371);
nand U7734 (N_7734,N_7428,N_7210);
xor U7735 (N_7735,N_7430,N_7251);
or U7736 (N_7736,N_7341,N_7012);
nand U7737 (N_7737,N_7116,N_7370);
nand U7738 (N_7738,N_7166,N_7420);
nand U7739 (N_7739,N_7011,N_7469);
xnor U7740 (N_7740,N_7460,N_7448);
and U7741 (N_7741,N_7330,N_7293);
or U7742 (N_7742,N_7462,N_7235);
and U7743 (N_7743,N_7087,N_7162);
nand U7744 (N_7744,N_7164,N_7368);
or U7745 (N_7745,N_7289,N_7041);
nand U7746 (N_7746,N_7147,N_7313);
or U7747 (N_7747,N_7096,N_7301);
xor U7748 (N_7748,N_7180,N_7123);
xnor U7749 (N_7749,N_7418,N_7007);
xnor U7750 (N_7750,N_7066,N_7387);
nand U7751 (N_7751,N_7290,N_7489);
and U7752 (N_7752,N_7145,N_7225);
nor U7753 (N_7753,N_7468,N_7341);
or U7754 (N_7754,N_7073,N_7001);
xor U7755 (N_7755,N_7166,N_7202);
xnor U7756 (N_7756,N_7360,N_7112);
or U7757 (N_7757,N_7179,N_7265);
and U7758 (N_7758,N_7298,N_7141);
nand U7759 (N_7759,N_7382,N_7233);
nand U7760 (N_7760,N_7302,N_7414);
or U7761 (N_7761,N_7171,N_7228);
xnor U7762 (N_7762,N_7254,N_7374);
nor U7763 (N_7763,N_7019,N_7212);
nor U7764 (N_7764,N_7159,N_7173);
and U7765 (N_7765,N_7378,N_7211);
nand U7766 (N_7766,N_7295,N_7423);
and U7767 (N_7767,N_7453,N_7326);
and U7768 (N_7768,N_7387,N_7289);
xor U7769 (N_7769,N_7118,N_7079);
nor U7770 (N_7770,N_7037,N_7401);
nand U7771 (N_7771,N_7045,N_7047);
nand U7772 (N_7772,N_7428,N_7076);
xor U7773 (N_7773,N_7061,N_7476);
or U7774 (N_7774,N_7384,N_7128);
or U7775 (N_7775,N_7202,N_7011);
nor U7776 (N_7776,N_7062,N_7156);
and U7777 (N_7777,N_7308,N_7496);
or U7778 (N_7778,N_7110,N_7401);
and U7779 (N_7779,N_7496,N_7405);
and U7780 (N_7780,N_7428,N_7475);
xnor U7781 (N_7781,N_7376,N_7373);
or U7782 (N_7782,N_7250,N_7450);
nand U7783 (N_7783,N_7021,N_7285);
and U7784 (N_7784,N_7150,N_7215);
or U7785 (N_7785,N_7075,N_7492);
and U7786 (N_7786,N_7274,N_7082);
nor U7787 (N_7787,N_7094,N_7488);
and U7788 (N_7788,N_7130,N_7194);
xnor U7789 (N_7789,N_7279,N_7072);
or U7790 (N_7790,N_7105,N_7302);
nand U7791 (N_7791,N_7054,N_7202);
nor U7792 (N_7792,N_7471,N_7058);
nor U7793 (N_7793,N_7131,N_7494);
or U7794 (N_7794,N_7399,N_7482);
nor U7795 (N_7795,N_7133,N_7382);
or U7796 (N_7796,N_7073,N_7140);
nor U7797 (N_7797,N_7246,N_7115);
or U7798 (N_7798,N_7165,N_7327);
xor U7799 (N_7799,N_7019,N_7148);
or U7800 (N_7800,N_7249,N_7013);
xnor U7801 (N_7801,N_7305,N_7136);
nand U7802 (N_7802,N_7447,N_7194);
and U7803 (N_7803,N_7009,N_7213);
nand U7804 (N_7804,N_7274,N_7474);
and U7805 (N_7805,N_7430,N_7360);
nor U7806 (N_7806,N_7209,N_7279);
xor U7807 (N_7807,N_7460,N_7492);
xnor U7808 (N_7808,N_7496,N_7398);
nor U7809 (N_7809,N_7128,N_7155);
or U7810 (N_7810,N_7407,N_7317);
and U7811 (N_7811,N_7269,N_7165);
and U7812 (N_7812,N_7371,N_7432);
xnor U7813 (N_7813,N_7332,N_7174);
or U7814 (N_7814,N_7165,N_7191);
or U7815 (N_7815,N_7475,N_7058);
and U7816 (N_7816,N_7436,N_7464);
xor U7817 (N_7817,N_7160,N_7020);
and U7818 (N_7818,N_7261,N_7430);
nor U7819 (N_7819,N_7399,N_7192);
or U7820 (N_7820,N_7429,N_7434);
xnor U7821 (N_7821,N_7223,N_7283);
xor U7822 (N_7822,N_7057,N_7188);
and U7823 (N_7823,N_7094,N_7180);
or U7824 (N_7824,N_7379,N_7335);
or U7825 (N_7825,N_7439,N_7122);
nor U7826 (N_7826,N_7019,N_7072);
or U7827 (N_7827,N_7323,N_7477);
xnor U7828 (N_7828,N_7151,N_7393);
and U7829 (N_7829,N_7499,N_7313);
nand U7830 (N_7830,N_7444,N_7156);
nor U7831 (N_7831,N_7220,N_7112);
xor U7832 (N_7832,N_7222,N_7084);
and U7833 (N_7833,N_7266,N_7094);
nand U7834 (N_7834,N_7404,N_7073);
and U7835 (N_7835,N_7335,N_7499);
or U7836 (N_7836,N_7327,N_7133);
xnor U7837 (N_7837,N_7241,N_7113);
xnor U7838 (N_7838,N_7079,N_7237);
nor U7839 (N_7839,N_7371,N_7207);
xnor U7840 (N_7840,N_7346,N_7413);
nand U7841 (N_7841,N_7340,N_7124);
and U7842 (N_7842,N_7223,N_7204);
nor U7843 (N_7843,N_7313,N_7497);
and U7844 (N_7844,N_7339,N_7030);
nand U7845 (N_7845,N_7287,N_7100);
nand U7846 (N_7846,N_7041,N_7468);
nor U7847 (N_7847,N_7497,N_7292);
and U7848 (N_7848,N_7169,N_7343);
or U7849 (N_7849,N_7171,N_7191);
nand U7850 (N_7850,N_7215,N_7392);
and U7851 (N_7851,N_7495,N_7010);
nand U7852 (N_7852,N_7132,N_7192);
nand U7853 (N_7853,N_7260,N_7153);
nor U7854 (N_7854,N_7488,N_7019);
nand U7855 (N_7855,N_7352,N_7403);
nor U7856 (N_7856,N_7107,N_7222);
nand U7857 (N_7857,N_7334,N_7473);
nor U7858 (N_7858,N_7461,N_7256);
nand U7859 (N_7859,N_7360,N_7467);
nand U7860 (N_7860,N_7316,N_7436);
and U7861 (N_7861,N_7215,N_7425);
nor U7862 (N_7862,N_7437,N_7306);
or U7863 (N_7863,N_7124,N_7350);
and U7864 (N_7864,N_7459,N_7408);
and U7865 (N_7865,N_7401,N_7194);
xor U7866 (N_7866,N_7238,N_7169);
nor U7867 (N_7867,N_7478,N_7347);
nand U7868 (N_7868,N_7319,N_7242);
nor U7869 (N_7869,N_7317,N_7409);
xnor U7870 (N_7870,N_7357,N_7195);
and U7871 (N_7871,N_7424,N_7072);
xor U7872 (N_7872,N_7351,N_7117);
xor U7873 (N_7873,N_7445,N_7390);
nand U7874 (N_7874,N_7146,N_7017);
and U7875 (N_7875,N_7394,N_7416);
nand U7876 (N_7876,N_7300,N_7022);
nor U7877 (N_7877,N_7206,N_7271);
nor U7878 (N_7878,N_7323,N_7315);
nor U7879 (N_7879,N_7480,N_7000);
and U7880 (N_7880,N_7011,N_7179);
xnor U7881 (N_7881,N_7383,N_7072);
and U7882 (N_7882,N_7152,N_7399);
nor U7883 (N_7883,N_7214,N_7223);
nor U7884 (N_7884,N_7004,N_7273);
and U7885 (N_7885,N_7471,N_7094);
or U7886 (N_7886,N_7391,N_7332);
nor U7887 (N_7887,N_7441,N_7423);
and U7888 (N_7888,N_7146,N_7473);
xnor U7889 (N_7889,N_7276,N_7005);
nand U7890 (N_7890,N_7204,N_7050);
and U7891 (N_7891,N_7484,N_7299);
xnor U7892 (N_7892,N_7404,N_7147);
nand U7893 (N_7893,N_7077,N_7191);
and U7894 (N_7894,N_7061,N_7104);
and U7895 (N_7895,N_7000,N_7116);
nor U7896 (N_7896,N_7351,N_7277);
or U7897 (N_7897,N_7046,N_7068);
nand U7898 (N_7898,N_7408,N_7099);
nand U7899 (N_7899,N_7094,N_7415);
xnor U7900 (N_7900,N_7053,N_7179);
or U7901 (N_7901,N_7478,N_7264);
xnor U7902 (N_7902,N_7059,N_7284);
nand U7903 (N_7903,N_7495,N_7144);
nor U7904 (N_7904,N_7294,N_7173);
or U7905 (N_7905,N_7253,N_7056);
or U7906 (N_7906,N_7335,N_7103);
or U7907 (N_7907,N_7422,N_7423);
nand U7908 (N_7908,N_7452,N_7302);
nor U7909 (N_7909,N_7055,N_7155);
nand U7910 (N_7910,N_7106,N_7454);
or U7911 (N_7911,N_7308,N_7103);
or U7912 (N_7912,N_7140,N_7169);
nor U7913 (N_7913,N_7049,N_7279);
and U7914 (N_7914,N_7289,N_7148);
nor U7915 (N_7915,N_7165,N_7459);
and U7916 (N_7916,N_7100,N_7461);
xnor U7917 (N_7917,N_7372,N_7379);
nor U7918 (N_7918,N_7384,N_7118);
or U7919 (N_7919,N_7070,N_7355);
and U7920 (N_7920,N_7272,N_7471);
or U7921 (N_7921,N_7303,N_7431);
xnor U7922 (N_7922,N_7149,N_7075);
nand U7923 (N_7923,N_7406,N_7137);
and U7924 (N_7924,N_7158,N_7081);
nand U7925 (N_7925,N_7182,N_7419);
xor U7926 (N_7926,N_7449,N_7149);
nor U7927 (N_7927,N_7400,N_7410);
or U7928 (N_7928,N_7354,N_7011);
xnor U7929 (N_7929,N_7316,N_7428);
and U7930 (N_7930,N_7354,N_7107);
xnor U7931 (N_7931,N_7068,N_7403);
xnor U7932 (N_7932,N_7292,N_7042);
xor U7933 (N_7933,N_7019,N_7490);
nor U7934 (N_7934,N_7036,N_7431);
nor U7935 (N_7935,N_7222,N_7446);
or U7936 (N_7936,N_7016,N_7357);
xnor U7937 (N_7937,N_7199,N_7025);
xnor U7938 (N_7938,N_7289,N_7331);
xor U7939 (N_7939,N_7440,N_7117);
or U7940 (N_7940,N_7437,N_7351);
xnor U7941 (N_7941,N_7310,N_7413);
xnor U7942 (N_7942,N_7094,N_7001);
xor U7943 (N_7943,N_7088,N_7319);
or U7944 (N_7944,N_7413,N_7043);
nand U7945 (N_7945,N_7321,N_7325);
nand U7946 (N_7946,N_7100,N_7339);
nor U7947 (N_7947,N_7419,N_7298);
nand U7948 (N_7948,N_7172,N_7394);
nand U7949 (N_7949,N_7257,N_7098);
nor U7950 (N_7950,N_7212,N_7097);
or U7951 (N_7951,N_7172,N_7188);
nand U7952 (N_7952,N_7165,N_7178);
or U7953 (N_7953,N_7480,N_7373);
nand U7954 (N_7954,N_7333,N_7190);
nand U7955 (N_7955,N_7303,N_7404);
and U7956 (N_7956,N_7061,N_7402);
and U7957 (N_7957,N_7436,N_7468);
nand U7958 (N_7958,N_7279,N_7156);
nand U7959 (N_7959,N_7023,N_7301);
and U7960 (N_7960,N_7199,N_7365);
nor U7961 (N_7961,N_7037,N_7391);
nand U7962 (N_7962,N_7357,N_7375);
nand U7963 (N_7963,N_7341,N_7445);
and U7964 (N_7964,N_7219,N_7483);
xnor U7965 (N_7965,N_7268,N_7318);
nand U7966 (N_7966,N_7252,N_7422);
and U7967 (N_7967,N_7292,N_7437);
or U7968 (N_7968,N_7158,N_7214);
and U7969 (N_7969,N_7154,N_7181);
and U7970 (N_7970,N_7096,N_7425);
and U7971 (N_7971,N_7150,N_7008);
and U7972 (N_7972,N_7186,N_7207);
or U7973 (N_7973,N_7318,N_7192);
nand U7974 (N_7974,N_7139,N_7447);
xor U7975 (N_7975,N_7352,N_7239);
nand U7976 (N_7976,N_7219,N_7308);
and U7977 (N_7977,N_7024,N_7222);
nor U7978 (N_7978,N_7064,N_7114);
nor U7979 (N_7979,N_7329,N_7489);
nand U7980 (N_7980,N_7322,N_7146);
and U7981 (N_7981,N_7315,N_7236);
nor U7982 (N_7982,N_7384,N_7418);
nor U7983 (N_7983,N_7098,N_7248);
nor U7984 (N_7984,N_7093,N_7485);
or U7985 (N_7985,N_7041,N_7400);
and U7986 (N_7986,N_7337,N_7304);
nor U7987 (N_7987,N_7475,N_7387);
xnor U7988 (N_7988,N_7064,N_7028);
xnor U7989 (N_7989,N_7078,N_7156);
nor U7990 (N_7990,N_7398,N_7492);
or U7991 (N_7991,N_7294,N_7026);
nor U7992 (N_7992,N_7150,N_7458);
or U7993 (N_7993,N_7326,N_7175);
nor U7994 (N_7994,N_7369,N_7195);
and U7995 (N_7995,N_7403,N_7056);
xnor U7996 (N_7996,N_7193,N_7004);
nor U7997 (N_7997,N_7213,N_7066);
nor U7998 (N_7998,N_7061,N_7341);
or U7999 (N_7999,N_7234,N_7120);
nand U8000 (N_8000,N_7885,N_7875);
nor U8001 (N_8001,N_7751,N_7912);
nand U8002 (N_8002,N_7636,N_7720);
xor U8003 (N_8003,N_7818,N_7528);
and U8004 (N_8004,N_7508,N_7899);
xnor U8005 (N_8005,N_7650,N_7781);
and U8006 (N_8006,N_7570,N_7608);
nand U8007 (N_8007,N_7854,N_7647);
or U8008 (N_8008,N_7676,N_7759);
nand U8009 (N_8009,N_7567,N_7810);
xnor U8010 (N_8010,N_7744,N_7724);
and U8011 (N_8011,N_7832,N_7664);
and U8012 (N_8012,N_7597,N_7773);
nand U8013 (N_8013,N_7690,N_7671);
nor U8014 (N_8014,N_7628,N_7610);
or U8015 (N_8015,N_7856,N_7517);
nor U8016 (N_8016,N_7710,N_7822);
or U8017 (N_8017,N_7725,N_7891);
and U8018 (N_8018,N_7753,N_7577);
xnor U8019 (N_8019,N_7551,N_7794);
nand U8020 (N_8020,N_7967,N_7663);
nor U8021 (N_8021,N_7548,N_7541);
or U8022 (N_8022,N_7591,N_7749);
or U8023 (N_8023,N_7969,N_7809);
nand U8024 (N_8024,N_7898,N_7828);
or U8025 (N_8025,N_7711,N_7626);
or U8026 (N_8026,N_7826,N_7950);
or U8027 (N_8027,N_7585,N_7621);
or U8028 (N_8028,N_7732,N_7764);
xnor U8029 (N_8029,N_7827,N_7658);
and U8030 (N_8030,N_7735,N_7963);
and U8031 (N_8031,N_7736,N_7845);
nand U8032 (N_8032,N_7646,N_7503);
nand U8033 (N_8033,N_7986,N_7971);
nand U8034 (N_8034,N_7512,N_7807);
or U8035 (N_8035,N_7787,N_7961);
xor U8036 (N_8036,N_7775,N_7761);
nand U8037 (N_8037,N_7739,N_7993);
or U8038 (N_8038,N_7581,N_7640);
or U8039 (N_8039,N_7605,N_7678);
xnor U8040 (N_8040,N_7590,N_7976);
nor U8041 (N_8041,N_7682,N_7716);
nand U8042 (N_8042,N_7555,N_7842);
nand U8043 (N_8043,N_7660,N_7547);
nand U8044 (N_8044,N_7997,N_7858);
and U8045 (N_8045,N_7878,N_7959);
xnor U8046 (N_8046,N_7979,N_7755);
nor U8047 (N_8047,N_7587,N_7977);
xnor U8048 (N_8048,N_7593,N_7927);
nor U8049 (N_8049,N_7903,N_7533);
and U8050 (N_8050,N_7834,N_7728);
nor U8051 (N_8051,N_7844,N_7501);
xnor U8052 (N_8052,N_7520,N_7988);
or U8053 (N_8053,N_7507,N_7734);
and U8054 (N_8054,N_7576,N_7894);
and U8055 (N_8055,N_7670,N_7960);
xnor U8056 (N_8056,N_7887,N_7513);
or U8057 (N_8057,N_7872,N_7865);
or U8058 (N_8058,N_7880,N_7638);
and U8059 (N_8059,N_7905,N_7957);
or U8060 (N_8060,N_7830,N_7583);
and U8061 (N_8061,N_7730,N_7586);
nor U8062 (N_8062,N_7667,N_7805);
nor U8063 (N_8063,N_7552,N_7972);
nor U8064 (N_8064,N_7833,N_7841);
xnor U8065 (N_8065,N_7537,N_7648);
and U8066 (N_8066,N_7578,N_7633);
nor U8067 (N_8067,N_7651,N_7702);
nand U8068 (N_8068,N_7900,N_7549);
or U8069 (N_8069,N_7677,N_7619);
and U8070 (N_8070,N_7579,N_7847);
or U8071 (N_8071,N_7776,N_7708);
nor U8072 (N_8072,N_7820,N_7510);
nor U8073 (N_8073,N_7639,N_7746);
nor U8074 (N_8074,N_7584,N_7895);
nand U8075 (N_8075,N_7952,N_7985);
or U8076 (N_8076,N_7742,N_7851);
xor U8077 (N_8077,N_7799,N_7866);
or U8078 (N_8078,N_7796,N_7774);
or U8079 (N_8079,N_7554,N_7611);
and U8080 (N_8080,N_7915,N_7893);
or U8081 (N_8081,N_7877,N_7740);
and U8082 (N_8082,N_7712,N_7925);
nor U8083 (N_8083,N_7917,N_7791);
or U8084 (N_8084,N_7543,N_7522);
xor U8085 (N_8085,N_7763,N_7762);
xor U8086 (N_8086,N_7630,N_7978);
xor U8087 (N_8087,N_7813,N_7538);
xor U8088 (N_8088,N_7991,N_7815);
nand U8089 (N_8089,N_7792,N_7526);
nor U8090 (N_8090,N_7954,N_7693);
nand U8091 (N_8091,N_7598,N_7609);
nor U8092 (N_8092,N_7523,N_7754);
and U8093 (N_8093,N_7649,N_7758);
and U8094 (N_8094,N_7989,N_7518);
nor U8095 (N_8095,N_7777,N_7916);
xnor U8096 (N_8096,N_7714,N_7596);
nor U8097 (N_8097,N_7862,N_7637);
or U8098 (N_8098,N_7808,N_7536);
or U8099 (N_8099,N_7784,N_7782);
or U8100 (N_8100,N_7629,N_7803);
and U8101 (N_8101,N_7902,N_7539);
nand U8102 (N_8102,N_7686,N_7652);
and U8103 (N_8103,N_7573,N_7766);
nand U8104 (N_8104,N_7962,N_7531);
nor U8105 (N_8105,N_7668,N_7980);
xor U8106 (N_8106,N_7814,N_7506);
and U8107 (N_8107,N_7550,N_7645);
xor U8108 (N_8108,N_7653,N_7857);
nor U8109 (N_8109,N_7515,N_7603);
nor U8110 (N_8110,N_7757,N_7624);
xnor U8111 (N_8111,N_7750,N_7882);
and U8112 (N_8112,N_7582,N_7929);
and U8113 (N_8113,N_7884,N_7798);
or U8114 (N_8114,N_7968,N_7945);
or U8115 (N_8115,N_7709,N_7530);
or U8116 (N_8116,N_7890,N_7729);
nor U8117 (N_8117,N_7500,N_7848);
or U8118 (N_8118,N_7502,N_7767);
and U8119 (N_8119,N_7564,N_7689);
xnor U8120 (N_8120,N_7731,N_7931);
nor U8121 (N_8121,N_7901,N_7535);
nand U8122 (N_8122,N_7718,N_7540);
or U8123 (N_8123,N_7569,N_7760);
or U8124 (N_8124,N_7935,N_7566);
nor U8125 (N_8125,N_7911,N_7553);
nand U8126 (N_8126,N_7701,N_7704);
nand U8127 (N_8127,N_7620,N_7839);
and U8128 (N_8128,N_7859,N_7680);
nand U8129 (N_8129,N_7723,N_7542);
nand U8130 (N_8130,N_7769,N_7521);
nand U8131 (N_8131,N_7713,N_7996);
and U8132 (N_8132,N_7559,N_7852);
nor U8133 (N_8133,N_7965,N_7788);
or U8134 (N_8134,N_7897,N_7756);
xor U8135 (N_8135,N_7688,N_7934);
xnor U8136 (N_8136,N_7726,N_7745);
nor U8137 (N_8137,N_7659,N_7793);
nor U8138 (N_8138,N_7821,N_7594);
nand U8139 (N_8139,N_7644,N_7837);
xor U8140 (N_8140,N_7703,N_7920);
nor U8141 (N_8141,N_7871,N_7705);
nor U8142 (N_8142,N_7944,N_7907);
nor U8143 (N_8143,N_7527,N_7800);
nor U8144 (N_8144,N_7879,N_7642);
nor U8145 (N_8145,N_7683,N_7942);
xnor U8146 (N_8146,N_7641,N_7982);
and U8147 (N_8147,N_7966,N_7511);
or U8148 (N_8148,N_7601,N_7904);
nand U8149 (N_8149,N_7816,N_7896);
nand U8150 (N_8150,N_7558,N_7707);
nor U8151 (N_8151,N_7881,N_7673);
and U8152 (N_8152,N_7943,N_7625);
xnor U8153 (N_8153,N_7823,N_7568);
nand U8154 (N_8154,N_7616,N_7618);
or U8155 (N_8155,N_7940,N_7635);
nand U8156 (N_8156,N_7797,N_7696);
or U8157 (N_8157,N_7679,N_7923);
and U8158 (N_8158,N_7752,N_7948);
or U8159 (N_8159,N_7717,N_7860);
nand U8160 (N_8160,N_7571,N_7995);
nor U8161 (N_8161,N_7574,N_7811);
or U8162 (N_8162,N_7994,N_7643);
xnor U8163 (N_8163,N_7909,N_7964);
nand U8164 (N_8164,N_7694,N_7906);
and U8165 (N_8165,N_7604,N_7937);
xor U8166 (N_8166,N_7956,N_7727);
xnor U8167 (N_8167,N_7765,N_7698);
nand U8168 (N_8168,N_7801,N_7778);
and U8169 (N_8169,N_7806,N_7665);
xnor U8170 (N_8170,N_7958,N_7924);
xor U8171 (N_8171,N_7771,N_7886);
and U8172 (N_8172,N_7666,N_7974);
nor U8173 (N_8173,N_7721,N_7657);
and U8174 (N_8174,N_7910,N_7932);
xnor U8175 (N_8175,N_7662,N_7692);
nor U8176 (N_8176,N_7947,N_7853);
xnor U8177 (N_8177,N_7654,N_7747);
and U8178 (N_8178,N_7623,N_7595);
and U8179 (N_8179,N_7873,N_7614);
xnor U8180 (N_8180,N_7699,N_7908);
nand U8181 (N_8181,N_7840,N_7933);
or U8182 (N_8182,N_7748,N_7634);
nor U8183 (N_8183,N_7846,N_7804);
and U8184 (N_8184,N_7975,N_7913);
or U8185 (N_8185,N_7922,N_7615);
xor U8186 (N_8186,N_7743,N_7722);
and U8187 (N_8187,N_7999,N_7600);
nor U8188 (N_8188,N_7928,N_7733);
and U8189 (N_8189,N_7835,N_7612);
or U8190 (N_8190,N_7674,N_7602);
nand U8191 (N_8191,N_7560,N_7505);
nand U8192 (N_8192,N_7607,N_7921);
and U8193 (N_8193,N_7946,N_7829);
nor U8194 (N_8194,N_7627,N_7831);
nand U8195 (N_8195,N_7892,N_7883);
xor U8196 (N_8196,N_7919,N_7684);
and U8197 (N_8197,N_7783,N_7592);
nand U8198 (N_8198,N_7655,N_7867);
or U8199 (N_8199,N_7719,N_7785);
and U8200 (N_8200,N_7930,N_7545);
nor U8201 (N_8201,N_7516,N_7534);
and U8202 (N_8202,N_7557,N_7825);
nand U8203 (N_8203,N_7990,N_7795);
or U8204 (N_8204,N_7556,N_7812);
xnor U8205 (N_8205,N_7973,N_7855);
and U8206 (N_8206,N_7863,N_7669);
xnor U8207 (N_8207,N_7504,N_7706);
nand U8208 (N_8208,N_7589,N_7780);
nand U8209 (N_8209,N_7802,N_7779);
and U8210 (N_8210,N_7741,N_7563);
nand U8211 (N_8211,N_7697,N_7715);
nor U8212 (N_8212,N_7981,N_7687);
or U8213 (N_8213,N_7613,N_7889);
or U8214 (N_8214,N_7819,N_7532);
nand U8215 (N_8215,N_7983,N_7695);
or U8216 (N_8216,N_7838,N_7738);
nor U8217 (N_8217,N_7874,N_7580);
or U8218 (N_8218,N_7561,N_7984);
nor U8219 (N_8219,N_7770,N_7632);
or U8220 (N_8220,N_7588,N_7824);
and U8221 (N_8221,N_7768,N_7868);
or U8222 (N_8222,N_7606,N_7914);
nand U8223 (N_8223,N_7572,N_7938);
nand U8224 (N_8224,N_7786,N_7617);
or U8225 (N_8225,N_7941,N_7790);
and U8226 (N_8226,N_7939,N_7700);
xnor U8227 (N_8227,N_7575,N_7949);
and U8228 (N_8228,N_7524,N_7849);
and U8229 (N_8229,N_7876,N_7562);
xor U8230 (N_8230,N_7685,N_7737);
nand U8231 (N_8231,N_7864,N_7817);
or U8232 (N_8232,N_7525,N_7850);
nand U8233 (N_8233,N_7998,N_7529);
or U8234 (N_8234,N_7544,N_7869);
xnor U8235 (N_8235,N_7509,N_7951);
or U8236 (N_8236,N_7936,N_7970);
or U8237 (N_8237,N_7656,N_7622);
xnor U8238 (N_8238,N_7861,N_7992);
nor U8239 (N_8239,N_7870,N_7565);
nor U8240 (N_8240,N_7953,N_7631);
nand U8241 (N_8241,N_7926,N_7519);
or U8242 (N_8242,N_7675,N_7681);
or U8243 (N_8243,N_7918,N_7772);
and U8244 (N_8244,N_7836,N_7546);
nor U8245 (N_8245,N_7661,N_7599);
nand U8246 (N_8246,N_7514,N_7843);
nor U8247 (N_8247,N_7955,N_7691);
and U8248 (N_8248,N_7672,N_7987);
nand U8249 (N_8249,N_7888,N_7789);
nand U8250 (N_8250,N_7830,N_7928);
or U8251 (N_8251,N_7622,N_7985);
xnor U8252 (N_8252,N_7652,N_7762);
and U8253 (N_8253,N_7808,N_7845);
xor U8254 (N_8254,N_7502,N_7821);
or U8255 (N_8255,N_7563,N_7571);
nor U8256 (N_8256,N_7654,N_7690);
or U8257 (N_8257,N_7557,N_7909);
and U8258 (N_8258,N_7847,N_7845);
and U8259 (N_8259,N_7513,N_7583);
nand U8260 (N_8260,N_7814,N_7834);
nand U8261 (N_8261,N_7952,N_7676);
nor U8262 (N_8262,N_7985,N_7546);
and U8263 (N_8263,N_7754,N_7692);
nand U8264 (N_8264,N_7748,N_7678);
nor U8265 (N_8265,N_7841,N_7878);
and U8266 (N_8266,N_7752,N_7664);
and U8267 (N_8267,N_7593,N_7793);
nand U8268 (N_8268,N_7757,N_7822);
and U8269 (N_8269,N_7685,N_7504);
xnor U8270 (N_8270,N_7609,N_7994);
nor U8271 (N_8271,N_7739,N_7836);
or U8272 (N_8272,N_7567,N_7674);
nor U8273 (N_8273,N_7732,N_7521);
nand U8274 (N_8274,N_7733,N_7676);
xnor U8275 (N_8275,N_7568,N_7767);
or U8276 (N_8276,N_7650,N_7537);
nand U8277 (N_8277,N_7716,N_7885);
nor U8278 (N_8278,N_7706,N_7788);
and U8279 (N_8279,N_7663,N_7909);
nor U8280 (N_8280,N_7944,N_7574);
nand U8281 (N_8281,N_7703,N_7585);
nand U8282 (N_8282,N_7510,N_7736);
nor U8283 (N_8283,N_7708,N_7654);
or U8284 (N_8284,N_7800,N_7681);
and U8285 (N_8285,N_7665,N_7563);
nor U8286 (N_8286,N_7977,N_7796);
nor U8287 (N_8287,N_7609,N_7536);
and U8288 (N_8288,N_7895,N_7698);
and U8289 (N_8289,N_7574,N_7664);
xnor U8290 (N_8290,N_7664,N_7532);
nand U8291 (N_8291,N_7981,N_7500);
nor U8292 (N_8292,N_7933,N_7716);
nand U8293 (N_8293,N_7634,N_7598);
nand U8294 (N_8294,N_7507,N_7550);
and U8295 (N_8295,N_7664,N_7505);
xnor U8296 (N_8296,N_7507,N_7521);
or U8297 (N_8297,N_7667,N_7594);
nand U8298 (N_8298,N_7794,N_7558);
or U8299 (N_8299,N_7877,N_7744);
nor U8300 (N_8300,N_7631,N_7885);
nor U8301 (N_8301,N_7752,N_7609);
nand U8302 (N_8302,N_7625,N_7511);
or U8303 (N_8303,N_7776,N_7767);
nand U8304 (N_8304,N_7559,N_7566);
nor U8305 (N_8305,N_7523,N_7829);
or U8306 (N_8306,N_7568,N_7543);
xor U8307 (N_8307,N_7791,N_7588);
or U8308 (N_8308,N_7575,N_7769);
nand U8309 (N_8309,N_7714,N_7609);
and U8310 (N_8310,N_7890,N_7671);
xor U8311 (N_8311,N_7950,N_7867);
xnor U8312 (N_8312,N_7800,N_7945);
and U8313 (N_8313,N_7786,N_7753);
xnor U8314 (N_8314,N_7744,N_7954);
nand U8315 (N_8315,N_7525,N_7903);
xor U8316 (N_8316,N_7660,N_7969);
and U8317 (N_8317,N_7978,N_7968);
and U8318 (N_8318,N_7875,N_7546);
xnor U8319 (N_8319,N_7536,N_7931);
nor U8320 (N_8320,N_7585,N_7929);
or U8321 (N_8321,N_7986,N_7881);
nor U8322 (N_8322,N_7842,N_7876);
nand U8323 (N_8323,N_7725,N_7909);
nor U8324 (N_8324,N_7779,N_7820);
nand U8325 (N_8325,N_7597,N_7666);
and U8326 (N_8326,N_7618,N_7639);
nand U8327 (N_8327,N_7915,N_7720);
xor U8328 (N_8328,N_7964,N_7638);
nand U8329 (N_8329,N_7538,N_7967);
or U8330 (N_8330,N_7506,N_7688);
and U8331 (N_8331,N_7776,N_7806);
and U8332 (N_8332,N_7611,N_7511);
and U8333 (N_8333,N_7923,N_7797);
nor U8334 (N_8334,N_7575,N_7567);
nand U8335 (N_8335,N_7858,N_7958);
and U8336 (N_8336,N_7825,N_7595);
xor U8337 (N_8337,N_7980,N_7564);
nor U8338 (N_8338,N_7900,N_7502);
or U8339 (N_8339,N_7836,N_7834);
or U8340 (N_8340,N_7535,N_7758);
and U8341 (N_8341,N_7576,N_7594);
nor U8342 (N_8342,N_7524,N_7925);
and U8343 (N_8343,N_7778,N_7958);
and U8344 (N_8344,N_7952,N_7747);
nand U8345 (N_8345,N_7985,N_7806);
nor U8346 (N_8346,N_7935,N_7903);
nor U8347 (N_8347,N_7649,N_7856);
and U8348 (N_8348,N_7916,N_7653);
nor U8349 (N_8349,N_7573,N_7680);
xor U8350 (N_8350,N_7812,N_7521);
nor U8351 (N_8351,N_7594,N_7837);
xor U8352 (N_8352,N_7795,N_7669);
xor U8353 (N_8353,N_7872,N_7558);
xnor U8354 (N_8354,N_7961,N_7615);
nand U8355 (N_8355,N_7959,N_7966);
nand U8356 (N_8356,N_7692,N_7592);
or U8357 (N_8357,N_7592,N_7519);
and U8358 (N_8358,N_7929,N_7742);
nand U8359 (N_8359,N_7823,N_7791);
and U8360 (N_8360,N_7632,N_7602);
and U8361 (N_8361,N_7582,N_7606);
and U8362 (N_8362,N_7973,N_7629);
nor U8363 (N_8363,N_7852,N_7955);
and U8364 (N_8364,N_7555,N_7963);
nand U8365 (N_8365,N_7804,N_7893);
xnor U8366 (N_8366,N_7501,N_7826);
nand U8367 (N_8367,N_7978,N_7927);
and U8368 (N_8368,N_7723,N_7906);
or U8369 (N_8369,N_7862,N_7852);
nor U8370 (N_8370,N_7990,N_7528);
xnor U8371 (N_8371,N_7737,N_7857);
or U8372 (N_8372,N_7636,N_7618);
nor U8373 (N_8373,N_7768,N_7920);
nor U8374 (N_8374,N_7635,N_7835);
nand U8375 (N_8375,N_7877,N_7949);
and U8376 (N_8376,N_7820,N_7691);
and U8377 (N_8377,N_7654,N_7590);
or U8378 (N_8378,N_7916,N_7766);
xor U8379 (N_8379,N_7762,N_7539);
xor U8380 (N_8380,N_7873,N_7517);
or U8381 (N_8381,N_7892,N_7612);
xnor U8382 (N_8382,N_7848,N_7805);
xor U8383 (N_8383,N_7554,N_7534);
nand U8384 (N_8384,N_7598,N_7865);
xor U8385 (N_8385,N_7544,N_7604);
and U8386 (N_8386,N_7858,N_7621);
and U8387 (N_8387,N_7858,N_7991);
and U8388 (N_8388,N_7726,N_7908);
and U8389 (N_8389,N_7826,N_7539);
nor U8390 (N_8390,N_7600,N_7653);
nand U8391 (N_8391,N_7724,N_7864);
and U8392 (N_8392,N_7642,N_7731);
nor U8393 (N_8393,N_7587,N_7854);
or U8394 (N_8394,N_7752,N_7731);
or U8395 (N_8395,N_7937,N_7566);
xnor U8396 (N_8396,N_7751,N_7839);
xor U8397 (N_8397,N_7965,N_7667);
xor U8398 (N_8398,N_7590,N_7820);
nor U8399 (N_8399,N_7727,N_7602);
nand U8400 (N_8400,N_7746,N_7621);
xor U8401 (N_8401,N_7928,N_7778);
and U8402 (N_8402,N_7933,N_7638);
or U8403 (N_8403,N_7623,N_7660);
xor U8404 (N_8404,N_7668,N_7888);
or U8405 (N_8405,N_7502,N_7758);
xor U8406 (N_8406,N_7517,N_7985);
and U8407 (N_8407,N_7651,N_7832);
or U8408 (N_8408,N_7586,N_7644);
nor U8409 (N_8409,N_7997,N_7744);
xor U8410 (N_8410,N_7614,N_7700);
nand U8411 (N_8411,N_7671,N_7981);
nor U8412 (N_8412,N_7665,N_7876);
and U8413 (N_8413,N_7667,N_7691);
nand U8414 (N_8414,N_7918,N_7833);
nor U8415 (N_8415,N_7571,N_7993);
or U8416 (N_8416,N_7582,N_7629);
or U8417 (N_8417,N_7526,N_7599);
and U8418 (N_8418,N_7772,N_7936);
nand U8419 (N_8419,N_7727,N_7957);
or U8420 (N_8420,N_7590,N_7686);
and U8421 (N_8421,N_7578,N_7859);
and U8422 (N_8422,N_7542,N_7615);
nand U8423 (N_8423,N_7579,N_7941);
and U8424 (N_8424,N_7590,N_7814);
xor U8425 (N_8425,N_7747,N_7618);
or U8426 (N_8426,N_7609,N_7788);
nand U8427 (N_8427,N_7965,N_7518);
or U8428 (N_8428,N_7873,N_7523);
or U8429 (N_8429,N_7511,N_7708);
xor U8430 (N_8430,N_7870,N_7865);
xor U8431 (N_8431,N_7881,N_7639);
or U8432 (N_8432,N_7905,N_7629);
nor U8433 (N_8433,N_7732,N_7945);
or U8434 (N_8434,N_7943,N_7595);
nor U8435 (N_8435,N_7929,N_7736);
and U8436 (N_8436,N_7821,N_7954);
nor U8437 (N_8437,N_7861,N_7891);
and U8438 (N_8438,N_7568,N_7693);
or U8439 (N_8439,N_7718,N_7912);
or U8440 (N_8440,N_7551,N_7672);
and U8441 (N_8441,N_7543,N_7752);
xor U8442 (N_8442,N_7647,N_7919);
or U8443 (N_8443,N_7607,N_7939);
and U8444 (N_8444,N_7682,N_7857);
or U8445 (N_8445,N_7616,N_7760);
and U8446 (N_8446,N_7919,N_7593);
xnor U8447 (N_8447,N_7907,N_7735);
xor U8448 (N_8448,N_7576,N_7986);
nand U8449 (N_8449,N_7563,N_7846);
or U8450 (N_8450,N_7750,N_7669);
and U8451 (N_8451,N_7950,N_7564);
nand U8452 (N_8452,N_7895,N_7772);
and U8453 (N_8453,N_7872,N_7522);
xor U8454 (N_8454,N_7990,N_7631);
nand U8455 (N_8455,N_7542,N_7767);
nor U8456 (N_8456,N_7680,N_7589);
xor U8457 (N_8457,N_7893,N_7633);
and U8458 (N_8458,N_7677,N_7880);
and U8459 (N_8459,N_7587,N_7532);
or U8460 (N_8460,N_7837,N_7761);
nor U8461 (N_8461,N_7672,N_7535);
xor U8462 (N_8462,N_7824,N_7683);
nand U8463 (N_8463,N_7758,N_7916);
or U8464 (N_8464,N_7851,N_7990);
nand U8465 (N_8465,N_7774,N_7934);
and U8466 (N_8466,N_7878,N_7950);
and U8467 (N_8467,N_7920,N_7970);
xor U8468 (N_8468,N_7945,N_7550);
nor U8469 (N_8469,N_7639,N_7765);
xor U8470 (N_8470,N_7651,N_7584);
and U8471 (N_8471,N_7613,N_7725);
xor U8472 (N_8472,N_7662,N_7956);
xnor U8473 (N_8473,N_7836,N_7820);
and U8474 (N_8474,N_7573,N_7777);
or U8475 (N_8475,N_7811,N_7634);
or U8476 (N_8476,N_7790,N_7619);
nor U8477 (N_8477,N_7679,N_7960);
and U8478 (N_8478,N_7856,N_7970);
nor U8479 (N_8479,N_7608,N_7518);
xor U8480 (N_8480,N_7674,N_7711);
and U8481 (N_8481,N_7875,N_7581);
xnor U8482 (N_8482,N_7519,N_7758);
nand U8483 (N_8483,N_7716,N_7801);
nand U8484 (N_8484,N_7519,N_7779);
nand U8485 (N_8485,N_7677,N_7980);
or U8486 (N_8486,N_7511,N_7508);
nor U8487 (N_8487,N_7565,N_7755);
xor U8488 (N_8488,N_7521,N_7748);
or U8489 (N_8489,N_7599,N_7765);
nor U8490 (N_8490,N_7525,N_7993);
nor U8491 (N_8491,N_7788,N_7917);
nand U8492 (N_8492,N_7647,N_7644);
nor U8493 (N_8493,N_7693,N_7946);
and U8494 (N_8494,N_7748,N_7728);
or U8495 (N_8495,N_7696,N_7532);
nand U8496 (N_8496,N_7939,N_7819);
or U8497 (N_8497,N_7906,N_7774);
and U8498 (N_8498,N_7538,N_7689);
and U8499 (N_8499,N_7530,N_7649);
and U8500 (N_8500,N_8034,N_8233);
and U8501 (N_8501,N_8099,N_8307);
or U8502 (N_8502,N_8167,N_8050);
nor U8503 (N_8503,N_8132,N_8271);
or U8504 (N_8504,N_8181,N_8165);
or U8505 (N_8505,N_8096,N_8263);
or U8506 (N_8506,N_8362,N_8462);
or U8507 (N_8507,N_8429,N_8133);
nor U8508 (N_8508,N_8029,N_8045);
nor U8509 (N_8509,N_8182,N_8259);
or U8510 (N_8510,N_8152,N_8246);
and U8511 (N_8511,N_8423,N_8223);
and U8512 (N_8512,N_8146,N_8119);
and U8513 (N_8513,N_8469,N_8151);
nand U8514 (N_8514,N_8153,N_8476);
or U8515 (N_8515,N_8386,N_8170);
nor U8516 (N_8516,N_8248,N_8353);
nand U8517 (N_8517,N_8275,N_8496);
nand U8518 (N_8518,N_8474,N_8466);
xor U8519 (N_8519,N_8042,N_8304);
xor U8520 (N_8520,N_8201,N_8021);
and U8521 (N_8521,N_8380,N_8396);
nor U8522 (N_8522,N_8068,N_8158);
and U8523 (N_8523,N_8415,N_8063);
and U8524 (N_8524,N_8098,N_8150);
nor U8525 (N_8525,N_8094,N_8071);
nand U8526 (N_8526,N_8202,N_8406);
xor U8527 (N_8527,N_8349,N_8217);
and U8528 (N_8528,N_8377,N_8280);
xor U8529 (N_8529,N_8286,N_8001);
or U8530 (N_8530,N_8087,N_8114);
xor U8531 (N_8531,N_8055,N_8142);
and U8532 (N_8532,N_8149,N_8399);
or U8533 (N_8533,N_8011,N_8285);
nand U8534 (N_8534,N_8443,N_8434);
xnor U8535 (N_8535,N_8137,N_8076);
nand U8536 (N_8536,N_8230,N_8184);
xnor U8537 (N_8537,N_8141,N_8379);
or U8538 (N_8538,N_8446,N_8331);
or U8539 (N_8539,N_8097,N_8344);
nor U8540 (N_8540,N_8005,N_8420);
xnor U8541 (N_8541,N_8350,N_8252);
or U8542 (N_8542,N_8484,N_8456);
and U8543 (N_8543,N_8186,N_8166);
nor U8544 (N_8544,N_8053,N_8289);
and U8545 (N_8545,N_8266,N_8240);
or U8546 (N_8546,N_8010,N_8297);
xor U8547 (N_8547,N_8135,N_8337);
xnor U8548 (N_8548,N_8120,N_8065);
nor U8549 (N_8549,N_8100,N_8024);
nand U8550 (N_8550,N_8425,N_8140);
nor U8551 (N_8551,N_8499,N_8104);
nor U8552 (N_8552,N_8483,N_8421);
xor U8553 (N_8553,N_8007,N_8121);
nor U8554 (N_8554,N_8080,N_8258);
and U8555 (N_8555,N_8014,N_8113);
or U8556 (N_8556,N_8294,N_8361);
nand U8557 (N_8557,N_8162,N_8116);
xor U8558 (N_8558,N_8311,N_8332);
nand U8559 (N_8559,N_8083,N_8197);
or U8560 (N_8560,N_8126,N_8249);
nor U8561 (N_8561,N_8418,N_8487);
and U8562 (N_8562,N_8417,N_8288);
nand U8563 (N_8563,N_8461,N_8287);
xor U8564 (N_8564,N_8376,N_8416);
xor U8565 (N_8565,N_8205,N_8257);
xor U8566 (N_8566,N_8449,N_8025);
xnor U8567 (N_8567,N_8346,N_8348);
xnor U8568 (N_8568,N_8485,N_8039);
xnor U8569 (N_8569,N_8409,N_8327);
nor U8570 (N_8570,N_8281,N_8174);
nor U8571 (N_8571,N_8012,N_8452);
or U8572 (N_8572,N_8340,N_8195);
nor U8573 (N_8573,N_8437,N_8190);
xor U8574 (N_8574,N_8136,N_8156);
or U8575 (N_8575,N_8244,N_8352);
nand U8576 (N_8576,N_8306,N_8253);
or U8577 (N_8577,N_8325,N_8498);
nand U8578 (N_8578,N_8058,N_8370);
and U8579 (N_8579,N_8477,N_8060);
and U8580 (N_8580,N_8251,N_8033);
or U8581 (N_8581,N_8069,N_8389);
nand U8582 (N_8582,N_8118,N_8319);
nand U8583 (N_8583,N_8400,N_8216);
nor U8584 (N_8584,N_8375,N_8347);
xnor U8585 (N_8585,N_8108,N_8163);
xnor U8586 (N_8586,N_8122,N_8106);
xnor U8587 (N_8587,N_8075,N_8392);
or U8588 (N_8588,N_8084,N_8407);
nand U8589 (N_8589,N_8491,N_8459);
and U8590 (N_8590,N_8272,N_8191);
or U8591 (N_8591,N_8020,N_8478);
xor U8592 (N_8592,N_8131,N_8209);
nand U8593 (N_8593,N_8442,N_8435);
and U8594 (N_8594,N_8226,N_8358);
or U8595 (N_8595,N_8241,N_8291);
nand U8596 (N_8596,N_8200,N_8026);
xnor U8597 (N_8597,N_8277,N_8117);
or U8598 (N_8598,N_8388,N_8308);
xnor U8599 (N_8599,N_8061,N_8145);
nor U8600 (N_8600,N_8382,N_8293);
nor U8601 (N_8601,N_8189,N_8187);
xnor U8602 (N_8602,N_8221,N_8130);
and U8603 (N_8603,N_8073,N_8482);
nor U8604 (N_8604,N_8056,N_8427);
nand U8605 (N_8605,N_8105,N_8312);
and U8606 (N_8606,N_8188,N_8250);
nand U8607 (N_8607,N_8300,N_8225);
or U8608 (N_8608,N_8410,N_8237);
xor U8609 (N_8609,N_8198,N_8268);
nor U8610 (N_8610,N_8148,N_8101);
nor U8611 (N_8611,N_8044,N_8298);
or U8612 (N_8612,N_8016,N_8315);
nand U8613 (N_8613,N_8047,N_8214);
xor U8614 (N_8614,N_8243,N_8123);
nor U8615 (N_8615,N_8303,N_8036);
nand U8616 (N_8616,N_8004,N_8492);
and U8617 (N_8617,N_8090,N_8046);
and U8618 (N_8618,N_8179,N_8320);
xnor U8619 (N_8619,N_8404,N_8463);
xor U8620 (N_8620,N_8043,N_8364);
nand U8621 (N_8621,N_8138,N_8077);
xnor U8622 (N_8622,N_8003,N_8032);
xor U8623 (N_8623,N_8354,N_8430);
nor U8624 (N_8624,N_8472,N_8212);
xor U8625 (N_8625,N_8447,N_8481);
and U8626 (N_8626,N_8278,N_8206);
and U8627 (N_8627,N_8203,N_8147);
or U8628 (N_8628,N_8169,N_8035);
or U8629 (N_8629,N_8334,N_8305);
nand U8630 (N_8630,N_8092,N_8030);
nand U8631 (N_8631,N_8284,N_8115);
nand U8632 (N_8632,N_8448,N_8381);
and U8633 (N_8633,N_8345,N_8239);
and U8634 (N_8634,N_8144,N_8027);
nor U8635 (N_8635,N_8022,N_8048);
xnor U8636 (N_8636,N_8473,N_8321);
nand U8637 (N_8637,N_8454,N_8059);
nand U8638 (N_8638,N_8041,N_8196);
or U8639 (N_8639,N_8450,N_8091);
nor U8640 (N_8640,N_8103,N_8031);
or U8641 (N_8641,N_8316,N_8139);
and U8642 (N_8642,N_8438,N_8444);
nor U8643 (N_8643,N_8464,N_8424);
nor U8644 (N_8644,N_8222,N_8125);
and U8645 (N_8645,N_8038,N_8054);
or U8646 (N_8646,N_8018,N_8467);
and U8647 (N_8647,N_8265,N_8213);
or U8648 (N_8648,N_8372,N_8367);
and U8649 (N_8649,N_8339,N_8134);
nor U8650 (N_8650,N_8049,N_8220);
and U8651 (N_8651,N_8002,N_8299);
xor U8652 (N_8652,N_8460,N_8422);
nor U8653 (N_8653,N_8168,N_8269);
nor U8654 (N_8654,N_8095,N_8219);
nor U8655 (N_8655,N_8267,N_8072);
and U8656 (N_8656,N_8408,N_8365);
or U8657 (N_8657,N_8279,N_8317);
and U8658 (N_8658,N_8210,N_8211);
nor U8659 (N_8659,N_8235,N_8330);
and U8660 (N_8660,N_8255,N_8494);
xnor U8661 (N_8661,N_8078,N_8497);
nand U8662 (N_8662,N_8102,N_8155);
xnor U8663 (N_8663,N_8458,N_8490);
xor U8664 (N_8664,N_8451,N_8411);
xor U8665 (N_8665,N_8256,N_8176);
or U8666 (N_8666,N_8366,N_8276);
nor U8667 (N_8667,N_8470,N_8323);
nand U8668 (N_8668,N_8371,N_8242);
nor U8669 (N_8669,N_8391,N_8260);
and U8670 (N_8670,N_8081,N_8384);
nand U8671 (N_8671,N_8374,N_8394);
xnor U8672 (N_8672,N_8419,N_8015);
or U8673 (N_8673,N_8009,N_8160);
or U8674 (N_8674,N_8128,N_8088);
or U8675 (N_8675,N_8177,N_8397);
nor U8676 (N_8676,N_8273,N_8356);
or U8677 (N_8677,N_8234,N_8175);
or U8678 (N_8678,N_8171,N_8000);
and U8679 (N_8679,N_8052,N_8426);
nor U8680 (N_8680,N_8385,N_8343);
and U8681 (N_8681,N_8363,N_8161);
or U8682 (N_8682,N_8093,N_8431);
xnor U8683 (N_8683,N_8193,N_8432);
and U8684 (N_8684,N_8086,N_8199);
xor U8685 (N_8685,N_8207,N_8111);
nor U8686 (N_8686,N_8475,N_8479);
nand U8687 (N_8687,N_8359,N_8378);
and U8688 (N_8688,N_8236,N_8180);
and U8689 (N_8689,N_8082,N_8342);
nand U8690 (N_8690,N_8107,N_8274);
and U8691 (N_8691,N_8254,N_8290);
nor U8692 (N_8692,N_8395,N_8079);
or U8693 (N_8693,N_8428,N_8208);
nor U8694 (N_8694,N_8023,N_8070);
or U8695 (N_8695,N_8127,N_8393);
nand U8696 (N_8696,N_8282,N_8224);
nand U8697 (N_8697,N_8040,N_8445);
nand U8698 (N_8698,N_8231,N_8322);
nand U8699 (N_8699,N_8309,N_8390);
nand U8700 (N_8700,N_8338,N_8074);
nor U8701 (N_8701,N_8328,N_8245);
or U8702 (N_8702,N_8369,N_8159);
xnor U8703 (N_8703,N_8261,N_8164);
nor U8704 (N_8704,N_8313,N_8066);
nor U8705 (N_8705,N_8028,N_8489);
and U8706 (N_8706,N_8204,N_8112);
nor U8707 (N_8707,N_8192,N_8455);
nor U8708 (N_8708,N_8412,N_8318);
xnor U8709 (N_8709,N_8089,N_8008);
xnor U8710 (N_8710,N_8183,N_8302);
nand U8711 (N_8711,N_8129,N_8368);
or U8712 (N_8712,N_8468,N_8013);
nor U8713 (N_8713,N_8295,N_8486);
nor U8714 (N_8714,N_8247,N_8017);
nor U8715 (N_8715,N_8373,N_8301);
or U8716 (N_8716,N_8493,N_8414);
nand U8717 (N_8717,N_8310,N_8228);
xnor U8718 (N_8718,N_8057,N_8124);
xnor U8719 (N_8719,N_8062,N_8109);
nand U8720 (N_8720,N_8019,N_8173);
or U8721 (N_8721,N_8360,N_8324);
or U8722 (N_8722,N_8314,N_8405);
xnor U8723 (N_8723,N_8157,N_8227);
or U8724 (N_8724,N_8270,N_8292);
and U8725 (N_8725,N_8403,N_8283);
nor U8726 (N_8726,N_8215,N_8336);
xnor U8727 (N_8727,N_8441,N_8067);
xor U8728 (N_8728,N_8355,N_8433);
and U8729 (N_8729,N_8085,N_8185);
nor U8730 (N_8730,N_8296,N_8387);
and U8731 (N_8731,N_8439,N_8051);
or U8732 (N_8732,N_8154,N_8218);
nor U8733 (N_8733,N_8178,N_8495);
xor U8734 (N_8734,N_8333,N_8335);
and U8735 (N_8735,N_8357,N_8436);
nand U8736 (N_8736,N_8037,N_8465);
xnor U8737 (N_8737,N_8453,N_8471);
xor U8738 (N_8738,N_8143,N_8398);
nand U8739 (N_8739,N_8194,N_8264);
xor U8740 (N_8740,N_8238,N_8413);
and U8741 (N_8741,N_8440,N_8329);
xor U8742 (N_8742,N_8351,N_8172);
nand U8743 (N_8743,N_8262,N_8383);
nand U8744 (N_8744,N_8402,N_8480);
xnor U8745 (N_8745,N_8457,N_8341);
or U8746 (N_8746,N_8232,N_8229);
nor U8747 (N_8747,N_8064,N_8326);
nor U8748 (N_8748,N_8488,N_8401);
nand U8749 (N_8749,N_8110,N_8006);
nand U8750 (N_8750,N_8257,N_8197);
xnor U8751 (N_8751,N_8451,N_8241);
or U8752 (N_8752,N_8279,N_8154);
and U8753 (N_8753,N_8499,N_8287);
nand U8754 (N_8754,N_8178,N_8104);
or U8755 (N_8755,N_8442,N_8316);
and U8756 (N_8756,N_8199,N_8079);
and U8757 (N_8757,N_8282,N_8444);
and U8758 (N_8758,N_8019,N_8091);
and U8759 (N_8759,N_8490,N_8471);
nor U8760 (N_8760,N_8008,N_8481);
xor U8761 (N_8761,N_8282,N_8361);
xnor U8762 (N_8762,N_8158,N_8056);
and U8763 (N_8763,N_8236,N_8308);
or U8764 (N_8764,N_8071,N_8367);
nand U8765 (N_8765,N_8080,N_8403);
and U8766 (N_8766,N_8245,N_8217);
or U8767 (N_8767,N_8214,N_8328);
nor U8768 (N_8768,N_8145,N_8120);
nor U8769 (N_8769,N_8220,N_8105);
xnor U8770 (N_8770,N_8467,N_8399);
and U8771 (N_8771,N_8394,N_8481);
or U8772 (N_8772,N_8137,N_8485);
nor U8773 (N_8773,N_8368,N_8273);
nand U8774 (N_8774,N_8479,N_8411);
or U8775 (N_8775,N_8348,N_8424);
xnor U8776 (N_8776,N_8008,N_8345);
xor U8777 (N_8777,N_8245,N_8495);
xnor U8778 (N_8778,N_8379,N_8385);
nor U8779 (N_8779,N_8259,N_8269);
and U8780 (N_8780,N_8078,N_8343);
and U8781 (N_8781,N_8324,N_8416);
nand U8782 (N_8782,N_8235,N_8238);
nand U8783 (N_8783,N_8322,N_8401);
nand U8784 (N_8784,N_8338,N_8327);
or U8785 (N_8785,N_8443,N_8291);
nand U8786 (N_8786,N_8367,N_8027);
or U8787 (N_8787,N_8088,N_8031);
xnor U8788 (N_8788,N_8011,N_8448);
xnor U8789 (N_8789,N_8099,N_8398);
xor U8790 (N_8790,N_8400,N_8473);
and U8791 (N_8791,N_8475,N_8374);
nand U8792 (N_8792,N_8151,N_8480);
or U8793 (N_8793,N_8391,N_8437);
xnor U8794 (N_8794,N_8313,N_8276);
xor U8795 (N_8795,N_8095,N_8357);
nand U8796 (N_8796,N_8150,N_8494);
xor U8797 (N_8797,N_8087,N_8487);
xnor U8798 (N_8798,N_8345,N_8389);
and U8799 (N_8799,N_8068,N_8118);
or U8800 (N_8800,N_8103,N_8144);
nor U8801 (N_8801,N_8326,N_8076);
and U8802 (N_8802,N_8427,N_8401);
nor U8803 (N_8803,N_8406,N_8437);
xnor U8804 (N_8804,N_8051,N_8193);
nor U8805 (N_8805,N_8161,N_8191);
nand U8806 (N_8806,N_8315,N_8386);
nand U8807 (N_8807,N_8356,N_8301);
and U8808 (N_8808,N_8014,N_8069);
nand U8809 (N_8809,N_8450,N_8415);
or U8810 (N_8810,N_8461,N_8401);
nor U8811 (N_8811,N_8356,N_8280);
nand U8812 (N_8812,N_8414,N_8165);
nor U8813 (N_8813,N_8369,N_8024);
and U8814 (N_8814,N_8476,N_8218);
nand U8815 (N_8815,N_8106,N_8413);
xnor U8816 (N_8816,N_8263,N_8184);
nor U8817 (N_8817,N_8495,N_8342);
nor U8818 (N_8818,N_8263,N_8333);
and U8819 (N_8819,N_8253,N_8387);
nor U8820 (N_8820,N_8041,N_8448);
and U8821 (N_8821,N_8051,N_8352);
or U8822 (N_8822,N_8375,N_8408);
nor U8823 (N_8823,N_8137,N_8146);
nand U8824 (N_8824,N_8037,N_8375);
nand U8825 (N_8825,N_8103,N_8232);
nand U8826 (N_8826,N_8168,N_8220);
nor U8827 (N_8827,N_8499,N_8324);
nand U8828 (N_8828,N_8216,N_8435);
nor U8829 (N_8829,N_8153,N_8216);
or U8830 (N_8830,N_8409,N_8356);
nor U8831 (N_8831,N_8216,N_8486);
xnor U8832 (N_8832,N_8306,N_8015);
xnor U8833 (N_8833,N_8194,N_8305);
and U8834 (N_8834,N_8187,N_8105);
nor U8835 (N_8835,N_8305,N_8132);
or U8836 (N_8836,N_8314,N_8130);
nand U8837 (N_8837,N_8382,N_8072);
and U8838 (N_8838,N_8227,N_8494);
nand U8839 (N_8839,N_8330,N_8102);
xor U8840 (N_8840,N_8292,N_8333);
xor U8841 (N_8841,N_8360,N_8038);
xnor U8842 (N_8842,N_8113,N_8209);
nand U8843 (N_8843,N_8022,N_8374);
xnor U8844 (N_8844,N_8321,N_8250);
nor U8845 (N_8845,N_8069,N_8435);
nand U8846 (N_8846,N_8396,N_8086);
or U8847 (N_8847,N_8432,N_8292);
and U8848 (N_8848,N_8078,N_8459);
or U8849 (N_8849,N_8075,N_8270);
or U8850 (N_8850,N_8176,N_8279);
or U8851 (N_8851,N_8087,N_8495);
and U8852 (N_8852,N_8135,N_8044);
xor U8853 (N_8853,N_8169,N_8391);
xor U8854 (N_8854,N_8484,N_8482);
or U8855 (N_8855,N_8094,N_8341);
or U8856 (N_8856,N_8128,N_8353);
and U8857 (N_8857,N_8136,N_8272);
or U8858 (N_8858,N_8107,N_8371);
nor U8859 (N_8859,N_8247,N_8356);
xor U8860 (N_8860,N_8490,N_8018);
xnor U8861 (N_8861,N_8363,N_8395);
nand U8862 (N_8862,N_8157,N_8456);
xnor U8863 (N_8863,N_8370,N_8411);
and U8864 (N_8864,N_8035,N_8179);
xnor U8865 (N_8865,N_8189,N_8227);
nand U8866 (N_8866,N_8105,N_8027);
xor U8867 (N_8867,N_8410,N_8124);
xnor U8868 (N_8868,N_8247,N_8088);
nor U8869 (N_8869,N_8221,N_8379);
or U8870 (N_8870,N_8339,N_8165);
nor U8871 (N_8871,N_8274,N_8196);
nand U8872 (N_8872,N_8112,N_8471);
xnor U8873 (N_8873,N_8339,N_8283);
xor U8874 (N_8874,N_8070,N_8455);
xnor U8875 (N_8875,N_8196,N_8144);
and U8876 (N_8876,N_8358,N_8430);
nand U8877 (N_8877,N_8256,N_8306);
and U8878 (N_8878,N_8478,N_8049);
xnor U8879 (N_8879,N_8422,N_8263);
and U8880 (N_8880,N_8177,N_8206);
nand U8881 (N_8881,N_8036,N_8459);
nand U8882 (N_8882,N_8184,N_8086);
and U8883 (N_8883,N_8415,N_8490);
nand U8884 (N_8884,N_8461,N_8413);
or U8885 (N_8885,N_8320,N_8236);
and U8886 (N_8886,N_8349,N_8138);
nand U8887 (N_8887,N_8427,N_8364);
nand U8888 (N_8888,N_8252,N_8099);
nand U8889 (N_8889,N_8019,N_8171);
nor U8890 (N_8890,N_8234,N_8438);
or U8891 (N_8891,N_8094,N_8119);
or U8892 (N_8892,N_8392,N_8217);
xor U8893 (N_8893,N_8083,N_8246);
and U8894 (N_8894,N_8303,N_8107);
nand U8895 (N_8895,N_8185,N_8150);
xnor U8896 (N_8896,N_8277,N_8286);
xnor U8897 (N_8897,N_8184,N_8202);
xnor U8898 (N_8898,N_8389,N_8213);
or U8899 (N_8899,N_8105,N_8210);
nor U8900 (N_8900,N_8248,N_8245);
nor U8901 (N_8901,N_8018,N_8215);
nor U8902 (N_8902,N_8164,N_8117);
nand U8903 (N_8903,N_8016,N_8311);
nor U8904 (N_8904,N_8137,N_8467);
or U8905 (N_8905,N_8178,N_8003);
and U8906 (N_8906,N_8170,N_8018);
xor U8907 (N_8907,N_8426,N_8006);
and U8908 (N_8908,N_8414,N_8478);
nand U8909 (N_8909,N_8038,N_8309);
xnor U8910 (N_8910,N_8242,N_8162);
nor U8911 (N_8911,N_8032,N_8481);
nand U8912 (N_8912,N_8369,N_8451);
nand U8913 (N_8913,N_8319,N_8050);
nor U8914 (N_8914,N_8433,N_8204);
nor U8915 (N_8915,N_8202,N_8286);
xor U8916 (N_8916,N_8048,N_8425);
or U8917 (N_8917,N_8361,N_8008);
and U8918 (N_8918,N_8294,N_8376);
nor U8919 (N_8919,N_8268,N_8378);
nand U8920 (N_8920,N_8113,N_8399);
xor U8921 (N_8921,N_8225,N_8338);
nor U8922 (N_8922,N_8496,N_8050);
xnor U8923 (N_8923,N_8208,N_8331);
xnor U8924 (N_8924,N_8218,N_8484);
and U8925 (N_8925,N_8337,N_8051);
nand U8926 (N_8926,N_8099,N_8005);
or U8927 (N_8927,N_8075,N_8365);
xnor U8928 (N_8928,N_8182,N_8282);
nor U8929 (N_8929,N_8065,N_8138);
or U8930 (N_8930,N_8463,N_8104);
nand U8931 (N_8931,N_8301,N_8247);
nand U8932 (N_8932,N_8182,N_8050);
and U8933 (N_8933,N_8280,N_8148);
nand U8934 (N_8934,N_8321,N_8099);
and U8935 (N_8935,N_8237,N_8299);
and U8936 (N_8936,N_8053,N_8317);
xor U8937 (N_8937,N_8482,N_8449);
nand U8938 (N_8938,N_8061,N_8450);
or U8939 (N_8939,N_8030,N_8097);
xor U8940 (N_8940,N_8482,N_8188);
and U8941 (N_8941,N_8484,N_8325);
xor U8942 (N_8942,N_8109,N_8018);
nand U8943 (N_8943,N_8057,N_8066);
nor U8944 (N_8944,N_8313,N_8364);
nor U8945 (N_8945,N_8234,N_8182);
xor U8946 (N_8946,N_8019,N_8491);
nor U8947 (N_8947,N_8144,N_8299);
nor U8948 (N_8948,N_8075,N_8264);
or U8949 (N_8949,N_8151,N_8241);
and U8950 (N_8950,N_8163,N_8337);
or U8951 (N_8951,N_8428,N_8315);
nor U8952 (N_8952,N_8233,N_8170);
xnor U8953 (N_8953,N_8118,N_8131);
nor U8954 (N_8954,N_8002,N_8016);
and U8955 (N_8955,N_8078,N_8467);
and U8956 (N_8956,N_8354,N_8257);
nor U8957 (N_8957,N_8387,N_8135);
xor U8958 (N_8958,N_8201,N_8137);
nor U8959 (N_8959,N_8114,N_8149);
nor U8960 (N_8960,N_8271,N_8405);
or U8961 (N_8961,N_8108,N_8435);
nand U8962 (N_8962,N_8073,N_8304);
nor U8963 (N_8963,N_8391,N_8256);
nand U8964 (N_8964,N_8380,N_8492);
and U8965 (N_8965,N_8195,N_8467);
xnor U8966 (N_8966,N_8225,N_8322);
and U8967 (N_8967,N_8417,N_8331);
and U8968 (N_8968,N_8260,N_8034);
xor U8969 (N_8969,N_8293,N_8035);
or U8970 (N_8970,N_8400,N_8241);
or U8971 (N_8971,N_8006,N_8004);
nor U8972 (N_8972,N_8233,N_8017);
nor U8973 (N_8973,N_8007,N_8350);
xor U8974 (N_8974,N_8315,N_8232);
nand U8975 (N_8975,N_8269,N_8102);
and U8976 (N_8976,N_8266,N_8114);
or U8977 (N_8977,N_8274,N_8478);
nor U8978 (N_8978,N_8299,N_8288);
or U8979 (N_8979,N_8495,N_8113);
nand U8980 (N_8980,N_8044,N_8089);
xor U8981 (N_8981,N_8408,N_8202);
nor U8982 (N_8982,N_8276,N_8102);
nor U8983 (N_8983,N_8467,N_8254);
or U8984 (N_8984,N_8449,N_8304);
or U8985 (N_8985,N_8328,N_8443);
nand U8986 (N_8986,N_8146,N_8281);
or U8987 (N_8987,N_8272,N_8439);
xor U8988 (N_8988,N_8248,N_8232);
nor U8989 (N_8989,N_8250,N_8286);
xor U8990 (N_8990,N_8246,N_8457);
nor U8991 (N_8991,N_8363,N_8059);
nand U8992 (N_8992,N_8051,N_8461);
xor U8993 (N_8993,N_8089,N_8381);
or U8994 (N_8994,N_8126,N_8230);
or U8995 (N_8995,N_8002,N_8349);
and U8996 (N_8996,N_8124,N_8363);
and U8997 (N_8997,N_8493,N_8191);
and U8998 (N_8998,N_8268,N_8333);
and U8999 (N_8999,N_8182,N_8382);
nor U9000 (N_9000,N_8923,N_8959);
and U9001 (N_9001,N_8551,N_8518);
nor U9002 (N_9002,N_8787,N_8835);
or U9003 (N_9003,N_8912,N_8593);
nor U9004 (N_9004,N_8513,N_8503);
nor U9005 (N_9005,N_8798,N_8780);
nand U9006 (N_9006,N_8918,N_8693);
xor U9007 (N_9007,N_8872,N_8830);
nand U9008 (N_9008,N_8839,N_8633);
xor U9009 (N_9009,N_8816,N_8608);
nor U9010 (N_9010,N_8535,N_8519);
or U9011 (N_9011,N_8751,N_8699);
or U9012 (N_9012,N_8777,N_8901);
nand U9013 (N_9013,N_8555,N_8874);
nand U9014 (N_9014,N_8623,N_8612);
nand U9015 (N_9015,N_8720,N_8865);
or U9016 (N_9016,N_8610,N_8711);
and U9017 (N_9017,N_8613,N_8997);
nor U9018 (N_9018,N_8685,N_8534);
and U9019 (N_9019,N_8909,N_8927);
or U9020 (N_9020,N_8667,N_8826);
nor U9021 (N_9021,N_8524,N_8804);
xnor U9022 (N_9022,N_8682,N_8646);
nor U9023 (N_9023,N_8680,N_8989);
and U9024 (N_9024,N_8955,N_8630);
nor U9025 (N_9025,N_8726,N_8974);
nand U9026 (N_9026,N_8553,N_8913);
xnor U9027 (N_9027,N_8779,N_8517);
nand U9028 (N_9028,N_8601,N_8728);
xor U9029 (N_9029,N_8893,N_8514);
or U9030 (N_9030,N_8984,N_8626);
xor U9031 (N_9031,N_8676,N_8960);
nand U9032 (N_9032,N_8812,N_8785);
nand U9033 (N_9033,N_8618,N_8578);
xnor U9034 (N_9034,N_8577,N_8669);
and U9035 (N_9035,N_8888,N_8745);
nor U9036 (N_9036,N_8597,N_8805);
nor U9037 (N_9037,N_8713,N_8515);
and U9038 (N_9038,N_8871,N_8908);
or U9039 (N_9039,N_8994,N_8749);
or U9040 (N_9040,N_8701,N_8627);
xnor U9041 (N_9041,N_8890,N_8940);
and U9042 (N_9042,N_8600,N_8584);
or U9043 (N_9043,N_8716,N_8860);
nor U9044 (N_9044,N_8684,N_8760);
nand U9045 (N_9045,N_8722,N_8536);
xnor U9046 (N_9046,N_8730,N_8828);
xnor U9047 (N_9047,N_8574,N_8567);
nand U9048 (N_9048,N_8710,N_8793);
xnor U9049 (N_9049,N_8928,N_8939);
nor U9050 (N_9050,N_8668,N_8500);
nand U9051 (N_9051,N_8796,N_8604);
nand U9052 (N_9052,N_8547,N_8573);
and U9053 (N_9053,N_8824,N_8752);
xnor U9054 (N_9054,N_8673,N_8857);
and U9055 (N_9055,N_8647,N_8588);
nand U9056 (N_9056,N_8958,N_8611);
and U9057 (N_9057,N_8837,N_8671);
nor U9058 (N_9058,N_8689,N_8823);
nand U9059 (N_9059,N_8877,N_8954);
nand U9060 (N_9060,N_8763,N_8818);
or U9061 (N_9061,N_8972,N_8995);
or U9062 (N_9062,N_8963,N_8851);
nor U9063 (N_9063,N_8964,N_8866);
nor U9064 (N_9064,N_8813,N_8821);
nand U9065 (N_9065,N_8664,N_8781);
xor U9066 (N_9066,N_8742,N_8841);
and U9067 (N_9067,N_8530,N_8541);
xnor U9068 (N_9068,N_8846,N_8655);
or U9069 (N_9069,N_8591,N_8596);
and U9070 (N_9070,N_8993,N_8863);
and U9071 (N_9071,N_8703,N_8592);
and U9072 (N_9072,N_8620,N_8714);
and U9073 (N_9073,N_8783,N_8854);
or U9074 (N_9074,N_8746,N_8768);
nor U9075 (N_9075,N_8543,N_8904);
or U9076 (N_9076,N_8665,N_8521);
xor U9077 (N_9077,N_8510,N_8786);
nand U9078 (N_9078,N_8843,N_8661);
nor U9079 (N_9079,N_8965,N_8905);
and U9080 (N_9080,N_8801,N_8979);
nor U9081 (N_9081,N_8545,N_8876);
xnor U9082 (N_9082,N_8643,N_8946);
or U9083 (N_9083,N_8625,N_8750);
xor U9084 (N_9084,N_8624,N_8791);
or U9085 (N_9085,N_8914,N_8753);
and U9086 (N_9086,N_8983,N_8629);
nand U9087 (N_9087,N_8886,N_8638);
and U9088 (N_9088,N_8687,N_8840);
nor U9089 (N_9089,N_8700,N_8968);
nand U9090 (N_9090,N_8557,N_8970);
nand U9091 (N_9091,N_8617,N_8819);
nor U9092 (N_9092,N_8986,N_8754);
nor U9093 (N_9093,N_8729,N_8867);
or U9094 (N_9094,N_8585,N_8660);
nor U9095 (N_9095,N_8774,N_8769);
xnor U9096 (N_9096,N_8540,N_8741);
nor U9097 (N_9097,N_8598,N_8898);
xor U9098 (N_9098,N_8602,N_8707);
nor U9099 (N_9099,N_8675,N_8885);
nand U9100 (N_9100,N_8506,N_8947);
or U9101 (N_9101,N_8508,N_8875);
or U9102 (N_9102,N_8672,N_8897);
or U9103 (N_9103,N_8653,N_8747);
or U9104 (N_9104,N_8827,N_8836);
nand U9105 (N_9105,N_8579,N_8896);
xnor U9106 (N_9106,N_8645,N_8926);
or U9107 (N_9107,N_8554,N_8686);
nor U9108 (N_9108,N_8695,N_8757);
nand U9109 (N_9109,N_8792,N_8847);
or U9110 (N_9110,N_8985,N_8528);
or U9111 (N_9111,N_8637,N_8802);
nand U9112 (N_9112,N_8771,N_8733);
nand U9113 (N_9113,N_8938,N_8723);
and U9114 (N_9114,N_8690,N_8657);
nand U9115 (N_9115,N_8527,N_8772);
or U9116 (N_9116,N_8520,N_8599);
nand U9117 (N_9117,N_8755,N_8920);
or U9118 (N_9118,N_8868,N_8916);
or U9119 (N_9119,N_8589,N_8762);
xor U9120 (N_9120,N_8734,N_8834);
nand U9121 (N_9121,N_8878,N_8869);
nand U9122 (N_9122,N_8539,N_8512);
nand U9123 (N_9123,N_8619,N_8971);
xnor U9124 (N_9124,N_8932,N_8586);
or U9125 (N_9125,N_8571,N_8632);
and U9126 (N_9126,N_8806,N_8580);
or U9127 (N_9127,N_8873,N_8815);
nand U9128 (N_9128,N_8855,N_8807);
nand U9129 (N_9129,N_8825,N_8859);
or U9130 (N_9130,N_8694,N_8709);
and U9131 (N_9131,N_8704,N_8744);
and U9132 (N_9132,N_8509,N_8894);
or U9133 (N_9133,N_8556,N_8563);
or U9134 (N_9134,N_8537,N_8737);
xnor U9135 (N_9135,N_8910,N_8950);
xnor U9136 (N_9136,N_8549,N_8935);
nand U9137 (N_9137,N_8583,N_8882);
nor U9138 (N_9138,N_8507,N_8548);
xnor U9139 (N_9139,N_8748,N_8969);
xor U9140 (N_9140,N_8799,N_8849);
and U9141 (N_9141,N_8558,N_8915);
xnor U9142 (N_9142,N_8953,N_8797);
or U9143 (N_9143,N_8727,N_8856);
nand U9144 (N_9144,N_8505,N_8991);
nor U9145 (N_9145,N_8999,N_8952);
nor U9146 (N_9146,N_8560,N_8717);
xor U9147 (N_9147,N_8765,N_8666);
xnor U9148 (N_9148,N_8538,N_8990);
nor U9149 (N_9149,N_8654,N_8688);
xor U9150 (N_9150,N_8870,N_8708);
xnor U9151 (N_9151,N_8622,N_8973);
and U9152 (N_9152,N_8758,N_8670);
or U9153 (N_9153,N_8552,N_8853);
xnor U9154 (N_9154,N_8697,N_8766);
and U9155 (N_9155,N_8956,N_8924);
nand U9156 (N_9156,N_8649,N_8790);
or U9157 (N_9157,N_8844,N_8523);
nor U9158 (N_9158,N_8677,N_8606);
xnor U9159 (N_9159,N_8966,N_8941);
or U9160 (N_9160,N_8900,N_8712);
or U9161 (N_9161,N_8715,N_8581);
and U9162 (N_9162,N_8800,N_8982);
or U9163 (N_9163,N_8562,N_8767);
nor U9164 (N_9164,N_8842,N_8829);
and U9165 (N_9165,N_8858,N_8702);
xor U9166 (N_9166,N_8569,N_8681);
nand U9167 (N_9167,N_8850,N_8788);
and U9168 (N_9168,N_8895,N_8852);
nand U9169 (N_9169,N_8761,N_8811);
nand U9170 (N_9170,N_8822,N_8561);
xnor U9171 (N_9171,N_8921,N_8810);
or U9172 (N_9172,N_8595,N_8731);
nand U9173 (N_9173,N_8683,N_8609);
nand U9174 (N_9174,N_8678,N_8582);
nor U9175 (N_9175,N_8902,N_8640);
nand U9176 (N_9176,N_8962,N_8568);
xnor U9177 (N_9177,N_8881,N_8501);
and U9178 (N_9178,N_8735,N_8725);
nand U9179 (N_9179,N_8739,N_8906);
and U9180 (N_9180,N_8542,N_8516);
or U9181 (N_9181,N_8884,N_8502);
or U9182 (N_9182,N_8566,N_8845);
and U9183 (N_9183,N_8831,N_8559);
nand U9184 (N_9184,N_8736,N_8706);
xor U9185 (N_9185,N_8838,N_8978);
nand U9186 (N_9186,N_8603,N_8719);
nand U9187 (N_9187,N_8764,N_8576);
and U9188 (N_9188,N_8980,N_8526);
xor U9189 (N_9189,N_8614,N_8705);
or U9190 (N_9190,N_8642,N_8948);
xor U9191 (N_9191,N_8773,N_8907);
or U9192 (N_9192,N_8756,N_8759);
xnor U9193 (N_9193,N_8943,N_8892);
nor U9194 (N_9194,N_8889,N_8644);
nor U9195 (N_9195,N_8981,N_8662);
xor U9196 (N_9196,N_8652,N_8778);
nand U9197 (N_9197,N_8891,N_8590);
and U9198 (N_9198,N_8658,N_8605);
nor U9199 (N_9199,N_8937,N_8532);
and U9200 (N_9200,N_8621,N_8833);
xnor U9201 (N_9201,N_8794,N_8951);
nand U9202 (N_9202,N_8988,N_8814);
and U9203 (N_9203,N_8529,N_8977);
or U9204 (N_9204,N_8817,N_8639);
and U9205 (N_9205,N_8848,N_8934);
nor U9206 (N_9206,N_8936,N_8957);
xor U9207 (N_9207,N_8674,N_8992);
or U9208 (N_9208,N_8533,N_8911);
or U9209 (N_9209,N_8740,N_8930);
nand U9210 (N_9210,N_8925,N_8864);
and U9211 (N_9211,N_8546,N_8987);
and U9212 (N_9212,N_8975,N_8775);
nor U9213 (N_9213,N_8564,N_8522);
nor U9214 (N_9214,N_8732,N_8616);
nor U9215 (N_9215,N_8883,N_8572);
or U9216 (N_9216,N_8663,N_8743);
and U9217 (N_9217,N_8967,N_8656);
nor U9218 (N_9218,N_8650,N_8544);
nand U9219 (N_9219,N_8679,N_8776);
and U9220 (N_9220,N_8789,N_8721);
nand U9221 (N_9221,N_8738,N_8651);
or U9222 (N_9222,N_8659,N_8724);
and U9223 (N_9223,N_8628,N_8770);
nand U9224 (N_9224,N_8976,N_8696);
and U9225 (N_9225,N_8615,N_8820);
nor U9226 (N_9226,N_8784,N_8698);
nor U9227 (N_9227,N_8795,N_8631);
nor U9228 (N_9228,N_8504,N_8903);
nand U9229 (N_9229,N_8525,N_8899);
or U9230 (N_9230,N_8917,N_8691);
nor U9231 (N_9231,N_8949,N_8587);
nand U9232 (N_9232,N_8945,N_8692);
or U9233 (N_9233,N_8648,N_8636);
nor U9234 (N_9234,N_8998,N_8861);
nand U9235 (N_9235,N_8607,N_8880);
or U9236 (N_9236,N_8570,N_8511);
xor U9237 (N_9237,N_8565,N_8635);
and U9238 (N_9238,N_8996,N_8550);
and U9239 (N_9239,N_8919,N_8808);
nand U9240 (N_9240,N_8809,N_8887);
or U9241 (N_9241,N_8832,N_8931);
xor U9242 (N_9242,N_8933,N_8942);
nor U9243 (N_9243,N_8922,N_8594);
nand U9244 (N_9244,N_8944,N_8782);
or U9245 (N_9245,N_8718,N_8641);
xor U9246 (N_9246,N_8634,N_8961);
and U9247 (N_9247,N_8929,N_8575);
and U9248 (N_9248,N_8879,N_8803);
nand U9249 (N_9249,N_8862,N_8531);
nor U9250 (N_9250,N_8634,N_8898);
nor U9251 (N_9251,N_8921,N_8733);
xor U9252 (N_9252,N_8921,N_8804);
nand U9253 (N_9253,N_8736,N_8658);
or U9254 (N_9254,N_8655,N_8943);
nand U9255 (N_9255,N_8728,N_8696);
xnor U9256 (N_9256,N_8960,N_8581);
xnor U9257 (N_9257,N_8859,N_8641);
nor U9258 (N_9258,N_8991,N_8572);
xor U9259 (N_9259,N_8891,N_8933);
nand U9260 (N_9260,N_8650,N_8566);
or U9261 (N_9261,N_8662,N_8728);
xor U9262 (N_9262,N_8527,N_8523);
nor U9263 (N_9263,N_8676,N_8596);
or U9264 (N_9264,N_8715,N_8604);
nand U9265 (N_9265,N_8795,N_8512);
nand U9266 (N_9266,N_8830,N_8960);
nor U9267 (N_9267,N_8944,N_8931);
nor U9268 (N_9268,N_8828,N_8723);
nand U9269 (N_9269,N_8818,N_8568);
nand U9270 (N_9270,N_8771,N_8748);
nor U9271 (N_9271,N_8585,N_8978);
xnor U9272 (N_9272,N_8593,N_8730);
and U9273 (N_9273,N_8703,N_8887);
or U9274 (N_9274,N_8807,N_8695);
and U9275 (N_9275,N_8957,N_8800);
nand U9276 (N_9276,N_8902,N_8992);
or U9277 (N_9277,N_8906,N_8911);
and U9278 (N_9278,N_8826,N_8938);
xor U9279 (N_9279,N_8622,N_8905);
xor U9280 (N_9280,N_8629,N_8690);
xor U9281 (N_9281,N_8811,N_8841);
and U9282 (N_9282,N_8741,N_8574);
xor U9283 (N_9283,N_8991,N_8730);
nand U9284 (N_9284,N_8781,N_8603);
xor U9285 (N_9285,N_8775,N_8579);
or U9286 (N_9286,N_8998,N_8589);
nor U9287 (N_9287,N_8684,N_8732);
xor U9288 (N_9288,N_8986,N_8708);
or U9289 (N_9289,N_8613,N_8773);
xor U9290 (N_9290,N_8509,N_8767);
nor U9291 (N_9291,N_8875,N_8796);
xnor U9292 (N_9292,N_8749,N_8730);
nand U9293 (N_9293,N_8900,N_8776);
and U9294 (N_9294,N_8830,N_8524);
and U9295 (N_9295,N_8977,N_8973);
nand U9296 (N_9296,N_8582,N_8982);
xnor U9297 (N_9297,N_8971,N_8875);
nor U9298 (N_9298,N_8672,N_8766);
and U9299 (N_9299,N_8754,N_8663);
nand U9300 (N_9300,N_8642,N_8994);
and U9301 (N_9301,N_8771,N_8863);
or U9302 (N_9302,N_8547,N_8579);
and U9303 (N_9303,N_8897,N_8777);
nor U9304 (N_9304,N_8678,N_8834);
nand U9305 (N_9305,N_8548,N_8534);
and U9306 (N_9306,N_8855,N_8628);
and U9307 (N_9307,N_8534,N_8561);
or U9308 (N_9308,N_8714,N_8616);
or U9309 (N_9309,N_8644,N_8987);
and U9310 (N_9310,N_8654,N_8702);
nor U9311 (N_9311,N_8942,N_8842);
nor U9312 (N_9312,N_8546,N_8953);
nand U9313 (N_9313,N_8891,N_8529);
and U9314 (N_9314,N_8684,N_8902);
nand U9315 (N_9315,N_8753,N_8585);
and U9316 (N_9316,N_8912,N_8837);
xnor U9317 (N_9317,N_8638,N_8579);
nand U9318 (N_9318,N_8648,N_8723);
xnor U9319 (N_9319,N_8993,N_8576);
or U9320 (N_9320,N_8751,N_8566);
and U9321 (N_9321,N_8622,N_8593);
and U9322 (N_9322,N_8562,N_8902);
and U9323 (N_9323,N_8738,N_8868);
or U9324 (N_9324,N_8571,N_8830);
nor U9325 (N_9325,N_8983,N_8787);
nor U9326 (N_9326,N_8976,N_8902);
nand U9327 (N_9327,N_8958,N_8924);
or U9328 (N_9328,N_8821,N_8996);
nand U9329 (N_9329,N_8679,N_8617);
nand U9330 (N_9330,N_8574,N_8808);
or U9331 (N_9331,N_8991,N_8839);
nand U9332 (N_9332,N_8891,N_8987);
xnor U9333 (N_9333,N_8879,N_8801);
or U9334 (N_9334,N_8612,N_8726);
or U9335 (N_9335,N_8654,N_8758);
nand U9336 (N_9336,N_8943,N_8726);
nor U9337 (N_9337,N_8894,N_8734);
nor U9338 (N_9338,N_8863,N_8638);
nor U9339 (N_9339,N_8947,N_8655);
or U9340 (N_9340,N_8888,N_8785);
nand U9341 (N_9341,N_8579,N_8825);
or U9342 (N_9342,N_8809,N_8591);
and U9343 (N_9343,N_8655,N_8735);
or U9344 (N_9344,N_8769,N_8842);
nor U9345 (N_9345,N_8566,N_8909);
nor U9346 (N_9346,N_8681,N_8891);
nand U9347 (N_9347,N_8555,N_8648);
or U9348 (N_9348,N_8870,N_8649);
nor U9349 (N_9349,N_8509,N_8884);
xor U9350 (N_9350,N_8574,N_8674);
nor U9351 (N_9351,N_8677,N_8538);
nor U9352 (N_9352,N_8999,N_8548);
nor U9353 (N_9353,N_8517,N_8974);
xor U9354 (N_9354,N_8816,N_8615);
xnor U9355 (N_9355,N_8560,N_8882);
or U9356 (N_9356,N_8636,N_8559);
nor U9357 (N_9357,N_8788,N_8775);
nor U9358 (N_9358,N_8666,N_8533);
nor U9359 (N_9359,N_8736,N_8525);
xnor U9360 (N_9360,N_8812,N_8578);
and U9361 (N_9361,N_8932,N_8864);
nor U9362 (N_9362,N_8931,N_8967);
and U9363 (N_9363,N_8568,N_8718);
xor U9364 (N_9364,N_8511,N_8905);
or U9365 (N_9365,N_8729,N_8922);
or U9366 (N_9366,N_8960,N_8568);
nand U9367 (N_9367,N_8954,N_8911);
nand U9368 (N_9368,N_8893,N_8934);
xor U9369 (N_9369,N_8750,N_8985);
and U9370 (N_9370,N_8865,N_8664);
and U9371 (N_9371,N_8978,N_8733);
nand U9372 (N_9372,N_8798,N_8501);
and U9373 (N_9373,N_8857,N_8692);
and U9374 (N_9374,N_8707,N_8970);
xor U9375 (N_9375,N_8749,N_8693);
xor U9376 (N_9376,N_8931,N_8732);
nor U9377 (N_9377,N_8649,N_8513);
nand U9378 (N_9378,N_8559,N_8627);
or U9379 (N_9379,N_8976,N_8720);
nor U9380 (N_9380,N_8747,N_8836);
nand U9381 (N_9381,N_8603,N_8547);
and U9382 (N_9382,N_8994,N_8986);
nor U9383 (N_9383,N_8904,N_8844);
xor U9384 (N_9384,N_8865,N_8881);
nor U9385 (N_9385,N_8504,N_8820);
nor U9386 (N_9386,N_8906,N_8596);
xor U9387 (N_9387,N_8719,N_8988);
nand U9388 (N_9388,N_8758,N_8835);
nor U9389 (N_9389,N_8712,N_8793);
nor U9390 (N_9390,N_8860,N_8588);
xor U9391 (N_9391,N_8830,N_8889);
xor U9392 (N_9392,N_8734,N_8887);
or U9393 (N_9393,N_8663,N_8506);
and U9394 (N_9394,N_8712,N_8855);
and U9395 (N_9395,N_8785,N_8958);
and U9396 (N_9396,N_8668,N_8845);
or U9397 (N_9397,N_8948,N_8555);
or U9398 (N_9398,N_8940,N_8963);
or U9399 (N_9399,N_8749,N_8544);
or U9400 (N_9400,N_8675,N_8737);
and U9401 (N_9401,N_8652,N_8934);
nand U9402 (N_9402,N_8822,N_8632);
nand U9403 (N_9403,N_8878,N_8695);
xor U9404 (N_9404,N_8979,N_8929);
nand U9405 (N_9405,N_8518,N_8829);
nand U9406 (N_9406,N_8575,N_8716);
nor U9407 (N_9407,N_8537,N_8820);
or U9408 (N_9408,N_8766,N_8838);
and U9409 (N_9409,N_8853,N_8630);
xnor U9410 (N_9410,N_8870,N_8534);
nand U9411 (N_9411,N_8809,N_8909);
xnor U9412 (N_9412,N_8976,N_8762);
or U9413 (N_9413,N_8768,N_8690);
and U9414 (N_9414,N_8678,N_8863);
nor U9415 (N_9415,N_8575,N_8712);
nand U9416 (N_9416,N_8534,N_8746);
xor U9417 (N_9417,N_8680,N_8964);
xor U9418 (N_9418,N_8646,N_8538);
xor U9419 (N_9419,N_8966,N_8744);
nor U9420 (N_9420,N_8740,N_8516);
and U9421 (N_9421,N_8855,N_8738);
xor U9422 (N_9422,N_8908,N_8955);
xor U9423 (N_9423,N_8911,N_8541);
and U9424 (N_9424,N_8976,N_8512);
xor U9425 (N_9425,N_8871,N_8581);
nand U9426 (N_9426,N_8896,N_8936);
or U9427 (N_9427,N_8897,N_8669);
nor U9428 (N_9428,N_8693,N_8630);
nand U9429 (N_9429,N_8837,N_8758);
and U9430 (N_9430,N_8866,N_8911);
xnor U9431 (N_9431,N_8916,N_8706);
nand U9432 (N_9432,N_8972,N_8575);
xnor U9433 (N_9433,N_8768,N_8844);
nand U9434 (N_9434,N_8819,N_8702);
and U9435 (N_9435,N_8789,N_8684);
xnor U9436 (N_9436,N_8575,N_8702);
nor U9437 (N_9437,N_8648,N_8890);
and U9438 (N_9438,N_8795,N_8937);
nand U9439 (N_9439,N_8875,N_8664);
nor U9440 (N_9440,N_8879,N_8818);
or U9441 (N_9441,N_8995,N_8504);
and U9442 (N_9442,N_8779,N_8530);
and U9443 (N_9443,N_8683,N_8875);
nand U9444 (N_9444,N_8708,N_8928);
nand U9445 (N_9445,N_8534,N_8539);
or U9446 (N_9446,N_8632,N_8607);
nand U9447 (N_9447,N_8650,N_8886);
nand U9448 (N_9448,N_8501,N_8879);
or U9449 (N_9449,N_8692,N_8988);
nor U9450 (N_9450,N_8788,N_8765);
or U9451 (N_9451,N_8818,N_8683);
or U9452 (N_9452,N_8917,N_8722);
or U9453 (N_9453,N_8949,N_8803);
or U9454 (N_9454,N_8967,N_8677);
or U9455 (N_9455,N_8753,N_8968);
nand U9456 (N_9456,N_8597,N_8817);
and U9457 (N_9457,N_8531,N_8897);
nor U9458 (N_9458,N_8637,N_8573);
and U9459 (N_9459,N_8673,N_8578);
xor U9460 (N_9460,N_8931,N_8938);
or U9461 (N_9461,N_8849,N_8905);
nor U9462 (N_9462,N_8642,N_8645);
or U9463 (N_9463,N_8934,N_8518);
nand U9464 (N_9464,N_8645,N_8605);
nand U9465 (N_9465,N_8959,N_8976);
and U9466 (N_9466,N_8984,N_8700);
or U9467 (N_9467,N_8740,N_8582);
nand U9468 (N_9468,N_8598,N_8536);
xor U9469 (N_9469,N_8511,N_8526);
xnor U9470 (N_9470,N_8501,N_8651);
and U9471 (N_9471,N_8517,N_8579);
or U9472 (N_9472,N_8745,N_8563);
xnor U9473 (N_9473,N_8912,N_8544);
nand U9474 (N_9474,N_8506,N_8633);
xor U9475 (N_9475,N_8612,N_8937);
or U9476 (N_9476,N_8971,N_8615);
nand U9477 (N_9477,N_8949,N_8628);
nor U9478 (N_9478,N_8509,N_8588);
or U9479 (N_9479,N_8622,N_8743);
nor U9480 (N_9480,N_8637,N_8635);
xnor U9481 (N_9481,N_8714,N_8736);
nor U9482 (N_9482,N_8592,N_8682);
nor U9483 (N_9483,N_8680,N_8891);
and U9484 (N_9484,N_8739,N_8508);
and U9485 (N_9485,N_8756,N_8623);
nor U9486 (N_9486,N_8591,N_8699);
nor U9487 (N_9487,N_8937,N_8871);
or U9488 (N_9488,N_8612,N_8927);
or U9489 (N_9489,N_8976,N_8813);
nor U9490 (N_9490,N_8914,N_8895);
xnor U9491 (N_9491,N_8937,N_8753);
nand U9492 (N_9492,N_8900,N_8626);
nor U9493 (N_9493,N_8862,N_8829);
nor U9494 (N_9494,N_8996,N_8771);
nand U9495 (N_9495,N_8843,N_8627);
and U9496 (N_9496,N_8883,N_8992);
nor U9497 (N_9497,N_8876,N_8991);
xnor U9498 (N_9498,N_8840,N_8634);
or U9499 (N_9499,N_8983,N_8669);
nor U9500 (N_9500,N_9076,N_9451);
or U9501 (N_9501,N_9067,N_9004);
xnor U9502 (N_9502,N_9392,N_9255);
and U9503 (N_9503,N_9213,N_9128);
nand U9504 (N_9504,N_9352,N_9404);
or U9505 (N_9505,N_9216,N_9252);
nor U9506 (N_9506,N_9228,N_9242);
xnor U9507 (N_9507,N_9139,N_9312);
nor U9508 (N_9508,N_9092,N_9140);
nand U9509 (N_9509,N_9165,N_9401);
xor U9510 (N_9510,N_9259,N_9211);
and U9511 (N_9511,N_9097,N_9008);
nand U9512 (N_9512,N_9298,N_9224);
xnor U9513 (N_9513,N_9390,N_9247);
and U9514 (N_9514,N_9494,N_9210);
nand U9515 (N_9515,N_9031,N_9305);
nor U9516 (N_9516,N_9274,N_9275);
xor U9517 (N_9517,N_9053,N_9142);
xnor U9518 (N_9518,N_9409,N_9283);
and U9519 (N_9519,N_9360,N_9416);
nand U9520 (N_9520,N_9129,N_9127);
xor U9521 (N_9521,N_9002,N_9119);
xor U9522 (N_9522,N_9383,N_9443);
xnor U9523 (N_9523,N_9108,N_9209);
xor U9524 (N_9524,N_9282,N_9445);
or U9525 (N_9525,N_9019,N_9174);
nand U9526 (N_9526,N_9368,N_9233);
or U9527 (N_9527,N_9199,N_9299);
and U9528 (N_9528,N_9302,N_9171);
or U9529 (N_9529,N_9057,N_9315);
xnor U9530 (N_9530,N_9395,N_9001);
or U9531 (N_9531,N_9332,N_9202);
nand U9532 (N_9532,N_9162,N_9191);
or U9533 (N_9533,N_9079,N_9195);
xor U9534 (N_9534,N_9354,N_9058);
or U9535 (N_9535,N_9487,N_9015);
nand U9536 (N_9536,N_9263,N_9101);
or U9537 (N_9537,N_9267,N_9133);
or U9538 (N_9538,N_9449,N_9313);
nor U9539 (N_9539,N_9178,N_9244);
nand U9540 (N_9540,N_9326,N_9388);
nor U9541 (N_9541,N_9272,N_9007);
nand U9542 (N_9542,N_9033,N_9422);
or U9543 (N_9543,N_9251,N_9218);
nand U9544 (N_9544,N_9406,N_9116);
or U9545 (N_9545,N_9304,N_9175);
xor U9546 (N_9546,N_9037,N_9464);
or U9547 (N_9547,N_9232,N_9093);
or U9548 (N_9548,N_9417,N_9363);
and U9549 (N_9549,N_9027,N_9441);
nor U9550 (N_9550,N_9324,N_9215);
or U9551 (N_9551,N_9163,N_9415);
nor U9552 (N_9552,N_9138,N_9353);
xnor U9553 (N_9553,N_9488,N_9229);
and U9554 (N_9554,N_9239,N_9080);
or U9555 (N_9555,N_9009,N_9351);
nand U9556 (N_9556,N_9219,N_9125);
xnor U9557 (N_9557,N_9427,N_9414);
or U9558 (N_9558,N_9480,N_9072);
xnor U9559 (N_9559,N_9418,N_9468);
nor U9560 (N_9560,N_9230,N_9316);
nand U9561 (N_9561,N_9448,N_9447);
or U9562 (N_9562,N_9115,N_9379);
xnor U9563 (N_9563,N_9311,N_9056);
nor U9564 (N_9564,N_9087,N_9065);
and U9565 (N_9565,N_9021,N_9350);
and U9566 (N_9566,N_9490,N_9234);
nor U9567 (N_9567,N_9336,N_9075);
xnor U9568 (N_9568,N_9003,N_9329);
or U9569 (N_9569,N_9039,N_9457);
xor U9570 (N_9570,N_9249,N_9179);
nand U9571 (N_9571,N_9044,N_9107);
and U9572 (N_9572,N_9201,N_9187);
nand U9573 (N_9573,N_9170,N_9277);
nor U9574 (N_9574,N_9279,N_9258);
and U9575 (N_9575,N_9069,N_9439);
xnor U9576 (N_9576,N_9180,N_9126);
or U9577 (N_9577,N_9102,N_9454);
xnor U9578 (N_9578,N_9483,N_9032);
and U9579 (N_9579,N_9325,N_9048);
nand U9580 (N_9580,N_9161,N_9430);
and U9581 (N_9581,N_9182,N_9131);
and U9582 (N_9582,N_9014,N_9356);
nor U9583 (N_9583,N_9297,N_9212);
or U9584 (N_9584,N_9264,N_9113);
or U9585 (N_9585,N_9309,N_9099);
nand U9586 (N_9586,N_9321,N_9123);
nand U9587 (N_9587,N_9347,N_9030);
nand U9588 (N_9588,N_9331,N_9035);
xor U9589 (N_9589,N_9143,N_9456);
nand U9590 (N_9590,N_9185,N_9022);
and U9591 (N_9591,N_9398,N_9340);
and U9592 (N_9592,N_9444,N_9085);
or U9593 (N_9593,N_9100,N_9446);
nand U9594 (N_9594,N_9137,N_9168);
nor U9595 (N_9595,N_9296,N_9288);
nand U9596 (N_9596,N_9074,N_9177);
nor U9597 (N_9597,N_9424,N_9018);
and U9598 (N_9598,N_9411,N_9105);
and U9599 (N_9599,N_9405,N_9337);
or U9600 (N_9600,N_9235,N_9156);
xnor U9601 (N_9601,N_9290,N_9475);
nand U9602 (N_9602,N_9465,N_9203);
nor U9603 (N_9603,N_9429,N_9358);
nand U9604 (N_9604,N_9381,N_9471);
or U9605 (N_9605,N_9476,N_9342);
nand U9606 (N_9606,N_9064,N_9090);
nor U9607 (N_9607,N_9106,N_9073);
nor U9608 (N_9608,N_9359,N_9261);
and U9609 (N_9609,N_9120,N_9148);
and U9610 (N_9610,N_9440,N_9042);
and U9611 (N_9611,N_9121,N_9472);
nand U9612 (N_9612,N_9110,N_9364);
and U9613 (N_9613,N_9425,N_9034);
nand U9614 (N_9614,N_9206,N_9083);
nor U9615 (N_9615,N_9135,N_9349);
or U9616 (N_9616,N_9481,N_9291);
nor U9617 (N_9617,N_9433,N_9208);
or U9618 (N_9618,N_9280,N_9150);
and U9619 (N_9619,N_9068,N_9478);
nor U9620 (N_9620,N_9276,N_9450);
nand U9621 (N_9621,N_9489,N_9196);
and U9622 (N_9622,N_9183,N_9144);
nand U9623 (N_9623,N_9253,N_9306);
nand U9624 (N_9624,N_9491,N_9286);
nand U9625 (N_9625,N_9245,N_9438);
nand U9626 (N_9626,N_9285,N_9289);
xnor U9627 (N_9627,N_9339,N_9348);
nand U9628 (N_9628,N_9086,N_9455);
and U9629 (N_9629,N_9496,N_9492);
and U9630 (N_9630,N_9378,N_9301);
and U9631 (N_9631,N_9365,N_9375);
xor U9632 (N_9632,N_9469,N_9393);
nor U9633 (N_9633,N_9256,N_9112);
nor U9634 (N_9634,N_9338,N_9154);
and U9635 (N_9635,N_9169,N_9373);
xnor U9636 (N_9636,N_9371,N_9151);
or U9637 (N_9637,N_9486,N_9343);
nand U9638 (N_9638,N_9372,N_9246);
nor U9639 (N_9639,N_9382,N_9153);
and U9640 (N_9640,N_9071,N_9400);
xnor U9641 (N_9641,N_9374,N_9361);
xor U9642 (N_9642,N_9096,N_9493);
and U9643 (N_9643,N_9062,N_9281);
xor U9644 (N_9644,N_9017,N_9010);
xnor U9645 (N_9645,N_9149,N_9222);
nor U9646 (N_9646,N_9434,N_9453);
or U9647 (N_9647,N_9376,N_9172);
and U9648 (N_9648,N_9497,N_9117);
nand U9649 (N_9649,N_9498,N_9432);
and U9650 (N_9650,N_9197,N_9081);
nor U9651 (N_9651,N_9084,N_9463);
nor U9652 (N_9652,N_9026,N_9420);
nand U9653 (N_9653,N_9000,N_9270);
xor U9654 (N_9654,N_9314,N_9370);
and U9655 (N_9655,N_9426,N_9303);
nor U9656 (N_9656,N_9460,N_9060);
nor U9657 (N_9657,N_9470,N_9158);
xor U9658 (N_9658,N_9095,N_9467);
nor U9659 (N_9659,N_9173,N_9189);
xor U9660 (N_9660,N_9052,N_9070);
xor U9661 (N_9661,N_9059,N_9380);
nor U9662 (N_9662,N_9317,N_9367);
xnor U9663 (N_9663,N_9396,N_9435);
xnor U9664 (N_9664,N_9413,N_9190);
or U9665 (N_9665,N_9181,N_9243);
xnor U9666 (N_9666,N_9442,N_9366);
nand U9667 (N_9667,N_9221,N_9369);
xnor U9668 (N_9668,N_9205,N_9082);
and U9669 (N_9669,N_9050,N_9308);
nor U9670 (N_9670,N_9094,N_9051);
nand U9671 (N_9671,N_9028,N_9262);
nand U9672 (N_9672,N_9198,N_9236);
xnor U9673 (N_9673,N_9260,N_9477);
or U9674 (N_9674,N_9319,N_9389);
xnor U9675 (N_9675,N_9452,N_9346);
xnor U9676 (N_9676,N_9407,N_9167);
and U9677 (N_9677,N_9330,N_9066);
nor U9678 (N_9678,N_9385,N_9155);
nand U9679 (N_9679,N_9054,N_9226);
nor U9680 (N_9680,N_9238,N_9227);
xor U9681 (N_9681,N_9461,N_9046);
nand U9682 (N_9682,N_9005,N_9334);
or U9683 (N_9683,N_9192,N_9152);
and U9684 (N_9684,N_9482,N_9287);
and U9685 (N_9685,N_9357,N_9147);
xnor U9686 (N_9686,N_9204,N_9333);
and U9687 (N_9687,N_9013,N_9271);
xor U9688 (N_9688,N_9327,N_9024);
xor U9689 (N_9689,N_9320,N_9436);
and U9690 (N_9690,N_9421,N_9335);
xnor U9691 (N_9691,N_9164,N_9310);
or U9692 (N_9692,N_9223,N_9266);
nand U9693 (N_9693,N_9045,N_9278);
nand U9694 (N_9694,N_9495,N_9055);
nand U9695 (N_9695,N_9250,N_9193);
or U9696 (N_9696,N_9166,N_9402);
nor U9697 (N_9697,N_9437,N_9294);
nand U9698 (N_9698,N_9265,N_9078);
and U9699 (N_9699,N_9394,N_9114);
nand U9700 (N_9700,N_9462,N_9295);
or U9701 (N_9701,N_9328,N_9061);
xor U9702 (N_9702,N_9207,N_9038);
nor U9703 (N_9703,N_9040,N_9362);
nand U9704 (N_9704,N_9016,N_9184);
nor U9705 (N_9705,N_9186,N_9176);
xor U9706 (N_9706,N_9023,N_9043);
nand U9707 (N_9707,N_9254,N_9091);
nand U9708 (N_9708,N_9466,N_9089);
or U9709 (N_9709,N_9323,N_9322);
and U9710 (N_9710,N_9269,N_9292);
nand U9711 (N_9711,N_9047,N_9403);
and U9712 (N_9712,N_9225,N_9474);
nor U9713 (N_9713,N_9231,N_9109);
nand U9714 (N_9714,N_9423,N_9077);
nand U9715 (N_9715,N_9111,N_9134);
or U9716 (N_9716,N_9006,N_9200);
and U9717 (N_9717,N_9020,N_9011);
and U9718 (N_9718,N_9300,N_9408);
or U9719 (N_9719,N_9025,N_9458);
xor U9720 (N_9720,N_9036,N_9473);
and U9721 (N_9721,N_9419,N_9132);
xor U9722 (N_9722,N_9194,N_9220);
or U9723 (N_9723,N_9088,N_9397);
and U9724 (N_9724,N_9041,N_9049);
xnor U9725 (N_9725,N_9237,N_9484);
nand U9726 (N_9726,N_9159,N_9241);
and U9727 (N_9727,N_9098,N_9248);
nand U9728 (N_9728,N_9214,N_9377);
nand U9729 (N_9729,N_9479,N_9399);
xor U9730 (N_9730,N_9257,N_9391);
xnor U9731 (N_9731,N_9387,N_9188);
nor U9732 (N_9732,N_9318,N_9217);
and U9733 (N_9733,N_9063,N_9240);
xnor U9734 (N_9734,N_9029,N_9341);
nor U9735 (N_9735,N_9130,N_9160);
or U9736 (N_9736,N_9459,N_9122);
and U9737 (N_9737,N_9345,N_9499);
xnor U9738 (N_9738,N_9268,N_9307);
nor U9739 (N_9739,N_9104,N_9284);
and U9740 (N_9740,N_9386,N_9293);
xnor U9741 (N_9741,N_9136,N_9431);
and U9742 (N_9742,N_9355,N_9344);
nor U9743 (N_9743,N_9146,N_9273);
nor U9744 (N_9744,N_9124,N_9412);
and U9745 (N_9745,N_9410,N_9103);
xnor U9746 (N_9746,N_9428,N_9485);
xnor U9747 (N_9747,N_9157,N_9145);
or U9748 (N_9748,N_9384,N_9012);
nand U9749 (N_9749,N_9141,N_9118);
and U9750 (N_9750,N_9499,N_9215);
nor U9751 (N_9751,N_9453,N_9194);
nor U9752 (N_9752,N_9070,N_9077);
or U9753 (N_9753,N_9284,N_9264);
nand U9754 (N_9754,N_9414,N_9043);
xor U9755 (N_9755,N_9212,N_9181);
nand U9756 (N_9756,N_9036,N_9463);
or U9757 (N_9757,N_9087,N_9487);
xnor U9758 (N_9758,N_9197,N_9432);
and U9759 (N_9759,N_9235,N_9299);
nor U9760 (N_9760,N_9316,N_9174);
nand U9761 (N_9761,N_9036,N_9486);
nor U9762 (N_9762,N_9469,N_9332);
xnor U9763 (N_9763,N_9377,N_9437);
or U9764 (N_9764,N_9054,N_9352);
nand U9765 (N_9765,N_9435,N_9120);
xnor U9766 (N_9766,N_9236,N_9177);
nand U9767 (N_9767,N_9289,N_9468);
nand U9768 (N_9768,N_9143,N_9253);
nor U9769 (N_9769,N_9270,N_9038);
nor U9770 (N_9770,N_9474,N_9330);
xnor U9771 (N_9771,N_9266,N_9475);
xnor U9772 (N_9772,N_9227,N_9383);
xnor U9773 (N_9773,N_9445,N_9287);
or U9774 (N_9774,N_9069,N_9492);
and U9775 (N_9775,N_9123,N_9337);
nand U9776 (N_9776,N_9330,N_9254);
xnor U9777 (N_9777,N_9492,N_9088);
or U9778 (N_9778,N_9017,N_9306);
nor U9779 (N_9779,N_9036,N_9050);
xor U9780 (N_9780,N_9135,N_9488);
and U9781 (N_9781,N_9310,N_9183);
xnor U9782 (N_9782,N_9102,N_9420);
nand U9783 (N_9783,N_9136,N_9377);
nand U9784 (N_9784,N_9055,N_9076);
nor U9785 (N_9785,N_9095,N_9082);
nor U9786 (N_9786,N_9442,N_9113);
nor U9787 (N_9787,N_9269,N_9058);
and U9788 (N_9788,N_9023,N_9237);
nor U9789 (N_9789,N_9397,N_9314);
xor U9790 (N_9790,N_9055,N_9437);
and U9791 (N_9791,N_9138,N_9052);
or U9792 (N_9792,N_9222,N_9123);
nand U9793 (N_9793,N_9365,N_9172);
nand U9794 (N_9794,N_9065,N_9001);
or U9795 (N_9795,N_9006,N_9013);
xor U9796 (N_9796,N_9414,N_9098);
and U9797 (N_9797,N_9082,N_9404);
nor U9798 (N_9798,N_9352,N_9314);
nor U9799 (N_9799,N_9456,N_9175);
nand U9800 (N_9800,N_9199,N_9020);
nor U9801 (N_9801,N_9279,N_9057);
and U9802 (N_9802,N_9325,N_9436);
nor U9803 (N_9803,N_9176,N_9062);
and U9804 (N_9804,N_9023,N_9180);
or U9805 (N_9805,N_9370,N_9497);
and U9806 (N_9806,N_9344,N_9218);
and U9807 (N_9807,N_9448,N_9158);
or U9808 (N_9808,N_9260,N_9045);
xor U9809 (N_9809,N_9460,N_9342);
nand U9810 (N_9810,N_9304,N_9428);
or U9811 (N_9811,N_9151,N_9269);
nor U9812 (N_9812,N_9392,N_9194);
nor U9813 (N_9813,N_9364,N_9438);
and U9814 (N_9814,N_9272,N_9126);
xor U9815 (N_9815,N_9150,N_9438);
nor U9816 (N_9816,N_9111,N_9428);
xnor U9817 (N_9817,N_9426,N_9494);
nor U9818 (N_9818,N_9093,N_9020);
nor U9819 (N_9819,N_9042,N_9496);
nor U9820 (N_9820,N_9443,N_9439);
nor U9821 (N_9821,N_9427,N_9370);
nor U9822 (N_9822,N_9214,N_9085);
or U9823 (N_9823,N_9460,N_9081);
nor U9824 (N_9824,N_9384,N_9079);
xor U9825 (N_9825,N_9101,N_9253);
or U9826 (N_9826,N_9180,N_9042);
or U9827 (N_9827,N_9370,N_9307);
or U9828 (N_9828,N_9061,N_9327);
xor U9829 (N_9829,N_9325,N_9084);
or U9830 (N_9830,N_9496,N_9406);
nor U9831 (N_9831,N_9222,N_9157);
nor U9832 (N_9832,N_9098,N_9200);
xnor U9833 (N_9833,N_9384,N_9316);
or U9834 (N_9834,N_9111,N_9439);
nand U9835 (N_9835,N_9176,N_9001);
or U9836 (N_9836,N_9256,N_9484);
xor U9837 (N_9837,N_9128,N_9004);
nor U9838 (N_9838,N_9299,N_9019);
xor U9839 (N_9839,N_9426,N_9432);
nor U9840 (N_9840,N_9238,N_9178);
nor U9841 (N_9841,N_9454,N_9005);
xor U9842 (N_9842,N_9026,N_9304);
xnor U9843 (N_9843,N_9086,N_9493);
and U9844 (N_9844,N_9221,N_9000);
or U9845 (N_9845,N_9373,N_9142);
or U9846 (N_9846,N_9052,N_9072);
or U9847 (N_9847,N_9093,N_9479);
nand U9848 (N_9848,N_9384,N_9399);
nor U9849 (N_9849,N_9306,N_9093);
and U9850 (N_9850,N_9055,N_9113);
nand U9851 (N_9851,N_9108,N_9395);
or U9852 (N_9852,N_9382,N_9210);
xnor U9853 (N_9853,N_9226,N_9089);
nand U9854 (N_9854,N_9069,N_9460);
xnor U9855 (N_9855,N_9303,N_9386);
and U9856 (N_9856,N_9446,N_9470);
xnor U9857 (N_9857,N_9324,N_9166);
or U9858 (N_9858,N_9113,N_9298);
or U9859 (N_9859,N_9428,N_9259);
or U9860 (N_9860,N_9443,N_9159);
and U9861 (N_9861,N_9139,N_9047);
and U9862 (N_9862,N_9212,N_9337);
or U9863 (N_9863,N_9117,N_9080);
nor U9864 (N_9864,N_9004,N_9193);
and U9865 (N_9865,N_9086,N_9332);
nor U9866 (N_9866,N_9133,N_9324);
or U9867 (N_9867,N_9376,N_9409);
nor U9868 (N_9868,N_9012,N_9186);
or U9869 (N_9869,N_9244,N_9418);
or U9870 (N_9870,N_9419,N_9381);
nand U9871 (N_9871,N_9106,N_9352);
and U9872 (N_9872,N_9244,N_9142);
or U9873 (N_9873,N_9104,N_9444);
xor U9874 (N_9874,N_9456,N_9203);
nand U9875 (N_9875,N_9367,N_9074);
or U9876 (N_9876,N_9408,N_9113);
or U9877 (N_9877,N_9338,N_9174);
xor U9878 (N_9878,N_9489,N_9261);
nor U9879 (N_9879,N_9131,N_9072);
xor U9880 (N_9880,N_9464,N_9476);
xor U9881 (N_9881,N_9309,N_9181);
nand U9882 (N_9882,N_9082,N_9375);
nor U9883 (N_9883,N_9361,N_9219);
and U9884 (N_9884,N_9431,N_9327);
and U9885 (N_9885,N_9231,N_9473);
xor U9886 (N_9886,N_9215,N_9060);
or U9887 (N_9887,N_9282,N_9411);
and U9888 (N_9888,N_9078,N_9230);
and U9889 (N_9889,N_9280,N_9113);
xnor U9890 (N_9890,N_9317,N_9231);
xnor U9891 (N_9891,N_9077,N_9029);
or U9892 (N_9892,N_9345,N_9257);
nor U9893 (N_9893,N_9439,N_9358);
and U9894 (N_9894,N_9082,N_9299);
nand U9895 (N_9895,N_9494,N_9422);
or U9896 (N_9896,N_9302,N_9306);
or U9897 (N_9897,N_9434,N_9439);
nand U9898 (N_9898,N_9116,N_9095);
or U9899 (N_9899,N_9089,N_9361);
nand U9900 (N_9900,N_9417,N_9153);
nor U9901 (N_9901,N_9063,N_9332);
and U9902 (N_9902,N_9198,N_9340);
nor U9903 (N_9903,N_9166,N_9359);
nor U9904 (N_9904,N_9100,N_9076);
nand U9905 (N_9905,N_9268,N_9220);
nor U9906 (N_9906,N_9189,N_9005);
nor U9907 (N_9907,N_9229,N_9149);
nor U9908 (N_9908,N_9163,N_9271);
or U9909 (N_9909,N_9135,N_9023);
nand U9910 (N_9910,N_9114,N_9343);
or U9911 (N_9911,N_9124,N_9377);
nand U9912 (N_9912,N_9124,N_9048);
or U9913 (N_9913,N_9239,N_9308);
nand U9914 (N_9914,N_9230,N_9348);
and U9915 (N_9915,N_9447,N_9327);
nor U9916 (N_9916,N_9269,N_9305);
xor U9917 (N_9917,N_9330,N_9160);
xnor U9918 (N_9918,N_9486,N_9018);
or U9919 (N_9919,N_9232,N_9347);
nor U9920 (N_9920,N_9424,N_9264);
and U9921 (N_9921,N_9494,N_9104);
nand U9922 (N_9922,N_9100,N_9485);
xnor U9923 (N_9923,N_9219,N_9294);
or U9924 (N_9924,N_9169,N_9337);
and U9925 (N_9925,N_9351,N_9496);
nor U9926 (N_9926,N_9306,N_9471);
xor U9927 (N_9927,N_9065,N_9162);
or U9928 (N_9928,N_9398,N_9120);
nor U9929 (N_9929,N_9338,N_9171);
nor U9930 (N_9930,N_9069,N_9061);
and U9931 (N_9931,N_9443,N_9459);
nand U9932 (N_9932,N_9256,N_9197);
nand U9933 (N_9933,N_9237,N_9160);
nor U9934 (N_9934,N_9052,N_9046);
or U9935 (N_9935,N_9256,N_9267);
xor U9936 (N_9936,N_9202,N_9012);
or U9937 (N_9937,N_9428,N_9366);
xnor U9938 (N_9938,N_9398,N_9416);
nor U9939 (N_9939,N_9167,N_9362);
nand U9940 (N_9940,N_9030,N_9396);
xor U9941 (N_9941,N_9420,N_9147);
or U9942 (N_9942,N_9209,N_9324);
xor U9943 (N_9943,N_9255,N_9146);
xor U9944 (N_9944,N_9322,N_9195);
nand U9945 (N_9945,N_9334,N_9045);
or U9946 (N_9946,N_9029,N_9198);
nand U9947 (N_9947,N_9400,N_9275);
nand U9948 (N_9948,N_9186,N_9054);
nand U9949 (N_9949,N_9290,N_9393);
or U9950 (N_9950,N_9235,N_9124);
nand U9951 (N_9951,N_9201,N_9240);
xor U9952 (N_9952,N_9314,N_9244);
nor U9953 (N_9953,N_9198,N_9246);
nor U9954 (N_9954,N_9150,N_9453);
xnor U9955 (N_9955,N_9346,N_9394);
nor U9956 (N_9956,N_9384,N_9430);
nor U9957 (N_9957,N_9141,N_9180);
nor U9958 (N_9958,N_9159,N_9376);
xor U9959 (N_9959,N_9124,N_9360);
nand U9960 (N_9960,N_9124,N_9271);
xnor U9961 (N_9961,N_9443,N_9264);
and U9962 (N_9962,N_9134,N_9191);
nor U9963 (N_9963,N_9189,N_9444);
nor U9964 (N_9964,N_9315,N_9477);
nor U9965 (N_9965,N_9316,N_9351);
or U9966 (N_9966,N_9076,N_9220);
and U9967 (N_9967,N_9132,N_9198);
and U9968 (N_9968,N_9463,N_9489);
and U9969 (N_9969,N_9352,N_9071);
or U9970 (N_9970,N_9174,N_9175);
nand U9971 (N_9971,N_9020,N_9284);
nand U9972 (N_9972,N_9372,N_9089);
nor U9973 (N_9973,N_9332,N_9175);
nor U9974 (N_9974,N_9450,N_9391);
nand U9975 (N_9975,N_9244,N_9101);
or U9976 (N_9976,N_9328,N_9010);
nand U9977 (N_9977,N_9263,N_9470);
nand U9978 (N_9978,N_9393,N_9351);
or U9979 (N_9979,N_9390,N_9215);
or U9980 (N_9980,N_9343,N_9215);
or U9981 (N_9981,N_9269,N_9165);
xnor U9982 (N_9982,N_9343,N_9321);
xnor U9983 (N_9983,N_9474,N_9422);
xor U9984 (N_9984,N_9163,N_9160);
nor U9985 (N_9985,N_9147,N_9119);
or U9986 (N_9986,N_9027,N_9068);
nor U9987 (N_9987,N_9027,N_9122);
nor U9988 (N_9988,N_9301,N_9450);
nor U9989 (N_9989,N_9422,N_9256);
xnor U9990 (N_9990,N_9416,N_9450);
nand U9991 (N_9991,N_9201,N_9166);
and U9992 (N_9992,N_9057,N_9184);
nor U9993 (N_9993,N_9257,N_9095);
or U9994 (N_9994,N_9119,N_9117);
or U9995 (N_9995,N_9235,N_9021);
nand U9996 (N_9996,N_9284,N_9488);
and U9997 (N_9997,N_9164,N_9237);
and U9998 (N_9998,N_9000,N_9212);
or U9999 (N_9999,N_9223,N_9478);
and U10000 (N_10000,N_9506,N_9517);
nor U10001 (N_10001,N_9588,N_9872);
xor U10002 (N_10002,N_9554,N_9541);
nand U10003 (N_10003,N_9654,N_9746);
nand U10004 (N_10004,N_9794,N_9714);
nand U10005 (N_10005,N_9800,N_9835);
nand U10006 (N_10006,N_9724,N_9860);
or U10007 (N_10007,N_9734,N_9676);
xnor U10008 (N_10008,N_9905,N_9834);
and U10009 (N_10009,N_9888,N_9942);
or U10010 (N_10010,N_9780,N_9957);
xor U10011 (N_10011,N_9883,N_9509);
xor U10012 (N_10012,N_9770,N_9947);
and U10013 (N_10013,N_9903,N_9900);
xor U10014 (N_10014,N_9821,N_9784);
or U10015 (N_10015,N_9817,N_9820);
and U10016 (N_10016,N_9890,N_9980);
nand U10017 (N_10017,N_9582,N_9832);
and U10018 (N_10018,N_9624,N_9635);
nor U10019 (N_10019,N_9776,N_9544);
xnor U10020 (N_10020,N_9553,N_9906);
xnor U10021 (N_10021,N_9859,N_9687);
or U10022 (N_10022,N_9975,N_9722);
xnor U10023 (N_10023,N_9916,N_9801);
xnor U10024 (N_10024,N_9809,N_9973);
nand U10025 (N_10025,N_9774,N_9732);
nor U10026 (N_10026,N_9962,N_9640);
or U10027 (N_10027,N_9502,N_9937);
and U10028 (N_10028,N_9529,N_9637);
xor U10029 (N_10029,N_9857,N_9824);
or U10030 (N_10030,N_9984,N_9717);
nand U10031 (N_10031,N_9601,N_9775);
nand U10032 (N_10032,N_9713,N_9871);
nor U10033 (N_10033,N_9852,N_9546);
or U10034 (N_10034,N_9828,N_9799);
nor U10035 (N_10035,N_9989,N_9694);
or U10036 (N_10036,N_9970,N_9995);
nor U10037 (N_10037,N_9666,N_9864);
nand U10038 (N_10038,N_9585,N_9966);
nor U10039 (N_10039,N_9881,N_9510);
or U10040 (N_10040,N_9846,N_9758);
xnor U10041 (N_10041,N_9662,N_9699);
nor U10042 (N_10042,N_9551,N_9878);
xor U10043 (N_10043,N_9511,N_9867);
nor U10044 (N_10044,N_9697,N_9983);
xor U10045 (N_10045,N_9682,N_9545);
nor U10046 (N_10046,N_9623,N_9849);
or U10047 (N_10047,N_9706,N_9939);
xnor U10048 (N_10048,N_9547,N_9610);
and U10049 (N_10049,N_9708,N_9723);
or U10050 (N_10050,N_9972,N_9994);
and U10051 (N_10051,N_9715,N_9744);
xor U10052 (N_10052,N_9752,N_9653);
nor U10053 (N_10053,N_9842,N_9954);
nor U10054 (N_10054,N_9534,N_9894);
nand U10055 (N_10055,N_9643,N_9761);
nor U10056 (N_10056,N_9673,N_9971);
and U10057 (N_10057,N_9961,N_9967);
or U10058 (N_10058,N_9677,N_9868);
nor U10059 (N_10059,N_9663,N_9721);
nor U10060 (N_10060,N_9802,N_9571);
xor U10061 (N_10061,N_9630,N_9874);
nor U10062 (N_10062,N_9922,N_9825);
nand U10063 (N_10063,N_9908,N_9921);
or U10064 (N_10064,N_9865,N_9923);
nor U10065 (N_10065,N_9965,N_9591);
nand U10066 (N_10066,N_9512,N_9577);
nand U10067 (N_10067,N_9990,N_9958);
xor U10068 (N_10068,N_9827,N_9614);
nand U10069 (N_10069,N_9831,N_9870);
nand U10070 (N_10070,N_9685,N_9669);
and U10071 (N_10071,N_9552,N_9538);
nor U10072 (N_10072,N_9597,N_9934);
nand U10073 (N_10073,N_9963,N_9838);
xnor U10074 (N_10074,N_9543,N_9559);
or U10075 (N_10075,N_9913,N_9897);
or U10076 (N_10076,N_9701,N_9932);
nand U10077 (N_10077,N_9636,N_9690);
nor U10078 (N_10078,N_9675,N_9818);
nor U10079 (N_10079,N_9814,N_9747);
nand U10080 (N_10080,N_9592,N_9866);
nand U10081 (N_10081,N_9986,N_9647);
or U10082 (N_10082,N_9626,N_9729);
nor U10083 (N_10083,N_9889,N_9741);
or U10084 (N_10084,N_9648,N_9556);
and U10085 (N_10085,N_9508,N_9596);
and U10086 (N_10086,N_9974,N_9524);
or U10087 (N_10087,N_9615,N_9887);
and U10088 (N_10088,N_9912,N_9940);
nor U10089 (N_10089,N_9791,N_9884);
and U10090 (N_10090,N_9960,N_9514);
and U10091 (N_10091,N_9798,N_9847);
nand U10092 (N_10092,N_9700,N_9593);
nand U10093 (N_10093,N_9790,N_9924);
and U10094 (N_10094,N_9855,N_9943);
or U10095 (N_10095,N_9539,N_9679);
xnor U10096 (N_10096,N_9667,N_9787);
xor U10097 (N_10097,N_9627,N_9815);
and U10098 (N_10098,N_9763,N_9902);
nand U10099 (N_10099,N_9745,N_9590);
xor U10100 (N_10100,N_9914,N_9767);
nor U10101 (N_10101,N_9642,N_9816);
nor U10102 (N_10102,N_9657,N_9688);
nand U10103 (N_10103,N_9656,N_9788);
and U10104 (N_10104,N_9580,N_9594);
or U10105 (N_10105,N_9629,N_9562);
xnor U10106 (N_10106,N_9581,N_9993);
nor U10107 (N_10107,N_9606,N_9985);
or U10108 (N_10108,N_9751,N_9773);
nor U10109 (N_10109,N_9613,N_9503);
and U10110 (N_10110,N_9698,N_9768);
nand U10111 (N_10111,N_9600,N_9987);
or U10112 (N_10112,N_9756,N_9716);
nand U10113 (N_10113,N_9952,N_9991);
xnor U10114 (N_10114,N_9956,N_9726);
or U10115 (N_10115,N_9599,N_9813);
and U10116 (N_10116,N_9665,N_9583);
xor U10117 (N_10117,N_9584,N_9725);
and U10118 (N_10118,N_9576,N_9574);
xnor U10119 (N_10119,N_9605,N_9655);
or U10120 (N_10120,N_9733,N_9786);
xor U10121 (N_10121,N_9612,N_9705);
nand U10122 (N_10122,N_9856,N_9759);
and U10123 (N_10123,N_9836,N_9822);
xor U10124 (N_10124,N_9650,N_9862);
or U10125 (N_10125,N_9941,N_9720);
or U10126 (N_10126,N_9777,N_9548);
nor U10127 (N_10127,N_9896,N_9804);
and U10128 (N_10128,N_9739,N_9981);
and U10129 (N_10129,N_9919,N_9826);
and U10130 (N_10130,N_9707,N_9792);
nor U10131 (N_10131,N_9819,N_9712);
nor U10132 (N_10132,N_9785,N_9660);
or U10133 (N_10133,N_9945,N_9621);
or U10134 (N_10134,N_9565,N_9737);
or U10135 (N_10135,N_9535,N_9608);
and U10136 (N_10136,N_9587,N_9840);
and U10137 (N_10137,N_9651,N_9589);
xor U10138 (N_10138,N_9964,N_9797);
xnor U10139 (N_10139,N_9812,N_9928);
nor U10140 (N_10140,N_9772,N_9978);
xnor U10141 (N_10141,N_9572,N_9749);
or U10142 (N_10142,N_9644,N_9740);
nand U10143 (N_10143,N_9550,N_9769);
or U10144 (N_10144,N_9979,N_9728);
and U10145 (N_10145,N_9936,N_9880);
nor U10146 (N_10146,N_9771,N_9638);
xor U10147 (N_10147,N_9528,N_9803);
nand U10148 (N_10148,N_9992,N_9680);
and U10149 (N_10149,N_9575,N_9861);
and U10150 (N_10150,N_9968,N_9639);
xnor U10151 (N_10151,N_9918,N_9689);
xor U10152 (N_10152,N_9750,N_9661);
nor U10153 (N_10153,N_9757,N_9730);
nand U10154 (N_10154,N_9891,N_9873);
and U10155 (N_10155,N_9904,N_9693);
xnor U10156 (N_10156,N_9837,N_9781);
or U10157 (N_10157,N_9931,N_9920);
xor U10158 (N_10158,N_9999,N_9805);
xor U10159 (N_10159,N_9731,N_9927);
nor U10160 (N_10160,N_9568,N_9531);
and U10161 (N_10161,N_9504,N_9537);
nand U10162 (N_10162,N_9844,N_9877);
xnor U10163 (N_10163,N_9930,N_9808);
or U10164 (N_10164,N_9631,N_9901);
and U10165 (N_10165,N_9507,N_9807);
nor U10166 (N_10166,N_9632,N_9998);
nor U10167 (N_10167,N_9823,N_9540);
nor U10168 (N_10168,N_9634,N_9762);
xnor U10169 (N_10169,N_9564,N_9926);
nand U10170 (N_10170,N_9738,N_9782);
xor U10171 (N_10171,N_9793,N_9619);
or U10172 (N_10172,N_9858,N_9727);
nor U10173 (N_10173,N_9779,N_9670);
or U10174 (N_10174,N_9607,N_9778);
and U10175 (N_10175,N_9611,N_9748);
xor U10176 (N_10176,N_9863,N_9501);
and U10177 (N_10177,N_9953,N_9684);
xor U10178 (N_10178,N_9710,N_9915);
nand U10179 (N_10179,N_9625,N_9946);
and U10180 (N_10180,N_9951,N_9555);
nand U10181 (N_10181,N_9711,N_9703);
and U10182 (N_10182,N_9959,N_9850);
xor U10183 (N_10183,N_9950,N_9753);
xnor U10184 (N_10184,N_9518,N_9505);
or U10185 (N_10185,N_9843,N_9641);
and U10186 (N_10186,N_9696,N_9526);
xnor U10187 (N_10187,N_9851,N_9602);
and U10188 (N_10188,N_9718,N_9875);
nor U10189 (N_10189,N_9911,N_9649);
and U10190 (N_10190,N_9841,N_9530);
or U10191 (N_10191,N_9743,N_9977);
xor U10192 (N_10192,N_9542,N_9882);
or U10193 (N_10193,N_9810,N_9899);
or U10194 (N_10194,N_9892,N_9532);
nand U10195 (N_10195,N_9567,N_9754);
and U10196 (N_10196,N_9944,N_9628);
nand U10197 (N_10197,N_9566,N_9969);
xnor U10198 (N_10198,N_9755,N_9789);
nor U10199 (N_10199,N_9885,N_9811);
and U10200 (N_10200,N_9617,N_9549);
and U10201 (N_10201,N_9795,N_9520);
nor U10202 (N_10202,N_9742,N_9833);
or U10203 (N_10203,N_9695,N_9598);
or U10204 (N_10204,N_9949,N_9622);
or U10205 (N_10205,N_9516,N_9735);
or U10206 (N_10206,N_9521,N_9691);
xnor U10207 (N_10207,N_9879,N_9845);
or U10208 (N_10208,N_9560,N_9603);
or U10209 (N_10209,N_9925,N_9573);
nand U10210 (N_10210,N_9681,N_9830);
or U10211 (N_10211,N_9561,N_9869);
or U10212 (N_10212,N_9853,N_9683);
xnor U10213 (N_10213,N_9909,N_9525);
nand U10214 (N_10214,N_9570,N_9563);
nor U10215 (N_10215,N_9736,N_9806);
or U10216 (N_10216,N_9578,N_9618);
and U10217 (N_10217,N_9783,N_9659);
or U10218 (N_10218,N_9558,N_9616);
and U10219 (N_10219,N_9766,N_9586);
or U10220 (N_10220,N_9886,N_9895);
xnor U10221 (N_10221,N_9664,N_9917);
or U10222 (N_10222,N_9876,N_9686);
or U10223 (N_10223,N_9609,N_9848);
nor U10224 (N_10224,N_9839,N_9523);
nor U10225 (N_10225,N_9658,N_9604);
xor U10226 (N_10226,N_9702,N_9645);
or U10227 (N_10227,N_9672,N_9527);
xor U10228 (N_10228,N_9907,N_9829);
nand U10229 (N_10229,N_9620,N_9652);
nor U10230 (N_10230,N_9893,N_9595);
and U10231 (N_10231,N_9709,N_9938);
xor U10232 (N_10232,N_9955,N_9500);
nand U10233 (N_10233,N_9579,N_9522);
nand U10234 (N_10234,N_9704,N_9996);
and U10235 (N_10235,N_9674,N_9646);
xor U10236 (N_10236,N_9764,N_9513);
nand U10237 (N_10237,N_9519,N_9948);
or U10238 (N_10238,N_9536,N_9678);
xnor U10239 (N_10239,N_9765,N_9719);
nor U10240 (N_10240,N_9910,N_9557);
nor U10241 (N_10241,N_9935,N_9760);
xnor U10242 (N_10242,N_9898,N_9997);
nand U10243 (N_10243,N_9982,N_9854);
and U10244 (N_10244,N_9933,N_9692);
and U10245 (N_10245,N_9988,N_9533);
nand U10246 (N_10246,N_9515,N_9929);
nor U10247 (N_10247,N_9976,N_9569);
and U10248 (N_10248,N_9668,N_9671);
nand U10249 (N_10249,N_9633,N_9796);
nand U10250 (N_10250,N_9528,N_9968);
nor U10251 (N_10251,N_9980,N_9642);
xor U10252 (N_10252,N_9928,N_9951);
nand U10253 (N_10253,N_9783,N_9613);
xnor U10254 (N_10254,N_9973,N_9909);
and U10255 (N_10255,N_9705,N_9848);
and U10256 (N_10256,N_9545,N_9578);
nand U10257 (N_10257,N_9801,N_9787);
nand U10258 (N_10258,N_9796,N_9945);
and U10259 (N_10259,N_9615,N_9933);
nand U10260 (N_10260,N_9587,N_9984);
nand U10261 (N_10261,N_9589,N_9639);
and U10262 (N_10262,N_9717,N_9706);
and U10263 (N_10263,N_9533,N_9924);
or U10264 (N_10264,N_9978,N_9586);
nor U10265 (N_10265,N_9709,N_9760);
or U10266 (N_10266,N_9792,N_9769);
xnor U10267 (N_10267,N_9808,N_9879);
xor U10268 (N_10268,N_9891,N_9994);
xnor U10269 (N_10269,N_9660,N_9804);
xor U10270 (N_10270,N_9560,N_9944);
xor U10271 (N_10271,N_9659,N_9979);
nor U10272 (N_10272,N_9979,N_9636);
nor U10273 (N_10273,N_9870,N_9648);
nand U10274 (N_10274,N_9637,N_9754);
and U10275 (N_10275,N_9788,N_9854);
xnor U10276 (N_10276,N_9735,N_9697);
xor U10277 (N_10277,N_9716,N_9762);
nor U10278 (N_10278,N_9942,N_9646);
nor U10279 (N_10279,N_9768,N_9586);
or U10280 (N_10280,N_9721,N_9706);
nor U10281 (N_10281,N_9772,N_9929);
and U10282 (N_10282,N_9837,N_9591);
xor U10283 (N_10283,N_9716,N_9636);
xnor U10284 (N_10284,N_9917,N_9854);
and U10285 (N_10285,N_9713,N_9695);
or U10286 (N_10286,N_9900,N_9775);
nand U10287 (N_10287,N_9958,N_9986);
xnor U10288 (N_10288,N_9969,N_9517);
or U10289 (N_10289,N_9605,N_9904);
nand U10290 (N_10290,N_9606,N_9724);
xnor U10291 (N_10291,N_9773,N_9657);
nand U10292 (N_10292,N_9938,N_9725);
nor U10293 (N_10293,N_9882,N_9618);
xor U10294 (N_10294,N_9832,N_9960);
nand U10295 (N_10295,N_9521,N_9999);
nand U10296 (N_10296,N_9649,N_9548);
xnor U10297 (N_10297,N_9717,N_9863);
and U10298 (N_10298,N_9794,N_9704);
nand U10299 (N_10299,N_9867,N_9632);
xor U10300 (N_10300,N_9857,N_9658);
or U10301 (N_10301,N_9836,N_9883);
xor U10302 (N_10302,N_9785,N_9682);
nor U10303 (N_10303,N_9780,N_9528);
or U10304 (N_10304,N_9784,N_9985);
and U10305 (N_10305,N_9524,N_9549);
and U10306 (N_10306,N_9630,N_9584);
or U10307 (N_10307,N_9647,N_9595);
xnor U10308 (N_10308,N_9618,N_9681);
nor U10309 (N_10309,N_9800,N_9589);
and U10310 (N_10310,N_9965,N_9511);
or U10311 (N_10311,N_9519,N_9847);
or U10312 (N_10312,N_9533,N_9594);
nand U10313 (N_10313,N_9940,N_9934);
or U10314 (N_10314,N_9555,N_9775);
nand U10315 (N_10315,N_9750,N_9856);
nand U10316 (N_10316,N_9703,N_9835);
nor U10317 (N_10317,N_9650,N_9978);
nor U10318 (N_10318,N_9702,N_9680);
xor U10319 (N_10319,N_9932,N_9577);
xor U10320 (N_10320,N_9955,N_9682);
nand U10321 (N_10321,N_9595,N_9843);
xnor U10322 (N_10322,N_9716,N_9789);
nor U10323 (N_10323,N_9598,N_9755);
nand U10324 (N_10324,N_9544,N_9848);
xor U10325 (N_10325,N_9626,N_9718);
nor U10326 (N_10326,N_9693,N_9862);
nor U10327 (N_10327,N_9625,N_9728);
nor U10328 (N_10328,N_9734,N_9627);
or U10329 (N_10329,N_9945,N_9863);
nand U10330 (N_10330,N_9761,N_9845);
nor U10331 (N_10331,N_9525,N_9841);
xor U10332 (N_10332,N_9967,N_9600);
nor U10333 (N_10333,N_9893,N_9787);
or U10334 (N_10334,N_9826,N_9812);
and U10335 (N_10335,N_9925,N_9621);
or U10336 (N_10336,N_9503,N_9780);
or U10337 (N_10337,N_9706,N_9887);
nand U10338 (N_10338,N_9648,N_9753);
xor U10339 (N_10339,N_9955,N_9600);
nor U10340 (N_10340,N_9592,N_9720);
nand U10341 (N_10341,N_9978,N_9938);
xor U10342 (N_10342,N_9616,N_9929);
or U10343 (N_10343,N_9617,N_9773);
nor U10344 (N_10344,N_9729,N_9785);
xnor U10345 (N_10345,N_9937,N_9567);
xnor U10346 (N_10346,N_9704,N_9702);
nand U10347 (N_10347,N_9713,N_9610);
nor U10348 (N_10348,N_9634,N_9654);
nor U10349 (N_10349,N_9572,N_9590);
or U10350 (N_10350,N_9555,N_9584);
or U10351 (N_10351,N_9585,N_9735);
nand U10352 (N_10352,N_9718,N_9798);
nand U10353 (N_10353,N_9556,N_9680);
or U10354 (N_10354,N_9613,N_9843);
and U10355 (N_10355,N_9809,N_9943);
and U10356 (N_10356,N_9983,N_9660);
nand U10357 (N_10357,N_9848,N_9679);
or U10358 (N_10358,N_9844,N_9881);
nand U10359 (N_10359,N_9658,N_9983);
and U10360 (N_10360,N_9993,N_9851);
nor U10361 (N_10361,N_9868,N_9578);
or U10362 (N_10362,N_9520,N_9717);
nor U10363 (N_10363,N_9532,N_9792);
xnor U10364 (N_10364,N_9613,N_9625);
or U10365 (N_10365,N_9885,N_9691);
nor U10366 (N_10366,N_9646,N_9862);
xor U10367 (N_10367,N_9856,N_9506);
or U10368 (N_10368,N_9679,N_9913);
and U10369 (N_10369,N_9776,N_9656);
nor U10370 (N_10370,N_9539,N_9902);
xor U10371 (N_10371,N_9970,N_9941);
nand U10372 (N_10372,N_9599,N_9943);
or U10373 (N_10373,N_9739,N_9988);
or U10374 (N_10374,N_9656,N_9951);
and U10375 (N_10375,N_9626,N_9516);
nand U10376 (N_10376,N_9678,N_9586);
nand U10377 (N_10377,N_9988,N_9710);
nor U10378 (N_10378,N_9543,N_9985);
or U10379 (N_10379,N_9625,N_9599);
and U10380 (N_10380,N_9656,N_9635);
or U10381 (N_10381,N_9963,N_9886);
xnor U10382 (N_10382,N_9723,N_9682);
xor U10383 (N_10383,N_9625,N_9846);
and U10384 (N_10384,N_9891,N_9550);
and U10385 (N_10385,N_9971,N_9512);
or U10386 (N_10386,N_9963,N_9541);
nor U10387 (N_10387,N_9970,N_9809);
nor U10388 (N_10388,N_9805,N_9774);
and U10389 (N_10389,N_9814,N_9926);
xor U10390 (N_10390,N_9991,N_9733);
nor U10391 (N_10391,N_9724,N_9761);
and U10392 (N_10392,N_9639,N_9618);
xnor U10393 (N_10393,N_9579,N_9889);
and U10394 (N_10394,N_9792,N_9510);
nand U10395 (N_10395,N_9635,N_9969);
nor U10396 (N_10396,N_9535,N_9590);
nand U10397 (N_10397,N_9695,N_9679);
nor U10398 (N_10398,N_9608,N_9804);
xnor U10399 (N_10399,N_9805,N_9891);
xor U10400 (N_10400,N_9848,N_9663);
nand U10401 (N_10401,N_9676,N_9668);
nand U10402 (N_10402,N_9635,N_9678);
nand U10403 (N_10403,N_9892,N_9705);
and U10404 (N_10404,N_9903,N_9766);
nand U10405 (N_10405,N_9953,N_9628);
nor U10406 (N_10406,N_9953,N_9812);
nor U10407 (N_10407,N_9522,N_9716);
xnor U10408 (N_10408,N_9552,N_9568);
and U10409 (N_10409,N_9758,N_9624);
nand U10410 (N_10410,N_9910,N_9768);
or U10411 (N_10411,N_9698,N_9687);
nor U10412 (N_10412,N_9505,N_9749);
or U10413 (N_10413,N_9963,N_9528);
and U10414 (N_10414,N_9939,N_9771);
nand U10415 (N_10415,N_9614,N_9896);
or U10416 (N_10416,N_9600,N_9934);
nand U10417 (N_10417,N_9585,N_9640);
nor U10418 (N_10418,N_9800,N_9727);
or U10419 (N_10419,N_9577,N_9797);
nand U10420 (N_10420,N_9630,N_9738);
or U10421 (N_10421,N_9769,N_9650);
xor U10422 (N_10422,N_9894,N_9943);
nor U10423 (N_10423,N_9790,N_9596);
nor U10424 (N_10424,N_9716,N_9846);
nor U10425 (N_10425,N_9941,N_9706);
nand U10426 (N_10426,N_9602,N_9642);
nor U10427 (N_10427,N_9701,N_9973);
nand U10428 (N_10428,N_9807,N_9542);
nor U10429 (N_10429,N_9576,N_9681);
or U10430 (N_10430,N_9738,N_9648);
xor U10431 (N_10431,N_9543,N_9628);
xnor U10432 (N_10432,N_9802,N_9865);
or U10433 (N_10433,N_9954,N_9646);
and U10434 (N_10434,N_9743,N_9939);
xnor U10435 (N_10435,N_9968,N_9653);
nor U10436 (N_10436,N_9862,N_9873);
nor U10437 (N_10437,N_9711,N_9919);
nor U10438 (N_10438,N_9993,N_9916);
and U10439 (N_10439,N_9962,N_9992);
nor U10440 (N_10440,N_9696,N_9900);
nor U10441 (N_10441,N_9615,N_9703);
nor U10442 (N_10442,N_9910,N_9915);
xnor U10443 (N_10443,N_9614,N_9509);
xnor U10444 (N_10444,N_9614,N_9580);
and U10445 (N_10445,N_9605,N_9619);
or U10446 (N_10446,N_9983,N_9885);
nand U10447 (N_10447,N_9616,N_9969);
or U10448 (N_10448,N_9924,N_9910);
xor U10449 (N_10449,N_9593,N_9971);
and U10450 (N_10450,N_9792,N_9788);
or U10451 (N_10451,N_9721,N_9731);
and U10452 (N_10452,N_9987,N_9813);
and U10453 (N_10453,N_9514,N_9562);
nand U10454 (N_10454,N_9858,N_9908);
xor U10455 (N_10455,N_9855,N_9740);
nand U10456 (N_10456,N_9891,N_9688);
xor U10457 (N_10457,N_9751,N_9984);
nor U10458 (N_10458,N_9781,N_9611);
and U10459 (N_10459,N_9507,N_9919);
and U10460 (N_10460,N_9885,N_9680);
or U10461 (N_10461,N_9594,N_9529);
xnor U10462 (N_10462,N_9881,N_9999);
and U10463 (N_10463,N_9970,N_9729);
and U10464 (N_10464,N_9924,N_9654);
xnor U10465 (N_10465,N_9687,N_9722);
nor U10466 (N_10466,N_9531,N_9960);
and U10467 (N_10467,N_9642,N_9542);
or U10468 (N_10468,N_9626,N_9617);
and U10469 (N_10469,N_9556,N_9662);
xnor U10470 (N_10470,N_9956,N_9816);
xnor U10471 (N_10471,N_9797,N_9678);
and U10472 (N_10472,N_9968,N_9663);
nor U10473 (N_10473,N_9849,N_9505);
nor U10474 (N_10474,N_9771,N_9538);
nand U10475 (N_10475,N_9532,N_9534);
or U10476 (N_10476,N_9587,N_9635);
nor U10477 (N_10477,N_9937,N_9776);
and U10478 (N_10478,N_9551,N_9500);
nor U10479 (N_10479,N_9902,N_9610);
xor U10480 (N_10480,N_9882,N_9885);
xnor U10481 (N_10481,N_9669,N_9761);
nand U10482 (N_10482,N_9860,N_9787);
nand U10483 (N_10483,N_9934,N_9850);
nor U10484 (N_10484,N_9630,N_9696);
xor U10485 (N_10485,N_9579,N_9837);
xnor U10486 (N_10486,N_9508,N_9536);
and U10487 (N_10487,N_9683,N_9545);
nor U10488 (N_10488,N_9605,N_9722);
nor U10489 (N_10489,N_9875,N_9763);
nand U10490 (N_10490,N_9630,N_9779);
nand U10491 (N_10491,N_9661,N_9527);
xnor U10492 (N_10492,N_9800,N_9733);
xnor U10493 (N_10493,N_9563,N_9847);
and U10494 (N_10494,N_9912,N_9780);
xor U10495 (N_10495,N_9541,N_9681);
nand U10496 (N_10496,N_9778,N_9596);
nor U10497 (N_10497,N_9525,N_9645);
xnor U10498 (N_10498,N_9915,N_9737);
and U10499 (N_10499,N_9818,N_9964);
xor U10500 (N_10500,N_10013,N_10286);
xnor U10501 (N_10501,N_10300,N_10329);
xor U10502 (N_10502,N_10238,N_10402);
xor U10503 (N_10503,N_10061,N_10060);
nor U10504 (N_10504,N_10012,N_10084);
nand U10505 (N_10505,N_10222,N_10324);
xnor U10506 (N_10506,N_10073,N_10299);
nand U10507 (N_10507,N_10235,N_10115);
nor U10508 (N_10508,N_10215,N_10129);
nor U10509 (N_10509,N_10043,N_10425);
or U10510 (N_10510,N_10135,N_10263);
or U10511 (N_10511,N_10323,N_10478);
or U10512 (N_10512,N_10080,N_10394);
nor U10513 (N_10513,N_10275,N_10145);
xnor U10514 (N_10514,N_10024,N_10033);
xor U10515 (N_10515,N_10314,N_10270);
nand U10516 (N_10516,N_10347,N_10441);
nand U10517 (N_10517,N_10313,N_10417);
xnor U10518 (N_10518,N_10422,N_10220);
xor U10519 (N_10519,N_10136,N_10202);
or U10520 (N_10520,N_10316,N_10130);
nand U10521 (N_10521,N_10030,N_10373);
or U10522 (N_10522,N_10387,N_10424);
xor U10523 (N_10523,N_10230,N_10361);
and U10524 (N_10524,N_10171,N_10332);
nand U10525 (N_10525,N_10040,N_10000);
or U10526 (N_10526,N_10053,N_10267);
or U10527 (N_10527,N_10277,N_10272);
xor U10528 (N_10528,N_10414,N_10208);
nor U10529 (N_10529,N_10365,N_10231);
or U10530 (N_10530,N_10320,N_10391);
and U10531 (N_10531,N_10307,N_10127);
xnor U10532 (N_10532,N_10091,N_10253);
or U10533 (N_10533,N_10195,N_10146);
and U10534 (N_10534,N_10438,N_10315);
and U10535 (N_10535,N_10229,N_10151);
xor U10536 (N_10536,N_10062,N_10183);
and U10537 (N_10537,N_10252,N_10104);
nand U10538 (N_10538,N_10206,N_10047);
xor U10539 (N_10539,N_10228,N_10492);
xor U10540 (N_10540,N_10003,N_10363);
nand U10541 (N_10541,N_10490,N_10039);
and U10542 (N_10542,N_10125,N_10095);
and U10543 (N_10543,N_10430,N_10261);
or U10544 (N_10544,N_10432,N_10065);
nand U10545 (N_10545,N_10297,N_10102);
nand U10546 (N_10546,N_10008,N_10219);
nor U10547 (N_10547,N_10377,N_10395);
and U10548 (N_10548,N_10379,N_10437);
nand U10549 (N_10549,N_10048,N_10167);
nand U10550 (N_10550,N_10243,N_10015);
and U10551 (N_10551,N_10192,N_10173);
nand U10552 (N_10552,N_10210,N_10240);
or U10553 (N_10553,N_10006,N_10093);
and U10554 (N_10554,N_10434,N_10049);
nor U10555 (N_10555,N_10453,N_10353);
nand U10556 (N_10556,N_10152,N_10227);
nand U10557 (N_10557,N_10085,N_10029);
nor U10558 (N_10558,N_10205,N_10489);
or U10559 (N_10559,N_10132,N_10260);
xnor U10560 (N_10560,N_10165,N_10038);
xor U10561 (N_10561,N_10465,N_10462);
nor U10562 (N_10562,N_10249,N_10471);
xor U10563 (N_10563,N_10203,N_10393);
and U10564 (N_10564,N_10472,N_10100);
nor U10565 (N_10565,N_10440,N_10481);
xnor U10566 (N_10566,N_10218,N_10103);
and U10567 (N_10567,N_10367,N_10287);
nand U10568 (N_10568,N_10181,N_10056);
or U10569 (N_10569,N_10058,N_10483);
nor U10570 (N_10570,N_10486,N_10211);
nand U10571 (N_10571,N_10009,N_10431);
and U10572 (N_10572,N_10426,N_10196);
nand U10573 (N_10573,N_10098,N_10031);
nand U10574 (N_10574,N_10390,N_10303);
or U10575 (N_10575,N_10351,N_10294);
and U10576 (N_10576,N_10140,N_10160);
or U10577 (N_10577,N_10467,N_10023);
xor U10578 (N_10578,N_10474,N_10435);
nand U10579 (N_10579,N_10011,N_10381);
nor U10580 (N_10580,N_10449,N_10087);
nor U10581 (N_10581,N_10150,N_10198);
xnor U10582 (N_10582,N_10330,N_10312);
nand U10583 (N_10583,N_10411,N_10439);
nor U10584 (N_10584,N_10289,N_10116);
nor U10585 (N_10585,N_10075,N_10461);
nand U10586 (N_10586,N_10090,N_10068);
and U10587 (N_10587,N_10477,N_10273);
nor U10588 (N_10588,N_10371,N_10427);
nor U10589 (N_10589,N_10027,N_10339);
nand U10590 (N_10590,N_10082,N_10112);
or U10591 (N_10591,N_10436,N_10348);
and U10592 (N_10592,N_10050,N_10178);
nand U10593 (N_10593,N_10405,N_10456);
nor U10594 (N_10594,N_10443,N_10157);
xor U10595 (N_10595,N_10284,N_10460);
nand U10596 (N_10596,N_10185,N_10175);
nand U10597 (N_10597,N_10120,N_10259);
nor U10598 (N_10598,N_10176,N_10199);
xor U10599 (N_10599,N_10459,N_10002);
or U10600 (N_10600,N_10457,N_10473);
or U10601 (N_10601,N_10141,N_10292);
nor U10602 (N_10602,N_10071,N_10366);
and U10603 (N_10603,N_10164,N_10239);
xor U10604 (N_10604,N_10423,N_10233);
and U10605 (N_10605,N_10334,N_10433);
nor U10606 (N_10606,N_10242,N_10020);
or U10607 (N_10607,N_10291,N_10362);
xnor U10608 (N_10608,N_10311,N_10350);
nor U10609 (N_10609,N_10386,N_10126);
nand U10610 (N_10610,N_10216,N_10221);
nor U10611 (N_10611,N_10005,N_10418);
and U10612 (N_10612,N_10207,N_10279);
nor U10613 (N_10613,N_10335,N_10236);
and U10614 (N_10614,N_10118,N_10448);
nor U10615 (N_10615,N_10389,N_10399);
or U10616 (N_10616,N_10293,N_10042);
and U10617 (N_10617,N_10321,N_10147);
and U10618 (N_10618,N_10110,N_10139);
and U10619 (N_10619,N_10026,N_10217);
xnor U10620 (N_10620,N_10143,N_10131);
xnor U10621 (N_10621,N_10213,N_10487);
nor U10622 (N_10622,N_10066,N_10070);
xnor U10623 (N_10623,N_10288,N_10428);
or U10624 (N_10624,N_10370,N_10097);
or U10625 (N_10625,N_10099,N_10072);
nand U10626 (N_10626,N_10480,N_10153);
xnor U10627 (N_10627,N_10336,N_10105);
xor U10628 (N_10628,N_10148,N_10154);
or U10629 (N_10629,N_10309,N_10484);
xor U10630 (N_10630,N_10122,N_10349);
nor U10631 (N_10631,N_10142,N_10032);
or U10632 (N_10632,N_10470,N_10296);
or U10633 (N_10633,N_10283,N_10224);
and U10634 (N_10634,N_10302,N_10276);
or U10635 (N_10635,N_10264,N_10017);
nor U10636 (N_10636,N_10204,N_10114);
and U10637 (N_10637,N_10214,N_10246);
nand U10638 (N_10638,N_10034,N_10403);
xnor U10639 (N_10639,N_10193,N_10086);
and U10640 (N_10640,N_10343,N_10344);
nor U10641 (N_10641,N_10188,N_10451);
nand U10642 (N_10642,N_10016,N_10452);
nor U10643 (N_10643,N_10357,N_10341);
nand U10644 (N_10644,N_10466,N_10212);
and U10645 (N_10645,N_10269,N_10245);
xnor U10646 (N_10646,N_10079,N_10498);
and U10647 (N_10647,N_10191,N_10310);
or U10648 (N_10648,N_10400,N_10375);
nor U10649 (N_10649,N_10429,N_10069);
xor U10650 (N_10650,N_10124,N_10385);
nand U10651 (N_10651,N_10179,N_10159);
and U10652 (N_10652,N_10369,N_10201);
or U10653 (N_10653,N_10162,N_10200);
nor U10654 (N_10654,N_10025,N_10265);
xor U10655 (N_10655,N_10019,N_10244);
and U10656 (N_10656,N_10352,N_10442);
nand U10657 (N_10657,N_10088,N_10223);
xnor U10658 (N_10658,N_10306,N_10144);
or U10659 (N_10659,N_10416,N_10055);
nor U10660 (N_10660,N_10354,N_10186);
nand U10661 (N_10661,N_10010,N_10407);
nand U10662 (N_10662,N_10137,N_10355);
xor U10663 (N_10663,N_10290,N_10446);
and U10664 (N_10664,N_10067,N_10494);
xor U10665 (N_10665,N_10406,N_10096);
or U10666 (N_10666,N_10155,N_10117);
nand U10667 (N_10667,N_10123,N_10057);
nand U10668 (N_10668,N_10014,N_10396);
nand U10669 (N_10669,N_10319,N_10172);
nor U10670 (N_10670,N_10081,N_10021);
nor U10671 (N_10671,N_10378,N_10052);
nor U10672 (N_10672,N_10454,N_10111);
xor U10673 (N_10673,N_10074,N_10078);
or U10674 (N_10674,N_10190,N_10476);
or U10675 (N_10675,N_10168,N_10397);
or U10676 (N_10676,N_10479,N_10285);
xor U10677 (N_10677,N_10464,N_10046);
or U10678 (N_10678,N_10298,N_10359);
nor U10679 (N_10679,N_10475,N_10388);
xnor U10680 (N_10680,N_10237,N_10257);
nand U10681 (N_10681,N_10234,N_10256);
nor U10682 (N_10682,N_10182,N_10495);
xnor U10683 (N_10683,N_10226,N_10333);
nor U10684 (N_10684,N_10189,N_10083);
nor U10685 (N_10685,N_10121,N_10413);
and U10686 (N_10686,N_10419,N_10415);
xnor U10687 (N_10687,N_10404,N_10281);
xnor U10688 (N_10688,N_10177,N_10169);
or U10689 (N_10689,N_10282,N_10001);
and U10690 (N_10690,N_10368,N_10274);
xnor U10691 (N_10691,N_10197,N_10410);
nand U10692 (N_10692,N_10278,N_10251);
nand U10693 (N_10693,N_10496,N_10271);
nor U10694 (N_10694,N_10063,N_10374);
nor U10695 (N_10695,N_10035,N_10345);
xnor U10696 (N_10696,N_10119,N_10308);
nand U10697 (N_10697,N_10163,N_10036);
and U10698 (N_10698,N_10304,N_10051);
and U10699 (N_10699,N_10037,N_10360);
and U10700 (N_10700,N_10340,N_10018);
nand U10701 (N_10701,N_10497,N_10326);
xnor U10702 (N_10702,N_10022,N_10248);
and U10703 (N_10703,N_10262,N_10225);
nor U10704 (N_10704,N_10383,N_10089);
xor U10705 (N_10705,N_10028,N_10392);
nand U10706 (N_10706,N_10187,N_10109);
and U10707 (N_10707,N_10113,N_10158);
nand U10708 (N_10708,N_10133,N_10401);
nand U10709 (N_10709,N_10376,N_10044);
nand U10710 (N_10710,N_10108,N_10134);
nand U10711 (N_10711,N_10059,N_10128);
nor U10712 (N_10712,N_10305,N_10408);
nor U10713 (N_10713,N_10106,N_10325);
nor U10714 (N_10714,N_10255,N_10232);
xor U10715 (N_10715,N_10364,N_10041);
nor U10716 (N_10716,N_10485,N_10076);
nor U10717 (N_10717,N_10170,N_10209);
or U10718 (N_10718,N_10412,N_10382);
nand U10719 (N_10719,N_10444,N_10174);
xor U10720 (N_10720,N_10380,N_10094);
nor U10721 (N_10721,N_10358,N_10346);
nand U10722 (N_10722,N_10101,N_10493);
nand U10723 (N_10723,N_10295,N_10488);
and U10724 (N_10724,N_10447,N_10092);
nor U10725 (N_10725,N_10064,N_10491);
xor U10726 (N_10726,N_10180,N_10445);
nand U10727 (N_10727,N_10337,N_10328);
nor U10728 (N_10728,N_10254,N_10194);
nand U10729 (N_10729,N_10007,N_10482);
or U10730 (N_10730,N_10420,N_10463);
and U10731 (N_10731,N_10469,N_10384);
and U10732 (N_10732,N_10342,N_10054);
nand U10733 (N_10733,N_10327,N_10322);
nand U10734 (N_10734,N_10372,N_10149);
or U10735 (N_10735,N_10184,N_10107);
nor U10736 (N_10736,N_10156,N_10166);
nor U10737 (N_10737,N_10468,N_10356);
nor U10738 (N_10738,N_10077,N_10045);
xnor U10739 (N_10739,N_10318,N_10004);
xnor U10740 (N_10740,N_10250,N_10338);
xnor U10741 (N_10741,N_10421,N_10409);
and U10742 (N_10742,N_10268,N_10450);
nand U10743 (N_10743,N_10398,N_10499);
nor U10744 (N_10744,N_10138,N_10258);
or U10745 (N_10745,N_10331,N_10280);
and U10746 (N_10746,N_10301,N_10458);
nand U10747 (N_10747,N_10455,N_10317);
xnor U10748 (N_10748,N_10161,N_10266);
or U10749 (N_10749,N_10247,N_10241);
nor U10750 (N_10750,N_10036,N_10044);
and U10751 (N_10751,N_10398,N_10016);
nor U10752 (N_10752,N_10388,N_10272);
xnor U10753 (N_10753,N_10061,N_10032);
xor U10754 (N_10754,N_10071,N_10241);
nor U10755 (N_10755,N_10139,N_10232);
and U10756 (N_10756,N_10157,N_10133);
or U10757 (N_10757,N_10319,N_10473);
and U10758 (N_10758,N_10331,N_10337);
nor U10759 (N_10759,N_10371,N_10454);
nor U10760 (N_10760,N_10405,N_10082);
xnor U10761 (N_10761,N_10289,N_10349);
nor U10762 (N_10762,N_10069,N_10321);
nor U10763 (N_10763,N_10064,N_10017);
and U10764 (N_10764,N_10130,N_10126);
and U10765 (N_10765,N_10249,N_10494);
nand U10766 (N_10766,N_10238,N_10214);
or U10767 (N_10767,N_10202,N_10454);
and U10768 (N_10768,N_10059,N_10488);
or U10769 (N_10769,N_10348,N_10075);
xor U10770 (N_10770,N_10012,N_10144);
and U10771 (N_10771,N_10091,N_10172);
xnor U10772 (N_10772,N_10469,N_10256);
nor U10773 (N_10773,N_10312,N_10447);
or U10774 (N_10774,N_10443,N_10299);
nand U10775 (N_10775,N_10404,N_10069);
or U10776 (N_10776,N_10339,N_10153);
nand U10777 (N_10777,N_10158,N_10078);
or U10778 (N_10778,N_10041,N_10291);
and U10779 (N_10779,N_10146,N_10455);
xnor U10780 (N_10780,N_10010,N_10331);
nor U10781 (N_10781,N_10444,N_10134);
and U10782 (N_10782,N_10098,N_10226);
and U10783 (N_10783,N_10344,N_10467);
nor U10784 (N_10784,N_10197,N_10213);
nand U10785 (N_10785,N_10015,N_10113);
nor U10786 (N_10786,N_10135,N_10331);
nand U10787 (N_10787,N_10047,N_10109);
xor U10788 (N_10788,N_10414,N_10127);
and U10789 (N_10789,N_10104,N_10130);
nand U10790 (N_10790,N_10233,N_10231);
and U10791 (N_10791,N_10137,N_10461);
and U10792 (N_10792,N_10490,N_10325);
or U10793 (N_10793,N_10479,N_10343);
nand U10794 (N_10794,N_10047,N_10082);
nand U10795 (N_10795,N_10304,N_10310);
nor U10796 (N_10796,N_10093,N_10427);
xor U10797 (N_10797,N_10163,N_10469);
nor U10798 (N_10798,N_10194,N_10221);
and U10799 (N_10799,N_10138,N_10024);
xor U10800 (N_10800,N_10136,N_10194);
xor U10801 (N_10801,N_10206,N_10413);
or U10802 (N_10802,N_10239,N_10038);
nand U10803 (N_10803,N_10073,N_10489);
or U10804 (N_10804,N_10055,N_10038);
xnor U10805 (N_10805,N_10084,N_10190);
nand U10806 (N_10806,N_10407,N_10372);
nor U10807 (N_10807,N_10184,N_10415);
and U10808 (N_10808,N_10487,N_10291);
xor U10809 (N_10809,N_10156,N_10486);
nor U10810 (N_10810,N_10002,N_10195);
and U10811 (N_10811,N_10340,N_10077);
or U10812 (N_10812,N_10260,N_10141);
nor U10813 (N_10813,N_10196,N_10458);
nor U10814 (N_10814,N_10065,N_10472);
nand U10815 (N_10815,N_10242,N_10481);
and U10816 (N_10816,N_10054,N_10170);
or U10817 (N_10817,N_10468,N_10091);
nand U10818 (N_10818,N_10353,N_10397);
or U10819 (N_10819,N_10008,N_10022);
or U10820 (N_10820,N_10209,N_10155);
nor U10821 (N_10821,N_10172,N_10432);
xnor U10822 (N_10822,N_10092,N_10095);
and U10823 (N_10823,N_10354,N_10337);
or U10824 (N_10824,N_10316,N_10180);
nand U10825 (N_10825,N_10334,N_10171);
nor U10826 (N_10826,N_10092,N_10052);
nand U10827 (N_10827,N_10457,N_10463);
or U10828 (N_10828,N_10091,N_10030);
or U10829 (N_10829,N_10303,N_10009);
nor U10830 (N_10830,N_10156,N_10094);
nand U10831 (N_10831,N_10445,N_10245);
xnor U10832 (N_10832,N_10174,N_10272);
and U10833 (N_10833,N_10289,N_10210);
xor U10834 (N_10834,N_10276,N_10090);
or U10835 (N_10835,N_10209,N_10135);
xor U10836 (N_10836,N_10072,N_10261);
nand U10837 (N_10837,N_10118,N_10135);
and U10838 (N_10838,N_10392,N_10361);
xor U10839 (N_10839,N_10000,N_10484);
xnor U10840 (N_10840,N_10467,N_10012);
and U10841 (N_10841,N_10383,N_10092);
or U10842 (N_10842,N_10042,N_10410);
nand U10843 (N_10843,N_10034,N_10198);
and U10844 (N_10844,N_10373,N_10364);
nand U10845 (N_10845,N_10138,N_10190);
xnor U10846 (N_10846,N_10055,N_10123);
and U10847 (N_10847,N_10491,N_10094);
xor U10848 (N_10848,N_10463,N_10389);
and U10849 (N_10849,N_10372,N_10408);
or U10850 (N_10850,N_10372,N_10324);
and U10851 (N_10851,N_10240,N_10251);
and U10852 (N_10852,N_10103,N_10306);
xor U10853 (N_10853,N_10229,N_10066);
nor U10854 (N_10854,N_10289,N_10357);
and U10855 (N_10855,N_10208,N_10190);
nand U10856 (N_10856,N_10385,N_10402);
xor U10857 (N_10857,N_10215,N_10199);
and U10858 (N_10858,N_10038,N_10017);
and U10859 (N_10859,N_10298,N_10409);
or U10860 (N_10860,N_10330,N_10203);
and U10861 (N_10861,N_10152,N_10388);
nand U10862 (N_10862,N_10010,N_10374);
xnor U10863 (N_10863,N_10343,N_10250);
or U10864 (N_10864,N_10313,N_10422);
and U10865 (N_10865,N_10066,N_10402);
and U10866 (N_10866,N_10478,N_10488);
and U10867 (N_10867,N_10479,N_10421);
xor U10868 (N_10868,N_10418,N_10057);
or U10869 (N_10869,N_10117,N_10294);
or U10870 (N_10870,N_10379,N_10158);
nand U10871 (N_10871,N_10445,N_10008);
xnor U10872 (N_10872,N_10096,N_10421);
or U10873 (N_10873,N_10215,N_10184);
xnor U10874 (N_10874,N_10385,N_10367);
xor U10875 (N_10875,N_10004,N_10416);
nor U10876 (N_10876,N_10270,N_10416);
nor U10877 (N_10877,N_10337,N_10499);
nor U10878 (N_10878,N_10134,N_10095);
and U10879 (N_10879,N_10451,N_10398);
nor U10880 (N_10880,N_10486,N_10264);
xor U10881 (N_10881,N_10371,N_10363);
nor U10882 (N_10882,N_10201,N_10248);
nor U10883 (N_10883,N_10409,N_10053);
xor U10884 (N_10884,N_10329,N_10473);
nand U10885 (N_10885,N_10022,N_10157);
and U10886 (N_10886,N_10461,N_10497);
and U10887 (N_10887,N_10477,N_10225);
or U10888 (N_10888,N_10346,N_10232);
or U10889 (N_10889,N_10098,N_10329);
nor U10890 (N_10890,N_10153,N_10295);
xor U10891 (N_10891,N_10490,N_10487);
nor U10892 (N_10892,N_10012,N_10026);
and U10893 (N_10893,N_10112,N_10345);
nand U10894 (N_10894,N_10119,N_10462);
nor U10895 (N_10895,N_10119,N_10314);
and U10896 (N_10896,N_10469,N_10102);
and U10897 (N_10897,N_10137,N_10425);
and U10898 (N_10898,N_10355,N_10237);
xnor U10899 (N_10899,N_10075,N_10016);
xnor U10900 (N_10900,N_10199,N_10226);
and U10901 (N_10901,N_10335,N_10162);
and U10902 (N_10902,N_10179,N_10385);
xnor U10903 (N_10903,N_10284,N_10088);
nand U10904 (N_10904,N_10011,N_10480);
xnor U10905 (N_10905,N_10199,N_10127);
or U10906 (N_10906,N_10308,N_10186);
and U10907 (N_10907,N_10138,N_10240);
and U10908 (N_10908,N_10342,N_10049);
or U10909 (N_10909,N_10283,N_10209);
nand U10910 (N_10910,N_10315,N_10261);
and U10911 (N_10911,N_10023,N_10448);
xnor U10912 (N_10912,N_10157,N_10281);
and U10913 (N_10913,N_10454,N_10429);
and U10914 (N_10914,N_10266,N_10013);
and U10915 (N_10915,N_10161,N_10271);
and U10916 (N_10916,N_10366,N_10369);
or U10917 (N_10917,N_10410,N_10232);
or U10918 (N_10918,N_10269,N_10274);
or U10919 (N_10919,N_10395,N_10364);
nor U10920 (N_10920,N_10337,N_10358);
xor U10921 (N_10921,N_10369,N_10060);
nand U10922 (N_10922,N_10025,N_10165);
and U10923 (N_10923,N_10286,N_10233);
nor U10924 (N_10924,N_10049,N_10099);
or U10925 (N_10925,N_10052,N_10104);
xnor U10926 (N_10926,N_10109,N_10340);
xnor U10927 (N_10927,N_10281,N_10495);
nor U10928 (N_10928,N_10301,N_10426);
and U10929 (N_10929,N_10220,N_10395);
xor U10930 (N_10930,N_10183,N_10040);
or U10931 (N_10931,N_10166,N_10349);
and U10932 (N_10932,N_10467,N_10392);
xnor U10933 (N_10933,N_10238,N_10045);
or U10934 (N_10934,N_10498,N_10367);
nor U10935 (N_10935,N_10269,N_10256);
nand U10936 (N_10936,N_10092,N_10264);
or U10937 (N_10937,N_10000,N_10261);
nand U10938 (N_10938,N_10265,N_10339);
nor U10939 (N_10939,N_10255,N_10003);
and U10940 (N_10940,N_10219,N_10320);
or U10941 (N_10941,N_10435,N_10128);
nor U10942 (N_10942,N_10402,N_10455);
and U10943 (N_10943,N_10341,N_10258);
xor U10944 (N_10944,N_10339,N_10379);
and U10945 (N_10945,N_10411,N_10004);
and U10946 (N_10946,N_10439,N_10019);
and U10947 (N_10947,N_10236,N_10009);
and U10948 (N_10948,N_10406,N_10421);
and U10949 (N_10949,N_10293,N_10405);
nor U10950 (N_10950,N_10271,N_10343);
or U10951 (N_10951,N_10128,N_10208);
and U10952 (N_10952,N_10450,N_10430);
or U10953 (N_10953,N_10304,N_10176);
nand U10954 (N_10954,N_10369,N_10154);
or U10955 (N_10955,N_10383,N_10309);
xnor U10956 (N_10956,N_10215,N_10494);
or U10957 (N_10957,N_10125,N_10356);
xor U10958 (N_10958,N_10482,N_10460);
nand U10959 (N_10959,N_10039,N_10323);
or U10960 (N_10960,N_10406,N_10015);
xnor U10961 (N_10961,N_10316,N_10007);
and U10962 (N_10962,N_10266,N_10301);
and U10963 (N_10963,N_10114,N_10412);
xor U10964 (N_10964,N_10478,N_10076);
nor U10965 (N_10965,N_10460,N_10262);
nor U10966 (N_10966,N_10173,N_10229);
and U10967 (N_10967,N_10067,N_10377);
and U10968 (N_10968,N_10236,N_10392);
or U10969 (N_10969,N_10276,N_10469);
or U10970 (N_10970,N_10385,N_10230);
nand U10971 (N_10971,N_10407,N_10062);
nor U10972 (N_10972,N_10320,N_10041);
or U10973 (N_10973,N_10376,N_10190);
nand U10974 (N_10974,N_10412,N_10060);
nand U10975 (N_10975,N_10416,N_10161);
nand U10976 (N_10976,N_10476,N_10108);
or U10977 (N_10977,N_10266,N_10327);
nor U10978 (N_10978,N_10412,N_10062);
nor U10979 (N_10979,N_10240,N_10454);
nand U10980 (N_10980,N_10250,N_10266);
nand U10981 (N_10981,N_10141,N_10484);
or U10982 (N_10982,N_10050,N_10439);
nor U10983 (N_10983,N_10041,N_10028);
nor U10984 (N_10984,N_10294,N_10480);
nand U10985 (N_10985,N_10199,N_10223);
xor U10986 (N_10986,N_10079,N_10162);
or U10987 (N_10987,N_10030,N_10385);
or U10988 (N_10988,N_10180,N_10273);
and U10989 (N_10989,N_10443,N_10045);
nor U10990 (N_10990,N_10025,N_10099);
or U10991 (N_10991,N_10028,N_10291);
and U10992 (N_10992,N_10119,N_10218);
or U10993 (N_10993,N_10252,N_10213);
nor U10994 (N_10994,N_10473,N_10301);
nor U10995 (N_10995,N_10273,N_10475);
nand U10996 (N_10996,N_10112,N_10460);
xor U10997 (N_10997,N_10342,N_10115);
nand U10998 (N_10998,N_10447,N_10473);
or U10999 (N_10999,N_10412,N_10046);
or U11000 (N_11000,N_10923,N_10886);
xnor U11001 (N_11001,N_10604,N_10813);
nand U11002 (N_11002,N_10748,N_10721);
xnor U11003 (N_11003,N_10883,N_10808);
or U11004 (N_11004,N_10908,N_10733);
or U11005 (N_11005,N_10595,N_10516);
nand U11006 (N_11006,N_10567,N_10824);
and U11007 (N_11007,N_10788,N_10834);
and U11008 (N_11008,N_10718,N_10769);
and U11009 (N_11009,N_10662,N_10511);
xnor U11010 (N_11010,N_10901,N_10587);
xnor U11011 (N_11011,N_10907,N_10905);
nor U11012 (N_11012,N_10720,N_10641);
nand U11013 (N_11013,N_10770,N_10805);
nand U11014 (N_11014,N_10759,N_10583);
nand U11015 (N_11015,N_10543,N_10727);
or U11016 (N_11016,N_10990,N_10958);
xnor U11017 (N_11017,N_10730,N_10609);
and U11018 (N_11018,N_10622,N_10625);
xor U11019 (N_11019,N_10779,N_10508);
xor U11020 (N_11020,N_10700,N_10763);
or U11021 (N_11021,N_10984,N_10957);
nand U11022 (N_11022,N_10650,N_10776);
xnor U11023 (N_11023,N_10585,N_10642);
and U11024 (N_11024,N_10894,N_10869);
or U11025 (N_11025,N_10684,N_10519);
or U11026 (N_11026,N_10986,N_10814);
and U11027 (N_11027,N_10826,N_10610);
and U11028 (N_11028,N_10971,N_10955);
nand U11029 (N_11029,N_10888,N_10688);
or U11030 (N_11030,N_10995,N_10784);
xnor U11031 (N_11031,N_10638,N_10956);
or U11032 (N_11032,N_10938,N_10945);
xnor U11033 (N_11033,N_10860,N_10649);
and U11034 (N_11034,N_10674,N_10941);
nand U11035 (N_11035,N_10676,N_10996);
and U11036 (N_11036,N_10829,N_10856);
and U11037 (N_11037,N_10812,N_10836);
and U11038 (N_11038,N_10513,N_10906);
and U11039 (N_11039,N_10879,N_10538);
nor U11040 (N_11040,N_10618,N_10589);
xor U11041 (N_11041,N_10600,N_10507);
nor U11042 (N_11042,N_10991,N_10821);
xor U11043 (N_11043,N_10789,N_10777);
and U11044 (N_11044,N_10708,N_10668);
nor U11045 (N_11045,N_10741,N_10503);
or U11046 (N_11046,N_10963,N_10531);
and U11047 (N_11047,N_10659,N_10796);
or U11048 (N_11048,N_10695,N_10505);
or U11049 (N_11049,N_10732,N_10870);
and U11050 (N_11050,N_10702,N_10540);
xor U11051 (N_11051,N_10847,N_10988);
xnor U11052 (N_11052,N_10564,N_10675);
nand U11053 (N_11053,N_10857,N_10555);
nand U11054 (N_11054,N_10500,N_10950);
nor U11055 (N_11055,N_10739,N_10672);
nor U11056 (N_11056,N_10933,N_10530);
or U11057 (N_11057,N_10736,N_10539);
or U11058 (N_11058,N_10939,N_10645);
xnor U11059 (N_11059,N_10717,N_10854);
and U11060 (N_11060,N_10707,N_10795);
or U11061 (N_11061,N_10782,N_10635);
or U11062 (N_11062,N_10900,N_10859);
nor U11063 (N_11063,N_10517,N_10831);
xnor U11064 (N_11064,N_10630,N_10999);
or U11065 (N_11065,N_10764,N_10877);
nand U11066 (N_11066,N_10837,N_10974);
or U11067 (N_11067,N_10897,N_10588);
nand U11068 (N_11068,N_10528,N_10937);
and U11069 (N_11069,N_10767,N_10623);
nor U11070 (N_11070,N_10822,N_10644);
and U11071 (N_11071,N_10802,N_10799);
and U11072 (N_11072,N_10863,N_10873);
and U11073 (N_11073,N_10801,N_10646);
or U11074 (N_11074,N_10929,N_10692);
or U11075 (N_11075,N_10534,N_10580);
nand U11076 (N_11076,N_10669,N_10994);
nand U11077 (N_11077,N_10792,N_10849);
nor U11078 (N_11078,N_10755,N_10568);
nor U11079 (N_11079,N_10554,N_10791);
or U11080 (N_11080,N_10798,N_10656);
and U11081 (N_11081,N_10615,N_10846);
xnor U11082 (N_11082,N_10576,N_10940);
or U11083 (N_11083,N_10689,N_10780);
nor U11084 (N_11084,N_10607,N_10880);
or U11085 (N_11085,N_10614,N_10872);
nor U11086 (N_11086,N_10713,N_10816);
and U11087 (N_11087,N_10734,N_10606);
or U11088 (N_11088,N_10603,N_10919);
nor U11089 (N_11089,N_10670,N_10922);
nor U11090 (N_11090,N_10616,N_10895);
and U11091 (N_11091,N_10552,N_10850);
or U11092 (N_11092,N_10876,N_10632);
and U11093 (N_11093,N_10914,N_10743);
xor U11094 (N_11094,N_10811,N_10778);
and U11095 (N_11095,N_10572,N_10740);
or U11096 (N_11096,N_10570,N_10673);
and U11097 (N_11097,N_10785,N_10989);
nor U11098 (N_11098,N_10709,N_10651);
or U11099 (N_11099,N_10865,N_10719);
and U11100 (N_11100,N_10557,N_10896);
nand U11101 (N_11101,N_10874,N_10648);
or U11102 (N_11102,N_10993,N_10611);
nor U11103 (N_11103,N_10680,N_10591);
and U11104 (N_11104,N_10526,N_10553);
and U11105 (N_11105,N_10928,N_10613);
or U11106 (N_11106,N_10547,N_10696);
nor U11107 (N_11107,N_10884,N_10504);
or U11108 (N_11108,N_10664,N_10890);
nor U11109 (N_11109,N_10620,N_10742);
xnor U11110 (N_11110,N_10828,N_10746);
nand U11111 (N_11111,N_10525,N_10545);
or U11112 (N_11112,N_10946,N_10617);
nor U11113 (N_11113,N_10965,N_10703);
nor U11114 (N_11114,N_10749,N_10571);
or U11115 (N_11115,N_10514,N_10934);
xor U11116 (N_11116,N_10686,N_10842);
xor U11117 (N_11117,N_10819,N_10601);
nor U11118 (N_11118,N_10992,N_10637);
nor U11119 (N_11119,N_10862,N_10705);
or U11120 (N_11120,N_10731,N_10775);
nor U11121 (N_11121,N_10577,N_10581);
xnor U11122 (N_11122,N_10747,N_10744);
and U11123 (N_11123,N_10925,N_10735);
xnor U11124 (N_11124,N_10579,N_10712);
xnor U11125 (N_11125,N_10520,N_10927);
nand U11126 (N_11126,N_10948,N_10685);
xnor U11127 (N_11127,N_10605,N_10726);
nand U11128 (N_11128,N_10771,N_10845);
and U11129 (N_11129,N_10871,N_10760);
or U11130 (N_11130,N_10930,N_10982);
nand U11131 (N_11131,N_10977,N_10521);
nand U11132 (N_11132,N_10921,N_10947);
xor U11133 (N_11133,N_10597,N_10682);
or U11134 (N_11134,N_10858,N_10599);
nor U11135 (N_11135,N_10536,N_10839);
and U11136 (N_11136,N_10754,N_10772);
nor U11137 (N_11137,N_10912,N_10657);
nor U11138 (N_11138,N_10586,N_10968);
or U11139 (N_11139,N_10810,N_10537);
nor U11140 (N_11140,N_10952,N_10745);
or U11141 (N_11141,N_10626,N_10882);
nand U11142 (N_11142,N_10911,N_10691);
nor U11143 (N_11143,N_10924,N_10833);
and U11144 (N_11144,N_10594,N_10851);
and U11145 (N_11145,N_10861,N_10962);
nor U11146 (N_11146,N_10885,N_10729);
nand U11147 (N_11147,N_10596,N_10843);
and U11148 (N_11148,N_10830,N_10578);
xor U11149 (N_11149,N_10681,N_10752);
nand U11150 (N_11150,N_10631,N_10502);
nand U11151 (N_11151,N_10926,N_10844);
and U11152 (N_11152,N_10690,N_10960);
xnor U11153 (N_11153,N_10549,N_10660);
nand U11154 (N_11154,N_10898,N_10711);
and U11155 (N_11155,N_10766,N_10809);
xnor U11156 (N_11156,N_10509,N_10817);
nor U11157 (N_11157,N_10550,N_10556);
xor U11158 (N_11158,N_10679,N_10935);
and U11159 (N_11159,N_10698,N_10797);
nor U11160 (N_11160,N_10751,N_10942);
xnor U11161 (N_11161,N_10997,N_10574);
nor U11162 (N_11162,N_10533,N_10909);
and U11163 (N_11163,N_10697,N_10608);
nor U11164 (N_11164,N_10541,N_10501);
or U11165 (N_11165,N_10762,N_10818);
nand U11166 (N_11166,N_10915,N_10665);
nor U11167 (N_11167,N_10820,N_10724);
and U11168 (N_11168,N_10979,N_10667);
nor U11169 (N_11169,N_10619,N_10584);
xor U11170 (N_11170,N_10804,N_10640);
nand U11171 (N_11171,N_10853,N_10881);
xor U11172 (N_11172,N_10978,N_10867);
nor U11173 (N_11173,N_10967,N_10949);
or U11174 (N_11174,N_10562,N_10918);
xor U11175 (N_11175,N_10983,N_10544);
and U11176 (N_11176,N_10633,N_10981);
nor U11177 (N_11177,N_10756,N_10786);
xor U11178 (N_11178,N_10551,N_10980);
or U11179 (N_11179,N_10823,N_10899);
xnor U11180 (N_11180,N_10987,N_10563);
or U11181 (N_11181,N_10694,N_10548);
and U11182 (N_11182,N_10728,N_10561);
nor U11183 (N_11183,N_10639,N_10806);
xor U11184 (N_11184,N_10781,N_10913);
nor U11185 (N_11185,N_10868,N_10566);
xnor U11186 (N_11186,N_10864,N_10532);
xor U11187 (N_11187,N_10893,N_10838);
and U11188 (N_11188,N_10954,N_10904);
nor U11189 (N_11189,N_10590,N_10943);
nand U11190 (N_11190,N_10953,N_10753);
or U11191 (N_11191,N_10969,N_10598);
nand U11192 (N_11192,N_10663,N_10790);
and U11193 (N_11193,N_10661,N_10787);
or U11194 (N_11194,N_10774,N_10693);
nand U11195 (N_11195,N_10931,N_10524);
nor U11196 (N_11196,N_10973,N_10917);
and U11197 (N_11197,N_10757,N_10621);
xor U11198 (N_11198,N_10783,N_10624);
or U11199 (N_11199,N_10527,N_10878);
xnor U11200 (N_11200,N_10773,N_10506);
nor U11201 (N_11201,N_10737,N_10723);
and U11202 (N_11202,N_10964,N_10841);
and U11203 (N_11203,N_10903,N_10518);
nand U11204 (N_11204,N_10529,N_10951);
xnor U11205 (N_11205,N_10800,N_10510);
and U11206 (N_11206,N_10875,N_10891);
nand U11207 (N_11207,N_10629,N_10835);
nand U11208 (N_11208,N_10827,N_10815);
nor U11209 (N_11209,N_10592,N_10636);
nand U11210 (N_11210,N_10654,N_10716);
xor U11211 (N_11211,N_10569,N_10852);
or U11212 (N_11212,N_10612,N_10655);
xor U11213 (N_11213,N_10546,N_10683);
and U11214 (N_11214,N_10765,N_10643);
and U11215 (N_11215,N_10560,N_10970);
or U11216 (N_11216,N_10565,N_10704);
nand U11217 (N_11217,N_10701,N_10807);
xor U11218 (N_11218,N_10866,N_10558);
nor U11219 (N_11219,N_10602,N_10722);
nand U11220 (N_11220,N_10593,N_10658);
xnor U11221 (N_11221,N_10710,N_10768);
and U11222 (N_11222,N_10523,N_10961);
xnor U11223 (N_11223,N_10535,N_10634);
nand U11224 (N_11224,N_10855,N_10515);
and U11225 (N_11225,N_10892,N_10666);
nand U11226 (N_11226,N_10738,N_10652);
or U11227 (N_11227,N_10944,N_10976);
xnor U11228 (N_11228,N_10832,N_10889);
nor U11229 (N_11229,N_10542,N_10932);
and U11230 (N_11230,N_10653,N_10575);
and U11231 (N_11231,N_10936,N_10975);
nor U11232 (N_11232,N_10920,N_10761);
or U11233 (N_11233,N_10627,N_10825);
and U11234 (N_11234,N_10910,N_10793);
xor U11235 (N_11235,N_10750,N_10706);
nand U11236 (N_11236,N_10671,N_10902);
or U11237 (N_11237,N_10559,N_10998);
nand U11238 (N_11238,N_10522,N_10887);
or U11239 (N_11239,N_10715,N_10972);
nor U11240 (N_11240,N_10840,N_10699);
xnor U11241 (N_11241,N_10916,N_10966);
xor U11242 (N_11242,N_10512,N_10758);
and U11243 (N_11243,N_10628,N_10803);
nand U11244 (N_11244,N_10714,N_10725);
and U11245 (N_11245,N_10794,N_10985);
xnor U11246 (N_11246,N_10573,N_10678);
nand U11247 (N_11247,N_10848,N_10959);
or U11248 (N_11248,N_10647,N_10687);
or U11249 (N_11249,N_10582,N_10677);
nand U11250 (N_11250,N_10897,N_10965);
or U11251 (N_11251,N_10596,N_10640);
nand U11252 (N_11252,N_10610,N_10531);
nor U11253 (N_11253,N_10582,N_10735);
xor U11254 (N_11254,N_10889,N_10534);
and U11255 (N_11255,N_10924,N_10915);
xor U11256 (N_11256,N_10863,N_10588);
or U11257 (N_11257,N_10853,N_10900);
or U11258 (N_11258,N_10801,N_10549);
or U11259 (N_11259,N_10688,N_10713);
and U11260 (N_11260,N_10962,N_10707);
and U11261 (N_11261,N_10955,N_10802);
and U11262 (N_11262,N_10893,N_10515);
or U11263 (N_11263,N_10960,N_10905);
and U11264 (N_11264,N_10766,N_10732);
and U11265 (N_11265,N_10907,N_10856);
xor U11266 (N_11266,N_10871,N_10777);
or U11267 (N_11267,N_10634,N_10868);
or U11268 (N_11268,N_10535,N_10587);
xnor U11269 (N_11269,N_10552,N_10963);
or U11270 (N_11270,N_10504,N_10690);
or U11271 (N_11271,N_10611,N_10864);
nor U11272 (N_11272,N_10642,N_10524);
and U11273 (N_11273,N_10536,N_10539);
nand U11274 (N_11274,N_10733,N_10835);
and U11275 (N_11275,N_10629,N_10610);
nor U11276 (N_11276,N_10903,N_10557);
nand U11277 (N_11277,N_10995,N_10947);
and U11278 (N_11278,N_10567,N_10751);
nand U11279 (N_11279,N_10697,N_10675);
xnor U11280 (N_11280,N_10756,N_10864);
nand U11281 (N_11281,N_10537,N_10964);
or U11282 (N_11282,N_10916,N_10700);
nor U11283 (N_11283,N_10566,N_10786);
and U11284 (N_11284,N_10950,N_10551);
and U11285 (N_11285,N_10690,N_10516);
nand U11286 (N_11286,N_10668,N_10684);
and U11287 (N_11287,N_10546,N_10605);
nand U11288 (N_11288,N_10907,N_10792);
xor U11289 (N_11289,N_10511,N_10805);
nand U11290 (N_11290,N_10502,N_10519);
nand U11291 (N_11291,N_10677,N_10970);
or U11292 (N_11292,N_10704,N_10787);
xnor U11293 (N_11293,N_10906,N_10864);
and U11294 (N_11294,N_10840,N_10918);
xnor U11295 (N_11295,N_10988,N_10969);
or U11296 (N_11296,N_10993,N_10737);
or U11297 (N_11297,N_10578,N_10832);
or U11298 (N_11298,N_10788,N_10847);
or U11299 (N_11299,N_10914,N_10823);
nor U11300 (N_11300,N_10758,N_10935);
xnor U11301 (N_11301,N_10611,N_10667);
or U11302 (N_11302,N_10811,N_10542);
and U11303 (N_11303,N_10543,N_10924);
xor U11304 (N_11304,N_10707,N_10984);
nor U11305 (N_11305,N_10794,N_10619);
xnor U11306 (N_11306,N_10555,N_10915);
nand U11307 (N_11307,N_10834,N_10509);
nand U11308 (N_11308,N_10526,N_10814);
nor U11309 (N_11309,N_10803,N_10749);
xor U11310 (N_11310,N_10574,N_10528);
nor U11311 (N_11311,N_10584,N_10568);
nor U11312 (N_11312,N_10683,N_10650);
or U11313 (N_11313,N_10577,N_10939);
or U11314 (N_11314,N_10680,N_10961);
or U11315 (N_11315,N_10981,N_10864);
xnor U11316 (N_11316,N_10891,N_10872);
or U11317 (N_11317,N_10636,N_10818);
or U11318 (N_11318,N_10992,N_10639);
or U11319 (N_11319,N_10607,N_10873);
or U11320 (N_11320,N_10862,N_10993);
or U11321 (N_11321,N_10746,N_10538);
nor U11322 (N_11322,N_10525,N_10860);
and U11323 (N_11323,N_10517,N_10923);
and U11324 (N_11324,N_10813,N_10643);
and U11325 (N_11325,N_10761,N_10818);
nor U11326 (N_11326,N_10759,N_10808);
and U11327 (N_11327,N_10963,N_10797);
and U11328 (N_11328,N_10567,N_10995);
xor U11329 (N_11329,N_10759,N_10713);
xor U11330 (N_11330,N_10691,N_10920);
or U11331 (N_11331,N_10504,N_10836);
or U11332 (N_11332,N_10977,N_10687);
nor U11333 (N_11333,N_10530,N_10765);
xnor U11334 (N_11334,N_10678,N_10749);
and U11335 (N_11335,N_10854,N_10572);
xor U11336 (N_11336,N_10660,N_10760);
and U11337 (N_11337,N_10976,N_10685);
xor U11338 (N_11338,N_10711,N_10988);
nand U11339 (N_11339,N_10890,N_10513);
nor U11340 (N_11340,N_10579,N_10525);
or U11341 (N_11341,N_10982,N_10634);
nand U11342 (N_11342,N_10927,N_10733);
nor U11343 (N_11343,N_10692,N_10630);
xnor U11344 (N_11344,N_10540,N_10899);
xor U11345 (N_11345,N_10685,N_10917);
and U11346 (N_11346,N_10716,N_10506);
nand U11347 (N_11347,N_10793,N_10549);
and U11348 (N_11348,N_10897,N_10740);
or U11349 (N_11349,N_10546,N_10725);
xnor U11350 (N_11350,N_10509,N_10516);
or U11351 (N_11351,N_10889,N_10660);
and U11352 (N_11352,N_10908,N_10725);
and U11353 (N_11353,N_10549,N_10671);
xor U11354 (N_11354,N_10845,N_10858);
or U11355 (N_11355,N_10529,N_10727);
and U11356 (N_11356,N_10852,N_10720);
or U11357 (N_11357,N_10690,N_10981);
nor U11358 (N_11358,N_10908,N_10827);
nor U11359 (N_11359,N_10501,N_10890);
or U11360 (N_11360,N_10703,N_10577);
nand U11361 (N_11361,N_10584,N_10670);
nand U11362 (N_11362,N_10962,N_10677);
xnor U11363 (N_11363,N_10801,N_10940);
nand U11364 (N_11364,N_10525,N_10741);
xnor U11365 (N_11365,N_10855,N_10825);
nand U11366 (N_11366,N_10843,N_10963);
nand U11367 (N_11367,N_10807,N_10659);
xor U11368 (N_11368,N_10805,N_10582);
nor U11369 (N_11369,N_10783,N_10656);
nor U11370 (N_11370,N_10950,N_10577);
nor U11371 (N_11371,N_10731,N_10726);
or U11372 (N_11372,N_10758,N_10814);
nor U11373 (N_11373,N_10513,N_10951);
nor U11374 (N_11374,N_10870,N_10646);
xnor U11375 (N_11375,N_10759,N_10928);
and U11376 (N_11376,N_10670,N_10673);
nor U11377 (N_11377,N_10515,N_10781);
or U11378 (N_11378,N_10881,N_10855);
nand U11379 (N_11379,N_10813,N_10883);
nand U11380 (N_11380,N_10924,N_10769);
xor U11381 (N_11381,N_10927,N_10512);
xor U11382 (N_11382,N_10599,N_10959);
xor U11383 (N_11383,N_10761,N_10815);
and U11384 (N_11384,N_10502,N_10671);
nand U11385 (N_11385,N_10689,N_10700);
nand U11386 (N_11386,N_10644,N_10800);
and U11387 (N_11387,N_10748,N_10907);
nor U11388 (N_11388,N_10720,N_10526);
xor U11389 (N_11389,N_10641,N_10725);
nor U11390 (N_11390,N_10645,N_10921);
nand U11391 (N_11391,N_10735,N_10623);
nand U11392 (N_11392,N_10979,N_10799);
nand U11393 (N_11393,N_10875,N_10709);
and U11394 (N_11394,N_10849,N_10521);
and U11395 (N_11395,N_10862,N_10516);
and U11396 (N_11396,N_10957,N_10530);
and U11397 (N_11397,N_10535,N_10719);
nor U11398 (N_11398,N_10726,N_10517);
nor U11399 (N_11399,N_10564,N_10723);
xnor U11400 (N_11400,N_10723,N_10642);
nor U11401 (N_11401,N_10612,N_10784);
nand U11402 (N_11402,N_10522,N_10909);
nor U11403 (N_11403,N_10687,N_10950);
nand U11404 (N_11404,N_10641,N_10920);
xnor U11405 (N_11405,N_10615,N_10790);
nand U11406 (N_11406,N_10519,N_10552);
nor U11407 (N_11407,N_10521,N_10736);
or U11408 (N_11408,N_10909,N_10776);
nand U11409 (N_11409,N_10690,N_10587);
xor U11410 (N_11410,N_10758,N_10718);
xnor U11411 (N_11411,N_10651,N_10603);
nor U11412 (N_11412,N_10707,N_10783);
nand U11413 (N_11413,N_10874,N_10944);
nor U11414 (N_11414,N_10802,N_10916);
and U11415 (N_11415,N_10647,N_10759);
and U11416 (N_11416,N_10748,N_10706);
and U11417 (N_11417,N_10899,N_10908);
and U11418 (N_11418,N_10525,N_10856);
nor U11419 (N_11419,N_10799,N_10789);
nand U11420 (N_11420,N_10513,N_10519);
xnor U11421 (N_11421,N_10787,N_10531);
xnor U11422 (N_11422,N_10822,N_10582);
nand U11423 (N_11423,N_10661,N_10591);
nor U11424 (N_11424,N_10878,N_10787);
nor U11425 (N_11425,N_10718,N_10689);
nor U11426 (N_11426,N_10801,N_10928);
nand U11427 (N_11427,N_10891,N_10758);
and U11428 (N_11428,N_10790,N_10986);
or U11429 (N_11429,N_10975,N_10522);
nor U11430 (N_11430,N_10559,N_10671);
nor U11431 (N_11431,N_10664,N_10821);
and U11432 (N_11432,N_10548,N_10910);
xnor U11433 (N_11433,N_10626,N_10726);
xor U11434 (N_11434,N_10667,N_10735);
and U11435 (N_11435,N_10923,N_10530);
and U11436 (N_11436,N_10766,N_10762);
nand U11437 (N_11437,N_10750,N_10858);
nand U11438 (N_11438,N_10965,N_10544);
or U11439 (N_11439,N_10950,N_10931);
or U11440 (N_11440,N_10982,N_10539);
nand U11441 (N_11441,N_10725,N_10699);
and U11442 (N_11442,N_10678,N_10775);
and U11443 (N_11443,N_10873,N_10593);
nand U11444 (N_11444,N_10738,N_10987);
nor U11445 (N_11445,N_10642,N_10768);
or U11446 (N_11446,N_10747,N_10599);
or U11447 (N_11447,N_10862,N_10572);
nand U11448 (N_11448,N_10863,N_10691);
or U11449 (N_11449,N_10567,N_10538);
nand U11450 (N_11450,N_10958,N_10694);
xor U11451 (N_11451,N_10907,N_10718);
nor U11452 (N_11452,N_10599,N_10907);
and U11453 (N_11453,N_10549,N_10658);
xnor U11454 (N_11454,N_10503,N_10591);
xnor U11455 (N_11455,N_10923,N_10573);
nand U11456 (N_11456,N_10839,N_10654);
nand U11457 (N_11457,N_10756,N_10510);
nand U11458 (N_11458,N_10907,N_10732);
nand U11459 (N_11459,N_10968,N_10685);
and U11460 (N_11460,N_10840,N_10994);
or U11461 (N_11461,N_10649,N_10811);
or U11462 (N_11462,N_10705,N_10960);
and U11463 (N_11463,N_10661,N_10877);
nand U11464 (N_11464,N_10533,N_10558);
nand U11465 (N_11465,N_10544,N_10609);
xnor U11466 (N_11466,N_10843,N_10732);
or U11467 (N_11467,N_10861,N_10904);
or U11468 (N_11468,N_10944,N_10661);
and U11469 (N_11469,N_10753,N_10831);
nor U11470 (N_11470,N_10855,N_10999);
nor U11471 (N_11471,N_10920,N_10646);
nor U11472 (N_11472,N_10518,N_10500);
and U11473 (N_11473,N_10550,N_10571);
nand U11474 (N_11474,N_10527,N_10510);
nand U11475 (N_11475,N_10680,N_10744);
and U11476 (N_11476,N_10802,N_10772);
nand U11477 (N_11477,N_10775,N_10894);
nand U11478 (N_11478,N_10971,N_10761);
xor U11479 (N_11479,N_10598,N_10611);
xnor U11480 (N_11480,N_10910,N_10530);
nand U11481 (N_11481,N_10962,N_10910);
xor U11482 (N_11482,N_10680,N_10702);
and U11483 (N_11483,N_10972,N_10622);
and U11484 (N_11484,N_10666,N_10567);
and U11485 (N_11485,N_10582,N_10511);
and U11486 (N_11486,N_10838,N_10909);
or U11487 (N_11487,N_10879,N_10795);
and U11488 (N_11488,N_10914,N_10549);
xnor U11489 (N_11489,N_10951,N_10850);
nand U11490 (N_11490,N_10527,N_10542);
nor U11491 (N_11491,N_10919,N_10932);
or U11492 (N_11492,N_10686,N_10858);
xnor U11493 (N_11493,N_10840,N_10830);
nand U11494 (N_11494,N_10692,N_10715);
or U11495 (N_11495,N_10858,N_10567);
nor U11496 (N_11496,N_10531,N_10598);
nand U11497 (N_11497,N_10851,N_10868);
nand U11498 (N_11498,N_10865,N_10650);
and U11499 (N_11499,N_10776,N_10898);
and U11500 (N_11500,N_11408,N_11322);
and U11501 (N_11501,N_11496,N_11034);
nor U11502 (N_11502,N_11354,N_11285);
nand U11503 (N_11503,N_11280,N_11314);
or U11504 (N_11504,N_11021,N_11129);
or U11505 (N_11505,N_11168,N_11458);
nand U11506 (N_11506,N_11371,N_11307);
xnor U11507 (N_11507,N_11015,N_11214);
and U11508 (N_11508,N_11238,N_11392);
nand U11509 (N_11509,N_11378,N_11036);
or U11510 (N_11510,N_11135,N_11389);
xnor U11511 (N_11511,N_11023,N_11001);
xor U11512 (N_11512,N_11289,N_11117);
nor U11513 (N_11513,N_11278,N_11063);
nand U11514 (N_11514,N_11412,N_11002);
nand U11515 (N_11515,N_11213,N_11096);
and U11516 (N_11516,N_11283,N_11252);
nand U11517 (N_11517,N_11288,N_11317);
nor U11518 (N_11518,N_11120,N_11026);
or U11519 (N_11519,N_11027,N_11234);
and U11520 (N_11520,N_11179,N_11123);
xor U11521 (N_11521,N_11480,N_11147);
nor U11522 (N_11522,N_11401,N_11483);
nand U11523 (N_11523,N_11399,N_11196);
or U11524 (N_11524,N_11164,N_11498);
or U11525 (N_11525,N_11300,N_11353);
or U11526 (N_11526,N_11381,N_11270);
or U11527 (N_11527,N_11070,N_11228);
nor U11528 (N_11528,N_11057,N_11390);
or U11529 (N_11529,N_11441,N_11106);
xnor U11530 (N_11530,N_11360,N_11165);
or U11531 (N_11531,N_11031,N_11160);
nand U11532 (N_11532,N_11019,N_11330);
or U11533 (N_11533,N_11052,N_11009);
nand U11534 (N_11534,N_11351,N_11373);
xnor U11535 (N_11535,N_11454,N_11246);
xor U11536 (N_11536,N_11258,N_11451);
or U11537 (N_11537,N_11124,N_11247);
xor U11538 (N_11538,N_11079,N_11460);
xnor U11539 (N_11539,N_11199,N_11302);
and U11540 (N_11540,N_11253,N_11215);
xor U11541 (N_11541,N_11207,N_11103);
nor U11542 (N_11542,N_11184,N_11490);
xnor U11543 (N_11543,N_11464,N_11411);
and U11544 (N_11544,N_11418,N_11339);
or U11545 (N_11545,N_11011,N_11427);
and U11546 (N_11546,N_11139,N_11175);
nor U11547 (N_11547,N_11433,N_11447);
xnor U11548 (N_11548,N_11173,N_11294);
nand U11549 (N_11549,N_11193,N_11054);
and U11550 (N_11550,N_11102,N_11166);
nand U11551 (N_11551,N_11405,N_11449);
xor U11552 (N_11552,N_11315,N_11035);
or U11553 (N_11553,N_11340,N_11384);
and U11554 (N_11554,N_11051,N_11479);
nand U11555 (N_11555,N_11276,N_11254);
and U11556 (N_11556,N_11167,N_11347);
nand U11557 (N_11557,N_11355,N_11066);
nand U11558 (N_11558,N_11010,N_11398);
xnor U11559 (N_11559,N_11180,N_11113);
nor U11560 (N_11560,N_11368,N_11251);
and U11561 (N_11561,N_11041,N_11383);
and U11562 (N_11562,N_11331,N_11342);
nand U11563 (N_11563,N_11499,N_11363);
or U11564 (N_11564,N_11150,N_11305);
or U11565 (N_11565,N_11438,N_11277);
and U11566 (N_11566,N_11260,N_11459);
nand U11567 (N_11567,N_11461,N_11329);
nor U11568 (N_11568,N_11341,N_11145);
xor U11569 (N_11569,N_11194,N_11221);
nand U11570 (N_11570,N_11003,N_11245);
and U11571 (N_11571,N_11092,N_11064);
or U11572 (N_11572,N_11171,N_11059);
xor U11573 (N_11573,N_11078,N_11348);
nand U11574 (N_11574,N_11039,N_11290);
and U11575 (N_11575,N_11308,N_11328);
xnor U11576 (N_11576,N_11430,N_11095);
xor U11577 (N_11577,N_11144,N_11127);
xor U11578 (N_11578,N_11379,N_11295);
xor U11579 (N_11579,N_11361,N_11432);
xor U11580 (N_11580,N_11022,N_11343);
xor U11581 (N_11581,N_11249,N_11088);
nor U11582 (N_11582,N_11481,N_11386);
xor U11583 (N_11583,N_11471,N_11143);
nand U11584 (N_11584,N_11200,N_11385);
nor U11585 (N_11585,N_11201,N_11191);
xor U11586 (N_11586,N_11197,N_11058);
and U11587 (N_11587,N_11219,N_11017);
nor U11588 (N_11588,N_11000,N_11446);
xnor U11589 (N_11589,N_11416,N_11190);
and U11590 (N_11590,N_11099,N_11350);
and U11591 (N_11591,N_11272,N_11257);
and U11592 (N_11592,N_11216,N_11138);
and U11593 (N_11593,N_11437,N_11131);
xor U11594 (N_11594,N_11151,N_11387);
or U11595 (N_11595,N_11268,N_11032);
nand U11596 (N_11596,N_11406,N_11267);
nor U11597 (N_11597,N_11377,N_11409);
nand U11598 (N_11598,N_11134,N_11085);
and U11599 (N_11599,N_11466,N_11309);
nand U11600 (N_11600,N_11467,N_11485);
nor U11601 (N_11601,N_11158,N_11489);
nand U11602 (N_11602,N_11203,N_11133);
or U11603 (N_11603,N_11273,N_11028);
xnor U11604 (N_11604,N_11357,N_11428);
nor U11605 (N_11605,N_11205,N_11156);
nor U11606 (N_11606,N_11029,N_11271);
nor U11607 (N_11607,N_11045,N_11025);
nor U11608 (N_11608,N_11419,N_11125);
nand U11609 (N_11609,N_11198,N_11185);
nand U11610 (N_11610,N_11421,N_11349);
nand U11611 (N_11611,N_11013,N_11475);
nand U11612 (N_11612,N_11209,N_11382);
or U11613 (N_11613,N_11006,N_11132);
nand U11614 (N_11614,N_11301,N_11231);
and U11615 (N_11615,N_11202,N_11274);
nor U11616 (N_11616,N_11286,N_11181);
and U11617 (N_11617,N_11468,N_11072);
xnor U11618 (N_11618,N_11242,N_11004);
nor U11619 (N_11619,N_11323,N_11100);
and U11620 (N_11620,N_11391,N_11204);
or U11621 (N_11621,N_11415,N_11093);
nor U11622 (N_11622,N_11239,N_11080);
and U11623 (N_11623,N_11312,N_11410);
nand U11624 (N_11624,N_11320,N_11044);
xor U11625 (N_11625,N_11452,N_11376);
xnor U11626 (N_11626,N_11413,N_11388);
and U11627 (N_11627,N_11208,N_11366);
nor U11628 (N_11628,N_11121,N_11014);
nor U11629 (N_11629,N_11488,N_11060);
xnor U11630 (N_11630,N_11367,N_11108);
or U11631 (N_11631,N_11334,N_11319);
or U11632 (N_11632,N_11352,N_11082);
and U11633 (N_11633,N_11287,N_11259);
or U11634 (N_11634,N_11243,N_11462);
nor U11635 (N_11635,N_11112,N_11395);
or U11636 (N_11636,N_11225,N_11358);
nand U11637 (N_11637,N_11050,N_11470);
or U11638 (N_11638,N_11291,N_11310);
nand U11639 (N_11639,N_11033,N_11443);
xnor U11640 (N_11640,N_11492,N_11071);
nand U11641 (N_11641,N_11299,N_11222);
or U11642 (N_11642,N_11473,N_11126);
nand U11643 (N_11643,N_11316,N_11226);
xnor U11644 (N_11644,N_11397,N_11332);
and U11645 (N_11645,N_11154,N_11296);
nor U11646 (N_11646,N_11115,N_11061);
nand U11647 (N_11647,N_11148,N_11486);
xnor U11648 (N_11648,N_11414,N_11012);
nand U11649 (N_11649,N_11256,N_11420);
nor U11650 (N_11650,N_11469,N_11396);
and U11651 (N_11651,N_11229,N_11403);
or U11652 (N_11652,N_11359,N_11210);
xnor U11653 (N_11653,N_11069,N_11345);
nand U11654 (N_11654,N_11176,N_11264);
and U11655 (N_11655,N_11338,N_11174);
and U11656 (N_11656,N_11476,N_11062);
and U11657 (N_11657,N_11495,N_11195);
and U11658 (N_11658,N_11116,N_11233);
nand U11659 (N_11659,N_11083,N_11105);
and U11660 (N_11660,N_11074,N_11370);
nor U11661 (N_11661,N_11232,N_11212);
nand U11662 (N_11662,N_11436,N_11261);
and U11663 (N_11663,N_11220,N_11374);
nand U11664 (N_11664,N_11068,N_11086);
and U11665 (N_11665,N_11162,N_11038);
xnor U11666 (N_11666,N_11056,N_11426);
or U11667 (N_11667,N_11043,N_11335);
nor U11668 (N_11668,N_11442,N_11110);
xor U11669 (N_11669,N_11404,N_11217);
nand U11670 (N_11670,N_11097,N_11472);
nor U11671 (N_11671,N_11337,N_11255);
nor U11672 (N_11672,N_11048,N_11107);
nor U11673 (N_11673,N_11393,N_11163);
and U11674 (N_11674,N_11444,N_11297);
and U11675 (N_11675,N_11047,N_11281);
xnor U11676 (N_11676,N_11077,N_11478);
nor U11677 (N_11677,N_11087,N_11450);
or U11678 (N_11678,N_11321,N_11445);
or U11679 (N_11679,N_11230,N_11439);
and U11680 (N_11680,N_11333,N_11474);
xor U11681 (N_11681,N_11188,N_11098);
and U11682 (N_11682,N_11081,N_11326);
or U11683 (N_11683,N_11407,N_11380);
or U11684 (N_11684,N_11109,N_11206);
nand U11685 (N_11685,N_11402,N_11153);
nand U11686 (N_11686,N_11269,N_11084);
nand U11687 (N_11687,N_11292,N_11020);
and U11688 (N_11688,N_11311,N_11037);
or U11689 (N_11689,N_11211,N_11152);
nor U11690 (N_11690,N_11130,N_11182);
nand U11691 (N_11691,N_11146,N_11170);
nand U11692 (N_11692,N_11227,N_11089);
xor U11693 (N_11693,N_11266,N_11075);
nor U11694 (N_11694,N_11298,N_11018);
nor U11695 (N_11695,N_11394,N_11055);
or U11696 (N_11696,N_11375,N_11073);
and U11697 (N_11697,N_11187,N_11453);
nor U11698 (N_11698,N_11094,N_11076);
and U11699 (N_11699,N_11046,N_11365);
and U11700 (N_11700,N_11159,N_11030);
nor U11701 (N_11701,N_11284,N_11024);
xor U11702 (N_11702,N_11128,N_11356);
nand U11703 (N_11703,N_11157,N_11429);
xor U11704 (N_11704,N_11183,N_11325);
nor U11705 (N_11705,N_11118,N_11065);
or U11706 (N_11706,N_11318,N_11434);
xnor U11707 (N_11707,N_11161,N_11040);
nand U11708 (N_11708,N_11275,N_11007);
nor U11709 (N_11709,N_11346,N_11484);
or U11710 (N_11710,N_11306,N_11431);
nand U11711 (N_11711,N_11090,N_11304);
nand U11712 (N_11712,N_11101,N_11440);
nand U11713 (N_11713,N_11293,N_11465);
nor U11714 (N_11714,N_11425,N_11424);
or U11715 (N_11715,N_11364,N_11423);
or U11716 (N_11716,N_11477,N_11303);
nor U11717 (N_11717,N_11049,N_11119);
nand U11718 (N_11718,N_11223,N_11111);
nand U11719 (N_11719,N_11177,N_11497);
nor U11720 (N_11720,N_11456,N_11487);
nor U11721 (N_11721,N_11178,N_11236);
nor U11722 (N_11722,N_11136,N_11493);
xor U11723 (N_11723,N_11448,N_11482);
xor U11724 (N_11724,N_11362,N_11224);
nand U11725 (N_11725,N_11248,N_11455);
or U11726 (N_11726,N_11091,N_11067);
or U11727 (N_11727,N_11140,N_11141);
nand U11728 (N_11728,N_11008,N_11491);
or U11729 (N_11729,N_11463,N_11189);
xnor U11730 (N_11730,N_11169,N_11457);
and U11731 (N_11731,N_11327,N_11324);
or U11732 (N_11732,N_11313,N_11282);
nor U11733 (N_11733,N_11053,N_11155);
or U11734 (N_11734,N_11172,N_11400);
and U11735 (N_11735,N_11137,N_11149);
nor U11736 (N_11736,N_11369,N_11235);
or U11737 (N_11737,N_11435,N_11005);
and U11738 (N_11738,N_11142,N_11422);
xnor U11739 (N_11739,N_11279,N_11417);
or U11740 (N_11740,N_11241,N_11237);
nor U11741 (N_11741,N_11240,N_11104);
xor U11742 (N_11742,N_11250,N_11336);
nand U11743 (N_11743,N_11016,N_11494);
xnor U11744 (N_11744,N_11344,N_11265);
xor U11745 (N_11745,N_11114,N_11372);
and U11746 (N_11746,N_11192,N_11218);
or U11747 (N_11747,N_11262,N_11042);
and U11748 (N_11748,N_11122,N_11263);
nor U11749 (N_11749,N_11186,N_11244);
and U11750 (N_11750,N_11066,N_11210);
and U11751 (N_11751,N_11028,N_11003);
nand U11752 (N_11752,N_11076,N_11064);
or U11753 (N_11753,N_11338,N_11323);
nor U11754 (N_11754,N_11177,N_11215);
and U11755 (N_11755,N_11201,N_11047);
and U11756 (N_11756,N_11176,N_11144);
nand U11757 (N_11757,N_11006,N_11274);
nor U11758 (N_11758,N_11346,N_11403);
nand U11759 (N_11759,N_11068,N_11452);
nand U11760 (N_11760,N_11489,N_11483);
and U11761 (N_11761,N_11089,N_11121);
nor U11762 (N_11762,N_11224,N_11459);
nand U11763 (N_11763,N_11471,N_11079);
xor U11764 (N_11764,N_11062,N_11350);
or U11765 (N_11765,N_11023,N_11257);
nor U11766 (N_11766,N_11152,N_11417);
and U11767 (N_11767,N_11134,N_11240);
nand U11768 (N_11768,N_11202,N_11172);
and U11769 (N_11769,N_11381,N_11398);
or U11770 (N_11770,N_11357,N_11236);
and U11771 (N_11771,N_11012,N_11370);
and U11772 (N_11772,N_11337,N_11257);
nand U11773 (N_11773,N_11329,N_11276);
and U11774 (N_11774,N_11424,N_11172);
xor U11775 (N_11775,N_11151,N_11159);
or U11776 (N_11776,N_11266,N_11130);
and U11777 (N_11777,N_11451,N_11482);
or U11778 (N_11778,N_11325,N_11413);
xor U11779 (N_11779,N_11024,N_11321);
xnor U11780 (N_11780,N_11102,N_11173);
or U11781 (N_11781,N_11240,N_11060);
nor U11782 (N_11782,N_11224,N_11372);
or U11783 (N_11783,N_11065,N_11080);
and U11784 (N_11784,N_11282,N_11396);
nor U11785 (N_11785,N_11388,N_11376);
xnor U11786 (N_11786,N_11115,N_11173);
nor U11787 (N_11787,N_11124,N_11112);
or U11788 (N_11788,N_11029,N_11212);
and U11789 (N_11789,N_11491,N_11043);
and U11790 (N_11790,N_11165,N_11470);
and U11791 (N_11791,N_11058,N_11212);
nand U11792 (N_11792,N_11316,N_11492);
or U11793 (N_11793,N_11061,N_11025);
xor U11794 (N_11794,N_11028,N_11123);
nand U11795 (N_11795,N_11130,N_11078);
xnor U11796 (N_11796,N_11168,N_11182);
nor U11797 (N_11797,N_11212,N_11272);
xor U11798 (N_11798,N_11375,N_11055);
nor U11799 (N_11799,N_11411,N_11320);
xor U11800 (N_11800,N_11419,N_11438);
or U11801 (N_11801,N_11482,N_11221);
xnor U11802 (N_11802,N_11152,N_11139);
xnor U11803 (N_11803,N_11290,N_11226);
or U11804 (N_11804,N_11340,N_11126);
or U11805 (N_11805,N_11428,N_11192);
or U11806 (N_11806,N_11489,N_11299);
nand U11807 (N_11807,N_11379,N_11436);
xnor U11808 (N_11808,N_11336,N_11042);
nor U11809 (N_11809,N_11420,N_11250);
xor U11810 (N_11810,N_11339,N_11136);
nor U11811 (N_11811,N_11320,N_11151);
nor U11812 (N_11812,N_11041,N_11057);
nand U11813 (N_11813,N_11259,N_11319);
or U11814 (N_11814,N_11071,N_11161);
nand U11815 (N_11815,N_11404,N_11464);
nor U11816 (N_11816,N_11298,N_11394);
and U11817 (N_11817,N_11236,N_11473);
xnor U11818 (N_11818,N_11231,N_11361);
or U11819 (N_11819,N_11037,N_11158);
nand U11820 (N_11820,N_11011,N_11444);
and U11821 (N_11821,N_11306,N_11396);
and U11822 (N_11822,N_11483,N_11097);
and U11823 (N_11823,N_11276,N_11312);
nor U11824 (N_11824,N_11077,N_11393);
nor U11825 (N_11825,N_11129,N_11304);
nor U11826 (N_11826,N_11271,N_11005);
and U11827 (N_11827,N_11149,N_11134);
or U11828 (N_11828,N_11417,N_11048);
xnor U11829 (N_11829,N_11118,N_11359);
nand U11830 (N_11830,N_11074,N_11042);
xor U11831 (N_11831,N_11129,N_11015);
xnor U11832 (N_11832,N_11323,N_11397);
and U11833 (N_11833,N_11163,N_11287);
nand U11834 (N_11834,N_11039,N_11013);
xnor U11835 (N_11835,N_11233,N_11455);
or U11836 (N_11836,N_11024,N_11407);
and U11837 (N_11837,N_11048,N_11206);
and U11838 (N_11838,N_11248,N_11394);
nor U11839 (N_11839,N_11246,N_11257);
or U11840 (N_11840,N_11089,N_11079);
nor U11841 (N_11841,N_11158,N_11287);
xnor U11842 (N_11842,N_11147,N_11078);
nor U11843 (N_11843,N_11397,N_11092);
nor U11844 (N_11844,N_11089,N_11195);
nand U11845 (N_11845,N_11041,N_11253);
nor U11846 (N_11846,N_11023,N_11116);
or U11847 (N_11847,N_11287,N_11171);
or U11848 (N_11848,N_11124,N_11238);
nor U11849 (N_11849,N_11375,N_11230);
and U11850 (N_11850,N_11283,N_11074);
nand U11851 (N_11851,N_11388,N_11328);
nand U11852 (N_11852,N_11364,N_11324);
nand U11853 (N_11853,N_11325,N_11232);
xor U11854 (N_11854,N_11232,N_11143);
and U11855 (N_11855,N_11057,N_11248);
nor U11856 (N_11856,N_11461,N_11438);
and U11857 (N_11857,N_11347,N_11262);
nor U11858 (N_11858,N_11091,N_11309);
nor U11859 (N_11859,N_11136,N_11041);
xnor U11860 (N_11860,N_11454,N_11416);
and U11861 (N_11861,N_11464,N_11107);
or U11862 (N_11862,N_11068,N_11419);
nand U11863 (N_11863,N_11393,N_11434);
nand U11864 (N_11864,N_11455,N_11019);
or U11865 (N_11865,N_11091,N_11464);
nand U11866 (N_11866,N_11171,N_11322);
or U11867 (N_11867,N_11205,N_11385);
nor U11868 (N_11868,N_11034,N_11051);
nand U11869 (N_11869,N_11158,N_11141);
or U11870 (N_11870,N_11399,N_11336);
or U11871 (N_11871,N_11378,N_11090);
or U11872 (N_11872,N_11017,N_11476);
and U11873 (N_11873,N_11423,N_11080);
nand U11874 (N_11874,N_11016,N_11258);
or U11875 (N_11875,N_11197,N_11300);
xnor U11876 (N_11876,N_11361,N_11060);
xnor U11877 (N_11877,N_11355,N_11015);
or U11878 (N_11878,N_11092,N_11200);
xnor U11879 (N_11879,N_11157,N_11364);
nand U11880 (N_11880,N_11299,N_11074);
xnor U11881 (N_11881,N_11082,N_11175);
or U11882 (N_11882,N_11264,N_11111);
and U11883 (N_11883,N_11489,N_11400);
nand U11884 (N_11884,N_11431,N_11459);
xnor U11885 (N_11885,N_11046,N_11106);
or U11886 (N_11886,N_11205,N_11118);
nand U11887 (N_11887,N_11354,N_11235);
and U11888 (N_11888,N_11499,N_11315);
nor U11889 (N_11889,N_11313,N_11070);
and U11890 (N_11890,N_11252,N_11399);
xnor U11891 (N_11891,N_11047,N_11175);
and U11892 (N_11892,N_11284,N_11351);
nor U11893 (N_11893,N_11388,N_11457);
and U11894 (N_11894,N_11032,N_11031);
nand U11895 (N_11895,N_11435,N_11378);
and U11896 (N_11896,N_11179,N_11453);
and U11897 (N_11897,N_11465,N_11125);
nor U11898 (N_11898,N_11145,N_11357);
nor U11899 (N_11899,N_11454,N_11448);
or U11900 (N_11900,N_11317,N_11491);
and U11901 (N_11901,N_11411,N_11101);
nand U11902 (N_11902,N_11119,N_11333);
and U11903 (N_11903,N_11463,N_11236);
xor U11904 (N_11904,N_11477,N_11387);
or U11905 (N_11905,N_11330,N_11195);
xor U11906 (N_11906,N_11228,N_11142);
nor U11907 (N_11907,N_11149,N_11361);
xor U11908 (N_11908,N_11485,N_11072);
nand U11909 (N_11909,N_11227,N_11405);
and U11910 (N_11910,N_11286,N_11299);
nor U11911 (N_11911,N_11049,N_11363);
or U11912 (N_11912,N_11157,N_11218);
and U11913 (N_11913,N_11172,N_11017);
and U11914 (N_11914,N_11126,N_11341);
nand U11915 (N_11915,N_11054,N_11128);
nor U11916 (N_11916,N_11286,N_11472);
and U11917 (N_11917,N_11360,N_11080);
nand U11918 (N_11918,N_11125,N_11113);
nand U11919 (N_11919,N_11376,N_11422);
xnor U11920 (N_11920,N_11108,N_11498);
nor U11921 (N_11921,N_11398,N_11178);
nor U11922 (N_11922,N_11222,N_11436);
nand U11923 (N_11923,N_11475,N_11313);
xnor U11924 (N_11924,N_11486,N_11048);
nand U11925 (N_11925,N_11010,N_11458);
nor U11926 (N_11926,N_11042,N_11309);
nand U11927 (N_11927,N_11395,N_11203);
or U11928 (N_11928,N_11480,N_11441);
nand U11929 (N_11929,N_11218,N_11360);
xnor U11930 (N_11930,N_11324,N_11232);
nand U11931 (N_11931,N_11285,N_11001);
nor U11932 (N_11932,N_11311,N_11348);
and U11933 (N_11933,N_11414,N_11486);
or U11934 (N_11934,N_11160,N_11201);
nand U11935 (N_11935,N_11295,N_11444);
nor U11936 (N_11936,N_11436,N_11423);
and U11937 (N_11937,N_11113,N_11332);
nand U11938 (N_11938,N_11485,N_11000);
or U11939 (N_11939,N_11121,N_11274);
xor U11940 (N_11940,N_11042,N_11207);
nand U11941 (N_11941,N_11196,N_11138);
or U11942 (N_11942,N_11470,N_11281);
and U11943 (N_11943,N_11207,N_11131);
xor U11944 (N_11944,N_11221,N_11392);
and U11945 (N_11945,N_11286,N_11255);
and U11946 (N_11946,N_11156,N_11413);
and U11947 (N_11947,N_11222,N_11381);
and U11948 (N_11948,N_11197,N_11117);
and U11949 (N_11949,N_11294,N_11407);
nand U11950 (N_11950,N_11245,N_11351);
and U11951 (N_11951,N_11184,N_11325);
nor U11952 (N_11952,N_11092,N_11193);
or U11953 (N_11953,N_11197,N_11383);
or U11954 (N_11954,N_11013,N_11470);
xor U11955 (N_11955,N_11305,N_11274);
and U11956 (N_11956,N_11378,N_11328);
xnor U11957 (N_11957,N_11304,N_11097);
xor U11958 (N_11958,N_11113,N_11419);
nand U11959 (N_11959,N_11472,N_11101);
nand U11960 (N_11960,N_11437,N_11353);
or U11961 (N_11961,N_11064,N_11140);
or U11962 (N_11962,N_11312,N_11114);
nand U11963 (N_11963,N_11247,N_11117);
xor U11964 (N_11964,N_11290,N_11050);
nor U11965 (N_11965,N_11350,N_11408);
and U11966 (N_11966,N_11118,N_11104);
xor U11967 (N_11967,N_11479,N_11141);
xor U11968 (N_11968,N_11445,N_11369);
nor U11969 (N_11969,N_11321,N_11230);
and U11970 (N_11970,N_11150,N_11324);
or U11971 (N_11971,N_11092,N_11390);
and U11972 (N_11972,N_11275,N_11418);
nor U11973 (N_11973,N_11404,N_11191);
or U11974 (N_11974,N_11451,N_11325);
nor U11975 (N_11975,N_11146,N_11364);
nor U11976 (N_11976,N_11053,N_11233);
or U11977 (N_11977,N_11411,N_11375);
or U11978 (N_11978,N_11155,N_11224);
nand U11979 (N_11979,N_11495,N_11258);
xnor U11980 (N_11980,N_11081,N_11242);
xor U11981 (N_11981,N_11032,N_11301);
or U11982 (N_11982,N_11302,N_11241);
and U11983 (N_11983,N_11272,N_11274);
or U11984 (N_11984,N_11048,N_11146);
and U11985 (N_11985,N_11204,N_11147);
nand U11986 (N_11986,N_11366,N_11459);
nor U11987 (N_11987,N_11261,N_11294);
nor U11988 (N_11988,N_11289,N_11025);
xnor U11989 (N_11989,N_11089,N_11366);
nor U11990 (N_11990,N_11054,N_11320);
nor U11991 (N_11991,N_11019,N_11300);
nor U11992 (N_11992,N_11422,N_11479);
or U11993 (N_11993,N_11107,N_11262);
and U11994 (N_11994,N_11225,N_11325);
nor U11995 (N_11995,N_11213,N_11252);
or U11996 (N_11996,N_11499,N_11488);
nor U11997 (N_11997,N_11049,N_11071);
nand U11998 (N_11998,N_11050,N_11077);
and U11999 (N_11999,N_11177,N_11241);
and U12000 (N_12000,N_11997,N_11644);
xor U12001 (N_12001,N_11990,N_11963);
and U12002 (N_12002,N_11941,N_11846);
xor U12003 (N_12003,N_11934,N_11769);
nand U12004 (N_12004,N_11547,N_11514);
or U12005 (N_12005,N_11950,N_11542);
or U12006 (N_12006,N_11745,N_11894);
or U12007 (N_12007,N_11903,N_11961);
nand U12008 (N_12008,N_11541,N_11840);
or U12009 (N_12009,N_11975,N_11838);
and U12010 (N_12010,N_11749,N_11931);
xor U12011 (N_12011,N_11982,N_11864);
nand U12012 (N_12012,N_11517,N_11955);
xor U12013 (N_12013,N_11669,N_11591);
or U12014 (N_12014,N_11713,N_11582);
and U12015 (N_12015,N_11536,N_11815);
nand U12016 (N_12016,N_11897,N_11549);
and U12017 (N_12017,N_11730,N_11970);
xor U12018 (N_12018,N_11759,N_11562);
or U12019 (N_12019,N_11622,N_11831);
nor U12020 (N_12020,N_11988,N_11723);
nand U12021 (N_12021,N_11510,N_11910);
xor U12022 (N_12022,N_11810,N_11889);
or U12023 (N_12023,N_11584,N_11866);
or U12024 (N_12024,N_11893,N_11556);
xor U12025 (N_12025,N_11671,N_11594);
xor U12026 (N_12026,N_11835,N_11758);
nor U12027 (N_12027,N_11693,N_11719);
nor U12028 (N_12028,N_11887,N_11827);
or U12029 (N_12029,N_11919,N_11617);
xor U12030 (N_12030,N_11691,N_11874);
or U12031 (N_12031,N_11848,N_11552);
xnor U12032 (N_12032,N_11626,N_11881);
or U12033 (N_12033,N_11969,N_11611);
nand U12034 (N_12034,N_11511,N_11711);
or U12035 (N_12035,N_11906,N_11638);
nand U12036 (N_12036,N_11686,N_11861);
and U12037 (N_12037,N_11725,N_11603);
xnor U12038 (N_12038,N_11625,N_11872);
and U12039 (N_12039,N_11663,N_11800);
or U12040 (N_12040,N_11976,N_11994);
and U12041 (N_12041,N_11731,N_11890);
xor U12042 (N_12042,N_11736,N_11916);
xor U12043 (N_12043,N_11520,N_11544);
nand U12044 (N_12044,N_11804,N_11847);
nand U12045 (N_12045,N_11540,N_11981);
and U12046 (N_12046,N_11998,N_11940);
or U12047 (N_12047,N_11704,N_11643);
nand U12048 (N_12048,N_11798,N_11937);
nand U12049 (N_12049,N_11606,N_11968);
nand U12050 (N_12050,N_11949,N_11886);
nor U12051 (N_12051,N_11646,N_11645);
or U12052 (N_12052,N_11647,N_11882);
xnor U12053 (N_12053,N_11590,N_11634);
and U12054 (N_12054,N_11561,N_11688);
nand U12055 (N_12055,N_11913,N_11853);
or U12056 (N_12056,N_11935,N_11554);
or U12057 (N_12057,N_11533,N_11574);
nand U12058 (N_12058,N_11777,N_11608);
nor U12059 (N_12059,N_11926,N_11885);
nor U12060 (N_12060,N_11539,N_11709);
nor U12061 (N_12061,N_11966,N_11991);
and U12062 (N_12062,N_11813,N_11604);
or U12063 (N_12063,N_11525,N_11986);
nand U12064 (N_12064,N_11631,N_11766);
xnor U12065 (N_12065,N_11965,N_11971);
and U12066 (N_12066,N_11828,N_11860);
and U12067 (N_12067,N_11649,N_11555);
nand U12068 (N_12068,N_11805,N_11901);
nand U12069 (N_12069,N_11871,N_11942);
nor U12070 (N_12070,N_11844,N_11746);
xor U12071 (N_12071,N_11548,N_11714);
and U12072 (N_12072,N_11795,N_11773);
or U12073 (N_12073,N_11858,N_11535);
nor U12074 (N_12074,N_11879,N_11782);
and U12075 (N_12075,N_11505,N_11789);
xor U12076 (N_12076,N_11595,N_11863);
nor U12077 (N_12077,N_11924,N_11953);
or U12078 (N_12078,N_11569,N_11902);
or U12079 (N_12079,N_11697,N_11735);
and U12080 (N_12080,N_11642,N_11748);
and U12081 (N_12081,N_11531,N_11873);
xor U12082 (N_12082,N_11637,N_11618);
or U12083 (N_12083,N_11756,N_11527);
nor U12084 (N_12084,N_11808,N_11980);
and U12085 (N_12085,N_11785,N_11564);
and U12086 (N_12086,N_11502,N_11772);
and U12087 (N_12087,N_11571,N_11673);
xnor U12088 (N_12088,N_11705,N_11509);
nor U12089 (N_12089,N_11712,N_11557);
and U12090 (N_12090,N_11972,N_11764);
nor U12091 (N_12091,N_11678,N_11674);
nor U12092 (N_12092,N_11951,N_11737);
nor U12093 (N_12093,N_11726,N_11918);
xor U12094 (N_12094,N_11899,N_11884);
nand U12095 (N_12095,N_11654,N_11753);
xnor U12096 (N_12096,N_11812,N_11996);
and U12097 (N_12097,N_11932,N_11927);
nand U12098 (N_12098,N_11818,N_11834);
and U12099 (N_12099,N_11706,N_11661);
nor U12100 (N_12100,N_11743,N_11898);
nand U12101 (N_12101,N_11629,N_11823);
nand U12102 (N_12102,N_11911,N_11985);
and U12103 (N_12103,N_11515,N_11601);
and U12104 (N_12104,N_11778,N_11679);
xor U12105 (N_12105,N_11630,N_11639);
and U12106 (N_12106,N_11776,N_11685);
xor U12107 (N_12107,N_11522,N_11702);
nor U12108 (N_12108,N_11904,N_11716);
xor U12109 (N_12109,N_11666,N_11754);
nor U12110 (N_12110,N_11786,N_11665);
xnor U12111 (N_12111,N_11944,N_11814);
nor U12112 (N_12112,N_11765,N_11851);
and U12113 (N_12113,N_11974,N_11788);
xor U12114 (N_12114,N_11938,N_11751);
nor U12115 (N_12115,N_11526,N_11843);
nand U12116 (N_12116,N_11842,N_11816);
nor U12117 (N_12117,N_11558,N_11833);
and U12118 (N_12118,N_11640,N_11537);
or U12119 (N_12119,N_11727,N_11523);
nor U12120 (N_12120,N_11599,N_11581);
nand U12121 (N_12121,N_11662,N_11891);
nand U12122 (N_12122,N_11930,N_11849);
and U12123 (N_12123,N_11605,N_11774);
xnor U12124 (N_12124,N_11832,N_11578);
nand U12125 (N_12125,N_11580,N_11614);
nor U12126 (N_12126,N_11803,N_11781);
or U12127 (N_12127,N_11920,N_11793);
nand U12128 (N_12128,N_11621,N_11682);
and U12129 (N_12129,N_11690,N_11952);
nand U12130 (N_12130,N_11587,N_11729);
and U12131 (N_12131,N_11780,N_11825);
xnor U12132 (N_12132,N_11947,N_11612);
nand U12133 (N_12133,N_11545,N_11633);
nand U12134 (N_12134,N_11912,N_11768);
and U12135 (N_12135,N_11909,N_11850);
and U12136 (N_12136,N_11992,N_11512);
nand U12137 (N_12137,N_11984,N_11876);
and U12138 (N_12138,N_11597,N_11859);
or U12139 (N_12139,N_11794,N_11914);
or U12140 (N_12140,N_11720,N_11946);
nand U12141 (N_12141,N_11747,N_11752);
nand U12142 (N_12142,N_11967,N_11869);
or U12143 (N_12143,N_11917,N_11960);
or U12144 (N_12144,N_11762,N_11892);
nand U12145 (N_12145,N_11895,N_11676);
xnor U12146 (N_12146,N_11733,N_11770);
or U12147 (N_12147,N_11610,N_11822);
xnor U12148 (N_12148,N_11824,N_11734);
or U12149 (N_12149,N_11579,N_11732);
nor U12150 (N_12150,N_11623,N_11632);
xor U12151 (N_12151,N_11880,N_11757);
nand U12152 (N_12152,N_11503,N_11560);
and U12153 (N_12153,N_11703,N_11698);
or U12154 (N_12154,N_11677,N_11896);
and U12155 (N_12155,N_11551,N_11915);
nand U12156 (N_12156,N_11925,N_11799);
nor U12157 (N_12157,N_11738,N_11576);
and U12158 (N_12158,N_11664,N_11907);
nand U12159 (N_12159,N_11783,N_11829);
or U12160 (N_12160,N_11583,N_11839);
nor U12161 (N_12161,N_11928,N_11741);
xnor U12162 (N_12162,N_11806,N_11636);
nand U12163 (N_12163,N_11979,N_11763);
and U12164 (N_12164,N_11855,N_11641);
or U12165 (N_12165,N_11628,N_11694);
or U12166 (N_12166,N_11856,N_11857);
or U12167 (N_12167,N_11607,N_11801);
or U12168 (N_12168,N_11989,N_11532);
nand U12169 (N_12169,N_11648,N_11696);
and U12170 (N_12170,N_11667,N_11900);
or U12171 (N_12171,N_11627,N_11521);
and U12172 (N_12172,N_11883,N_11593);
and U12173 (N_12173,N_11775,N_11784);
nand U12174 (N_12174,N_11715,N_11945);
xor U12175 (N_12175,N_11513,N_11739);
or U12176 (N_12176,N_11655,N_11750);
and U12177 (N_12177,N_11659,N_11820);
nand U12178 (N_12178,N_11566,N_11797);
nor U12179 (N_12179,N_11596,N_11936);
nor U12180 (N_12180,N_11506,N_11699);
nand U12181 (N_12181,N_11660,N_11650);
nand U12182 (N_12182,N_11819,N_11787);
nand U12183 (N_12183,N_11613,N_11616);
xnor U12184 (N_12184,N_11836,N_11958);
nand U12185 (N_12185,N_11534,N_11957);
nand U12186 (N_12186,N_11658,N_11933);
or U12187 (N_12187,N_11519,N_11609);
xnor U12188 (N_12188,N_11575,N_11852);
or U12189 (N_12189,N_11742,N_11817);
or U12190 (N_12190,N_11837,N_11572);
xor U12191 (N_12191,N_11538,N_11672);
xor U12192 (N_12192,N_11589,N_11959);
and U12193 (N_12193,N_11995,N_11518);
nor U12194 (N_12194,N_11954,N_11588);
or U12195 (N_12195,N_11692,N_11707);
nand U12196 (N_12196,N_11543,N_11761);
nor U12197 (N_12197,N_11948,N_11718);
nand U12198 (N_12198,N_11867,N_11500);
nor U12199 (N_12199,N_11722,N_11568);
and U12200 (N_12200,N_11598,N_11570);
and U12201 (N_12201,N_11675,N_11683);
or U12202 (N_12202,N_11651,N_11983);
or U12203 (N_12203,N_11508,N_11550);
nand U12204 (N_12204,N_11653,N_11792);
or U12205 (N_12205,N_11977,N_11865);
nand U12206 (N_12206,N_11740,N_11721);
nor U12207 (N_12207,N_11921,N_11565);
nand U12208 (N_12208,N_11767,N_11755);
and U12209 (N_12209,N_11962,N_11668);
xor U12210 (N_12210,N_11602,N_11524);
or U12211 (N_12211,N_11529,N_11504);
nor U12212 (N_12212,N_11680,N_11585);
xnor U12213 (N_12213,N_11875,N_11956);
xnor U12214 (N_12214,N_11717,N_11701);
or U12215 (N_12215,N_11790,N_11929);
xnor U12216 (N_12216,N_11615,N_11624);
xnor U12217 (N_12217,N_11681,N_11695);
or U12218 (N_12218,N_11744,N_11826);
nand U12219 (N_12219,N_11973,N_11687);
nand U12220 (N_12220,N_11563,N_11652);
nor U12221 (N_12221,N_11700,N_11845);
or U12222 (N_12222,N_11501,N_11710);
or U12223 (N_12223,N_11868,N_11619);
and U12224 (N_12224,N_11978,N_11943);
nand U12225 (N_12225,N_11516,N_11553);
or U12226 (N_12226,N_11656,N_11796);
nor U12227 (N_12227,N_11530,N_11728);
nand U12228 (N_12228,N_11600,N_11807);
nand U12229 (N_12229,N_11507,N_11993);
xnor U12230 (N_12230,N_11771,N_11546);
and U12231 (N_12231,N_11791,N_11586);
nor U12232 (N_12232,N_11878,N_11760);
and U12233 (N_12233,N_11573,N_11841);
nor U12234 (N_12234,N_11999,N_11559);
and U12235 (N_12235,N_11802,N_11908);
nand U12236 (N_12236,N_11635,N_11854);
nand U12237 (N_12237,N_11888,N_11657);
or U12238 (N_12238,N_11684,N_11670);
nor U12239 (N_12239,N_11964,N_11779);
nand U12240 (N_12240,N_11870,N_11724);
nand U12241 (N_12241,N_11987,N_11862);
or U12242 (N_12242,N_11830,N_11567);
nor U12243 (N_12243,N_11905,N_11592);
or U12244 (N_12244,N_11922,N_11923);
nand U12245 (N_12245,N_11708,N_11620);
nor U12246 (N_12246,N_11877,N_11689);
and U12247 (N_12247,N_11809,N_11821);
nand U12248 (N_12248,N_11528,N_11939);
and U12249 (N_12249,N_11811,N_11577);
nor U12250 (N_12250,N_11546,N_11809);
nor U12251 (N_12251,N_11500,N_11761);
or U12252 (N_12252,N_11751,N_11816);
nor U12253 (N_12253,N_11554,N_11780);
xor U12254 (N_12254,N_11802,N_11512);
xnor U12255 (N_12255,N_11804,N_11748);
or U12256 (N_12256,N_11701,N_11531);
nand U12257 (N_12257,N_11613,N_11721);
nand U12258 (N_12258,N_11799,N_11754);
nor U12259 (N_12259,N_11886,N_11903);
nor U12260 (N_12260,N_11880,N_11748);
and U12261 (N_12261,N_11701,N_11605);
nand U12262 (N_12262,N_11714,N_11725);
nor U12263 (N_12263,N_11800,N_11649);
nand U12264 (N_12264,N_11692,N_11838);
or U12265 (N_12265,N_11636,N_11591);
nor U12266 (N_12266,N_11942,N_11681);
and U12267 (N_12267,N_11999,N_11736);
xnor U12268 (N_12268,N_11526,N_11978);
nor U12269 (N_12269,N_11708,N_11686);
and U12270 (N_12270,N_11761,N_11726);
or U12271 (N_12271,N_11995,N_11746);
or U12272 (N_12272,N_11708,N_11678);
xnor U12273 (N_12273,N_11711,N_11926);
nor U12274 (N_12274,N_11861,N_11851);
or U12275 (N_12275,N_11503,N_11713);
nor U12276 (N_12276,N_11605,N_11720);
xor U12277 (N_12277,N_11743,N_11729);
and U12278 (N_12278,N_11694,N_11978);
and U12279 (N_12279,N_11676,N_11712);
xor U12280 (N_12280,N_11857,N_11833);
nor U12281 (N_12281,N_11941,N_11849);
xor U12282 (N_12282,N_11826,N_11967);
and U12283 (N_12283,N_11863,N_11914);
xor U12284 (N_12284,N_11965,N_11601);
nor U12285 (N_12285,N_11541,N_11926);
nor U12286 (N_12286,N_11894,N_11701);
or U12287 (N_12287,N_11542,N_11836);
and U12288 (N_12288,N_11640,N_11550);
and U12289 (N_12289,N_11591,N_11951);
xor U12290 (N_12290,N_11653,N_11634);
xor U12291 (N_12291,N_11802,N_11928);
or U12292 (N_12292,N_11796,N_11615);
nand U12293 (N_12293,N_11557,N_11788);
and U12294 (N_12294,N_11746,N_11617);
xnor U12295 (N_12295,N_11890,N_11696);
nand U12296 (N_12296,N_11814,N_11870);
xor U12297 (N_12297,N_11592,N_11658);
and U12298 (N_12298,N_11828,N_11976);
or U12299 (N_12299,N_11570,N_11959);
nor U12300 (N_12300,N_11778,N_11518);
nand U12301 (N_12301,N_11742,N_11950);
and U12302 (N_12302,N_11502,N_11643);
nand U12303 (N_12303,N_11864,N_11813);
or U12304 (N_12304,N_11816,N_11664);
or U12305 (N_12305,N_11594,N_11793);
nor U12306 (N_12306,N_11660,N_11802);
nand U12307 (N_12307,N_11519,N_11542);
or U12308 (N_12308,N_11954,N_11668);
nor U12309 (N_12309,N_11926,N_11538);
nand U12310 (N_12310,N_11706,N_11827);
nand U12311 (N_12311,N_11581,N_11741);
and U12312 (N_12312,N_11724,N_11921);
xnor U12313 (N_12313,N_11698,N_11682);
nor U12314 (N_12314,N_11930,N_11728);
xnor U12315 (N_12315,N_11962,N_11867);
nor U12316 (N_12316,N_11790,N_11827);
or U12317 (N_12317,N_11972,N_11963);
nand U12318 (N_12318,N_11993,N_11900);
or U12319 (N_12319,N_11610,N_11661);
or U12320 (N_12320,N_11658,N_11680);
nand U12321 (N_12321,N_11989,N_11829);
xor U12322 (N_12322,N_11718,N_11821);
nand U12323 (N_12323,N_11834,N_11524);
and U12324 (N_12324,N_11786,N_11658);
or U12325 (N_12325,N_11852,N_11628);
nor U12326 (N_12326,N_11561,N_11885);
xnor U12327 (N_12327,N_11655,N_11803);
nor U12328 (N_12328,N_11831,N_11507);
nor U12329 (N_12329,N_11572,N_11963);
xnor U12330 (N_12330,N_11854,N_11614);
nor U12331 (N_12331,N_11643,N_11532);
nor U12332 (N_12332,N_11990,N_11953);
xor U12333 (N_12333,N_11728,N_11803);
nand U12334 (N_12334,N_11953,N_11850);
nand U12335 (N_12335,N_11737,N_11939);
or U12336 (N_12336,N_11509,N_11881);
or U12337 (N_12337,N_11745,N_11597);
nand U12338 (N_12338,N_11755,N_11510);
or U12339 (N_12339,N_11705,N_11961);
and U12340 (N_12340,N_11719,N_11786);
or U12341 (N_12341,N_11576,N_11605);
and U12342 (N_12342,N_11675,N_11705);
and U12343 (N_12343,N_11930,N_11878);
and U12344 (N_12344,N_11870,N_11957);
nand U12345 (N_12345,N_11840,N_11524);
or U12346 (N_12346,N_11944,N_11882);
nand U12347 (N_12347,N_11931,N_11972);
and U12348 (N_12348,N_11741,N_11582);
nand U12349 (N_12349,N_11738,N_11681);
or U12350 (N_12350,N_11723,N_11666);
nor U12351 (N_12351,N_11874,N_11985);
nor U12352 (N_12352,N_11914,N_11658);
xnor U12353 (N_12353,N_11538,N_11569);
or U12354 (N_12354,N_11863,N_11861);
or U12355 (N_12355,N_11970,N_11500);
and U12356 (N_12356,N_11893,N_11658);
nor U12357 (N_12357,N_11693,N_11694);
nor U12358 (N_12358,N_11912,N_11818);
xor U12359 (N_12359,N_11579,N_11651);
xor U12360 (N_12360,N_11911,N_11830);
and U12361 (N_12361,N_11753,N_11812);
nor U12362 (N_12362,N_11723,N_11641);
and U12363 (N_12363,N_11806,N_11768);
nand U12364 (N_12364,N_11850,N_11903);
nand U12365 (N_12365,N_11826,N_11626);
xnor U12366 (N_12366,N_11540,N_11977);
nor U12367 (N_12367,N_11830,N_11845);
or U12368 (N_12368,N_11536,N_11704);
nor U12369 (N_12369,N_11640,N_11960);
and U12370 (N_12370,N_11662,N_11966);
xor U12371 (N_12371,N_11824,N_11543);
nor U12372 (N_12372,N_11995,N_11915);
nor U12373 (N_12373,N_11501,N_11968);
or U12374 (N_12374,N_11987,N_11808);
or U12375 (N_12375,N_11907,N_11565);
xnor U12376 (N_12376,N_11671,N_11740);
nand U12377 (N_12377,N_11772,N_11967);
nand U12378 (N_12378,N_11664,N_11580);
xor U12379 (N_12379,N_11551,N_11577);
or U12380 (N_12380,N_11500,N_11617);
nand U12381 (N_12381,N_11638,N_11616);
nand U12382 (N_12382,N_11516,N_11845);
nor U12383 (N_12383,N_11518,N_11768);
nand U12384 (N_12384,N_11975,N_11718);
nand U12385 (N_12385,N_11520,N_11730);
or U12386 (N_12386,N_11933,N_11887);
nor U12387 (N_12387,N_11932,N_11930);
and U12388 (N_12388,N_11964,N_11688);
or U12389 (N_12389,N_11644,N_11542);
nor U12390 (N_12390,N_11745,N_11828);
nor U12391 (N_12391,N_11504,N_11707);
or U12392 (N_12392,N_11767,N_11632);
xor U12393 (N_12393,N_11955,N_11606);
and U12394 (N_12394,N_11552,N_11943);
or U12395 (N_12395,N_11852,N_11826);
xor U12396 (N_12396,N_11824,N_11572);
or U12397 (N_12397,N_11612,N_11708);
nor U12398 (N_12398,N_11978,N_11649);
xor U12399 (N_12399,N_11847,N_11527);
nand U12400 (N_12400,N_11976,N_11829);
nor U12401 (N_12401,N_11641,N_11512);
and U12402 (N_12402,N_11677,N_11627);
or U12403 (N_12403,N_11602,N_11585);
xor U12404 (N_12404,N_11786,N_11664);
and U12405 (N_12405,N_11874,N_11976);
nor U12406 (N_12406,N_11883,N_11527);
nor U12407 (N_12407,N_11861,N_11621);
or U12408 (N_12408,N_11570,N_11848);
xor U12409 (N_12409,N_11556,N_11942);
and U12410 (N_12410,N_11632,N_11750);
xnor U12411 (N_12411,N_11528,N_11889);
and U12412 (N_12412,N_11517,N_11543);
xnor U12413 (N_12413,N_11637,N_11586);
or U12414 (N_12414,N_11932,N_11670);
nor U12415 (N_12415,N_11703,N_11511);
xnor U12416 (N_12416,N_11631,N_11907);
or U12417 (N_12417,N_11769,N_11612);
nor U12418 (N_12418,N_11593,N_11643);
and U12419 (N_12419,N_11930,N_11974);
nor U12420 (N_12420,N_11672,N_11995);
and U12421 (N_12421,N_11904,N_11985);
and U12422 (N_12422,N_11732,N_11934);
and U12423 (N_12423,N_11683,N_11863);
and U12424 (N_12424,N_11721,N_11811);
and U12425 (N_12425,N_11937,N_11644);
or U12426 (N_12426,N_11934,N_11658);
xor U12427 (N_12427,N_11909,N_11937);
or U12428 (N_12428,N_11503,N_11869);
and U12429 (N_12429,N_11706,N_11649);
nand U12430 (N_12430,N_11948,N_11850);
nand U12431 (N_12431,N_11781,N_11742);
xor U12432 (N_12432,N_11853,N_11796);
xor U12433 (N_12433,N_11611,N_11749);
nor U12434 (N_12434,N_11784,N_11560);
or U12435 (N_12435,N_11549,N_11691);
xnor U12436 (N_12436,N_11734,N_11986);
or U12437 (N_12437,N_11716,N_11760);
and U12438 (N_12438,N_11523,N_11953);
and U12439 (N_12439,N_11765,N_11516);
or U12440 (N_12440,N_11729,N_11768);
and U12441 (N_12441,N_11623,N_11852);
nand U12442 (N_12442,N_11958,N_11982);
and U12443 (N_12443,N_11772,N_11997);
nand U12444 (N_12444,N_11929,N_11818);
and U12445 (N_12445,N_11838,N_11742);
nand U12446 (N_12446,N_11687,N_11527);
and U12447 (N_12447,N_11716,N_11631);
xor U12448 (N_12448,N_11702,N_11966);
nor U12449 (N_12449,N_11618,N_11856);
xnor U12450 (N_12450,N_11556,N_11681);
xor U12451 (N_12451,N_11520,N_11617);
nand U12452 (N_12452,N_11518,N_11668);
nor U12453 (N_12453,N_11741,N_11857);
and U12454 (N_12454,N_11596,N_11597);
xnor U12455 (N_12455,N_11962,N_11618);
xnor U12456 (N_12456,N_11817,N_11847);
or U12457 (N_12457,N_11926,N_11600);
xor U12458 (N_12458,N_11623,N_11692);
and U12459 (N_12459,N_11842,N_11802);
xnor U12460 (N_12460,N_11567,N_11806);
nor U12461 (N_12461,N_11646,N_11693);
nand U12462 (N_12462,N_11574,N_11830);
xor U12463 (N_12463,N_11580,N_11691);
nor U12464 (N_12464,N_11564,N_11774);
or U12465 (N_12465,N_11705,N_11654);
nor U12466 (N_12466,N_11800,N_11554);
or U12467 (N_12467,N_11707,N_11988);
and U12468 (N_12468,N_11680,N_11755);
nand U12469 (N_12469,N_11620,N_11733);
xor U12470 (N_12470,N_11945,N_11703);
xor U12471 (N_12471,N_11675,N_11797);
xnor U12472 (N_12472,N_11963,N_11685);
and U12473 (N_12473,N_11606,N_11820);
or U12474 (N_12474,N_11734,N_11611);
or U12475 (N_12475,N_11505,N_11640);
nand U12476 (N_12476,N_11548,N_11967);
and U12477 (N_12477,N_11900,N_11795);
nand U12478 (N_12478,N_11960,N_11851);
and U12479 (N_12479,N_11561,N_11645);
or U12480 (N_12480,N_11836,N_11810);
or U12481 (N_12481,N_11749,N_11988);
nand U12482 (N_12482,N_11927,N_11502);
xnor U12483 (N_12483,N_11554,N_11576);
xnor U12484 (N_12484,N_11601,N_11967);
and U12485 (N_12485,N_11574,N_11519);
nand U12486 (N_12486,N_11714,N_11582);
nand U12487 (N_12487,N_11789,N_11674);
nor U12488 (N_12488,N_11864,N_11734);
or U12489 (N_12489,N_11558,N_11987);
or U12490 (N_12490,N_11814,N_11984);
and U12491 (N_12491,N_11745,N_11727);
nand U12492 (N_12492,N_11812,N_11624);
xor U12493 (N_12493,N_11519,N_11580);
and U12494 (N_12494,N_11914,N_11599);
and U12495 (N_12495,N_11600,N_11860);
and U12496 (N_12496,N_11606,N_11581);
or U12497 (N_12497,N_11644,N_11536);
or U12498 (N_12498,N_11770,N_11693);
and U12499 (N_12499,N_11880,N_11945);
or U12500 (N_12500,N_12333,N_12180);
xor U12501 (N_12501,N_12392,N_12441);
or U12502 (N_12502,N_12257,N_12395);
and U12503 (N_12503,N_12237,N_12393);
nand U12504 (N_12504,N_12286,N_12461);
nand U12505 (N_12505,N_12326,N_12493);
nor U12506 (N_12506,N_12018,N_12303);
and U12507 (N_12507,N_12318,N_12118);
xnor U12508 (N_12508,N_12101,N_12036);
and U12509 (N_12509,N_12131,N_12008);
and U12510 (N_12510,N_12343,N_12099);
and U12511 (N_12511,N_12438,N_12109);
nand U12512 (N_12512,N_12142,N_12121);
xnor U12513 (N_12513,N_12342,N_12273);
nor U12514 (N_12514,N_12351,N_12011);
or U12515 (N_12515,N_12282,N_12113);
nand U12516 (N_12516,N_12136,N_12074);
nor U12517 (N_12517,N_12266,N_12458);
xor U12518 (N_12518,N_12433,N_12375);
nor U12519 (N_12519,N_12495,N_12419);
and U12520 (N_12520,N_12256,N_12041);
xor U12521 (N_12521,N_12298,N_12184);
nor U12522 (N_12522,N_12323,N_12373);
or U12523 (N_12523,N_12030,N_12394);
nor U12524 (N_12524,N_12396,N_12426);
or U12525 (N_12525,N_12353,N_12094);
nand U12526 (N_12526,N_12452,N_12324);
nand U12527 (N_12527,N_12383,N_12022);
nor U12528 (N_12528,N_12001,N_12029);
xor U12529 (N_12529,N_12081,N_12049);
nand U12530 (N_12530,N_12454,N_12100);
or U12531 (N_12531,N_12183,N_12005);
or U12532 (N_12532,N_12095,N_12223);
nand U12533 (N_12533,N_12299,N_12388);
nor U12534 (N_12534,N_12337,N_12155);
xnor U12535 (N_12535,N_12272,N_12037);
and U12536 (N_12536,N_12439,N_12133);
xnor U12537 (N_12537,N_12243,N_12413);
nor U12538 (N_12538,N_12028,N_12140);
nand U12539 (N_12539,N_12235,N_12412);
or U12540 (N_12540,N_12479,N_12489);
or U12541 (N_12541,N_12411,N_12431);
or U12542 (N_12542,N_12244,N_12238);
or U12543 (N_12543,N_12421,N_12027);
and U12544 (N_12544,N_12080,N_12156);
xnor U12545 (N_12545,N_12170,N_12260);
nand U12546 (N_12546,N_12367,N_12089);
xnor U12547 (N_12547,N_12076,N_12124);
or U12548 (N_12548,N_12350,N_12130);
xor U12549 (N_12549,N_12239,N_12263);
nand U12550 (N_12550,N_12402,N_12294);
xnor U12551 (N_12551,N_12204,N_12186);
or U12552 (N_12552,N_12306,N_12476);
xnor U12553 (N_12553,N_12152,N_12195);
nor U12554 (N_12554,N_12056,N_12250);
xor U12555 (N_12555,N_12447,N_12295);
nor U12556 (N_12556,N_12006,N_12290);
xnor U12557 (N_12557,N_12415,N_12026);
or U12558 (N_12558,N_12078,N_12219);
or U12559 (N_12559,N_12482,N_12445);
nand U12560 (N_12560,N_12144,N_12284);
xnor U12561 (N_12561,N_12221,N_12448);
xnor U12562 (N_12562,N_12498,N_12356);
and U12563 (N_12563,N_12103,N_12416);
nand U12564 (N_12564,N_12134,N_12414);
nor U12565 (N_12565,N_12088,N_12400);
and U12566 (N_12566,N_12125,N_12405);
nand U12567 (N_12567,N_12443,N_12330);
or U12568 (N_12568,N_12399,N_12197);
nor U12569 (N_12569,N_12092,N_12168);
nor U12570 (N_12570,N_12345,N_12021);
or U12571 (N_12571,N_12382,N_12222);
or U12572 (N_12572,N_12214,N_12055);
or U12573 (N_12573,N_12348,N_12228);
xnor U12574 (N_12574,N_12010,N_12434);
nor U12575 (N_12575,N_12065,N_12230);
nor U12576 (N_12576,N_12391,N_12398);
xor U12577 (N_12577,N_12363,N_12457);
xnor U12578 (N_12578,N_12128,N_12016);
and U12579 (N_12579,N_12397,N_12496);
nand U12580 (N_12580,N_12096,N_12236);
and U12581 (N_12581,N_12034,N_12480);
and U12582 (N_12582,N_12329,N_12465);
and U12583 (N_12583,N_12310,N_12240);
or U12584 (N_12584,N_12174,N_12097);
xor U12585 (N_12585,N_12205,N_12473);
or U12586 (N_12586,N_12377,N_12090);
and U12587 (N_12587,N_12114,N_12105);
nand U12588 (N_12588,N_12060,N_12316);
nor U12589 (N_12589,N_12190,N_12147);
xnor U12590 (N_12590,N_12409,N_12360);
nand U12591 (N_12591,N_12317,N_12358);
nor U12592 (N_12592,N_12357,N_12137);
and U12593 (N_12593,N_12247,N_12213);
and U12594 (N_12594,N_12425,N_12064);
or U12595 (N_12595,N_12436,N_12371);
nand U12596 (N_12596,N_12442,N_12073);
xor U12597 (N_12597,N_12201,N_12004);
nand U12598 (N_12598,N_12051,N_12115);
or U12599 (N_12599,N_12408,N_12013);
nand U12600 (N_12600,N_12427,N_12252);
xnor U12601 (N_12601,N_12104,N_12313);
nor U12602 (N_12602,N_12403,N_12264);
or U12603 (N_12603,N_12162,N_12216);
and U12604 (N_12604,N_12042,N_12048);
nand U12605 (N_12605,N_12297,N_12422);
and U12606 (N_12606,N_12176,N_12093);
or U12607 (N_12607,N_12179,N_12429);
and U12608 (N_12608,N_12208,N_12420);
or U12609 (N_12609,N_12232,N_12366);
nor U12610 (N_12610,N_12033,N_12132);
and U12611 (N_12611,N_12122,N_12401);
or U12612 (N_12612,N_12325,N_12054);
or U12613 (N_12613,N_12296,N_12437);
xor U12614 (N_12614,N_12374,N_12492);
xnor U12615 (N_12615,N_12309,N_12475);
nand U12616 (N_12616,N_12069,N_12287);
xnor U12617 (N_12617,N_12261,N_12281);
nand U12618 (N_12618,N_12038,N_12071);
nor U12619 (N_12619,N_12206,N_12246);
nand U12620 (N_12620,N_12107,N_12117);
nand U12621 (N_12621,N_12462,N_12091);
nand U12622 (N_12622,N_12171,N_12161);
nor U12623 (N_12623,N_12410,N_12274);
and U12624 (N_12624,N_12423,N_12328);
nor U12625 (N_12625,N_12271,N_12307);
or U12626 (N_12626,N_12450,N_12052);
xnor U12627 (N_12627,N_12212,N_12196);
or U12628 (N_12628,N_12320,N_12334);
and U12629 (N_12629,N_12385,N_12300);
xnor U12630 (N_12630,N_12259,N_12058);
nand U12631 (N_12631,N_12165,N_12040);
and U12632 (N_12632,N_12460,N_12159);
xnor U12633 (N_12633,N_12157,N_12207);
nor U12634 (N_12634,N_12304,N_12477);
or U12635 (N_12635,N_12139,N_12389);
nor U12636 (N_12636,N_12308,N_12187);
and U12637 (N_12637,N_12497,N_12210);
nor U12638 (N_12638,N_12467,N_12311);
or U12639 (N_12639,N_12135,N_12061);
nor U12640 (N_12640,N_12209,N_12119);
nor U12641 (N_12641,N_12166,N_12087);
and U12642 (N_12642,N_12043,N_12446);
nor U12643 (N_12643,N_12149,N_12368);
nor U12644 (N_12644,N_12146,N_12319);
and U12645 (N_12645,N_12332,N_12015);
and U12646 (N_12646,N_12167,N_12478);
xnor U12647 (N_12647,N_12082,N_12490);
or U12648 (N_12648,N_12241,N_12491);
nand U12649 (N_12649,N_12127,N_12067);
nor U12650 (N_12650,N_12172,N_12075);
and U12651 (N_12651,N_12116,N_12032);
xor U12652 (N_12652,N_12321,N_12341);
nand U12653 (N_12653,N_12085,N_12463);
xor U12654 (N_12654,N_12083,N_12181);
nand U12655 (N_12655,N_12062,N_12203);
nand U12656 (N_12656,N_12023,N_12003);
and U12657 (N_12657,N_12251,N_12148);
xnor U12658 (N_12658,N_12380,N_12154);
and U12659 (N_12659,N_12077,N_12253);
nand U12660 (N_12660,N_12352,N_12488);
or U12661 (N_12661,N_12070,N_12111);
xor U12662 (N_12662,N_12215,N_12435);
nand U12663 (N_12663,N_12110,N_12378);
nor U12664 (N_12664,N_12002,N_12456);
or U12665 (N_12665,N_12007,N_12164);
xor U12666 (N_12666,N_12469,N_12258);
and U12667 (N_12667,N_12276,N_12163);
or U12668 (N_12668,N_12200,N_12072);
nand U12669 (N_12669,N_12384,N_12102);
nand U12670 (N_12670,N_12283,N_12335);
nand U12671 (N_12671,N_12193,N_12292);
or U12672 (N_12672,N_12362,N_12084);
nand U12673 (N_12673,N_12312,N_12047);
and U12674 (N_12674,N_12354,N_12305);
and U12675 (N_12675,N_12059,N_12270);
nor U12676 (N_12676,N_12129,N_12098);
nand U12677 (N_12677,N_12262,N_12359);
xor U12678 (N_12678,N_12227,N_12381);
nor U12679 (N_12679,N_12012,N_12444);
xor U12680 (N_12680,N_12050,N_12280);
nand U12681 (N_12681,N_12106,N_12024);
nor U12682 (N_12682,N_12202,N_12035);
or U12683 (N_12683,N_12386,N_12485);
nor U12684 (N_12684,N_12277,N_12123);
nor U12685 (N_12685,N_12379,N_12112);
or U12686 (N_12686,N_12406,N_12173);
or U12687 (N_12687,N_12301,N_12369);
xor U12688 (N_12688,N_12182,N_12459);
or U12689 (N_12689,N_12233,N_12349);
nor U12690 (N_12690,N_12407,N_12453);
nand U12691 (N_12691,N_12339,N_12249);
nand U12692 (N_12692,N_12269,N_12428);
or U12693 (N_12693,N_12120,N_12364);
nor U12694 (N_12694,N_12279,N_12019);
xnor U12695 (N_12695,N_12472,N_12199);
nand U12696 (N_12696,N_12372,N_12242);
nand U12697 (N_12697,N_12017,N_12229);
xor U12698 (N_12698,N_12254,N_12417);
nor U12699 (N_12699,N_12255,N_12045);
xor U12700 (N_12700,N_12178,N_12248);
nor U12701 (N_12701,N_12086,N_12177);
nor U12702 (N_12702,N_12265,N_12494);
xnor U12703 (N_12703,N_12138,N_12194);
or U12704 (N_12704,N_12151,N_12025);
nand U12705 (N_12705,N_12158,N_12031);
nand U12706 (N_12706,N_12145,N_12150);
nand U12707 (N_12707,N_12340,N_12390);
or U12708 (N_12708,N_12430,N_12474);
nand U12709 (N_12709,N_12291,N_12225);
nand U12710 (N_12710,N_12315,N_12484);
or U12711 (N_12711,N_12068,N_12169);
nand U12712 (N_12712,N_12486,N_12338);
nand U12713 (N_12713,N_12267,N_12314);
xnor U12714 (N_12714,N_12432,N_12376);
xor U12715 (N_12715,N_12000,N_12063);
nor U12716 (N_12716,N_12355,N_12387);
or U12717 (N_12717,N_12302,N_12499);
and U12718 (N_12718,N_12468,N_12039);
and U12719 (N_12719,N_12331,N_12141);
or U12720 (N_12720,N_12189,N_12175);
nor U12721 (N_12721,N_12451,N_12234);
or U12722 (N_12722,N_12275,N_12198);
or U12723 (N_12723,N_12231,N_12327);
and U12724 (N_12724,N_12336,N_12466);
nor U12725 (N_12725,N_12344,N_12226);
nand U12726 (N_12726,N_12185,N_12191);
xor U12727 (N_12727,N_12404,N_12218);
and U12728 (N_12728,N_12220,N_12470);
or U12729 (N_12729,N_12066,N_12365);
or U12730 (N_12730,N_12440,N_12449);
nand U12731 (N_12731,N_12285,N_12044);
or U12732 (N_12732,N_12293,N_12245);
nor U12733 (N_12733,N_12418,N_12160);
or U12734 (N_12734,N_12424,N_12211);
and U12735 (N_12735,N_12143,N_12217);
and U12736 (N_12736,N_12053,N_12046);
and U12737 (N_12737,N_12079,N_12153);
and U12738 (N_12738,N_12464,N_12126);
xnor U12739 (N_12739,N_12009,N_12289);
or U12740 (N_12740,N_12361,N_12322);
or U12741 (N_12741,N_12020,N_12455);
and U12742 (N_12742,N_12481,N_12471);
nor U12743 (N_12743,N_12014,N_12347);
or U12744 (N_12744,N_12057,N_12268);
and U12745 (N_12745,N_12108,N_12346);
nand U12746 (N_12746,N_12370,N_12288);
nand U12747 (N_12747,N_12487,N_12224);
nand U12748 (N_12748,N_12483,N_12192);
or U12749 (N_12749,N_12278,N_12188);
or U12750 (N_12750,N_12042,N_12090);
xnor U12751 (N_12751,N_12403,N_12304);
nand U12752 (N_12752,N_12189,N_12048);
nand U12753 (N_12753,N_12440,N_12040);
nand U12754 (N_12754,N_12475,N_12202);
xor U12755 (N_12755,N_12193,N_12375);
and U12756 (N_12756,N_12031,N_12345);
and U12757 (N_12757,N_12470,N_12465);
nor U12758 (N_12758,N_12040,N_12075);
xor U12759 (N_12759,N_12499,N_12495);
nand U12760 (N_12760,N_12193,N_12444);
and U12761 (N_12761,N_12342,N_12393);
or U12762 (N_12762,N_12075,N_12416);
xor U12763 (N_12763,N_12275,N_12017);
nor U12764 (N_12764,N_12003,N_12226);
nand U12765 (N_12765,N_12099,N_12158);
xnor U12766 (N_12766,N_12491,N_12331);
or U12767 (N_12767,N_12315,N_12301);
and U12768 (N_12768,N_12317,N_12150);
and U12769 (N_12769,N_12202,N_12369);
or U12770 (N_12770,N_12142,N_12242);
nand U12771 (N_12771,N_12232,N_12168);
nor U12772 (N_12772,N_12465,N_12011);
xor U12773 (N_12773,N_12355,N_12277);
and U12774 (N_12774,N_12198,N_12300);
nand U12775 (N_12775,N_12024,N_12134);
or U12776 (N_12776,N_12297,N_12250);
xnor U12777 (N_12777,N_12125,N_12346);
nand U12778 (N_12778,N_12037,N_12327);
or U12779 (N_12779,N_12105,N_12243);
nand U12780 (N_12780,N_12278,N_12013);
nor U12781 (N_12781,N_12480,N_12105);
nor U12782 (N_12782,N_12126,N_12477);
xnor U12783 (N_12783,N_12364,N_12496);
and U12784 (N_12784,N_12417,N_12400);
xnor U12785 (N_12785,N_12145,N_12186);
nand U12786 (N_12786,N_12433,N_12408);
nand U12787 (N_12787,N_12071,N_12049);
xor U12788 (N_12788,N_12029,N_12338);
or U12789 (N_12789,N_12077,N_12170);
or U12790 (N_12790,N_12027,N_12146);
and U12791 (N_12791,N_12433,N_12428);
nor U12792 (N_12792,N_12390,N_12214);
xnor U12793 (N_12793,N_12035,N_12495);
and U12794 (N_12794,N_12130,N_12116);
nand U12795 (N_12795,N_12167,N_12463);
nor U12796 (N_12796,N_12469,N_12041);
nand U12797 (N_12797,N_12376,N_12023);
nor U12798 (N_12798,N_12445,N_12497);
and U12799 (N_12799,N_12353,N_12338);
or U12800 (N_12800,N_12284,N_12365);
nor U12801 (N_12801,N_12365,N_12479);
and U12802 (N_12802,N_12319,N_12428);
and U12803 (N_12803,N_12160,N_12129);
xnor U12804 (N_12804,N_12431,N_12338);
or U12805 (N_12805,N_12313,N_12063);
nor U12806 (N_12806,N_12437,N_12081);
nor U12807 (N_12807,N_12092,N_12444);
or U12808 (N_12808,N_12156,N_12343);
nand U12809 (N_12809,N_12069,N_12005);
xnor U12810 (N_12810,N_12031,N_12169);
or U12811 (N_12811,N_12246,N_12274);
nand U12812 (N_12812,N_12223,N_12479);
and U12813 (N_12813,N_12276,N_12370);
or U12814 (N_12814,N_12104,N_12161);
xnor U12815 (N_12815,N_12363,N_12099);
nor U12816 (N_12816,N_12290,N_12340);
or U12817 (N_12817,N_12351,N_12109);
and U12818 (N_12818,N_12059,N_12368);
nor U12819 (N_12819,N_12239,N_12175);
nor U12820 (N_12820,N_12497,N_12094);
or U12821 (N_12821,N_12207,N_12052);
and U12822 (N_12822,N_12405,N_12058);
nor U12823 (N_12823,N_12206,N_12323);
nor U12824 (N_12824,N_12218,N_12466);
nand U12825 (N_12825,N_12087,N_12285);
or U12826 (N_12826,N_12324,N_12137);
nand U12827 (N_12827,N_12058,N_12389);
nand U12828 (N_12828,N_12383,N_12483);
xor U12829 (N_12829,N_12315,N_12284);
nand U12830 (N_12830,N_12389,N_12217);
nor U12831 (N_12831,N_12282,N_12314);
and U12832 (N_12832,N_12233,N_12390);
xnor U12833 (N_12833,N_12298,N_12329);
nor U12834 (N_12834,N_12165,N_12459);
xor U12835 (N_12835,N_12020,N_12194);
nor U12836 (N_12836,N_12356,N_12043);
or U12837 (N_12837,N_12046,N_12223);
and U12838 (N_12838,N_12160,N_12278);
xor U12839 (N_12839,N_12199,N_12253);
nand U12840 (N_12840,N_12343,N_12015);
and U12841 (N_12841,N_12435,N_12397);
or U12842 (N_12842,N_12179,N_12424);
nor U12843 (N_12843,N_12286,N_12462);
nor U12844 (N_12844,N_12008,N_12046);
nor U12845 (N_12845,N_12055,N_12257);
nand U12846 (N_12846,N_12487,N_12237);
xnor U12847 (N_12847,N_12078,N_12096);
nor U12848 (N_12848,N_12194,N_12385);
or U12849 (N_12849,N_12269,N_12173);
and U12850 (N_12850,N_12293,N_12271);
and U12851 (N_12851,N_12393,N_12125);
or U12852 (N_12852,N_12216,N_12420);
nand U12853 (N_12853,N_12132,N_12157);
nand U12854 (N_12854,N_12353,N_12388);
or U12855 (N_12855,N_12256,N_12152);
or U12856 (N_12856,N_12389,N_12435);
and U12857 (N_12857,N_12253,N_12168);
and U12858 (N_12858,N_12101,N_12006);
nand U12859 (N_12859,N_12397,N_12212);
nor U12860 (N_12860,N_12019,N_12112);
and U12861 (N_12861,N_12306,N_12178);
xnor U12862 (N_12862,N_12073,N_12485);
and U12863 (N_12863,N_12308,N_12320);
nand U12864 (N_12864,N_12298,N_12368);
nor U12865 (N_12865,N_12061,N_12431);
and U12866 (N_12866,N_12122,N_12402);
xnor U12867 (N_12867,N_12151,N_12437);
xnor U12868 (N_12868,N_12102,N_12092);
nand U12869 (N_12869,N_12056,N_12130);
and U12870 (N_12870,N_12395,N_12354);
and U12871 (N_12871,N_12003,N_12225);
xor U12872 (N_12872,N_12368,N_12171);
xor U12873 (N_12873,N_12117,N_12456);
or U12874 (N_12874,N_12180,N_12177);
and U12875 (N_12875,N_12031,N_12331);
nand U12876 (N_12876,N_12381,N_12232);
nor U12877 (N_12877,N_12328,N_12054);
xnor U12878 (N_12878,N_12124,N_12346);
nand U12879 (N_12879,N_12460,N_12310);
nand U12880 (N_12880,N_12061,N_12192);
nor U12881 (N_12881,N_12305,N_12120);
xnor U12882 (N_12882,N_12135,N_12284);
nor U12883 (N_12883,N_12038,N_12439);
or U12884 (N_12884,N_12053,N_12244);
xor U12885 (N_12885,N_12089,N_12285);
nor U12886 (N_12886,N_12454,N_12260);
or U12887 (N_12887,N_12098,N_12305);
nor U12888 (N_12888,N_12429,N_12146);
and U12889 (N_12889,N_12298,N_12058);
or U12890 (N_12890,N_12397,N_12330);
nor U12891 (N_12891,N_12497,N_12498);
nand U12892 (N_12892,N_12340,N_12036);
nand U12893 (N_12893,N_12178,N_12144);
nor U12894 (N_12894,N_12300,N_12102);
nor U12895 (N_12895,N_12498,N_12277);
or U12896 (N_12896,N_12194,N_12301);
xnor U12897 (N_12897,N_12255,N_12001);
xor U12898 (N_12898,N_12481,N_12255);
xnor U12899 (N_12899,N_12330,N_12260);
nor U12900 (N_12900,N_12030,N_12426);
or U12901 (N_12901,N_12196,N_12108);
and U12902 (N_12902,N_12325,N_12110);
nand U12903 (N_12903,N_12137,N_12376);
or U12904 (N_12904,N_12173,N_12293);
xnor U12905 (N_12905,N_12126,N_12223);
and U12906 (N_12906,N_12005,N_12151);
or U12907 (N_12907,N_12221,N_12198);
and U12908 (N_12908,N_12192,N_12263);
nor U12909 (N_12909,N_12331,N_12291);
and U12910 (N_12910,N_12268,N_12170);
and U12911 (N_12911,N_12325,N_12100);
nand U12912 (N_12912,N_12145,N_12406);
nand U12913 (N_12913,N_12275,N_12363);
xnor U12914 (N_12914,N_12124,N_12356);
xnor U12915 (N_12915,N_12386,N_12262);
xnor U12916 (N_12916,N_12368,N_12268);
xor U12917 (N_12917,N_12471,N_12341);
nor U12918 (N_12918,N_12060,N_12294);
or U12919 (N_12919,N_12081,N_12475);
or U12920 (N_12920,N_12180,N_12284);
nor U12921 (N_12921,N_12073,N_12272);
or U12922 (N_12922,N_12296,N_12112);
and U12923 (N_12923,N_12026,N_12429);
or U12924 (N_12924,N_12256,N_12158);
nand U12925 (N_12925,N_12299,N_12054);
or U12926 (N_12926,N_12468,N_12073);
or U12927 (N_12927,N_12300,N_12048);
nand U12928 (N_12928,N_12370,N_12496);
xor U12929 (N_12929,N_12086,N_12115);
nor U12930 (N_12930,N_12178,N_12230);
nand U12931 (N_12931,N_12353,N_12189);
nor U12932 (N_12932,N_12214,N_12174);
xnor U12933 (N_12933,N_12449,N_12415);
nor U12934 (N_12934,N_12496,N_12383);
or U12935 (N_12935,N_12338,N_12217);
xor U12936 (N_12936,N_12244,N_12007);
and U12937 (N_12937,N_12336,N_12373);
xnor U12938 (N_12938,N_12259,N_12235);
or U12939 (N_12939,N_12250,N_12174);
xnor U12940 (N_12940,N_12161,N_12017);
and U12941 (N_12941,N_12204,N_12166);
xnor U12942 (N_12942,N_12406,N_12274);
xor U12943 (N_12943,N_12017,N_12395);
nand U12944 (N_12944,N_12015,N_12116);
or U12945 (N_12945,N_12399,N_12168);
xor U12946 (N_12946,N_12056,N_12024);
nor U12947 (N_12947,N_12436,N_12206);
xor U12948 (N_12948,N_12349,N_12493);
or U12949 (N_12949,N_12159,N_12322);
or U12950 (N_12950,N_12262,N_12485);
xnor U12951 (N_12951,N_12278,N_12243);
nor U12952 (N_12952,N_12002,N_12090);
nand U12953 (N_12953,N_12057,N_12203);
nor U12954 (N_12954,N_12399,N_12228);
xnor U12955 (N_12955,N_12285,N_12300);
xor U12956 (N_12956,N_12394,N_12010);
xor U12957 (N_12957,N_12208,N_12281);
nand U12958 (N_12958,N_12207,N_12095);
nand U12959 (N_12959,N_12297,N_12029);
xnor U12960 (N_12960,N_12066,N_12018);
and U12961 (N_12961,N_12336,N_12455);
xor U12962 (N_12962,N_12004,N_12037);
nor U12963 (N_12963,N_12287,N_12138);
and U12964 (N_12964,N_12293,N_12455);
or U12965 (N_12965,N_12072,N_12112);
or U12966 (N_12966,N_12364,N_12046);
nor U12967 (N_12967,N_12024,N_12006);
nor U12968 (N_12968,N_12261,N_12260);
or U12969 (N_12969,N_12208,N_12144);
and U12970 (N_12970,N_12304,N_12361);
xor U12971 (N_12971,N_12007,N_12055);
nand U12972 (N_12972,N_12159,N_12468);
xnor U12973 (N_12973,N_12424,N_12439);
nor U12974 (N_12974,N_12174,N_12226);
and U12975 (N_12975,N_12261,N_12217);
xnor U12976 (N_12976,N_12367,N_12070);
nor U12977 (N_12977,N_12337,N_12499);
and U12978 (N_12978,N_12122,N_12029);
nor U12979 (N_12979,N_12327,N_12140);
xnor U12980 (N_12980,N_12436,N_12410);
nor U12981 (N_12981,N_12196,N_12001);
and U12982 (N_12982,N_12218,N_12306);
and U12983 (N_12983,N_12210,N_12165);
and U12984 (N_12984,N_12396,N_12152);
nand U12985 (N_12985,N_12091,N_12171);
or U12986 (N_12986,N_12372,N_12252);
nor U12987 (N_12987,N_12449,N_12469);
nor U12988 (N_12988,N_12281,N_12296);
and U12989 (N_12989,N_12465,N_12181);
and U12990 (N_12990,N_12231,N_12452);
or U12991 (N_12991,N_12428,N_12293);
xnor U12992 (N_12992,N_12225,N_12265);
and U12993 (N_12993,N_12014,N_12458);
xnor U12994 (N_12994,N_12388,N_12295);
nor U12995 (N_12995,N_12179,N_12371);
or U12996 (N_12996,N_12477,N_12109);
and U12997 (N_12997,N_12209,N_12101);
nand U12998 (N_12998,N_12089,N_12220);
and U12999 (N_12999,N_12425,N_12140);
or U13000 (N_13000,N_12958,N_12513);
nand U13001 (N_13001,N_12755,N_12758);
and U13002 (N_13002,N_12969,N_12874);
xnor U13003 (N_13003,N_12597,N_12771);
nand U13004 (N_13004,N_12650,N_12624);
xor U13005 (N_13005,N_12685,N_12670);
nor U13006 (N_13006,N_12655,N_12500);
nand U13007 (N_13007,N_12785,N_12636);
nor U13008 (N_13008,N_12551,N_12888);
and U13009 (N_13009,N_12817,N_12721);
and U13010 (N_13010,N_12664,N_12623);
nor U13011 (N_13011,N_12550,N_12825);
xor U13012 (N_13012,N_12812,N_12537);
nand U13013 (N_13013,N_12506,N_12644);
nand U13014 (N_13014,N_12704,N_12893);
nand U13015 (N_13015,N_12932,N_12764);
nand U13016 (N_13016,N_12991,N_12911);
xnor U13017 (N_13017,N_12663,N_12642);
nor U13018 (N_13018,N_12894,N_12542);
nor U13019 (N_13019,N_12973,N_12887);
and U13020 (N_13020,N_12773,N_12609);
nand U13021 (N_13021,N_12936,N_12787);
or U13022 (N_13022,N_12532,N_12892);
and U13023 (N_13023,N_12561,N_12846);
nor U13024 (N_13024,N_12985,N_12806);
nand U13025 (N_13025,N_12621,N_12730);
nand U13026 (N_13026,N_12614,N_12909);
nand U13027 (N_13027,N_12587,N_12610);
xor U13028 (N_13028,N_12805,N_12671);
xnor U13029 (N_13029,N_12914,N_12512);
nand U13030 (N_13030,N_12984,N_12800);
nand U13031 (N_13031,N_12856,N_12604);
xor U13032 (N_13032,N_12760,N_12665);
and U13033 (N_13033,N_12848,N_12908);
nor U13034 (N_13034,N_12601,N_12795);
nor U13035 (N_13035,N_12913,N_12545);
and U13036 (N_13036,N_12645,N_12835);
and U13037 (N_13037,N_12766,N_12581);
and U13038 (N_13038,N_12815,N_12699);
and U13039 (N_13039,N_12725,N_12631);
nor U13040 (N_13040,N_12682,N_12559);
nand U13041 (N_13041,N_12549,N_12741);
and U13042 (N_13042,N_12628,N_12865);
or U13043 (N_13043,N_12555,N_12576);
or U13044 (N_13044,N_12850,N_12625);
and U13045 (N_13045,N_12568,N_12728);
nor U13046 (N_13046,N_12627,N_12988);
and U13047 (N_13047,N_12578,N_12745);
nor U13048 (N_13048,N_12849,N_12620);
nand U13049 (N_13049,N_12509,N_12777);
nand U13050 (N_13050,N_12962,N_12851);
or U13051 (N_13051,N_12845,N_12928);
or U13052 (N_13052,N_12827,N_12789);
xor U13053 (N_13053,N_12660,N_12526);
nand U13054 (N_13054,N_12956,N_12823);
or U13055 (N_13055,N_12963,N_12633);
nand U13056 (N_13056,N_12582,N_12915);
xor U13057 (N_13057,N_12708,N_12743);
xor U13058 (N_13058,N_12612,N_12719);
nor U13059 (N_13059,N_12723,N_12592);
nor U13060 (N_13060,N_12989,N_12738);
xnor U13061 (N_13061,N_12536,N_12659);
xor U13062 (N_13062,N_12643,N_12674);
nor U13063 (N_13063,N_12905,N_12945);
xnor U13064 (N_13064,N_12733,N_12761);
and U13065 (N_13065,N_12554,N_12617);
xnor U13066 (N_13066,N_12833,N_12678);
nor U13067 (N_13067,N_12681,N_12540);
nor U13068 (N_13068,N_12531,N_12646);
nor U13069 (N_13069,N_12952,N_12838);
nor U13070 (N_13070,N_12781,N_12992);
and U13071 (N_13071,N_12747,N_12855);
and U13072 (N_13072,N_12565,N_12898);
nand U13073 (N_13073,N_12993,N_12955);
xor U13074 (N_13074,N_12701,N_12895);
xnor U13075 (N_13075,N_12979,N_12940);
nand U13076 (N_13076,N_12638,N_12960);
nor U13077 (N_13077,N_12837,N_12779);
nor U13078 (N_13078,N_12695,N_12971);
and U13079 (N_13079,N_12548,N_12890);
and U13080 (N_13080,N_12891,N_12954);
nor U13081 (N_13081,N_12784,N_12517);
and U13082 (N_13082,N_12937,N_12539);
xnor U13083 (N_13083,N_12949,N_12722);
or U13084 (N_13084,N_12982,N_12543);
nand U13085 (N_13085,N_12762,N_12921);
and U13086 (N_13086,N_12687,N_12753);
xnor U13087 (N_13087,N_12974,N_12562);
nor U13088 (N_13088,N_12804,N_12590);
xor U13089 (N_13089,N_12731,N_12616);
and U13090 (N_13090,N_12724,N_12713);
and U13091 (N_13091,N_12902,N_12712);
nand U13092 (N_13092,N_12515,N_12886);
or U13093 (N_13093,N_12688,N_12711);
nand U13094 (N_13094,N_12618,N_12756);
nor U13095 (N_13095,N_12875,N_12570);
or U13096 (N_13096,N_12818,N_12896);
xor U13097 (N_13097,N_12585,N_12705);
xor U13098 (N_13098,N_12808,N_12626);
xnor U13099 (N_13099,N_12706,N_12950);
or U13100 (N_13100,N_12700,N_12647);
xor U13101 (N_13101,N_12831,N_12683);
and U13102 (N_13102,N_12654,N_12709);
or U13103 (N_13103,N_12996,N_12727);
and U13104 (N_13104,N_12739,N_12853);
and U13105 (N_13105,N_12977,N_12630);
nand U13106 (N_13106,N_12583,N_12832);
nand U13107 (N_13107,N_12716,N_12944);
and U13108 (N_13108,N_12961,N_12652);
nand U13109 (N_13109,N_12596,N_12520);
xor U13110 (N_13110,N_12966,N_12686);
nand U13111 (N_13111,N_12946,N_12919);
xnor U13112 (N_13112,N_12567,N_12672);
nand U13113 (N_13113,N_12976,N_12514);
nor U13114 (N_13114,N_12829,N_12975);
xor U13115 (N_13115,N_12866,N_12553);
or U13116 (N_13116,N_12807,N_12508);
nor U13117 (N_13117,N_12987,N_12600);
nand U13118 (N_13118,N_12796,N_12676);
xor U13119 (N_13119,N_12953,N_12534);
xor U13120 (N_13120,N_12744,N_12883);
xnor U13121 (N_13121,N_12847,N_12603);
and U13122 (N_13122,N_12917,N_12613);
nor U13123 (N_13123,N_12792,N_12640);
nor U13124 (N_13124,N_12656,N_12941);
nor U13125 (N_13125,N_12588,N_12605);
or U13126 (N_13126,N_12729,N_12598);
xnor U13127 (N_13127,N_12813,N_12852);
nand U13128 (N_13128,N_12563,N_12594);
xor U13129 (N_13129,N_12589,N_12780);
nor U13130 (N_13130,N_12794,N_12697);
and U13131 (N_13131,N_12994,N_12591);
nand U13132 (N_13132,N_12965,N_12916);
and U13133 (N_13133,N_12602,N_12820);
or U13134 (N_13134,N_12749,N_12926);
nand U13135 (N_13135,N_12778,N_12673);
or U13136 (N_13136,N_12611,N_12740);
or U13137 (N_13137,N_12844,N_12521);
xnor U13138 (N_13138,N_12735,N_12879);
or U13139 (N_13139,N_12927,N_12912);
xor U13140 (N_13140,N_12904,N_12863);
nand U13141 (N_13141,N_12579,N_12821);
and U13142 (N_13142,N_12931,N_12751);
and U13143 (N_13143,N_12639,N_12869);
or U13144 (N_13144,N_12872,N_12742);
or U13145 (N_13145,N_12649,N_12797);
nand U13146 (N_13146,N_12897,N_12907);
nand U13147 (N_13147,N_12710,N_12607);
nor U13148 (N_13148,N_12586,N_12669);
xnor U13149 (N_13149,N_12910,N_12903);
nor U13150 (N_13150,N_12841,N_12861);
nand U13151 (N_13151,N_12803,N_12822);
xor U13152 (N_13152,N_12518,N_12703);
xor U13153 (N_13153,N_12889,N_12726);
and U13154 (N_13154,N_12791,N_12860);
and U13155 (N_13155,N_12793,N_12839);
nor U13156 (N_13156,N_12566,N_12775);
or U13157 (N_13157,N_12651,N_12957);
and U13158 (N_13158,N_12510,N_12843);
xor U13159 (N_13159,N_12533,N_12920);
nand U13160 (N_13160,N_12798,N_12680);
xnor U13161 (N_13161,N_12918,N_12980);
nor U13162 (N_13162,N_12877,N_12547);
and U13163 (N_13163,N_12560,N_12997);
and U13164 (N_13164,N_12629,N_12564);
and U13165 (N_13165,N_12575,N_12776);
nor U13166 (N_13166,N_12593,N_12767);
nor U13167 (N_13167,N_12868,N_12970);
or U13168 (N_13168,N_12720,N_12527);
and U13169 (N_13169,N_12675,N_12694);
nor U13170 (N_13170,N_12606,N_12964);
or U13171 (N_13171,N_12505,N_12943);
xnor U13172 (N_13172,N_12574,N_12535);
nand U13173 (N_13173,N_12774,N_12864);
or U13174 (N_13174,N_12939,N_12693);
xnor U13175 (N_13175,N_12922,N_12858);
and U13176 (N_13176,N_12502,N_12746);
and U13177 (N_13177,N_12859,N_12947);
nand U13178 (N_13178,N_12524,N_12689);
nor U13179 (N_13179,N_12811,N_12734);
nand U13180 (N_13180,N_12668,N_12923);
or U13181 (N_13181,N_12995,N_12990);
xnor U13182 (N_13182,N_12862,N_12632);
nor U13183 (N_13183,N_12790,N_12507);
nor U13184 (N_13184,N_12819,N_12615);
nand U13185 (N_13185,N_12986,N_12661);
or U13186 (N_13186,N_12692,N_12690);
and U13187 (N_13187,N_12679,N_12959);
xor U13188 (N_13188,N_12523,N_12836);
and U13189 (N_13189,N_12504,N_12881);
xor U13190 (N_13190,N_12658,N_12972);
or U13191 (N_13191,N_12870,N_12541);
or U13192 (N_13192,N_12840,N_12544);
nand U13193 (N_13193,N_12707,N_12934);
xor U13194 (N_13194,N_12769,N_12634);
xnor U13195 (N_13195,N_12653,N_12999);
or U13196 (N_13196,N_12906,N_12842);
and U13197 (N_13197,N_12801,N_12571);
xnor U13198 (N_13198,N_12828,N_12951);
nand U13199 (N_13199,N_12933,N_12608);
nor U13200 (N_13200,N_12691,N_12783);
and U13201 (N_13201,N_12718,N_12834);
nor U13202 (N_13202,N_12759,N_12648);
xnor U13203 (N_13203,N_12867,N_12511);
and U13204 (N_13204,N_12569,N_12935);
nand U13205 (N_13205,N_12657,N_12715);
xnor U13206 (N_13206,N_12599,N_12854);
nor U13207 (N_13207,N_12677,N_12750);
or U13208 (N_13208,N_12938,N_12814);
and U13209 (N_13209,N_12983,N_12768);
nor U13210 (N_13210,N_12667,N_12884);
nor U13211 (N_13211,N_12809,N_12871);
nor U13212 (N_13212,N_12885,N_12503);
or U13213 (N_13213,N_12876,N_12799);
xnor U13214 (N_13214,N_12595,N_12770);
or U13215 (N_13215,N_12528,N_12557);
nand U13216 (N_13216,N_12757,N_12763);
or U13217 (N_13217,N_12556,N_12998);
nor U13218 (N_13218,N_12516,N_12522);
nand U13219 (N_13219,N_12501,N_12529);
or U13220 (N_13220,N_12584,N_12978);
or U13221 (N_13221,N_12684,N_12873);
nand U13222 (N_13222,N_12622,N_12525);
xor U13223 (N_13223,N_12765,N_12830);
or U13224 (N_13224,N_12942,N_12802);
and U13225 (N_13225,N_12899,N_12748);
nand U13226 (N_13226,N_12857,N_12826);
xnor U13227 (N_13227,N_12737,N_12530);
xnor U13228 (N_13228,N_12732,N_12772);
nor U13229 (N_13229,N_12981,N_12878);
xnor U13230 (N_13230,N_12714,N_12968);
nor U13231 (N_13231,N_12538,N_12573);
xnor U13232 (N_13232,N_12782,N_12635);
and U13233 (N_13233,N_12948,N_12882);
xor U13234 (N_13234,N_12666,N_12572);
xnor U13235 (N_13235,N_12580,N_12519);
or U13236 (N_13236,N_12901,N_12925);
xnor U13237 (N_13237,N_12637,N_12641);
nand U13238 (N_13238,N_12702,N_12967);
and U13239 (N_13239,N_12717,N_12880);
nor U13240 (N_13240,N_12696,N_12754);
and U13241 (N_13241,N_12619,N_12924);
nor U13242 (N_13242,N_12929,N_12558);
nor U13243 (N_13243,N_12546,N_12752);
nor U13244 (N_13244,N_12698,N_12900);
and U13245 (N_13245,N_12930,N_12577);
and U13246 (N_13246,N_12816,N_12788);
and U13247 (N_13247,N_12786,N_12824);
and U13248 (N_13248,N_12736,N_12662);
xor U13249 (N_13249,N_12810,N_12552);
and U13250 (N_13250,N_12919,N_12887);
nor U13251 (N_13251,N_12678,N_12872);
and U13252 (N_13252,N_12868,N_12857);
nor U13253 (N_13253,N_12848,N_12598);
nor U13254 (N_13254,N_12616,N_12959);
nand U13255 (N_13255,N_12520,N_12605);
xnor U13256 (N_13256,N_12680,N_12672);
xnor U13257 (N_13257,N_12878,N_12911);
nor U13258 (N_13258,N_12578,N_12802);
or U13259 (N_13259,N_12570,N_12885);
xnor U13260 (N_13260,N_12732,N_12836);
or U13261 (N_13261,N_12911,N_12558);
nand U13262 (N_13262,N_12997,N_12533);
nand U13263 (N_13263,N_12678,N_12596);
xnor U13264 (N_13264,N_12735,N_12926);
or U13265 (N_13265,N_12883,N_12809);
nand U13266 (N_13266,N_12991,N_12563);
or U13267 (N_13267,N_12877,N_12918);
nand U13268 (N_13268,N_12810,N_12955);
and U13269 (N_13269,N_12553,N_12786);
nor U13270 (N_13270,N_12764,N_12590);
nand U13271 (N_13271,N_12690,N_12962);
xor U13272 (N_13272,N_12594,N_12848);
xor U13273 (N_13273,N_12518,N_12612);
and U13274 (N_13274,N_12803,N_12871);
nor U13275 (N_13275,N_12720,N_12552);
xor U13276 (N_13276,N_12558,N_12526);
nor U13277 (N_13277,N_12839,N_12904);
nand U13278 (N_13278,N_12659,N_12622);
nand U13279 (N_13279,N_12960,N_12695);
xor U13280 (N_13280,N_12693,N_12531);
nor U13281 (N_13281,N_12777,N_12719);
nand U13282 (N_13282,N_12590,N_12645);
nand U13283 (N_13283,N_12729,N_12508);
nor U13284 (N_13284,N_12590,N_12815);
xnor U13285 (N_13285,N_12864,N_12893);
nor U13286 (N_13286,N_12534,N_12656);
nand U13287 (N_13287,N_12943,N_12988);
nand U13288 (N_13288,N_12605,N_12537);
xor U13289 (N_13289,N_12947,N_12500);
xnor U13290 (N_13290,N_12830,N_12652);
nand U13291 (N_13291,N_12741,N_12506);
xnor U13292 (N_13292,N_12876,N_12915);
nor U13293 (N_13293,N_12822,N_12742);
xor U13294 (N_13294,N_12881,N_12957);
nand U13295 (N_13295,N_12799,N_12542);
and U13296 (N_13296,N_12646,N_12510);
and U13297 (N_13297,N_12644,N_12958);
xnor U13298 (N_13298,N_12751,N_12856);
and U13299 (N_13299,N_12564,N_12960);
xnor U13300 (N_13300,N_12622,N_12748);
nand U13301 (N_13301,N_12620,N_12505);
nand U13302 (N_13302,N_12931,N_12791);
xor U13303 (N_13303,N_12870,N_12989);
and U13304 (N_13304,N_12581,N_12604);
and U13305 (N_13305,N_12632,N_12600);
nand U13306 (N_13306,N_12631,N_12712);
or U13307 (N_13307,N_12985,N_12632);
xor U13308 (N_13308,N_12717,N_12584);
nor U13309 (N_13309,N_12724,N_12694);
or U13310 (N_13310,N_12956,N_12723);
nand U13311 (N_13311,N_12979,N_12959);
nor U13312 (N_13312,N_12734,N_12531);
and U13313 (N_13313,N_12882,N_12929);
and U13314 (N_13314,N_12965,N_12943);
and U13315 (N_13315,N_12895,N_12595);
xnor U13316 (N_13316,N_12850,N_12978);
nand U13317 (N_13317,N_12691,N_12906);
nor U13318 (N_13318,N_12641,N_12617);
xor U13319 (N_13319,N_12886,N_12586);
nor U13320 (N_13320,N_12593,N_12698);
nor U13321 (N_13321,N_12547,N_12988);
or U13322 (N_13322,N_12786,N_12604);
nor U13323 (N_13323,N_12702,N_12916);
or U13324 (N_13324,N_12576,N_12624);
nand U13325 (N_13325,N_12714,N_12864);
nor U13326 (N_13326,N_12946,N_12749);
and U13327 (N_13327,N_12508,N_12638);
or U13328 (N_13328,N_12675,N_12850);
and U13329 (N_13329,N_12766,N_12579);
xor U13330 (N_13330,N_12538,N_12957);
nor U13331 (N_13331,N_12899,N_12878);
xnor U13332 (N_13332,N_12707,N_12941);
and U13333 (N_13333,N_12582,N_12743);
xnor U13334 (N_13334,N_12790,N_12503);
nor U13335 (N_13335,N_12828,N_12814);
and U13336 (N_13336,N_12563,N_12567);
nor U13337 (N_13337,N_12556,N_12877);
and U13338 (N_13338,N_12715,N_12942);
nor U13339 (N_13339,N_12505,N_12584);
or U13340 (N_13340,N_12663,N_12900);
xor U13341 (N_13341,N_12798,N_12611);
xnor U13342 (N_13342,N_12624,N_12539);
nor U13343 (N_13343,N_12673,N_12660);
nor U13344 (N_13344,N_12870,N_12749);
and U13345 (N_13345,N_12950,N_12931);
or U13346 (N_13346,N_12733,N_12725);
nor U13347 (N_13347,N_12910,N_12866);
and U13348 (N_13348,N_12963,N_12608);
or U13349 (N_13349,N_12518,N_12903);
nor U13350 (N_13350,N_12886,N_12671);
nand U13351 (N_13351,N_12582,N_12754);
nor U13352 (N_13352,N_12838,N_12965);
or U13353 (N_13353,N_12866,N_12561);
nand U13354 (N_13354,N_12682,N_12545);
nor U13355 (N_13355,N_12720,N_12901);
or U13356 (N_13356,N_12698,N_12507);
nor U13357 (N_13357,N_12824,N_12552);
or U13358 (N_13358,N_12605,N_12895);
nor U13359 (N_13359,N_12915,N_12990);
nor U13360 (N_13360,N_12938,N_12909);
nand U13361 (N_13361,N_12834,N_12798);
nor U13362 (N_13362,N_12517,N_12752);
and U13363 (N_13363,N_12711,N_12704);
or U13364 (N_13364,N_12657,N_12926);
nand U13365 (N_13365,N_12939,N_12886);
or U13366 (N_13366,N_12655,N_12806);
xnor U13367 (N_13367,N_12661,N_12802);
xor U13368 (N_13368,N_12533,N_12519);
nor U13369 (N_13369,N_12825,N_12759);
nor U13370 (N_13370,N_12894,N_12645);
nor U13371 (N_13371,N_12664,N_12951);
xor U13372 (N_13372,N_12618,N_12923);
nor U13373 (N_13373,N_12731,N_12925);
nand U13374 (N_13374,N_12907,N_12874);
and U13375 (N_13375,N_12538,N_12887);
and U13376 (N_13376,N_12826,N_12618);
and U13377 (N_13377,N_12585,N_12736);
or U13378 (N_13378,N_12614,N_12731);
or U13379 (N_13379,N_12972,N_12629);
and U13380 (N_13380,N_12830,N_12519);
nor U13381 (N_13381,N_12778,N_12865);
or U13382 (N_13382,N_12880,N_12521);
nor U13383 (N_13383,N_12787,N_12833);
xnor U13384 (N_13384,N_12800,N_12612);
nor U13385 (N_13385,N_12914,N_12677);
nand U13386 (N_13386,N_12611,N_12781);
nor U13387 (N_13387,N_12637,N_12971);
nand U13388 (N_13388,N_12674,N_12641);
and U13389 (N_13389,N_12578,N_12637);
nor U13390 (N_13390,N_12520,N_12809);
or U13391 (N_13391,N_12505,N_12645);
xor U13392 (N_13392,N_12738,N_12882);
nand U13393 (N_13393,N_12789,N_12895);
nor U13394 (N_13394,N_12538,N_12563);
nor U13395 (N_13395,N_12992,N_12900);
xnor U13396 (N_13396,N_12681,N_12615);
nand U13397 (N_13397,N_12790,N_12509);
nor U13398 (N_13398,N_12589,N_12536);
nand U13399 (N_13399,N_12917,N_12646);
and U13400 (N_13400,N_12966,N_12691);
nand U13401 (N_13401,N_12528,N_12624);
and U13402 (N_13402,N_12556,N_12763);
nor U13403 (N_13403,N_12646,N_12979);
nand U13404 (N_13404,N_12509,N_12945);
xor U13405 (N_13405,N_12878,N_12640);
xnor U13406 (N_13406,N_12774,N_12733);
nand U13407 (N_13407,N_12704,N_12833);
nand U13408 (N_13408,N_12769,N_12930);
or U13409 (N_13409,N_12668,N_12682);
nor U13410 (N_13410,N_12734,N_12845);
or U13411 (N_13411,N_12784,N_12979);
and U13412 (N_13412,N_12556,N_12668);
nand U13413 (N_13413,N_12511,N_12694);
nor U13414 (N_13414,N_12719,N_12805);
and U13415 (N_13415,N_12778,N_12938);
nor U13416 (N_13416,N_12623,N_12541);
nand U13417 (N_13417,N_12576,N_12893);
or U13418 (N_13418,N_12692,N_12530);
or U13419 (N_13419,N_12508,N_12562);
xor U13420 (N_13420,N_12851,N_12974);
and U13421 (N_13421,N_12856,N_12940);
xor U13422 (N_13422,N_12712,N_12584);
and U13423 (N_13423,N_12635,N_12941);
or U13424 (N_13424,N_12907,N_12650);
nand U13425 (N_13425,N_12702,N_12818);
nand U13426 (N_13426,N_12726,N_12620);
and U13427 (N_13427,N_12574,N_12929);
and U13428 (N_13428,N_12651,N_12784);
nor U13429 (N_13429,N_12633,N_12899);
nor U13430 (N_13430,N_12781,N_12957);
nand U13431 (N_13431,N_12761,N_12547);
nand U13432 (N_13432,N_12691,N_12936);
xnor U13433 (N_13433,N_12544,N_12934);
xor U13434 (N_13434,N_12582,N_12824);
xor U13435 (N_13435,N_12515,N_12557);
nor U13436 (N_13436,N_12742,N_12679);
nor U13437 (N_13437,N_12698,N_12901);
and U13438 (N_13438,N_12807,N_12526);
nor U13439 (N_13439,N_12582,N_12584);
and U13440 (N_13440,N_12931,N_12822);
nor U13441 (N_13441,N_12772,N_12972);
xnor U13442 (N_13442,N_12882,N_12780);
nor U13443 (N_13443,N_12750,N_12972);
xnor U13444 (N_13444,N_12982,N_12869);
nand U13445 (N_13445,N_12832,N_12516);
xnor U13446 (N_13446,N_12868,N_12512);
xnor U13447 (N_13447,N_12796,N_12804);
and U13448 (N_13448,N_12734,N_12547);
nand U13449 (N_13449,N_12766,N_12623);
and U13450 (N_13450,N_12745,N_12877);
or U13451 (N_13451,N_12945,N_12995);
or U13452 (N_13452,N_12932,N_12885);
nor U13453 (N_13453,N_12691,N_12771);
xnor U13454 (N_13454,N_12648,N_12724);
nand U13455 (N_13455,N_12980,N_12508);
or U13456 (N_13456,N_12847,N_12842);
and U13457 (N_13457,N_12819,N_12664);
nor U13458 (N_13458,N_12956,N_12935);
nand U13459 (N_13459,N_12680,N_12561);
xor U13460 (N_13460,N_12712,N_12945);
and U13461 (N_13461,N_12953,N_12502);
or U13462 (N_13462,N_12815,N_12559);
and U13463 (N_13463,N_12711,N_12749);
and U13464 (N_13464,N_12586,N_12717);
nand U13465 (N_13465,N_12911,N_12562);
nor U13466 (N_13466,N_12523,N_12682);
or U13467 (N_13467,N_12533,N_12850);
xor U13468 (N_13468,N_12657,N_12859);
xor U13469 (N_13469,N_12842,N_12689);
and U13470 (N_13470,N_12672,N_12838);
xor U13471 (N_13471,N_12532,N_12859);
nor U13472 (N_13472,N_12708,N_12946);
xor U13473 (N_13473,N_12708,N_12721);
xor U13474 (N_13474,N_12732,N_12649);
or U13475 (N_13475,N_12717,N_12979);
or U13476 (N_13476,N_12802,N_12980);
or U13477 (N_13477,N_12568,N_12711);
nand U13478 (N_13478,N_12972,N_12979);
nand U13479 (N_13479,N_12558,N_12906);
nand U13480 (N_13480,N_12893,N_12792);
nor U13481 (N_13481,N_12970,N_12633);
nand U13482 (N_13482,N_12694,N_12561);
nand U13483 (N_13483,N_12878,N_12639);
nor U13484 (N_13484,N_12973,N_12503);
and U13485 (N_13485,N_12680,N_12772);
or U13486 (N_13486,N_12905,N_12823);
or U13487 (N_13487,N_12639,N_12652);
or U13488 (N_13488,N_12954,N_12783);
and U13489 (N_13489,N_12899,N_12733);
nor U13490 (N_13490,N_12629,N_12611);
nor U13491 (N_13491,N_12636,N_12614);
xnor U13492 (N_13492,N_12511,N_12888);
and U13493 (N_13493,N_12628,N_12738);
nand U13494 (N_13494,N_12902,N_12800);
and U13495 (N_13495,N_12842,N_12648);
nor U13496 (N_13496,N_12709,N_12766);
and U13497 (N_13497,N_12886,N_12717);
and U13498 (N_13498,N_12953,N_12750);
nor U13499 (N_13499,N_12935,N_12845);
xor U13500 (N_13500,N_13468,N_13248);
or U13501 (N_13501,N_13036,N_13095);
nand U13502 (N_13502,N_13480,N_13487);
nand U13503 (N_13503,N_13179,N_13329);
and U13504 (N_13504,N_13135,N_13301);
nand U13505 (N_13505,N_13255,N_13419);
and U13506 (N_13506,N_13281,N_13311);
and U13507 (N_13507,N_13396,N_13273);
or U13508 (N_13508,N_13360,N_13210);
or U13509 (N_13509,N_13139,N_13141);
and U13510 (N_13510,N_13312,N_13182);
nor U13511 (N_13511,N_13481,N_13336);
xnor U13512 (N_13512,N_13328,N_13047);
nand U13513 (N_13513,N_13226,N_13209);
nand U13514 (N_13514,N_13357,N_13298);
nand U13515 (N_13515,N_13362,N_13054);
or U13516 (N_13516,N_13014,N_13138);
and U13517 (N_13517,N_13451,N_13364);
nand U13518 (N_13518,N_13082,N_13458);
and U13519 (N_13519,N_13202,N_13446);
xor U13520 (N_13520,N_13274,N_13004);
nand U13521 (N_13521,N_13032,N_13253);
nor U13522 (N_13522,N_13296,N_13000);
or U13523 (N_13523,N_13476,N_13277);
nor U13524 (N_13524,N_13178,N_13087);
nor U13525 (N_13525,N_13031,N_13090);
nand U13526 (N_13526,N_13056,N_13465);
and U13527 (N_13527,N_13303,N_13279);
xnor U13528 (N_13528,N_13177,N_13350);
nand U13529 (N_13529,N_13400,N_13007);
and U13530 (N_13530,N_13453,N_13109);
or U13531 (N_13531,N_13028,N_13407);
nor U13532 (N_13532,N_13448,N_13349);
nand U13533 (N_13533,N_13211,N_13188);
or U13534 (N_13534,N_13406,N_13059);
nand U13535 (N_13535,N_13428,N_13409);
nand U13536 (N_13536,N_13471,N_13466);
and U13537 (N_13537,N_13333,N_13436);
nor U13538 (N_13538,N_13155,N_13467);
xnor U13539 (N_13539,N_13344,N_13153);
and U13540 (N_13540,N_13363,N_13175);
nand U13541 (N_13541,N_13143,N_13063);
nand U13542 (N_13542,N_13389,N_13170);
xnor U13543 (N_13543,N_13392,N_13072);
or U13544 (N_13544,N_13089,N_13067);
nor U13545 (N_13545,N_13173,N_13220);
xor U13546 (N_13546,N_13048,N_13423);
xor U13547 (N_13547,N_13245,N_13380);
and U13548 (N_13548,N_13447,N_13276);
nand U13549 (N_13549,N_13094,N_13314);
nor U13550 (N_13550,N_13099,N_13172);
and U13551 (N_13551,N_13140,N_13121);
nor U13552 (N_13552,N_13234,N_13215);
nor U13553 (N_13553,N_13294,N_13322);
and U13554 (N_13554,N_13414,N_13025);
nor U13555 (N_13555,N_13297,N_13435);
or U13556 (N_13556,N_13332,N_13093);
or U13557 (N_13557,N_13479,N_13079);
or U13558 (N_13558,N_13192,N_13161);
nand U13559 (N_13559,N_13433,N_13189);
or U13560 (N_13560,N_13216,N_13490);
and U13561 (N_13561,N_13424,N_13353);
nor U13562 (N_13562,N_13133,N_13163);
and U13563 (N_13563,N_13037,N_13417);
nand U13564 (N_13564,N_13271,N_13472);
nor U13565 (N_13565,N_13235,N_13038);
or U13566 (N_13566,N_13187,N_13016);
nor U13567 (N_13567,N_13387,N_13104);
or U13568 (N_13568,N_13391,N_13444);
and U13569 (N_13569,N_13002,N_13167);
and U13570 (N_13570,N_13009,N_13395);
nor U13571 (N_13571,N_13492,N_13237);
nor U13572 (N_13572,N_13158,N_13449);
or U13573 (N_13573,N_13431,N_13107);
xor U13574 (N_13574,N_13374,N_13377);
and U13575 (N_13575,N_13132,N_13166);
xor U13576 (N_13576,N_13434,N_13491);
and U13577 (N_13577,N_13223,N_13319);
or U13578 (N_13578,N_13194,N_13372);
nand U13579 (N_13579,N_13075,N_13205);
nor U13580 (N_13580,N_13217,N_13412);
or U13581 (N_13581,N_13200,N_13066);
xnor U13582 (N_13582,N_13097,N_13152);
or U13583 (N_13583,N_13219,N_13105);
xor U13584 (N_13584,N_13157,N_13456);
xor U13585 (N_13585,N_13213,N_13462);
nand U13586 (N_13586,N_13110,N_13044);
or U13587 (N_13587,N_13496,N_13069);
or U13588 (N_13588,N_13083,N_13484);
xor U13589 (N_13589,N_13488,N_13096);
and U13590 (N_13590,N_13231,N_13342);
nor U13591 (N_13591,N_13174,N_13345);
nand U13592 (N_13592,N_13136,N_13113);
nor U13593 (N_13593,N_13191,N_13003);
and U13594 (N_13594,N_13021,N_13290);
nor U13595 (N_13595,N_13498,N_13445);
or U13596 (N_13596,N_13247,N_13111);
or U13597 (N_13597,N_13049,N_13394);
nand U13598 (N_13598,N_13197,N_13416);
and U13599 (N_13599,N_13053,N_13493);
or U13600 (N_13600,N_13450,N_13029);
xor U13601 (N_13601,N_13088,N_13478);
or U13602 (N_13602,N_13365,N_13397);
nor U13603 (N_13603,N_13198,N_13461);
or U13604 (N_13604,N_13124,N_13227);
or U13605 (N_13605,N_13280,N_13061);
nand U13606 (N_13606,N_13454,N_13385);
nor U13607 (N_13607,N_13256,N_13199);
or U13608 (N_13608,N_13257,N_13159);
nor U13609 (N_13609,N_13258,N_13195);
or U13610 (N_13610,N_13183,N_13287);
nor U13611 (N_13611,N_13420,N_13052);
nand U13612 (N_13612,N_13373,N_13355);
xnor U13613 (N_13613,N_13438,N_13013);
xnor U13614 (N_13614,N_13019,N_13477);
nor U13615 (N_13615,N_13386,N_13230);
or U13616 (N_13616,N_13081,N_13410);
or U13617 (N_13617,N_13323,N_13078);
or U13618 (N_13618,N_13335,N_13254);
and U13619 (N_13619,N_13127,N_13317);
xnor U13620 (N_13620,N_13165,N_13125);
and U13621 (N_13621,N_13017,N_13015);
and U13622 (N_13622,N_13027,N_13086);
and U13623 (N_13623,N_13238,N_13370);
and U13624 (N_13624,N_13260,N_13318);
nor U13625 (N_13625,N_13084,N_13060);
xor U13626 (N_13626,N_13119,N_13232);
xor U13627 (N_13627,N_13250,N_13299);
xnor U13628 (N_13628,N_13288,N_13102);
and U13629 (N_13629,N_13313,N_13129);
xor U13630 (N_13630,N_13338,N_13282);
xnor U13631 (N_13631,N_13150,N_13413);
or U13632 (N_13632,N_13295,N_13265);
nand U13633 (N_13633,N_13270,N_13249);
and U13634 (N_13634,N_13243,N_13306);
nand U13635 (N_13635,N_13070,N_13405);
nor U13636 (N_13636,N_13128,N_13325);
and U13637 (N_13637,N_13246,N_13285);
or U13638 (N_13638,N_13429,N_13368);
xnor U13639 (N_13639,N_13421,N_13439);
nand U13640 (N_13640,N_13156,N_13452);
nor U13641 (N_13641,N_13310,N_13108);
and U13642 (N_13642,N_13092,N_13043);
nand U13643 (N_13643,N_13034,N_13403);
and U13644 (N_13644,N_13346,N_13040);
and U13645 (N_13645,N_13222,N_13278);
nand U13646 (N_13646,N_13304,N_13023);
and U13647 (N_13647,N_13240,N_13321);
nand U13648 (N_13648,N_13366,N_13390);
and U13649 (N_13649,N_13221,N_13154);
nor U13650 (N_13650,N_13340,N_13292);
and U13651 (N_13651,N_13184,N_13316);
nor U13652 (N_13652,N_13208,N_13418);
xnor U13653 (N_13653,N_13470,N_13206);
xnor U13654 (N_13654,N_13485,N_13196);
or U13655 (N_13655,N_13378,N_13399);
or U13656 (N_13656,N_13144,N_13126);
nor U13657 (N_13657,N_13148,N_13001);
nor U13658 (N_13658,N_13309,N_13051);
nor U13659 (N_13659,N_13176,N_13218);
and U13660 (N_13660,N_13459,N_13411);
nor U13661 (N_13661,N_13046,N_13171);
nand U13662 (N_13662,N_13062,N_13293);
and U13663 (N_13663,N_13499,N_13005);
xor U13664 (N_13664,N_13008,N_13214);
and U13665 (N_13665,N_13464,N_13057);
nand U13666 (N_13666,N_13455,N_13149);
or U13667 (N_13667,N_13489,N_13475);
nand U13668 (N_13668,N_13106,N_13358);
nand U13669 (N_13669,N_13112,N_13384);
xnor U13670 (N_13670,N_13033,N_13123);
nand U13671 (N_13671,N_13068,N_13229);
nand U13672 (N_13672,N_13151,N_13269);
xnor U13673 (N_13673,N_13483,N_13185);
and U13674 (N_13674,N_13233,N_13408);
or U13675 (N_13675,N_13204,N_13241);
and U13676 (N_13676,N_13065,N_13180);
or U13677 (N_13677,N_13207,N_13440);
nand U13678 (N_13678,N_13264,N_13193);
nand U13679 (N_13679,N_13291,N_13460);
nor U13680 (N_13680,N_13474,N_13118);
and U13681 (N_13681,N_13343,N_13324);
nor U13682 (N_13682,N_13388,N_13085);
xnor U13683 (N_13683,N_13259,N_13039);
xor U13684 (N_13684,N_13326,N_13283);
nor U13685 (N_13685,N_13441,N_13415);
nor U13686 (N_13686,N_13164,N_13045);
nor U13687 (N_13687,N_13361,N_13071);
nand U13688 (N_13688,N_13442,N_13263);
nor U13689 (N_13689,N_13073,N_13356);
and U13690 (N_13690,N_13236,N_13186);
or U13691 (N_13691,N_13116,N_13348);
xor U13692 (N_13692,N_13371,N_13120);
nand U13693 (N_13693,N_13076,N_13018);
or U13694 (N_13694,N_13268,N_13286);
and U13695 (N_13695,N_13103,N_13398);
or U13696 (N_13696,N_13382,N_13100);
nor U13697 (N_13697,N_13145,N_13266);
or U13698 (N_13698,N_13203,N_13341);
or U13699 (N_13699,N_13098,N_13181);
and U13700 (N_13700,N_13020,N_13275);
and U13701 (N_13701,N_13302,N_13327);
or U13702 (N_13702,N_13239,N_13042);
xnor U13703 (N_13703,N_13201,N_13427);
nand U13704 (N_13704,N_13212,N_13064);
nand U13705 (N_13705,N_13137,N_13284);
nor U13706 (N_13706,N_13339,N_13024);
nand U13707 (N_13707,N_13443,N_13463);
and U13708 (N_13708,N_13022,N_13228);
nor U13709 (N_13709,N_13315,N_13425);
and U13710 (N_13710,N_13404,N_13169);
nand U13711 (N_13711,N_13376,N_13430);
or U13712 (N_13712,N_13422,N_13012);
and U13713 (N_13713,N_13473,N_13077);
or U13714 (N_13714,N_13486,N_13162);
xor U13715 (N_13715,N_13101,N_13359);
nor U13716 (N_13716,N_13381,N_13224);
or U13717 (N_13717,N_13130,N_13331);
or U13718 (N_13718,N_13495,N_13337);
xor U13719 (N_13719,N_13334,N_13305);
nor U13720 (N_13720,N_13160,N_13497);
xnor U13721 (N_13721,N_13354,N_13190);
and U13722 (N_13722,N_13272,N_13330);
xor U13723 (N_13723,N_13383,N_13058);
or U13724 (N_13724,N_13026,N_13347);
and U13725 (N_13725,N_13437,N_13426);
nand U13726 (N_13726,N_13050,N_13494);
or U13727 (N_13727,N_13300,N_13351);
xnor U13728 (N_13728,N_13142,N_13035);
nor U13729 (N_13729,N_13369,N_13011);
xnor U13730 (N_13730,N_13080,N_13320);
nor U13731 (N_13731,N_13457,N_13393);
nor U13732 (N_13732,N_13352,N_13168);
or U13733 (N_13733,N_13401,N_13267);
or U13734 (N_13734,N_13030,N_13252);
or U13735 (N_13735,N_13402,N_13261);
nand U13736 (N_13736,N_13375,N_13482);
or U13737 (N_13737,N_13146,N_13469);
nor U13738 (N_13738,N_13147,N_13432);
or U13739 (N_13739,N_13041,N_13307);
or U13740 (N_13740,N_13117,N_13367);
or U13741 (N_13741,N_13379,N_13134);
or U13742 (N_13742,N_13242,N_13244);
nand U13743 (N_13743,N_13225,N_13114);
and U13744 (N_13744,N_13055,N_13289);
or U13745 (N_13745,N_13251,N_13115);
and U13746 (N_13746,N_13308,N_13006);
xor U13747 (N_13747,N_13131,N_13122);
and U13748 (N_13748,N_13262,N_13074);
and U13749 (N_13749,N_13091,N_13010);
or U13750 (N_13750,N_13106,N_13414);
or U13751 (N_13751,N_13168,N_13437);
and U13752 (N_13752,N_13340,N_13270);
or U13753 (N_13753,N_13096,N_13310);
nand U13754 (N_13754,N_13105,N_13411);
xor U13755 (N_13755,N_13313,N_13208);
and U13756 (N_13756,N_13035,N_13001);
nor U13757 (N_13757,N_13099,N_13465);
nand U13758 (N_13758,N_13083,N_13141);
or U13759 (N_13759,N_13496,N_13025);
and U13760 (N_13760,N_13114,N_13367);
nand U13761 (N_13761,N_13142,N_13474);
or U13762 (N_13762,N_13364,N_13450);
nor U13763 (N_13763,N_13122,N_13496);
nand U13764 (N_13764,N_13078,N_13032);
and U13765 (N_13765,N_13236,N_13238);
nor U13766 (N_13766,N_13107,N_13190);
or U13767 (N_13767,N_13385,N_13183);
nand U13768 (N_13768,N_13467,N_13143);
or U13769 (N_13769,N_13225,N_13398);
nor U13770 (N_13770,N_13133,N_13297);
nand U13771 (N_13771,N_13209,N_13218);
or U13772 (N_13772,N_13315,N_13279);
xnor U13773 (N_13773,N_13292,N_13131);
and U13774 (N_13774,N_13272,N_13171);
nor U13775 (N_13775,N_13310,N_13163);
nand U13776 (N_13776,N_13441,N_13290);
xor U13777 (N_13777,N_13442,N_13011);
nand U13778 (N_13778,N_13320,N_13462);
and U13779 (N_13779,N_13436,N_13117);
and U13780 (N_13780,N_13118,N_13004);
nand U13781 (N_13781,N_13417,N_13375);
nor U13782 (N_13782,N_13356,N_13227);
or U13783 (N_13783,N_13114,N_13109);
nand U13784 (N_13784,N_13323,N_13427);
nor U13785 (N_13785,N_13365,N_13255);
or U13786 (N_13786,N_13490,N_13230);
nand U13787 (N_13787,N_13323,N_13278);
nand U13788 (N_13788,N_13063,N_13249);
nand U13789 (N_13789,N_13155,N_13372);
nand U13790 (N_13790,N_13388,N_13071);
or U13791 (N_13791,N_13007,N_13419);
nand U13792 (N_13792,N_13148,N_13228);
nor U13793 (N_13793,N_13438,N_13003);
nor U13794 (N_13794,N_13423,N_13497);
nand U13795 (N_13795,N_13036,N_13334);
nand U13796 (N_13796,N_13070,N_13472);
nand U13797 (N_13797,N_13283,N_13205);
and U13798 (N_13798,N_13206,N_13245);
nor U13799 (N_13799,N_13272,N_13186);
and U13800 (N_13800,N_13473,N_13027);
xor U13801 (N_13801,N_13186,N_13191);
and U13802 (N_13802,N_13000,N_13462);
and U13803 (N_13803,N_13429,N_13444);
xnor U13804 (N_13804,N_13022,N_13208);
or U13805 (N_13805,N_13327,N_13296);
and U13806 (N_13806,N_13125,N_13231);
nor U13807 (N_13807,N_13311,N_13207);
or U13808 (N_13808,N_13433,N_13250);
nand U13809 (N_13809,N_13067,N_13076);
and U13810 (N_13810,N_13042,N_13376);
nor U13811 (N_13811,N_13393,N_13353);
or U13812 (N_13812,N_13305,N_13197);
xor U13813 (N_13813,N_13200,N_13382);
xor U13814 (N_13814,N_13435,N_13486);
and U13815 (N_13815,N_13418,N_13290);
xor U13816 (N_13816,N_13215,N_13495);
nor U13817 (N_13817,N_13312,N_13052);
xor U13818 (N_13818,N_13140,N_13489);
and U13819 (N_13819,N_13358,N_13185);
and U13820 (N_13820,N_13250,N_13453);
nor U13821 (N_13821,N_13409,N_13098);
nor U13822 (N_13822,N_13374,N_13264);
xor U13823 (N_13823,N_13112,N_13115);
or U13824 (N_13824,N_13202,N_13428);
xor U13825 (N_13825,N_13258,N_13159);
or U13826 (N_13826,N_13054,N_13408);
and U13827 (N_13827,N_13200,N_13073);
and U13828 (N_13828,N_13361,N_13259);
nor U13829 (N_13829,N_13322,N_13439);
and U13830 (N_13830,N_13120,N_13332);
nor U13831 (N_13831,N_13321,N_13257);
and U13832 (N_13832,N_13355,N_13045);
nor U13833 (N_13833,N_13124,N_13293);
nand U13834 (N_13834,N_13480,N_13105);
nand U13835 (N_13835,N_13084,N_13118);
and U13836 (N_13836,N_13000,N_13029);
nor U13837 (N_13837,N_13195,N_13317);
and U13838 (N_13838,N_13406,N_13375);
nand U13839 (N_13839,N_13231,N_13329);
nor U13840 (N_13840,N_13168,N_13303);
nor U13841 (N_13841,N_13085,N_13088);
and U13842 (N_13842,N_13265,N_13460);
xor U13843 (N_13843,N_13469,N_13192);
and U13844 (N_13844,N_13496,N_13187);
xor U13845 (N_13845,N_13229,N_13132);
or U13846 (N_13846,N_13440,N_13283);
and U13847 (N_13847,N_13040,N_13315);
nand U13848 (N_13848,N_13274,N_13343);
or U13849 (N_13849,N_13030,N_13159);
nor U13850 (N_13850,N_13051,N_13267);
nand U13851 (N_13851,N_13099,N_13343);
or U13852 (N_13852,N_13275,N_13018);
xor U13853 (N_13853,N_13359,N_13132);
or U13854 (N_13854,N_13049,N_13104);
xnor U13855 (N_13855,N_13236,N_13472);
nor U13856 (N_13856,N_13496,N_13323);
xnor U13857 (N_13857,N_13075,N_13161);
nand U13858 (N_13858,N_13025,N_13058);
or U13859 (N_13859,N_13341,N_13079);
and U13860 (N_13860,N_13337,N_13388);
nand U13861 (N_13861,N_13235,N_13322);
xnor U13862 (N_13862,N_13426,N_13250);
nand U13863 (N_13863,N_13118,N_13478);
or U13864 (N_13864,N_13192,N_13322);
or U13865 (N_13865,N_13415,N_13325);
nand U13866 (N_13866,N_13457,N_13054);
or U13867 (N_13867,N_13108,N_13447);
or U13868 (N_13868,N_13435,N_13343);
or U13869 (N_13869,N_13022,N_13145);
nor U13870 (N_13870,N_13349,N_13163);
nor U13871 (N_13871,N_13247,N_13160);
nor U13872 (N_13872,N_13280,N_13320);
xnor U13873 (N_13873,N_13489,N_13380);
nor U13874 (N_13874,N_13369,N_13178);
and U13875 (N_13875,N_13127,N_13177);
nand U13876 (N_13876,N_13035,N_13376);
nand U13877 (N_13877,N_13294,N_13173);
or U13878 (N_13878,N_13038,N_13118);
xnor U13879 (N_13879,N_13159,N_13106);
nand U13880 (N_13880,N_13359,N_13486);
or U13881 (N_13881,N_13148,N_13200);
and U13882 (N_13882,N_13254,N_13483);
or U13883 (N_13883,N_13396,N_13263);
xor U13884 (N_13884,N_13073,N_13354);
or U13885 (N_13885,N_13251,N_13279);
or U13886 (N_13886,N_13398,N_13471);
xnor U13887 (N_13887,N_13030,N_13175);
or U13888 (N_13888,N_13051,N_13108);
or U13889 (N_13889,N_13018,N_13321);
xor U13890 (N_13890,N_13092,N_13274);
and U13891 (N_13891,N_13218,N_13450);
and U13892 (N_13892,N_13340,N_13114);
xnor U13893 (N_13893,N_13025,N_13353);
and U13894 (N_13894,N_13024,N_13179);
nand U13895 (N_13895,N_13096,N_13108);
and U13896 (N_13896,N_13404,N_13271);
or U13897 (N_13897,N_13319,N_13453);
nor U13898 (N_13898,N_13162,N_13164);
nand U13899 (N_13899,N_13201,N_13006);
and U13900 (N_13900,N_13172,N_13425);
or U13901 (N_13901,N_13076,N_13102);
and U13902 (N_13902,N_13180,N_13186);
and U13903 (N_13903,N_13054,N_13145);
or U13904 (N_13904,N_13266,N_13146);
and U13905 (N_13905,N_13439,N_13362);
or U13906 (N_13906,N_13493,N_13255);
nand U13907 (N_13907,N_13085,N_13258);
nor U13908 (N_13908,N_13493,N_13432);
nand U13909 (N_13909,N_13267,N_13398);
xor U13910 (N_13910,N_13279,N_13232);
and U13911 (N_13911,N_13046,N_13160);
nor U13912 (N_13912,N_13294,N_13156);
nand U13913 (N_13913,N_13160,N_13315);
and U13914 (N_13914,N_13015,N_13135);
xor U13915 (N_13915,N_13479,N_13457);
xnor U13916 (N_13916,N_13267,N_13018);
or U13917 (N_13917,N_13236,N_13212);
xnor U13918 (N_13918,N_13349,N_13028);
xnor U13919 (N_13919,N_13195,N_13387);
nor U13920 (N_13920,N_13116,N_13272);
and U13921 (N_13921,N_13213,N_13396);
nand U13922 (N_13922,N_13056,N_13028);
nor U13923 (N_13923,N_13428,N_13016);
nand U13924 (N_13924,N_13191,N_13025);
and U13925 (N_13925,N_13362,N_13220);
or U13926 (N_13926,N_13060,N_13218);
xor U13927 (N_13927,N_13084,N_13337);
nor U13928 (N_13928,N_13459,N_13113);
nor U13929 (N_13929,N_13068,N_13326);
and U13930 (N_13930,N_13356,N_13196);
or U13931 (N_13931,N_13370,N_13341);
nor U13932 (N_13932,N_13336,N_13375);
and U13933 (N_13933,N_13050,N_13079);
xor U13934 (N_13934,N_13332,N_13351);
or U13935 (N_13935,N_13071,N_13341);
and U13936 (N_13936,N_13210,N_13393);
nand U13937 (N_13937,N_13289,N_13282);
nor U13938 (N_13938,N_13303,N_13325);
nand U13939 (N_13939,N_13283,N_13111);
nand U13940 (N_13940,N_13464,N_13268);
nor U13941 (N_13941,N_13273,N_13020);
and U13942 (N_13942,N_13320,N_13197);
and U13943 (N_13943,N_13190,N_13111);
or U13944 (N_13944,N_13136,N_13122);
xnor U13945 (N_13945,N_13386,N_13466);
or U13946 (N_13946,N_13290,N_13455);
nor U13947 (N_13947,N_13384,N_13162);
or U13948 (N_13948,N_13073,N_13079);
and U13949 (N_13949,N_13354,N_13357);
nand U13950 (N_13950,N_13045,N_13233);
nor U13951 (N_13951,N_13478,N_13465);
xor U13952 (N_13952,N_13468,N_13378);
and U13953 (N_13953,N_13077,N_13041);
xor U13954 (N_13954,N_13141,N_13075);
nand U13955 (N_13955,N_13298,N_13498);
or U13956 (N_13956,N_13339,N_13407);
or U13957 (N_13957,N_13310,N_13103);
and U13958 (N_13958,N_13278,N_13176);
nand U13959 (N_13959,N_13058,N_13181);
nand U13960 (N_13960,N_13090,N_13203);
or U13961 (N_13961,N_13138,N_13387);
nor U13962 (N_13962,N_13472,N_13150);
or U13963 (N_13963,N_13227,N_13165);
nor U13964 (N_13964,N_13341,N_13016);
and U13965 (N_13965,N_13106,N_13200);
xor U13966 (N_13966,N_13171,N_13137);
xnor U13967 (N_13967,N_13106,N_13267);
and U13968 (N_13968,N_13323,N_13371);
or U13969 (N_13969,N_13299,N_13009);
nor U13970 (N_13970,N_13458,N_13014);
xor U13971 (N_13971,N_13031,N_13386);
xnor U13972 (N_13972,N_13154,N_13437);
nand U13973 (N_13973,N_13334,N_13100);
or U13974 (N_13974,N_13085,N_13255);
xor U13975 (N_13975,N_13016,N_13171);
nor U13976 (N_13976,N_13006,N_13162);
xor U13977 (N_13977,N_13321,N_13141);
nor U13978 (N_13978,N_13449,N_13347);
or U13979 (N_13979,N_13169,N_13467);
nand U13980 (N_13980,N_13329,N_13133);
and U13981 (N_13981,N_13047,N_13074);
nand U13982 (N_13982,N_13035,N_13011);
xnor U13983 (N_13983,N_13461,N_13396);
nor U13984 (N_13984,N_13365,N_13492);
or U13985 (N_13985,N_13249,N_13205);
nand U13986 (N_13986,N_13215,N_13264);
or U13987 (N_13987,N_13195,N_13413);
and U13988 (N_13988,N_13330,N_13007);
nor U13989 (N_13989,N_13428,N_13257);
nor U13990 (N_13990,N_13163,N_13004);
xor U13991 (N_13991,N_13153,N_13190);
xnor U13992 (N_13992,N_13277,N_13118);
xor U13993 (N_13993,N_13255,N_13450);
xor U13994 (N_13994,N_13485,N_13310);
xor U13995 (N_13995,N_13144,N_13330);
nand U13996 (N_13996,N_13156,N_13453);
xnor U13997 (N_13997,N_13039,N_13254);
xnor U13998 (N_13998,N_13120,N_13244);
nor U13999 (N_13999,N_13481,N_13121);
nand U14000 (N_14000,N_13788,N_13760);
nand U14001 (N_14001,N_13609,N_13785);
nor U14002 (N_14002,N_13855,N_13852);
nor U14003 (N_14003,N_13822,N_13762);
or U14004 (N_14004,N_13794,N_13772);
nor U14005 (N_14005,N_13779,N_13702);
and U14006 (N_14006,N_13539,N_13726);
and U14007 (N_14007,N_13592,N_13918);
nor U14008 (N_14008,N_13747,N_13960);
xnor U14009 (N_14009,N_13645,N_13615);
nand U14010 (N_14010,N_13885,N_13742);
xnor U14011 (N_14011,N_13967,N_13781);
or U14012 (N_14012,N_13630,N_13571);
and U14013 (N_14013,N_13889,N_13997);
nand U14014 (N_14014,N_13533,N_13608);
and U14015 (N_14015,N_13984,N_13554);
nor U14016 (N_14016,N_13721,N_13530);
or U14017 (N_14017,N_13954,N_13665);
xnor U14018 (N_14018,N_13644,N_13986);
and U14019 (N_14019,N_13672,N_13769);
or U14020 (N_14020,N_13838,N_13687);
nor U14021 (N_14021,N_13866,N_13708);
nand U14022 (N_14022,N_13532,N_13707);
or U14023 (N_14023,N_13950,N_13650);
xnor U14024 (N_14024,N_13725,N_13836);
and U14025 (N_14025,N_13597,N_13992);
nand U14026 (N_14026,N_13511,N_13507);
and U14027 (N_14027,N_13872,N_13565);
xnor U14028 (N_14028,N_13913,N_13614);
or U14029 (N_14029,N_13828,N_13607);
xnor U14030 (N_14030,N_13655,N_13596);
or U14031 (N_14031,N_13955,N_13883);
and U14032 (N_14032,N_13520,N_13808);
or U14033 (N_14033,N_13518,N_13540);
and U14034 (N_14034,N_13865,N_13517);
and U14035 (N_14035,N_13504,N_13853);
nor U14036 (N_14036,N_13666,N_13871);
xor U14037 (N_14037,N_13776,N_13566);
nand U14038 (N_14038,N_13937,N_13935);
and U14039 (N_14039,N_13873,N_13682);
xnor U14040 (N_14040,N_13850,N_13624);
xor U14041 (N_14041,N_13878,N_13677);
or U14042 (N_14042,N_13928,N_13791);
nand U14043 (N_14043,N_13911,N_13800);
nand U14044 (N_14044,N_13670,N_13631);
nand U14045 (N_14045,N_13916,N_13629);
xnor U14046 (N_14046,N_13847,N_13861);
and U14047 (N_14047,N_13663,N_13538);
nand U14048 (N_14048,N_13844,N_13914);
or U14049 (N_14049,N_13525,N_13512);
xnor U14050 (N_14050,N_13896,N_13543);
xor U14051 (N_14051,N_13799,N_13733);
nand U14052 (N_14052,N_13719,N_13798);
xnor U14053 (N_14053,N_13537,N_13648);
xor U14054 (N_14054,N_13633,N_13999);
and U14055 (N_14055,N_13978,N_13612);
nand U14056 (N_14056,N_13976,N_13679);
nand U14057 (N_14057,N_13777,N_13970);
or U14058 (N_14058,N_13501,N_13859);
nand U14059 (N_14059,N_13979,N_13773);
xor U14060 (N_14060,N_13646,N_13958);
or U14061 (N_14061,N_13634,N_13793);
and U14062 (N_14062,N_13951,N_13635);
or U14063 (N_14063,N_13908,N_13524);
xnor U14064 (N_14064,N_13724,N_13503);
xor U14065 (N_14065,N_13647,N_13890);
or U14066 (N_14066,N_13681,N_13795);
xnor U14067 (N_14067,N_13548,N_13546);
and U14068 (N_14068,N_13764,N_13636);
and U14069 (N_14069,N_13660,N_13656);
and U14070 (N_14070,N_13673,N_13653);
and U14071 (N_14071,N_13741,N_13739);
nand U14072 (N_14072,N_13535,N_13750);
nor U14073 (N_14073,N_13903,N_13628);
and U14074 (N_14074,N_13796,N_13693);
nor U14075 (N_14075,N_13758,N_13744);
nand U14076 (N_14076,N_13829,N_13706);
and U14077 (N_14077,N_13560,N_13620);
nor U14078 (N_14078,N_13661,N_13920);
or U14079 (N_14079,N_13667,N_13998);
nand U14080 (N_14080,N_13917,N_13602);
nor U14081 (N_14081,N_13938,N_13782);
and U14082 (N_14082,N_13567,N_13731);
nand U14083 (N_14083,N_13888,N_13949);
nand U14084 (N_14084,N_13712,N_13572);
nand U14085 (N_14085,N_13601,N_13953);
and U14086 (N_14086,N_13519,N_13994);
or U14087 (N_14087,N_13698,N_13901);
or U14088 (N_14088,N_13618,N_13927);
nand U14089 (N_14089,N_13710,N_13716);
xnor U14090 (N_14090,N_13632,N_13505);
and U14091 (N_14091,N_13792,N_13689);
xnor U14092 (N_14092,N_13502,N_13743);
and U14093 (N_14093,N_13897,N_13522);
and U14094 (N_14094,N_13810,N_13685);
nand U14095 (N_14095,N_13748,N_13738);
or U14096 (N_14096,N_13649,N_13603);
nor U14097 (N_14097,N_13959,N_13995);
or U14098 (N_14098,N_13588,N_13867);
xnor U14099 (N_14099,N_13963,N_13893);
xor U14100 (N_14100,N_13616,N_13783);
nor U14101 (N_14101,N_13983,N_13876);
nor U14102 (N_14102,N_13766,N_13547);
nor U14103 (N_14103,N_13811,N_13541);
nand U14104 (N_14104,N_13837,N_13807);
and U14105 (N_14105,N_13912,N_13936);
or U14106 (N_14106,N_13559,N_13797);
xor U14107 (N_14107,N_13589,N_13642);
nand U14108 (N_14108,N_13723,N_13907);
or U14109 (N_14109,N_13858,N_13944);
nor U14110 (N_14110,N_13581,N_13801);
xnor U14111 (N_14111,N_13968,N_13513);
xor U14112 (N_14112,N_13638,N_13973);
nor U14113 (N_14113,N_13552,N_13771);
nor U14114 (N_14114,N_13851,N_13555);
nand U14115 (N_14115,N_13763,N_13942);
nand U14116 (N_14116,N_13842,N_13514);
nor U14117 (N_14117,N_13947,N_13508);
or U14118 (N_14118,N_13802,N_13599);
and U14119 (N_14119,N_13996,N_13722);
nor U14120 (N_14120,N_13606,N_13619);
and U14121 (N_14121,N_13678,N_13891);
or U14122 (N_14122,N_13803,N_13737);
nor U14123 (N_14123,N_13898,N_13544);
xnor U14124 (N_14124,N_13709,N_13759);
and U14125 (N_14125,N_13658,N_13860);
and U14126 (N_14126,N_13652,N_13510);
nand U14127 (N_14127,N_13985,N_13887);
nor U14128 (N_14128,N_13715,N_13840);
and U14129 (N_14129,N_13561,N_13969);
and U14130 (N_14130,N_13582,N_13923);
nor U14131 (N_14131,N_13946,N_13705);
nor U14132 (N_14132,N_13550,N_13965);
or U14133 (N_14133,N_13728,N_13730);
nand U14134 (N_14134,N_13906,N_13833);
nor U14135 (N_14135,N_13587,N_13882);
or U14136 (N_14136,N_13761,N_13961);
xor U14137 (N_14137,N_13506,N_13778);
nand U14138 (N_14138,N_13711,N_13956);
and U14139 (N_14139,N_13697,N_13880);
xnor U14140 (N_14140,N_13526,N_13557);
nor U14141 (N_14141,N_13625,N_13664);
xor U14142 (N_14142,N_13809,N_13659);
nand U14143 (N_14143,N_13831,N_13701);
or U14144 (N_14144,N_13734,N_13604);
nand U14145 (N_14145,N_13610,N_13875);
nor U14146 (N_14146,N_13804,N_13684);
and U14147 (N_14147,N_13825,N_13982);
nand U14148 (N_14148,N_13932,N_13749);
or U14149 (N_14149,N_13671,N_13756);
or U14150 (N_14150,N_13593,N_13720);
nor U14151 (N_14151,N_13639,N_13832);
xnor U14152 (N_14152,N_13848,N_13574);
nor U14153 (N_14153,N_13819,N_13700);
xor U14154 (N_14154,N_13899,N_13818);
nand U14155 (N_14155,N_13945,N_13590);
nand U14156 (N_14156,N_13657,N_13680);
or U14157 (N_14157,N_13521,N_13767);
nor U14158 (N_14158,N_13924,N_13516);
and U14159 (N_14159,N_13974,N_13562);
xor U14160 (N_14160,N_13688,N_13573);
xor U14161 (N_14161,N_13768,N_13790);
nor U14162 (N_14162,N_13568,N_13611);
and U14163 (N_14163,N_13886,N_13864);
or U14164 (N_14164,N_13922,N_13765);
and U14165 (N_14165,N_13643,N_13717);
and U14166 (N_14166,N_13905,N_13713);
or U14167 (N_14167,N_13839,N_13870);
or U14168 (N_14168,N_13826,N_13981);
or U14169 (N_14169,N_13570,N_13683);
and U14170 (N_14170,N_13988,N_13622);
and U14171 (N_14171,N_13740,N_13528);
and U14172 (N_14172,N_13919,N_13694);
xnor U14173 (N_14173,N_13784,N_13805);
or U14174 (N_14174,N_13676,N_13536);
nand U14175 (N_14175,N_13915,N_13894);
nand U14176 (N_14176,N_13929,N_13812);
nor U14177 (N_14177,N_13751,N_13754);
or U14178 (N_14178,N_13821,N_13863);
and U14179 (N_14179,N_13854,N_13736);
nor U14180 (N_14180,N_13626,N_13774);
nor U14181 (N_14181,N_13641,N_13962);
nor U14182 (N_14182,N_13904,N_13752);
and U14183 (N_14183,N_13987,N_13879);
or U14184 (N_14184,N_13869,N_13975);
xor U14185 (N_14185,N_13718,N_13827);
and U14186 (N_14186,N_13551,N_13627);
nand U14187 (N_14187,N_13699,N_13757);
nor U14188 (N_14188,N_13654,N_13993);
nor U14189 (N_14189,N_13835,N_13696);
nor U14190 (N_14190,N_13534,N_13934);
and U14191 (N_14191,N_13892,N_13753);
or U14192 (N_14192,N_13881,N_13745);
and U14193 (N_14193,N_13605,N_13991);
nand U14194 (N_14194,N_13529,N_13598);
or U14195 (N_14195,N_13877,N_13868);
nor U14196 (N_14196,N_13527,N_13775);
nand U14197 (N_14197,N_13563,N_13515);
nor U14198 (N_14198,N_13846,N_13553);
xor U14199 (N_14199,N_13841,N_13662);
nor U14200 (N_14200,N_13952,N_13637);
xnor U14201 (N_14201,N_13977,N_13930);
xor U14202 (N_14202,N_13780,N_13755);
and U14203 (N_14203,N_13948,N_13583);
xor U14204 (N_14204,N_13895,N_13824);
xnor U14205 (N_14205,N_13806,N_13813);
nand U14206 (N_14206,N_13910,N_13900);
or U14207 (N_14207,N_13558,N_13770);
or U14208 (N_14208,N_13786,N_13845);
nor U14209 (N_14209,N_13925,N_13675);
nor U14210 (N_14210,N_13823,N_13617);
nand U14211 (N_14211,N_13580,N_13690);
and U14212 (N_14212,N_13972,N_13816);
or U14213 (N_14213,N_13509,N_13549);
nand U14214 (N_14214,N_13692,N_13909);
nand U14215 (N_14215,N_13595,N_13523);
xor U14216 (N_14216,N_13669,N_13735);
nand U14217 (N_14217,N_13668,N_13817);
xnor U14218 (N_14218,N_13874,N_13989);
nor U14219 (N_14219,N_13862,N_13594);
and U14220 (N_14220,N_13542,N_13941);
nand U14221 (N_14221,N_13990,N_13545);
or U14222 (N_14222,N_13746,N_13815);
nor U14223 (N_14223,N_13814,N_13576);
nand U14224 (N_14224,N_13843,N_13964);
xor U14225 (N_14225,N_13933,N_13621);
nor U14226 (N_14226,N_13577,N_13695);
nor U14227 (N_14227,N_13940,N_13921);
xor U14228 (N_14228,N_13575,N_13789);
xor U14229 (N_14229,N_13727,N_13966);
or U14230 (N_14230,N_13600,N_13686);
nor U14231 (N_14231,N_13849,N_13787);
and U14232 (N_14232,N_13500,N_13926);
or U14233 (N_14233,N_13704,N_13586);
nor U14234 (N_14234,N_13830,N_13971);
nor U14235 (N_14235,N_13613,N_13591);
and U14236 (N_14236,N_13578,N_13584);
or U14237 (N_14237,N_13931,N_13556);
nor U14238 (N_14238,N_13691,N_13902);
xnor U14239 (N_14239,N_13857,N_13640);
or U14240 (N_14240,N_13856,N_13834);
nand U14241 (N_14241,N_13732,N_13585);
nand U14242 (N_14242,N_13579,N_13729);
nor U14243 (N_14243,N_13703,N_13884);
and U14244 (N_14244,N_13980,N_13651);
nand U14245 (N_14245,N_13564,N_13943);
xor U14246 (N_14246,N_13939,N_13623);
or U14247 (N_14247,N_13531,N_13569);
or U14248 (N_14248,N_13957,N_13674);
xor U14249 (N_14249,N_13820,N_13714);
or U14250 (N_14250,N_13975,N_13766);
nand U14251 (N_14251,N_13961,N_13890);
xor U14252 (N_14252,N_13636,N_13744);
nor U14253 (N_14253,N_13549,N_13728);
or U14254 (N_14254,N_13956,N_13542);
and U14255 (N_14255,N_13561,N_13626);
nor U14256 (N_14256,N_13618,N_13923);
xor U14257 (N_14257,N_13636,N_13844);
nor U14258 (N_14258,N_13842,N_13590);
nor U14259 (N_14259,N_13838,N_13981);
xnor U14260 (N_14260,N_13724,N_13685);
and U14261 (N_14261,N_13672,N_13878);
nand U14262 (N_14262,N_13878,N_13708);
and U14263 (N_14263,N_13584,N_13619);
and U14264 (N_14264,N_13770,N_13809);
nand U14265 (N_14265,N_13521,N_13516);
nand U14266 (N_14266,N_13700,N_13698);
nand U14267 (N_14267,N_13585,N_13834);
or U14268 (N_14268,N_13639,N_13576);
xor U14269 (N_14269,N_13956,N_13689);
xnor U14270 (N_14270,N_13975,N_13891);
and U14271 (N_14271,N_13668,N_13855);
and U14272 (N_14272,N_13942,N_13776);
nor U14273 (N_14273,N_13851,N_13814);
nor U14274 (N_14274,N_13763,N_13728);
xor U14275 (N_14275,N_13654,N_13531);
nor U14276 (N_14276,N_13607,N_13932);
nand U14277 (N_14277,N_13559,N_13693);
and U14278 (N_14278,N_13903,N_13850);
nor U14279 (N_14279,N_13917,N_13592);
xnor U14280 (N_14280,N_13776,N_13740);
or U14281 (N_14281,N_13954,N_13947);
nor U14282 (N_14282,N_13508,N_13818);
nand U14283 (N_14283,N_13609,N_13589);
nor U14284 (N_14284,N_13500,N_13540);
xor U14285 (N_14285,N_13565,N_13989);
and U14286 (N_14286,N_13580,N_13942);
nand U14287 (N_14287,N_13725,N_13828);
nand U14288 (N_14288,N_13932,N_13552);
or U14289 (N_14289,N_13515,N_13839);
or U14290 (N_14290,N_13623,N_13673);
and U14291 (N_14291,N_13766,N_13658);
and U14292 (N_14292,N_13748,N_13515);
or U14293 (N_14293,N_13775,N_13589);
xnor U14294 (N_14294,N_13870,N_13876);
nand U14295 (N_14295,N_13922,N_13722);
nand U14296 (N_14296,N_13694,N_13881);
xnor U14297 (N_14297,N_13528,N_13792);
nand U14298 (N_14298,N_13773,N_13945);
or U14299 (N_14299,N_13752,N_13746);
xor U14300 (N_14300,N_13978,N_13760);
nor U14301 (N_14301,N_13599,N_13775);
or U14302 (N_14302,N_13534,N_13634);
and U14303 (N_14303,N_13748,N_13910);
and U14304 (N_14304,N_13960,N_13711);
nor U14305 (N_14305,N_13760,N_13785);
xor U14306 (N_14306,N_13565,N_13995);
nand U14307 (N_14307,N_13624,N_13688);
and U14308 (N_14308,N_13850,N_13844);
nor U14309 (N_14309,N_13508,N_13793);
or U14310 (N_14310,N_13914,N_13949);
nand U14311 (N_14311,N_13861,N_13840);
xnor U14312 (N_14312,N_13836,N_13924);
xor U14313 (N_14313,N_13566,N_13808);
and U14314 (N_14314,N_13550,N_13880);
nand U14315 (N_14315,N_13968,N_13995);
and U14316 (N_14316,N_13925,N_13515);
xor U14317 (N_14317,N_13594,N_13696);
or U14318 (N_14318,N_13705,N_13667);
nor U14319 (N_14319,N_13808,N_13807);
nor U14320 (N_14320,N_13649,N_13897);
nor U14321 (N_14321,N_13537,N_13965);
or U14322 (N_14322,N_13776,N_13959);
or U14323 (N_14323,N_13562,N_13630);
or U14324 (N_14324,N_13706,N_13540);
nor U14325 (N_14325,N_13674,N_13971);
nand U14326 (N_14326,N_13611,N_13577);
nand U14327 (N_14327,N_13743,N_13558);
and U14328 (N_14328,N_13818,N_13706);
nor U14329 (N_14329,N_13647,N_13563);
nand U14330 (N_14330,N_13600,N_13985);
nand U14331 (N_14331,N_13672,N_13527);
or U14332 (N_14332,N_13751,N_13959);
and U14333 (N_14333,N_13955,N_13732);
and U14334 (N_14334,N_13915,N_13801);
xnor U14335 (N_14335,N_13556,N_13751);
nand U14336 (N_14336,N_13811,N_13635);
or U14337 (N_14337,N_13696,N_13752);
xor U14338 (N_14338,N_13818,N_13587);
nor U14339 (N_14339,N_13568,N_13614);
nor U14340 (N_14340,N_13926,N_13927);
xor U14341 (N_14341,N_13664,N_13855);
and U14342 (N_14342,N_13857,N_13911);
or U14343 (N_14343,N_13545,N_13725);
xnor U14344 (N_14344,N_13720,N_13979);
or U14345 (N_14345,N_13668,N_13736);
or U14346 (N_14346,N_13904,N_13896);
and U14347 (N_14347,N_13884,N_13755);
and U14348 (N_14348,N_13537,N_13628);
xnor U14349 (N_14349,N_13829,N_13618);
or U14350 (N_14350,N_13892,N_13739);
or U14351 (N_14351,N_13623,N_13831);
xor U14352 (N_14352,N_13642,N_13790);
or U14353 (N_14353,N_13901,N_13684);
or U14354 (N_14354,N_13982,N_13933);
and U14355 (N_14355,N_13676,N_13749);
and U14356 (N_14356,N_13783,N_13553);
nor U14357 (N_14357,N_13650,N_13598);
or U14358 (N_14358,N_13895,N_13643);
and U14359 (N_14359,N_13911,N_13718);
nor U14360 (N_14360,N_13854,N_13752);
nand U14361 (N_14361,N_13949,N_13699);
xnor U14362 (N_14362,N_13758,N_13747);
or U14363 (N_14363,N_13903,N_13834);
or U14364 (N_14364,N_13901,N_13511);
nor U14365 (N_14365,N_13876,N_13748);
and U14366 (N_14366,N_13525,N_13983);
xor U14367 (N_14367,N_13621,N_13583);
or U14368 (N_14368,N_13913,N_13557);
nor U14369 (N_14369,N_13503,N_13870);
and U14370 (N_14370,N_13920,N_13770);
nand U14371 (N_14371,N_13739,N_13507);
xor U14372 (N_14372,N_13870,N_13743);
nor U14373 (N_14373,N_13546,N_13514);
nor U14374 (N_14374,N_13795,N_13792);
or U14375 (N_14375,N_13611,N_13855);
xor U14376 (N_14376,N_13886,N_13512);
or U14377 (N_14377,N_13677,N_13792);
and U14378 (N_14378,N_13596,N_13928);
xnor U14379 (N_14379,N_13671,N_13539);
or U14380 (N_14380,N_13631,N_13789);
xnor U14381 (N_14381,N_13510,N_13675);
nand U14382 (N_14382,N_13685,N_13711);
xor U14383 (N_14383,N_13848,N_13714);
and U14384 (N_14384,N_13866,N_13693);
nor U14385 (N_14385,N_13878,N_13910);
or U14386 (N_14386,N_13906,N_13717);
nor U14387 (N_14387,N_13757,N_13758);
xor U14388 (N_14388,N_13877,N_13756);
or U14389 (N_14389,N_13831,N_13707);
or U14390 (N_14390,N_13568,N_13827);
xor U14391 (N_14391,N_13883,N_13989);
or U14392 (N_14392,N_13703,N_13702);
xnor U14393 (N_14393,N_13521,N_13713);
nor U14394 (N_14394,N_13943,N_13788);
xnor U14395 (N_14395,N_13764,N_13937);
and U14396 (N_14396,N_13702,N_13527);
xor U14397 (N_14397,N_13926,N_13778);
nand U14398 (N_14398,N_13511,N_13979);
xor U14399 (N_14399,N_13729,N_13971);
nor U14400 (N_14400,N_13785,N_13596);
xor U14401 (N_14401,N_13540,N_13834);
xnor U14402 (N_14402,N_13869,N_13723);
and U14403 (N_14403,N_13927,N_13674);
or U14404 (N_14404,N_13692,N_13555);
nor U14405 (N_14405,N_13746,N_13519);
or U14406 (N_14406,N_13641,N_13657);
nor U14407 (N_14407,N_13748,N_13535);
or U14408 (N_14408,N_13939,N_13646);
nand U14409 (N_14409,N_13945,N_13783);
and U14410 (N_14410,N_13945,N_13842);
nand U14411 (N_14411,N_13984,N_13883);
xnor U14412 (N_14412,N_13847,N_13588);
nor U14413 (N_14413,N_13724,N_13983);
xnor U14414 (N_14414,N_13918,N_13520);
nor U14415 (N_14415,N_13680,N_13949);
nand U14416 (N_14416,N_13644,N_13762);
and U14417 (N_14417,N_13919,N_13843);
nand U14418 (N_14418,N_13519,N_13613);
and U14419 (N_14419,N_13904,N_13792);
nand U14420 (N_14420,N_13934,N_13850);
and U14421 (N_14421,N_13708,N_13775);
nand U14422 (N_14422,N_13739,N_13774);
or U14423 (N_14423,N_13746,N_13888);
and U14424 (N_14424,N_13786,N_13595);
nor U14425 (N_14425,N_13777,N_13592);
and U14426 (N_14426,N_13883,N_13823);
and U14427 (N_14427,N_13509,N_13827);
and U14428 (N_14428,N_13869,N_13596);
and U14429 (N_14429,N_13575,N_13654);
nand U14430 (N_14430,N_13721,N_13960);
nand U14431 (N_14431,N_13519,N_13910);
and U14432 (N_14432,N_13855,N_13988);
or U14433 (N_14433,N_13895,N_13700);
nand U14434 (N_14434,N_13835,N_13736);
or U14435 (N_14435,N_13559,N_13788);
or U14436 (N_14436,N_13529,N_13961);
xor U14437 (N_14437,N_13694,N_13810);
and U14438 (N_14438,N_13963,N_13770);
and U14439 (N_14439,N_13645,N_13986);
or U14440 (N_14440,N_13858,N_13824);
xnor U14441 (N_14441,N_13762,N_13810);
nor U14442 (N_14442,N_13952,N_13552);
or U14443 (N_14443,N_13852,N_13749);
xor U14444 (N_14444,N_13542,N_13964);
and U14445 (N_14445,N_13648,N_13800);
nor U14446 (N_14446,N_13646,N_13692);
xnor U14447 (N_14447,N_13726,N_13740);
or U14448 (N_14448,N_13608,N_13787);
nand U14449 (N_14449,N_13948,N_13623);
xor U14450 (N_14450,N_13977,N_13564);
and U14451 (N_14451,N_13723,N_13722);
nand U14452 (N_14452,N_13517,N_13529);
or U14453 (N_14453,N_13677,N_13521);
nor U14454 (N_14454,N_13534,N_13683);
and U14455 (N_14455,N_13709,N_13638);
and U14456 (N_14456,N_13534,N_13931);
nand U14457 (N_14457,N_13844,N_13526);
xnor U14458 (N_14458,N_13644,N_13912);
nor U14459 (N_14459,N_13608,N_13621);
xor U14460 (N_14460,N_13542,N_13825);
xor U14461 (N_14461,N_13678,N_13593);
nand U14462 (N_14462,N_13981,N_13741);
nand U14463 (N_14463,N_13965,N_13954);
nand U14464 (N_14464,N_13806,N_13607);
or U14465 (N_14465,N_13634,N_13949);
xor U14466 (N_14466,N_13797,N_13737);
or U14467 (N_14467,N_13916,N_13965);
or U14468 (N_14468,N_13847,N_13590);
or U14469 (N_14469,N_13811,N_13928);
nor U14470 (N_14470,N_13855,N_13673);
nor U14471 (N_14471,N_13579,N_13722);
xor U14472 (N_14472,N_13919,N_13515);
nand U14473 (N_14473,N_13781,N_13859);
xor U14474 (N_14474,N_13659,N_13643);
xor U14475 (N_14475,N_13505,N_13877);
or U14476 (N_14476,N_13684,N_13572);
xor U14477 (N_14477,N_13863,N_13764);
nor U14478 (N_14478,N_13751,N_13707);
nor U14479 (N_14479,N_13634,N_13751);
nor U14480 (N_14480,N_13811,N_13917);
nand U14481 (N_14481,N_13626,N_13970);
and U14482 (N_14482,N_13709,N_13877);
nor U14483 (N_14483,N_13624,N_13555);
or U14484 (N_14484,N_13695,N_13859);
or U14485 (N_14485,N_13503,N_13703);
and U14486 (N_14486,N_13884,N_13650);
nor U14487 (N_14487,N_13608,N_13712);
xnor U14488 (N_14488,N_13811,N_13651);
or U14489 (N_14489,N_13707,N_13826);
nand U14490 (N_14490,N_13678,N_13841);
nor U14491 (N_14491,N_13714,N_13646);
nor U14492 (N_14492,N_13834,N_13715);
nor U14493 (N_14493,N_13682,N_13799);
and U14494 (N_14494,N_13630,N_13928);
and U14495 (N_14495,N_13565,N_13917);
or U14496 (N_14496,N_13898,N_13873);
nor U14497 (N_14497,N_13757,N_13505);
or U14498 (N_14498,N_13756,N_13732);
nand U14499 (N_14499,N_13526,N_13841);
xor U14500 (N_14500,N_14385,N_14279);
xor U14501 (N_14501,N_14335,N_14055);
xnor U14502 (N_14502,N_14021,N_14244);
nor U14503 (N_14503,N_14494,N_14280);
and U14504 (N_14504,N_14477,N_14082);
nor U14505 (N_14505,N_14475,N_14141);
nor U14506 (N_14506,N_14362,N_14234);
nand U14507 (N_14507,N_14427,N_14213);
nor U14508 (N_14508,N_14043,N_14194);
nor U14509 (N_14509,N_14386,N_14274);
xnor U14510 (N_14510,N_14446,N_14047);
or U14511 (N_14511,N_14139,N_14357);
nand U14512 (N_14512,N_14042,N_14358);
and U14513 (N_14513,N_14186,N_14014);
or U14514 (N_14514,N_14422,N_14191);
nor U14515 (N_14515,N_14078,N_14410);
nand U14516 (N_14516,N_14275,N_14440);
nor U14517 (N_14517,N_14005,N_14356);
nor U14518 (N_14518,N_14311,N_14355);
xnor U14519 (N_14519,N_14221,N_14322);
and U14520 (N_14520,N_14394,N_14432);
and U14521 (N_14521,N_14074,N_14188);
nor U14522 (N_14522,N_14392,N_14340);
or U14523 (N_14523,N_14418,N_14107);
or U14524 (N_14524,N_14415,N_14219);
or U14525 (N_14525,N_14041,N_14069);
nand U14526 (N_14526,N_14285,N_14384);
xor U14527 (N_14527,N_14298,N_14389);
nand U14528 (N_14528,N_14437,N_14169);
nand U14529 (N_14529,N_14129,N_14447);
and U14530 (N_14530,N_14474,N_14252);
or U14531 (N_14531,N_14250,N_14028);
xor U14532 (N_14532,N_14106,N_14488);
xnor U14533 (N_14533,N_14172,N_14202);
nand U14534 (N_14534,N_14443,N_14053);
nor U14535 (N_14535,N_14370,N_14148);
or U14536 (N_14536,N_14470,N_14299);
or U14537 (N_14537,N_14116,N_14154);
xor U14538 (N_14538,N_14426,N_14189);
nor U14539 (N_14539,N_14216,N_14227);
nor U14540 (N_14540,N_14282,N_14071);
or U14541 (N_14541,N_14400,N_14029);
nor U14542 (N_14542,N_14459,N_14336);
nand U14543 (N_14543,N_14088,N_14462);
and U14544 (N_14544,N_14246,N_14391);
or U14545 (N_14545,N_14050,N_14445);
nor U14546 (N_14546,N_14265,N_14425);
and U14547 (N_14547,N_14132,N_14058);
xnor U14548 (N_14548,N_14110,N_14038);
and U14549 (N_14549,N_14046,N_14348);
nand U14550 (N_14550,N_14395,N_14179);
and U14551 (N_14551,N_14196,N_14407);
or U14552 (N_14552,N_14433,N_14104);
nand U14553 (N_14553,N_14305,N_14127);
nor U14554 (N_14554,N_14167,N_14303);
xnor U14555 (N_14555,N_14192,N_14155);
and U14556 (N_14556,N_14093,N_14160);
nand U14557 (N_14557,N_14173,N_14396);
nand U14558 (N_14558,N_14486,N_14469);
nor U14559 (N_14559,N_14211,N_14487);
nor U14560 (N_14560,N_14214,N_14059);
and U14561 (N_14561,N_14151,N_14171);
and U14562 (N_14562,N_14091,N_14080);
nand U14563 (N_14563,N_14230,N_14268);
nor U14564 (N_14564,N_14312,N_14353);
nor U14565 (N_14565,N_14207,N_14119);
nand U14566 (N_14566,N_14347,N_14286);
and U14567 (N_14567,N_14332,N_14027);
or U14568 (N_14568,N_14452,N_14048);
nor U14569 (N_14569,N_14315,N_14424);
or U14570 (N_14570,N_14327,N_14181);
xor U14571 (N_14571,N_14263,N_14354);
nor U14572 (N_14572,N_14066,N_14455);
nor U14573 (N_14573,N_14254,N_14331);
and U14574 (N_14574,N_14460,N_14247);
nor U14575 (N_14575,N_14149,N_14086);
xnor U14576 (N_14576,N_14302,N_14098);
nor U14577 (N_14577,N_14032,N_14491);
nor U14578 (N_14578,N_14183,N_14320);
nor U14579 (N_14579,N_14372,N_14441);
and U14580 (N_14580,N_14077,N_14008);
nand U14581 (N_14581,N_14190,N_14031);
nand U14582 (N_14582,N_14283,N_14092);
xnor U14583 (N_14583,N_14476,N_14004);
nor U14584 (N_14584,N_14293,N_14136);
nand U14585 (N_14585,N_14444,N_14256);
nand U14586 (N_14586,N_14030,N_14481);
nand U14587 (N_14587,N_14325,N_14273);
and U14588 (N_14588,N_14065,N_14383);
xnor U14589 (N_14589,N_14212,N_14319);
xor U14590 (N_14590,N_14222,N_14430);
nor U14591 (N_14591,N_14420,N_14178);
nor U14592 (N_14592,N_14156,N_14090);
xor U14593 (N_14593,N_14024,N_14393);
and U14594 (N_14594,N_14133,N_14109);
nand U14595 (N_14595,N_14314,N_14350);
nand U14596 (N_14596,N_14084,N_14112);
nand U14597 (N_14597,N_14002,N_14471);
nand U14598 (N_14598,N_14295,N_14382);
nand U14599 (N_14599,N_14122,N_14316);
nand U14600 (N_14600,N_14208,N_14333);
nor U14601 (N_14601,N_14239,N_14158);
and U14602 (N_14602,N_14408,N_14342);
or U14603 (N_14603,N_14068,N_14205);
nand U14604 (N_14604,N_14210,N_14498);
xnor U14605 (N_14605,N_14397,N_14036);
or U14606 (N_14606,N_14180,N_14026);
or U14607 (N_14607,N_14419,N_14142);
or U14608 (N_14608,N_14060,N_14337);
nand U14609 (N_14609,N_14260,N_14379);
or U14610 (N_14610,N_14238,N_14094);
and U14611 (N_14611,N_14185,N_14233);
xnor U14612 (N_14612,N_14064,N_14095);
or U14613 (N_14613,N_14115,N_14170);
and U14614 (N_14614,N_14218,N_14224);
nand U14615 (N_14615,N_14496,N_14497);
or U14616 (N_14616,N_14016,N_14457);
nand U14617 (N_14617,N_14140,N_14478);
nand U14618 (N_14618,N_14304,N_14070);
nand U14619 (N_14619,N_14089,N_14429);
or U14620 (N_14620,N_14174,N_14226);
xnor U14621 (N_14621,N_14034,N_14329);
xor U14622 (N_14622,N_14468,N_14466);
nor U14623 (N_14623,N_14409,N_14241);
nand U14624 (N_14624,N_14007,N_14318);
or U14625 (N_14625,N_14037,N_14281);
and U14626 (N_14626,N_14472,N_14162);
nor U14627 (N_14627,N_14324,N_14063);
and U14628 (N_14628,N_14198,N_14414);
and U14629 (N_14629,N_14352,N_14017);
xor U14630 (N_14630,N_14204,N_14175);
xor U14631 (N_14631,N_14490,N_14360);
nand U14632 (N_14632,N_14144,N_14373);
xor U14633 (N_14633,N_14087,N_14366);
or U14634 (N_14634,N_14449,N_14482);
nor U14635 (N_14635,N_14334,N_14399);
nor U14636 (N_14636,N_14237,N_14276);
xnor U14637 (N_14637,N_14339,N_14495);
xor U14638 (N_14638,N_14294,N_14215);
nand U14639 (N_14639,N_14308,N_14165);
xnor U14640 (N_14640,N_14313,N_14269);
and U14641 (N_14641,N_14193,N_14448);
nand U14642 (N_14642,N_14292,N_14277);
nor U14643 (N_14643,N_14040,N_14184);
or U14644 (N_14644,N_14236,N_14376);
and U14645 (N_14645,N_14351,N_14417);
or U14646 (N_14646,N_14135,N_14010);
or U14647 (N_14647,N_14411,N_14051);
and U14648 (N_14648,N_14465,N_14442);
xnor U14649 (N_14649,N_14079,N_14012);
and U14650 (N_14650,N_14045,N_14461);
nor U14651 (N_14651,N_14159,N_14152);
xnor U14652 (N_14652,N_14330,N_14100);
and U14653 (N_14653,N_14272,N_14117);
xor U14654 (N_14654,N_14270,N_14105);
or U14655 (N_14655,N_14083,N_14401);
and U14656 (N_14656,N_14113,N_14343);
and U14657 (N_14657,N_14367,N_14365);
or U14658 (N_14658,N_14164,N_14076);
or U14659 (N_14659,N_14130,N_14242);
nand U14660 (N_14660,N_14439,N_14259);
nor U14661 (N_14661,N_14485,N_14266);
or U14662 (N_14662,N_14049,N_14387);
or U14663 (N_14663,N_14166,N_14232);
nor U14664 (N_14664,N_14229,N_14368);
or U14665 (N_14665,N_14006,N_14126);
xnor U14666 (N_14666,N_14288,N_14033);
and U14667 (N_14667,N_14450,N_14011);
or U14668 (N_14668,N_14398,N_14264);
or U14669 (N_14669,N_14454,N_14323);
nand U14670 (N_14670,N_14163,N_14145);
nor U14671 (N_14671,N_14072,N_14349);
or U14672 (N_14672,N_14492,N_14206);
nor U14673 (N_14673,N_14435,N_14085);
nor U14674 (N_14674,N_14103,N_14484);
or U14675 (N_14675,N_14489,N_14428);
and U14676 (N_14676,N_14378,N_14096);
xnor U14677 (N_14677,N_14346,N_14381);
and U14678 (N_14678,N_14168,N_14296);
nor U14679 (N_14679,N_14019,N_14153);
nor U14680 (N_14680,N_14035,N_14131);
nand U14681 (N_14681,N_14363,N_14257);
xor U14682 (N_14682,N_14251,N_14271);
nor U14683 (N_14683,N_14434,N_14297);
or U14684 (N_14684,N_14300,N_14483);
nand U14685 (N_14685,N_14499,N_14150);
and U14686 (N_14686,N_14310,N_14301);
or U14687 (N_14687,N_14118,N_14009);
nor U14688 (N_14688,N_14177,N_14328);
and U14689 (N_14689,N_14121,N_14000);
nand U14690 (N_14690,N_14405,N_14111);
and U14691 (N_14691,N_14464,N_14451);
or U14692 (N_14692,N_14431,N_14062);
and U14693 (N_14693,N_14138,N_14147);
nor U14694 (N_14694,N_14262,N_14480);
and U14695 (N_14695,N_14453,N_14013);
and U14696 (N_14696,N_14307,N_14228);
xor U14697 (N_14697,N_14404,N_14248);
or U14698 (N_14698,N_14120,N_14388);
xor U14699 (N_14699,N_14220,N_14493);
nand U14700 (N_14700,N_14341,N_14364);
xor U14701 (N_14701,N_14287,N_14161);
nor U14702 (N_14702,N_14406,N_14374);
nor U14703 (N_14703,N_14249,N_14436);
nand U14704 (N_14704,N_14197,N_14231);
or U14705 (N_14705,N_14317,N_14182);
nor U14706 (N_14706,N_14467,N_14416);
or U14707 (N_14707,N_14143,N_14423);
nand U14708 (N_14708,N_14099,N_14057);
or U14709 (N_14709,N_14023,N_14267);
and U14710 (N_14710,N_14201,N_14375);
nor U14711 (N_14711,N_14345,N_14081);
nand U14712 (N_14712,N_14235,N_14369);
or U14713 (N_14713,N_14052,N_14176);
xnor U14714 (N_14714,N_14458,N_14101);
xnor U14715 (N_14715,N_14245,N_14195);
xnor U14716 (N_14716,N_14015,N_14001);
xnor U14717 (N_14717,N_14371,N_14044);
xor U14718 (N_14718,N_14067,N_14438);
and U14719 (N_14719,N_14321,N_14217);
nor U14720 (N_14720,N_14003,N_14124);
nand U14721 (N_14721,N_14203,N_14413);
or U14722 (N_14722,N_14290,N_14309);
nand U14723 (N_14723,N_14018,N_14157);
nand U14724 (N_14724,N_14128,N_14403);
nand U14725 (N_14725,N_14056,N_14209);
xor U14726 (N_14726,N_14278,N_14097);
nor U14727 (N_14727,N_14025,N_14473);
or U14728 (N_14728,N_14338,N_14344);
nor U14729 (N_14729,N_14187,N_14075);
or U14730 (N_14730,N_14125,N_14061);
xor U14731 (N_14731,N_14102,N_14359);
nor U14732 (N_14732,N_14380,N_14253);
xor U14733 (N_14733,N_14306,N_14123);
or U14734 (N_14734,N_14421,N_14261);
nor U14735 (N_14735,N_14284,N_14020);
and U14736 (N_14736,N_14073,N_14326);
nand U14737 (N_14737,N_14361,N_14200);
nor U14738 (N_14738,N_14390,N_14108);
or U14739 (N_14739,N_14243,N_14225);
nand U14740 (N_14740,N_14240,N_14137);
nor U14741 (N_14741,N_14199,N_14377);
nand U14742 (N_14742,N_14289,N_14402);
and U14743 (N_14743,N_14039,N_14456);
nand U14744 (N_14744,N_14463,N_14134);
nand U14745 (N_14745,N_14114,N_14479);
or U14746 (N_14746,N_14258,N_14291);
nand U14747 (N_14747,N_14412,N_14146);
xnor U14748 (N_14748,N_14223,N_14022);
xnor U14749 (N_14749,N_14255,N_14054);
nand U14750 (N_14750,N_14201,N_14463);
xnor U14751 (N_14751,N_14400,N_14229);
xor U14752 (N_14752,N_14309,N_14464);
nor U14753 (N_14753,N_14307,N_14084);
nand U14754 (N_14754,N_14289,N_14407);
nand U14755 (N_14755,N_14158,N_14469);
or U14756 (N_14756,N_14078,N_14313);
nor U14757 (N_14757,N_14413,N_14162);
xnor U14758 (N_14758,N_14412,N_14495);
nor U14759 (N_14759,N_14105,N_14185);
and U14760 (N_14760,N_14311,N_14455);
nor U14761 (N_14761,N_14119,N_14263);
nor U14762 (N_14762,N_14233,N_14135);
or U14763 (N_14763,N_14143,N_14070);
nand U14764 (N_14764,N_14277,N_14446);
nand U14765 (N_14765,N_14032,N_14465);
nand U14766 (N_14766,N_14254,N_14001);
xnor U14767 (N_14767,N_14012,N_14483);
nand U14768 (N_14768,N_14057,N_14102);
nand U14769 (N_14769,N_14110,N_14216);
or U14770 (N_14770,N_14064,N_14112);
or U14771 (N_14771,N_14431,N_14171);
and U14772 (N_14772,N_14023,N_14461);
nor U14773 (N_14773,N_14220,N_14469);
and U14774 (N_14774,N_14462,N_14448);
xor U14775 (N_14775,N_14067,N_14418);
nor U14776 (N_14776,N_14284,N_14088);
xnor U14777 (N_14777,N_14001,N_14141);
nand U14778 (N_14778,N_14483,N_14158);
nand U14779 (N_14779,N_14122,N_14035);
nor U14780 (N_14780,N_14111,N_14150);
and U14781 (N_14781,N_14437,N_14338);
xnor U14782 (N_14782,N_14074,N_14456);
or U14783 (N_14783,N_14182,N_14295);
or U14784 (N_14784,N_14292,N_14246);
xor U14785 (N_14785,N_14010,N_14412);
xor U14786 (N_14786,N_14326,N_14397);
nor U14787 (N_14787,N_14280,N_14218);
nand U14788 (N_14788,N_14422,N_14146);
and U14789 (N_14789,N_14075,N_14292);
nand U14790 (N_14790,N_14338,N_14203);
nand U14791 (N_14791,N_14139,N_14133);
nand U14792 (N_14792,N_14320,N_14473);
nor U14793 (N_14793,N_14055,N_14131);
or U14794 (N_14794,N_14146,N_14339);
and U14795 (N_14795,N_14494,N_14224);
xor U14796 (N_14796,N_14230,N_14248);
and U14797 (N_14797,N_14490,N_14208);
xor U14798 (N_14798,N_14468,N_14062);
and U14799 (N_14799,N_14223,N_14455);
nand U14800 (N_14800,N_14106,N_14093);
nor U14801 (N_14801,N_14037,N_14109);
xor U14802 (N_14802,N_14169,N_14301);
or U14803 (N_14803,N_14183,N_14327);
and U14804 (N_14804,N_14471,N_14039);
or U14805 (N_14805,N_14351,N_14487);
xnor U14806 (N_14806,N_14119,N_14215);
or U14807 (N_14807,N_14362,N_14466);
and U14808 (N_14808,N_14090,N_14497);
nor U14809 (N_14809,N_14487,N_14486);
or U14810 (N_14810,N_14268,N_14169);
xnor U14811 (N_14811,N_14229,N_14304);
nand U14812 (N_14812,N_14457,N_14129);
or U14813 (N_14813,N_14376,N_14252);
nor U14814 (N_14814,N_14041,N_14321);
or U14815 (N_14815,N_14498,N_14365);
or U14816 (N_14816,N_14144,N_14345);
or U14817 (N_14817,N_14365,N_14366);
or U14818 (N_14818,N_14213,N_14109);
xnor U14819 (N_14819,N_14147,N_14142);
nor U14820 (N_14820,N_14231,N_14301);
nand U14821 (N_14821,N_14459,N_14072);
or U14822 (N_14822,N_14010,N_14005);
nand U14823 (N_14823,N_14022,N_14384);
nand U14824 (N_14824,N_14034,N_14448);
and U14825 (N_14825,N_14216,N_14340);
nor U14826 (N_14826,N_14401,N_14210);
nand U14827 (N_14827,N_14164,N_14131);
or U14828 (N_14828,N_14073,N_14249);
or U14829 (N_14829,N_14445,N_14173);
nand U14830 (N_14830,N_14066,N_14281);
nor U14831 (N_14831,N_14151,N_14160);
nor U14832 (N_14832,N_14021,N_14103);
and U14833 (N_14833,N_14475,N_14399);
or U14834 (N_14834,N_14176,N_14151);
nor U14835 (N_14835,N_14453,N_14298);
and U14836 (N_14836,N_14110,N_14046);
or U14837 (N_14837,N_14271,N_14234);
or U14838 (N_14838,N_14259,N_14002);
nor U14839 (N_14839,N_14233,N_14268);
and U14840 (N_14840,N_14286,N_14231);
xor U14841 (N_14841,N_14171,N_14350);
and U14842 (N_14842,N_14030,N_14284);
xor U14843 (N_14843,N_14171,N_14283);
and U14844 (N_14844,N_14223,N_14233);
xnor U14845 (N_14845,N_14440,N_14128);
xor U14846 (N_14846,N_14287,N_14061);
or U14847 (N_14847,N_14368,N_14344);
xor U14848 (N_14848,N_14141,N_14026);
and U14849 (N_14849,N_14097,N_14435);
or U14850 (N_14850,N_14018,N_14076);
nand U14851 (N_14851,N_14348,N_14171);
and U14852 (N_14852,N_14116,N_14482);
nor U14853 (N_14853,N_14162,N_14051);
xor U14854 (N_14854,N_14030,N_14172);
nor U14855 (N_14855,N_14487,N_14004);
nand U14856 (N_14856,N_14010,N_14123);
nor U14857 (N_14857,N_14242,N_14139);
or U14858 (N_14858,N_14399,N_14466);
xnor U14859 (N_14859,N_14312,N_14088);
or U14860 (N_14860,N_14146,N_14417);
and U14861 (N_14861,N_14369,N_14175);
nor U14862 (N_14862,N_14417,N_14422);
nand U14863 (N_14863,N_14077,N_14060);
and U14864 (N_14864,N_14166,N_14366);
nor U14865 (N_14865,N_14485,N_14103);
and U14866 (N_14866,N_14194,N_14054);
nor U14867 (N_14867,N_14371,N_14376);
nand U14868 (N_14868,N_14327,N_14326);
nor U14869 (N_14869,N_14311,N_14031);
or U14870 (N_14870,N_14126,N_14389);
nor U14871 (N_14871,N_14340,N_14123);
or U14872 (N_14872,N_14168,N_14498);
xnor U14873 (N_14873,N_14358,N_14127);
nor U14874 (N_14874,N_14137,N_14180);
and U14875 (N_14875,N_14124,N_14427);
xor U14876 (N_14876,N_14101,N_14336);
nor U14877 (N_14877,N_14050,N_14286);
nand U14878 (N_14878,N_14314,N_14187);
nor U14879 (N_14879,N_14111,N_14283);
and U14880 (N_14880,N_14033,N_14486);
or U14881 (N_14881,N_14336,N_14008);
nand U14882 (N_14882,N_14029,N_14085);
xnor U14883 (N_14883,N_14128,N_14489);
nor U14884 (N_14884,N_14011,N_14453);
and U14885 (N_14885,N_14242,N_14352);
and U14886 (N_14886,N_14412,N_14370);
and U14887 (N_14887,N_14189,N_14293);
and U14888 (N_14888,N_14329,N_14318);
and U14889 (N_14889,N_14240,N_14296);
xnor U14890 (N_14890,N_14351,N_14211);
nand U14891 (N_14891,N_14107,N_14448);
or U14892 (N_14892,N_14073,N_14295);
nand U14893 (N_14893,N_14013,N_14149);
xnor U14894 (N_14894,N_14357,N_14000);
and U14895 (N_14895,N_14215,N_14444);
nor U14896 (N_14896,N_14011,N_14411);
nor U14897 (N_14897,N_14292,N_14309);
nand U14898 (N_14898,N_14181,N_14342);
or U14899 (N_14899,N_14079,N_14084);
nand U14900 (N_14900,N_14249,N_14067);
or U14901 (N_14901,N_14158,N_14139);
or U14902 (N_14902,N_14063,N_14499);
nor U14903 (N_14903,N_14342,N_14410);
or U14904 (N_14904,N_14493,N_14307);
nor U14905 (N_14905,N_14180,N_14431);
or U14906 (N_14906,N_14130,N_14412);
or U14907 (N_14907,N_14274,N_14313);
xor U14908 (N_14908,N_14325,N_14102);
nor U14909 (N_14909,N_14311,N_14454);
and U14910 (N_14910,N_14383,N_14494);
and U14911 (N_14911,N_14388,N_14170);
nor U14912 (N_14912,N_14036,N_14268);
nor U14913 (N_14913,N_14246,N_14259);
and U14914 (N_14914,N_14369,N_14196);
nor U14915 (N_14915,N_14384,N_14386);
nand U14916 (N_14916,N_14329,N_14040);
nand U14917 (N_14917,N_14357,N_14197);
xnor U14918 (N_14918,N_14359,N_14320);
and U14919 (N_14919,N_14481,N_14156);
nand U14920 (N_14920,N_14241,N_14325);
nor U14921 (N_14921,N_14316,N_14136);
or U14922 (N_14922,N_14379,N_14070);
and U14923 (N_14923,N_14132,N_14067);
and U14924 (N_14924,N_14344,N_14372);
xnor U14925 (N_14925,N_14446,N_14034);
nand U14926 (N_14926,N_14354,N_14465);
nand U14927 (N_14927,N_14244,N_14163);
nor U14928 (N_14928,N_14189,N_14188);
or U14929 (N_14929,N_14235,N_14413);
nor U14930 (N_14930,N_14333,N_14292);
and U14931 (N_14931,N_14246,N_14194);
or U14932 (N_14932,N_14342,N_14182);
nand U14933 (N_14933,N_14234,N_14169);
nor U14934 (N_14934,N_14314,N_14183);
nand U14935 (N_14935,N_14305,N_14078);
nand U14936 (N_14936,N_14375,N_14226);
xor U14937 (N_14937,N_14012,N_14451);
nor U14938 (N_14938,N_14065,N_14424);
and U14939 (N_14939,N_14312,N_14243);
xnor U14940 (N_14940,N_14430,N_14354);
nor U14941 (N_14941,N_14155,N_14467);
nand U14942 (N_14942,N_14339,N_14112);
xor U14943 (N_14943,N_14393,N_14049);
nor U14944 (N_14944,N_14421,N_14355);
or U14945 (N_14945,N_14116,N_14129);
and U14946 (N_14946,N_14328,N_14341);
or U14947 (N_14947,N_14001,N_14026);
nor U14948 (N_14948,N_14411,N_14029);
xnor U14949 (N_14949,N_14041,N_14317);
xor U14950 (N_14950,N_14039,N_14360);
and U14951 (N_14951,N_14094,N_14249);
and U14952 (N_14952,N_14108,N_14469);
and U14953 (N_14953,N_14431,N_14101);
xor U14954 (N_14954,N_14373,N_14075);
or U14955 (N_14955,N_14066,N_14209);
nand U14956 (N_14956,N_14335,N_14428);
or U14957 (N_14957,N_14373,N_14099);
xnor U14958 (N_14958,N_14031,N_14310);
xnor U14959 (N_14959,N_14496,N_14442);
nand U14960 (N_14960,N_14278,N_14258);
or U14961 (N_14961,N_14375,N_14156);
or U14962 (N_14962,N_14131,N_14388);
nand U14963 (N_14963,N_14456,N_14453);
nand U14964 (N_14964,N_14422,N_14088);
xnor U14965 (N_14965,N_14465,N_14224);
nand U14966 (N_14966,N_14409,N_14021);
and U14967 (N_14967,N_14423,N_14285);
nand U14968 (N_14968,N_14401,N_14441);
nand U14969 (N_14969,N_14063,N_14211);
xor U14970 (N_14970,N_14281,N_14039);
xor U14971 (N_14971,N_14284,N_14469);
nor U14972 (N_14972,N_14024,N_14451);
or U14973 (N_14973,N_14275,N_14050);
nor U14974 (N_14974,N_14428,N_14474);
nor U14975 (N_14975,N_14193,N_14408);
and U14976 (N_14976,N_14191,N_14199);
xnor U14977 (N_14977,N_14474,N_14355);
or U14978 (N_14978,N_14481,N_14307);
or U14979 (N_14979,N_14377,N_14234);
nor U14980 (N_14980,N_14393,N_14337);
or U14981 (N_14981,N_14229,N_14253);
or U14982 (N_14982,N_14128,N_14300);
and U14983 (N_14983,N_14493,N_14249);
xnor U14984 (N_14984,N_14312,N_14473);
nand U14985 (N_14985,N_14386,N_14452);
xnor U14986 (N_14986,N_14406,N_14315);
and U14987 (N_14987,N_14365,N_14396);
or U14988 (N_14988,N_14063,N_14040);
nor U14989 (N_14989,N_14474,N_14360);
nand U14990 (N_14990,N_14139,N_14022);
or U14991 (N_14991,N_14293,N_14215);
or U14992 (N_14992,N_14475,N_14055);
and U14993 (N_14993,N_14245,N_14194);
nor U14994 (N_14994,N_14489,N_14038);
or U14995 (N_14995,N_14369,N_14421);
xnor U14996 (N_14996,N_14492,N_14185);
nand U14997 (N_14997,N_14132,N_14415);
xnor U14998 (N_14998,N_14225,N_14407);
nor U14999 (N_14999,N_14256,N_14198);
nand U15000 (N_15000,N_14847,N_14520);
nor U15001 (N_15001,N_14774,N_14818);
xor U15002 (N_15002,N_14738,N_14801);
xnor U15003 (N_15003,N_14620,N_14536);
xnor U15004 (N_15004,N_14976,N_14752);
xnor U15005 (N_15005,N_14585,N_14532);
xor U15006 (N_15006,N_14566,N_14875);
nand U15007 (N_15007,N_14761,N_14972);
nor U15008 (N_15008,N_14727,N_14991);
or U15009 (N_15009,N_14882,N_14552);
or U15010 (N_15010,N_14958,N_14911);
nor U15011 (N_15011,N_14680,N_14628);
nor U15012 (N_15012,N_14903,N_14515);
or U15013 (N_15013,N_14866,N_14583);
xnor U15014 (N_15014,N_14514,N_14768);
or U15015 (N_15015,N_14833,N_14975);
and U15016 (N_15016,N_14723,N_14849);
xor U15017 (N_15017,N_14516,N_14988);
or U15018 (N_15018,N_14509,N_14770);
nand U15019 (N_15019,N_14984,N_14610);
nand U15020 (N_15020,N_14923,N_14661);
nor U15021 (N_15021,N_14720,N_14672);
xor U15022 (N_15022,N_14852,N_14901);
and U15023 (N_15023,N_14960,N_14985);
xnor U15024 (N_15024,N_14600,N_14513);
xor U15025 (N_15025,N_14564,N_14613);
or U15026 (N_15026,N_14677,N_14538);
xor U15027 (N_15027,N_14953,N_14734);
nand U15028 (N_15028,N_14848,N_14922);
or U15029 (N_15029,N_14948,N_14612);
or U15030 (N_15030,N_14679,N_14952);
or U15031 (N_15031,N_14713,N_14842);
and U15032 (N_15032,N_14967,N_14799);
xor U15033 (N_15033,N_14886,N_14640);
and U15034 (N_15034,N_14835,N_14789);
nand U15035 (N_15035,N_14518,N_14887);
nand U15036 (N_15036,N_14986,N_14557);
and U15037 (N_15037,N_14556,N_14962);
and U15038 (N_15038,N_14646,N_14559);
or U15039 (N_15039,N_14541,N_14681);
xor U15040 (N_15040,N_14558,N_14531);
and U15041 (N_15041,N_14622,N_14634);
xnor U15042 (N_15042,N_14618,N_14917);
nor U15043 (N_15043,N_14696,N_14832);
or U15044 (N_15044,N_14932,N_14584);
or U15045 (N_15045,N_14678,N_14741);
and U15046 (N_15046,N_14873,N_14826);
or U15047 (N_15047,N_14876,N_14760);
nand U15048 (N_15048,N_14843,N_14632);
nand U15049 (N_15049,N_14937,N_14624);
nor U15050 (N_15050,N_14715,N_14825);
and U15051 (N_15051,N_14753,N_14820);
nand U15052 (N_15052,N_14663,N_14782);
nand U15053 (N_15053,N_14800,N_14551);
nor U15054 (N_15054,N_14872,N_14983);
nand U15055 (N_15055,N_14756,N_14511);
xnor U15056 (N_15056,N_14915,N_14951);
and U15057 (N_15057,N_14987,N_14897);
nand U15058 (N_15058,N_14945,N_14969);
nor U15059 (N_15059,N_14805,N_14865);
xor U15060 (N_15060,N_14750,N_14858);
xor U15061 (N_15061,N_14777,N_14808);
or U15062 (N_15062,N_14891,N_14638);
nor U15063 (N_15063,N_14929,N_14596);
or U15064 (N_15064,N_14836,N_14525);
or U15065 (N_15065,N_14565,N_14829);
or U15066 (N_15066,N_14528,N_14908);
and U15067 (N_15067,N_14587,N_14502);
and U15068 (N_15068,N_14659,N_14586);
nor U15069 (N_15069,N_14979,N_14883);
or U15070 (N_15070,N_14579,N_14535);
xor U15071 (N_15071,N_14605,N_14899);
or U15072 (N_15072,N_14860,N_14523);
and U15073 (N_15073,N_14740,N_14783);
nor U15074 (N_15074,N_14767,N_14582);
xor U15075 (N_15075,N_14621,N_14550);
or U15076 (N_15076,N_14614,N_14617);
xor U15077 (N_15077,N_14936,N_14772);
nor U15078 (N_15078,N_14717,N_14912);
nand U15079 (N_15079,N_14731,N_14700);
nand U15080 (N_15080,N_14934,N_14977);
xnor U15081 (N_15081,N_14931,N_14567);
nor U15082 (N_15082,N_14542,N_14841);
nor U15083 (N_15083,N_14803,N_14796);
and U15084 (N_15084,N_14759,N_14868);
or U15085 (N_15085,N_14593,N_14939);
and U15086 (N_15086,N_14812,N_14963);
xor U15087 (N_15087,N_14773,N_14674);
and U15088 (N_15088,N_14650,N_14645);
nor U15089 (N_15089,N_14685,N_14971);
or U15090 (N_15090,N_14973,N_14561);
nand U15091 (N_15091,N_14942,N_14735);
or U15092 (N_15092,N_14522,N_14993);
nand U15093 (N_15093,N_14869,N_14616);
nand U15094 (N_15094,N_14683,N_14743);
xnor U15095 (N_15095,N_14530,N_14888);
or U15096 (N_15096,N_14629,N_14545);
nand U15097 (N_15097,N_14742,N_14930);
xor U15098 (N_15098,N_14637,N_14701);
or U15099 (N_15099,N_14797,N_14606);
or U15100 (N_15100,N_14780,N_14980);
xor U15101 (N_15101,N_14935,N_14904);
nor U15102 (N_15102,N_14881,N_14840);
nor U15103 (N_15103,N_14537,N_14609);
or U15104 (N_15104,N_14686,N_14862);
and U15105 (N_15105,N_14655,N_14781);
nor U15106 (N_15106,N_14729,N_14652);
or U15107 (N_15107,N_14784,N_14776);
nor U15108 (N_15108,N_14692,N_14851);
or U15109 (N_15109,N_14505,N_14611);
xor U15110 (N_15110,N_14974,N_14944);
nor U15111 (N_15111,N_14758,N_14878);
nand U15112 (N_15112,N_14687,N_14806);
nand U15113 (N_15113,N_14795,N_14615);
or U15114 (N_15114,N_14941,N_14732);
and U15115 (N_15115,N_14570,N_14682);
nand U15116 (N_15116,N_14906,N_14639);
nand U15117 (N_15117,N_14867,N_14595);
and U15118 (N_15118,N_14625,N_14990);
and U15119 (N_15119,N_14746,N_14562);
and U15120 (N_15120,N_14745,N_14785);
nor U15121 (N_15121,N_14938,N_14708);
and U15122 (N_15122,N_14588,N_14668);
nand U15123 (N_15123,N_14943,N_14691);
and U15124 (N_15124,N_14627,N_14804);
nand U15125 (N_15125,N_14658,N_14712);
nand U15126 (N_15126,N_14794,N_14718);
nor U15127 (N_15127,N_14744,N_14693);
nand U15128 (N_15128,N_14819,N_14527);
xnor U15129 (N_15129,N_14589,N_14788);
xnor U15130 (N_15130,N_14762,N_14554);
and U15131 (N_15131,N_14529,N_14714);
nor U15132 (N_15132,N_14572,N_14998);
nor U15133 (N_15133,N_14790,N_14707);
nand U15134 (N_15134,N_14910,N_14623);
and U15135 (N_15135,N_14907,N_14747);
or U15136 (N_15136,N_14954,N_14893);
xor U15137 (N_15137,N_14940,N_14706);
nor U15138 (N_15138,N_14563,N_14709);
and U15139 (N_15139,N_14560,N_14539);
and U15140 (N_15140,N_14534,N_14657);
xnor U15141 (N_15141,N_14766,N_14879);
xor U15142 (N_15142,N_14870,N_14997);
and U15143 (N_15143,N_14857,N_14863);
and U15144 (N_15144,N_14591,N_14900);
nand U15145 (N_15145,N_14855,N_14555);
nand U15146 (N_15146,N_14633,N_14880);
or U15147 (N_15147,N_14512,N_14504);
nor U15148 (N_15148,N_14599,N_14684);
nand U15149 (N_15149,N_14636,N_14690);
or U15150 (N_15150,N_14946,N_14607);
or U15151 (N_15151,N_14547,N_14793);
xnor U15152 (N_15152,N_14726,N_14540);
nor U15153 (N_15153,N_14549,N_14918);
nand U15154 (N_15154,N_14665,N_14892);
nand U15155 (N_15155,N_14884,N_14926);
and U15156 (N_15156,N_14838,N_14533);
and U15157 (N_15157,N_14778,N_14861);
and U15158 (N_15158,N_14925,N_14856);
nand U15159 (N_15159,N_14755,N_14978);
nand U15160 (N_15160,N_14814,N_14846);
and U15161 (N_15161,N_14576,N_14698);
nor U15162 (N_15162,N_14653,N_14924);
and U15163 (N_15163,N_14581,N_14921);
xor U15164 (N_15164,N_14811,N_14580);
nand U15165 (N_15165,N_14575,N_14916);
xnor U15166 (N_15166,N_14786,N_14689);
and U15167 (N_15167,N_14568,N_14823);
nand U15168 (N_15168,N_14630,N_14982);
nor U15169 (N_15169,N_14577,N_14676);
xor U15170 (N_15170,N_14928,N_14635);
or U15171 (N_15171,N_14601,N_14524);
or U15172 (N_15172,N_14810,N_14598);
and U15173 (N_15173,N_14724,N_14507);
nand U15174 (N_15174,N_14837,N_14736);
or U15175 (N_15175,N_14737,N_14748);
nand U15176 (N_15176,N_14779,N_14824);
nand U15177 (N_15177,N_14574,N_14864);
or U15178 (N_15178,N_14839,N_14992);
xnor U15179 (N_15179,N_14673,N_14604);
xnor U15180 (N_15180,N_14895,N_14671);
nand U15181 (N_15181,N_14807,N_14754);
xnor U15182 (N_15182,N_14519,N_14651);
xor U15183 (N_15183,N_14765,N_14571);
or U15184 (N_15184,N_14521,N_14647);
xor U15185 (N_15185,N_14827,N_14961);
nand U15186 (N_15186,N_14970,N_14553);
nor U15187 (N_15187,N_14702,N_14592);
xor U15188 (N_15188,N_14859,N_14821);
xor U15189 (N_15189,N_14902,N_14695);
nor U15190 (N_15190,N_14844,N_14816);
xor U15191 (N_15191,N_14989,N_14894);
and U15192 (N_15192,N_14517,N_14968);
xnor U15193 (N_15193,N_14699,N_14578);
nor U15194 (N_15194,N_14890,N_14500);
and U15195 (N_15195,N_14947,N_14898);
xnor U15196 (N_15196,N_14526,N_14830);
nand U15197 (N_15197,N_14933,N_14644);
nor U15198 (N_15198,N_14854,N_14619);
nor U15199 (N_15199,N_14641,N_14791);
or U15200 (N_15200,N_14764,N_14956);
nor U15201 (N_15201,N_14763,N_14710);
and U15202 (N_15202,N_14669,N_14809);
xnor U15203 (N_15203,N_14733,N_14802);
xor U15204 (N_15204,N_14503,N_14728);
xnor U15205 (N_15205,N_14909,N_14817);
or U15206 (N_15206,N_14959,N_14654);
nand U15207 (N_15207,N_14667,N_14965);
xor U15208 (N_15208,N_14688,N_14649);
xnor U15209 (N_15209,N_14508,N_14853);
nand U15210 (N_15210,N_14885,N_14546);
or U15211 (N_15211,N_14642,N_14608);
or U15212 (N_15212,N_14874,N_14749);
nor U15213 (N_15213,N_14845,N_14771);
xnor U15214 (N_15214,N_14602,N_14999);
xor U15215 (N_15215,N_14662,N_14792);
nor U15216 (N_15216,N_14828,N_14834);
or U15217 (N_15217,N_14711,N_14927);
xor U15218 (N_15218,N_14914,N_14995);
and U15219 (N_15219,N_14751,N_14590);
xnor U15220 (N_15220,N_14648,N_14798);
nor U15221 (N_15221,N_14955,N_14739);
xor U15222 (N_15222,N_14594,N_14725);
xnor U15223 (N_15223,N_14775,N_14660);
or U15224 (N_15224,N_14719,N_14569);
nor U15225 (N_15225,N_14670,N_14787);
nand U15226 (N_15226,N_14905,N_14822);
nor U15227 (N_15227,N_14543,N_14631);
nor U15228 (N_15228,N_14544,N_14573);
xor U15229 (N_15229,N_14831,N_14694);
and U15230 (N_15230,N_14994,N_14964);
xnor U15231 (N_15231,N_14769,N_14548);
and U15232 (N_15232,N_14697,N_14981);
or U15233 (N_15233,N_14603,N_14815);
nand U15234 (N_15234,N_14716,N_14626);
xnor U15235 (N_15235,N_14919,N_14813);
and U15236 (N_15236,N_14877,N_14913);
or U15237 (N_15237,N_14643,N_14957);
and U15238 (N_15238,N_14889,N_14704);
or U15239 (N_15239,N_14675,N_14506);
and U15240 (N_15240,N_14896,N_14703);
xnor U15241 (N_15241,N_14757,N_14666);
and U15242 (N_15242,N_14597,N_14664);
or U15243 (N_15243,N_14705,N_14730);
xor U15244 (N_15244,N_14722,N_14949);
or U15245 (N_15245,N_14721,N_14510);
and U15246 (N_15246,N_14501,N_14920);
nand U15247 (N_15247,N_14950,N_14656);
and U15248 (N_15248,N_14850,N_14871);
or U15249 (N_15249,N_14966,N_14996);
or U15250 (N_15250,N_14719,N_14759);
xor U15251 (N_15251,N_14853,N_14554);
nand U15252 (N_15252,N_14850,N_14686);
and U15253 (N_15253,N_14636,N_14738);
xnor U15254 (N_15254,N_14622,N_14928);
xor U15255 (N_15255,N_14536,N_14871);
nor U15256 (N_15256,N_14652,N_14942);
nor U15257 (N_15257,N_14591,N_14984);
and U15258 (N_15258,N_14660,N_14590);
nor U15259 (N_15259,N_14792,N_14530);
nor U15260 (N_15260,N_14971,N_14836);
and U15261 (N_15261,N_14644,N_14842);
xnor U15262 (N_15262,N_14801,N_14722);
nor U15263 (N_15263,N_14937,N_14871);
nor U15264 (N_15264,N_14548,N_14748);
nand U15265 (N_15265,N_14739,N_14856);
and U15266 (N_15266,N_14641,N_14735);
nand U15267 (N_15267,N_14860,N_14557);
xor U15268 (N_15268,N_14600,N_14876);
and U15269 (N_15269,N_14910,N_14875);
or U15270 (N_15270,N_14528,N_14898);
nor U15271 (N_15271,N_14855,N_14523);
nor U15272 (N_15272,N_14787,N_14614);
and U15273 (N_15273,N_14801,N_14576);
nand U15274 (N_15274,N_14859,N_14512);
xor U15275 (N_15275,N_14876,N_14738);
or U15276 (N_15276,N_14550,N_14755);
nor U15277 (N_15277,N_14828,N_14763);
nor U15278 (N_15278,N_14567,N_14727);
and U15279 (N_15279,N_14905,N_14503);
xnor U15280 (N_15280,N_14776,N_14561);
nand U15281 (N_15281,N_14834,N_14607);
nand U15282 (N_15282,N_14742,N_14780);
xnor U15283 (N_15283,N_14739,N_14591);
nand U15284 (N_15284,N_14663,N_14690);
or U15285 (N_15285,N_14791,N_14805);
nand U15286 (N_15286,N_14794,N_14575);
and U15287 (N_15287,N_14860,N_14623);
or U15288 (N_15288,N_14871,N_14861);
or U15289 (N_15289,N_14876,N_14837);
nand U15290 (N_15290,N_14538,N_14582);
or U15291 (N_15291,N_14837,N_14500);
nor U15292 (N_15292,N_14872,N_14609);
xor U15293 (N_15293,N_14530,N_14716);
or U15294 (N_15294,N_14642,N_14606);
xnor U15295 (N_15295,N_14644,N_14646);
nand U15296 (N_15296,N_14598,N_14893);
xor U15297 (N_15297,N_14504,N_14550);
and U15298 (N_15298,N_14512,N_14913);
nand U15299 (N_15299,N_14753,N_14794);
nand U15300 (N_15300,N_14519,N_14807);
and U15301 (N_15301,N_14516,N_14964);
nor U15302 (N_15302,N_14642,N_14660);
or U15303 (N_15303,N_14664,N_14523);
nor U15304 (N_15304,N_14798,N_14654);
nor U15305 (N_15305,N_14623,N_14931);
or U15306 (N_15306,N_14767,N_14627);
and U15307 (N_15307,N_14979,N_14650);
or U15308 (N_15308,N_14736,N_14841);
nor U15309 (N_15309,N_14969,N_14812);
and U15310 (N_15310,N_14694,N_14548);
nand U15311 (N_15311,N_14798,N_14628);
or U15312 (N_15312,N_14535,N_14558);
nand U15313 (N_15313,N_14869,N_14737);
nor U15314 (N_15314,N_14636,N_14699);
or U15315 (N_15315,N_14665,N_14887);
nand U15316 (N_15316,N_14651,N_14510);
or U15317 (N_15317,N_14704,N_14951);
and U15318 (N_15318,N_14597,N_14790);
nor U15319 (N_15319,N_14688,N_14548);
nand U15320 (N_15320,N_14740,N_14512);
and U15321 (N_15321,N_14776,N_14984);
nand U15322 (N_15322,N_14575,N_14572);
and U15323 (N_15323,N_14662,N_14921);
nor U15324 (N_15324,N_14981,N_14769);
or U15325 (N_15325,N_14982,N_14799);
nor U15326 (N_15326,N_14778,N_14865);
nor U15327 (N_15327,N_14842,N_14538);
and U15328 (N_15328,N_14881,N_14891);
nand U15329 (N_15329,N_14824,N_14913);
and U15330 (N_15330,N_14928,N_14744);
xor U15331 (N_15331,N_14868,N_14973);
xor U15332 (N_15332,N_14517,N_14619);
and U15333 (N_15333,N_14941,N_14713);
xor U15334 (N_15334,N_14554,N_14815);
and U15335 (N_15335,N_14876,N_14970);
or U15336 (N_15336,N_14976,N_14918);
and U15337 (N_15337,N_14729,N_14681);
xor U15338 (N_15338,N_14711,N_14836);
xnor U15339 (N_15339,N_14838,N_14639);
nand U15340 (N_15340,N_14534,N_14582);
nor U15341 (N_15341,N_14842,N_14861);
nor U15342 (N_15342,N_14869,N_14893);
xor U15343 (N_15343,N_14962,N_14938);
and U15344 (N_15344,N_14541,N_14693);
and U15345 (N_15345,N_14521,N_14708);
nand U15346 (N_15346,N_14740,N_14638);
nand U15347 (N_15347,N_14908,N_14704);
nor U15348 (N_15348,N_14909,N_14826);
nor U15349 (N_15349,N_14691,N_14706);
nor U15350 (N_15350,N_14581,N_14514);
nand U15351 (N_15351,N_14726,N_14531);
or U15352 (N_15352,N_14715,N_14724);
xor U15353 (N_15353,N_14906,N_14526);
nand U15354 (N_15354,N_14865,N_14590);
or U15355 (N_15355,N_14677,N_14759);
and U15356 (N_15356,N_14628,N_14544);
or U15357 (N_15357,N_14687,N_14500);
and U15358 (N_15358,N_14971,N_14616);
and U15359 (N_15359,N_14760,N_14761);
and U15360 (N_15360,N_14841,N_14843);
nor U15361 (N_15361,N_14823,N_14911);
xor U15362 (N_15362,N_14600,N_14827);
xnor U15363 (N_15363,N_14958,N_14570);
xnor U15364 (N_15364,N_14502,N_14641);
or U15365 (N_15365,N_14870,N_14945);
nand U15366 (N_15366,N_14885,N_14791);
and U15367 (N_15367,N_14752,N_14779);
or U15368 (N_15368,N_14763,N_14509);
and U15369 (N_15369,N_14590,N_14762);
and U15370 (N_15370,N_14622,N_14602);
nor U15371 (N_15371,N_14978,N_14721);
nor U15372 (N_15372,N_14822,N_14974);
nor U15373 (N_15373,N_14896,N_14927);
or U15374 (N_15374,N_14958,N_14753);
nand U15375 (N_15375,N_14511,N_14753);
nand U15376 (N_15376,N_14837,N_14516);
or U15377 (N_15377,N_14611,N_14875);
nand U15378 (N_15378,N_14594,N_14616);
nor U15379 (N_15379,N_14529,N_14722);
and U15380 (N_15380,N_14767,N_14975);
nor U15381 (N_15381,N_14739,N_14665);
and U15382 (N_15382,N_14582,N_14725);
xnor U15383 (N_15383,N_14725,N_14939);
xnor U15384 (N_15384,N_14642,N_14941);
nand U15385 (N_15385,N_14900,N_14963);
nor U15386 (N_15386,N_14609,N_14974);
nor U15387 (N_15387,N_14960,N_14768);
nor U15388 (N_15388,N_14786,N_14971);
xor U15389 (N_15389,N_14638,N_14544);
or U15390 (N_15390,N_14562,N_14502);
and U15391 (N_15391,N_14855,N_14603);
and U15392 (N_15392,N_14888,N_14680);
nor U15393 (N_15393,N_14605,N_14856);
nand U15394 (N_15394,N_14876,N_14866);
and U15395 (N_15395,N_14555,N_14571);
and U15396 (N_15396,N_14611,N_14936);
nor U15397 (N_15397,N_14648,N_14962);
or U15398 (N_15398,N_14756,N_14643);
nor U15399 (N_15399,N_14846,N_14796);
nand U15400 (N_15400,N_14978,N_14797);
and U15401 (N_15401,N_14755,N_14955);
nor U15402 (N_15402,N_14805,N_14807);
nand U15403 (N_15403,N_14759,N_14756);
or U15404 (N_15404,N_14876,N_14617);
nor U15405 (N_15405,N_14689,N_14528);
nor U15406 (N_15406,N_14536,N_14578);
nand U15407 (N_15407,N_14626,N_14603);
xnor U15408 (N_15408,N_14996,N_14527);
and U15409 (N_15409,N_14705,N_14651);
nor U15410 (N_15410,N_14860,N_14574);
xnor U15411 (N_15411,N_14922,N_14983);
nand U15412 (N_15412,N_14798,N_14881);
xnor U15413 (N_15413,N_14958,N_14679);
and U15414 (N_15414,N_14725,N_14600);
or U15415 (N_15415,N_14597,N_14949);
and U15416 (N_15416,N_14746,N_14773);
and U15417 (N_15417,N_14966,N_14989);
or U15418 (N_15418,N_14715,N_14543);
nor U15419 (N_15419,N_14753,N_14670);
and U15420 (N_15420,N_14836,N_14699);
nor U15421 (N_15421,N_14917,N_14798);
nand U15422 (N_15422,N_14671,N_14561);
and U15423 (N_15423,N_14774,N_14725);
nand U15424 (N_15424,N_14640,N_14713);
nor U15425 (N_15425,N_14631,N_14839);
nand U15426 (N_15426,N_14669,N_14543);
xnor U15427 (N_15427,N_14561,N_14749);
nand U15428 (N_15428,N_14515,N_14748);
or U15429 (N_15429,N_14577,N_14959);
nor U15430 (N_15430,N_14502,N_14521);
or U15431 (N_15431,N_14685,N_14740);
and U15432 (N_15432,N_14607,N_14850);
nand U15433 (N_15433,N_14776,N_14549);
and U15434 (N_15434,N_14513,N_14889);
nor U15435 (N_15435,N_14949,N_14741);
nor U15436 (N_15436,N_14887,N_14634);
nand U15437 (N_15437,N_14631,N_14881);
or U15438 (N_15438,N_14960,N_14532);
and U15439 (N_15439,N_14910,N_14691);
nand U15440 (N_15440,N_14605,N_14934);
nand U15441 (N_15441,N_14634,N_14698);
or U15442 (N_15442,N_14736,N_14621);
xor U15443 (N_15443,N_14812,N_14802);
xor U15444 (N_15444,N_14775,N_14672);
nor U15445 (N_15445,N_14822,N_14659);
xnor U15446 (N_15446,N_14573,N_14748);
or U15447 (N_15447,N_14872,N_14848);
nand U15448 (N_15448,N_14750,N_14959);
xor U15449 (N_15449,N_14601,N_14831);
or U15450 (N_15450,N_14749,N_14701);
xor U15451 (N_15451,N_14886,N_14971);
or U15452 (N_15452,N_14604,N_14526);
nor U15453 (N_15453,N_14625,N_14653);
nor U15454 (N_15454,N_14529,N_14862);
and U15455 (N_15455,N_14506,N_14828);
xnor U15456 (N_15456,N_14666,N_14584);
nor U15457 (N_15457,N_14862,N_14797);
nand U15458 (N_15458,N_14610,N_14793);
nand U15459 (N_15459,N_14840,N_14660);
or U15460 (N_15460,N_14922,N_14540);
or U15461 (N_15461,N_14564,N_14676);
or U15462 (N_15462,N_14775,N_14622);
or U15463 (N_15463,N_14560,N_14958);
nor U15464 (N_15464,N_14879,N_14714);
nand U15465 (N_15465,N_14514,N_14787);
or U15466 (N_15466,N_14879,N_14701);
xor U15467 (N_15467,N_14513,N_14765);
nand U15468 (N_15468,N_14858,N_14743);
xor U15469 (N_15469,N_14724,N_14948);
and U15470 (N_15470,N_14727,N_14856);
or U15471 (N_15471,N_14770,N_14652);
nand U15472 (N_15472,N_14980,N_14603);
or U15473 (N_15473,N_14992,N_14874);
and U15474 (N_15474,N_14784,N_14841);
nand U15475 (N_15475,N_14746,N_14967);
nor U15476 (N_15476,N_14670,N_14684);
or U15477 (N_15477,N_14670,N_14956);
nand U15478 (N_15478,N_14703,N_14641);
xnor U15479 (N_15479,N_14756,N_14656);
nand U15480 (N_15480,N_14575,N_14890);
nand U15481 (N_15481,N_14963,N_14593);
nor U15482 (N_15482,N_14888,N_14772);
or U15483 (N_15483,N_14654,N_14976);
xnor U15484 (N_15484,N_14778,N_14926);
and U15485 (N_15485,N_14559,N_14851);
xnor U15486 (N_15486,N_14953,N_14808);
xor U15487 (N_15487,N_14847,N_14725);
or U15488 (N_15488,N_14614,N_14501);
nand U15489 (N_15489,N_14608,N_14792);
and U15490 (N_15490,N_14724,N_14689);
and U15491 (N_15491,N_14604,N_14706);
or U15492 (N_15492,N_14569,N_14614);
nand U15493 (N_15493,N_14534,N_14868);
and U15494 (N_15494,N_14872,N_14896);
xor U15495 (N_15495,N_14787,N_14599);
or U15496 (N_15496,N_14587,N_14676);
xnor U15497 (N_15497,N_14743,N_14725);
and U15498 (N_15498,N_14546,N_14789);
nor U15499 (N_15499,N_14824,N_14626);
and U15500 (N_15500,N_15101,N_15147);
or U15501 (N_15501,N_15045,N_15055);
and U15502 (N_15502,N_15091,N_15233);
xor U15503 (N_15503,N_15256,N_15088);
nor U15504 (N_15504,N_15223,N_15049);
xnor U15505 (N_15505,N_15203,N_15303);
nand U15506 (N_15506,N_15164,N_15335);
nor U15507 (N_15507,N_15375,N_15169);
or U15508 (N_15508,N_15085,N_15271);
xor U15509 (N_15509,N_15191,N_15136);
or U15510 (N_15510,N_15234,N_15311);
or U15511 (N_15511,N_15359,N_15298);
and U15512 (N_15512,N_15460,N_15369);
and U15513 (N_15513,N_15445,N_15035);
and U15514 (N_15514,N_15330,N_15202);
and U15515 (N_15515,N_15261,N_15137);
or U15516 (N_15516,N_15388,N_15038);
xor U15517 (N_15517,N_15441,N_15240);
nand U15518 (N_15518,N_15280,N_15022);
xnor U15519 (N_15519,N_15265,N_15396);
and U15520 (N_15520,N_15106,N_15392);
and U15521 (N_15521,N_15347,N_15186);
nor U15522 (N_15522,N_15353,N_15258);
or U15523 (N_15523,N_15173,N_15288);
nor U15524 (N_15524,N_15127,N_15414);
nand U15525 (N_15525,N_15366,N_15345);
xor U15526 (N_15526,N_15214,N_15105);
xnor U15527 (N_15527,N_15461,N_15430);
nand U15528 (N_15528,N_15170,N_15193);
and U15529 (N_15529,N_15005,N_15397);
nand U15530 (N_15530,N_15152,N_15423);
nor U15531 (N_15531,N_15301,N_15189);
xnor U15532 (N_15532,N_15046,N_15367);
or U15533 (N_15533,N_15245,N_15462);
xor U15534 (N_15534,N_15218,N_15268);
or U15535 (N_15535,N_15383,N_15458);
nor U15536 (N_15536,N_15207,N_15135);
nor U15537 (N_15537,N_15150,N_15482);
xor U15538 (N_15538,N_15490,N_15450);
nand U15539 (N_15539,N_15270,N_15086);
nor U15540 (N_15540,N_15184,N_15394);
xor U15541 (N_15541,N_15126,N_15432);
xnor U15542 (N_15542,N_15036,N_15011);
xor U15543 (N_15543,N_15165,N_15350);
nor U15544 (N_15544,N_15081,N_15130);
or U15545 (N_15545,N_15358,N_15179);
xor U15546 (N_15546,N_15419,N_15181);
or U15547 (N_15547,N_15365,N_15323);
xnor U15548 (N_15548,N_15324,N_15178);
or U15549 (N_15549,N_15077,N_15222);
nand U15550 (N_15550,N_15060,N_15144);
and U15551 (N_15551,N_15092,N_15031);
or U15552 (N_15552,N_15426,N_15442);
and U15553 (N_15553,N_15273,N_15448);
or U15554 (N_15554,N_15190,N_15420);
nor U15555 (N_15555,N_15058,N_15139);
or U15556 (N_15556,N_15128,N_15151);
xnor U15557 (N_15557,N_15197,N_15064);
nand U15558 (N_15558,N_15346,N_15318);
xor U15559 (N_15559,N_15332,N_15410);
or U15560 (N_15560,N_15242,N_15315);
and U15561 (N_15561,N_15006,N_15122);
xor U15562 (N_15562,N_15119,N_15230);
xnor U15563 (N_15563,N_15279,N_15103);
nand U15564 (N_15564,N_15390,N_15108);
nand U15565 (N_15565,N_15226,N_15090);
nand U15566 (N_15566,N_15386,N_15422);
nor U15567 (N_15567,N_15093,N_15095);
nand U15568 (N_15568,N_15219,N_15166);
and U15569 (N_15569,N_15489,N_15082);
xor U15570 (N_15570,N_15379,N_15019);
or U15571 (N_15571,N_15200,N_15304);
nor U15572 (N_15572,N_15043,N_15235);
and U15573 (N_15573,N_15444,N_15459);
xor U15574 (N_15574,N_15372,N_15014);
and U15575 (N_15575,N_15195,N_15282);
nor U15576 (N_15576,N_15163,N_15220);
nand U15577 (N_15577,N_15417,N_15037);
nor U15578 (N_15578,N_15326,N_15287);
and U15579 (N_15579,N_15308,N_15260);
and U15580 (N_15580,N_15352,N_15296);
nor U15581 (N_15581,N_15063,N_15452);
nand U15582 (N_15582,N_15246,N_15215);
and U15583 (N_15583,N_15297,N_15110);
nand U15584 (N_15584,N_15168,N_15355);
or U15585 (N_15585,N_15054,N_15340);
nor U15586 (N_15586,N_15041,N_15313);
nand U15587 (N_15587,N_15059,N_15427);
and U15588 (N_15588,N_15473,N_15062);
nor U15589 (N_15589,N_15157,N_15463);
nor U15590 (N_15590,N_15250,N_15053);
xor U15591 (N_15591,N_15149,N_15146);
and U15592 (N_15592,N_15125,N_15068);
and U15593 (N_15593,N_15252,N_15159);
nand U15594 (N_15594,N_15192,N_15385);
nand U15595 (N_15595,N_15034,N_15310);
xor U15596 (N_15596,N_15107,N_15455);
nor U15597 (N_15597,N_15325,N_15180);
nor U15598 (N_15598,N_15387,N_15209);
nor U15599 (N_15599,N_15408,N_15228);
xor U15600 (N_15600,N_15141,N_15247);
or U15601 (N_15601,N_15285,N_15348);
xor U15602 (N_15602,N_15351,N_15098);
nor U15603 (N_15603,N_15254,N_15469);
and U15604 (N_15604,N_15269,N_15000);
nor U15605 (N_15605,N_15494,N_15148);
nor U15606 (N_15606,N_15021,N_15156);
and U15607 (N_15607,N_15339,N_15020);
nor U15608 (N_15608,N_15134,N_15281);
xnor U15609 (N_15609,N_15231,N_15433);
and U15610 (N_15610,N_15371,N_15289);
nor U15611 (N_15611,N_15267,N_15485);
nand U15612 (N_15612,N_15470,N_15023);
nor U15613 (N_15613,N_15454,N_15073);
nor U15614 (N_15614,N_15336,N_15492);
nor U15615 (N_15615,N_15418,N_15290);
or U15616 (N_15616,N_15236,N_15381);
and U15617 (N_15617,N_15435,N_15145);
and U15618 (N_15618,N_15399,N_15016);
nor U15619 (N_15619,N_15050,N_15312);
or U15620 (N_15620,N_15251,N_15111);
xnor U15621 (N_15621,N_15116,N_15416);
and U15622 (N_15622,N_15115,N_15176);
and U15623 (N_15623,N_15133,N_15276);
xnor U15624 (N_15624,N_15465,N_15089);
nor U15625 (N_15625,N_15495,N_15362);
xnor U15626 (N_15626,N_15262,N_15124);
and U15627 (N_15627,N_15155,N_15319);
or U15628 (N_15628,N_15224,N_15074);
and U15629 (N_15629,N_15497,N_15177);
and U15630 (N_15630,N_15293,N_15140);
and U15631 (N_15631,N_15331,N_15275);
and U15632 (N_15632,N_15072,N_15158);
xnor U15633 (N_15633,N_15487,N_15118);
nand U15634 (N_15634,N_15208,N_15446);
nand U15635 (N_15635,N_15070,N_15027);
nand U15636 (N_15636,N_15206,N_15225);
or U15637 (N_15637,N_15097,N_15076);
nor U15638 (N_15638,N_15412,N_15406);
and U15639 (N_15639,N_15354,N_15259);
nand U15640 (N_15640,N_15316,N_15334);
or U15641 (N_15641,N_15198,N_15411);
nor U15642 (N_15642,N_15374,N_15025);
and U15643 (N_15643,N_15196,N_15322);
or U15644 (N_15644,N_15210,N_15464);
nor U15645 (N_15645,N_15314,N_15009);
or U15646 (N_15646,N_15428,N_15421);
nand U15647 (N_15647,N_15341,N_15447);
nor U15648 (N_15648,N_15183,N_15030);
xnor U15649 (N_15649,N_15257,N_15239);
or U15650 (N_15650,N_15160,N_15328);
nand U15651 (N_15651,N_15187,N_15439);
nand U15652 (N_15652,N_15129,N_15333);
or U15653 (N_15653,N_15204,N_15481);
nor U15654 (N_15654,N_15229,N_15211);
nor U15655 (N_15655,N_15398,N_15380);
and U15656 (N_15656,N_15425,N_15407);
nand U15657 (N_15657,N_15120,N_15466);
nand U15658 (N_15658,N_15018,N_15047);
and U15659 (N_15659,N_15468,N_15102);
and U15660 (N_15660,N_15138,N_15194);
xnor U15661 (N_15661,N_15302,N_15415);
nor U15662 (N_15662,N_15075,N_15429);
and U15663 (N_15663,N_15456,N_15478);
and U15664 (N_15664,N_15493,N_15278);
nor U15665 (N_15665,N_15363,N_15199);
or U15666 (N_15666,N_15498,N_15474);
or U15667 (N_15667,N_15434,N_15272);
xor U15668 (N_15668,N_15377,N_15401);
xnor U15669 (N_15669,N_15174,N_15044);
xnor U15670 (N_15670,N_15306,N_15232);
xor U15671 (N_15671,N_15389,N_15227);
nor U15672 (N_15672,N_15378,N_15449);
and U15673 (N_15673,N_15357,N_15087);
nand U15674 (N_15674,N_15475,N_15263);
nor U15675 (N_15675,N_15376,N_15373);
or U15676 (N_15676,N_15405,N_15286);
and U15677 (N_15677,N_15182,N_15026);
and U15678 (N_15678,N_15080,N_15013);
or U15679 (N_15679,N_15142,N_15061);
and U15680 (N_15680,N_15438,N_15069);
or U15681 (N_15681,N_15338,N_15042);
xor U15682 (N_15682,N_15007,N_15112);
nor U15683 (N_15683,N_15342,N_15395);
xor U15684 (N_15684,N_15364,N_15453);
xor U15685 (N_15685,N_15457,N_15431);
nor U15686 (N_15686,N_15066,N_15283);
xor U15687 (N_15687,N_15057,N_15004);
nand U15688 (N_15688,N_15451,N_15361);
or U15689 (N_15689,N_15188,N_15015);
nor U15690 (N_15690,N_15294,N_15477);
and U15691 (N_15691,N_15382,N_15033);
xnor U15692 (N_15692,N_15123,N_15266);
and U15693 (N_15693,N_15329,N_15321);
or U15694 (N_15694,N_15402,N_15003);
or U15695 (N_15695,N_15029,N_15132);
nand U15696 (N_15696,N_15213,N_15205);
or U15697 (N_15697,N_15424,N_15284);
nand U15698 (N_15698,N_15244,N_15305);
or U15699 (N_15699,N_15201,N_15216);
nand U15700 (N_15700,N_15488,N_15360);
nor U15701 (N_15701,N_15113,N_15143);
or U15702 (N_15702,N_15017,N_15307);
nand U15703 (N_15703,N_15171,N_15096);
nand U15704 (N_15704,N_15471,N_15309);
nand U15705 (N_15705,N_15343,N_15114);
and U15706 (N_15706,N_15499,N_15409);
nand U15707 (N_15707,N_15217,N_15368);
nand U15708 (N_15708,N_15277,N_15079);
xor U15709 (N_15709,N_15436,N_15052);
or U15710 (N_15710,N_15467,N_15243);
or U15711 (N_15711,N_15356,N_15221);
or U15712 (N_15712,N_15249,N_15264);
nand U15713 (N_15713,N_15344,N_15337);
xor U15714 (N_15714,N_15404,N_15131);
nor U15715 (N_15715,N_15083,N_15024);
xor U15716 (N_15716,N_15032,N_15008);
xor U15717 (N_15717,N_15300,N_15100);
or U15718 (N_15718,N_15048,N_15153);
and U15719 (N_15719,N_15291,N_15001);
xor U15720 (N_15720,N_15167,N_15400);
xnor U15721 (N_15721,N_15472,N_15486);
nor U15722 (N_15722,N_15028,N_15094);
and U15723 (N_15723,N_15010,N_15491);
or U15724 (N_15724,N_15109,N_15012);
or U15725 (N_15725,N_15248,N_15403);
and U15726 (N_15726,N_15117,N_15440);
nor U15727 (N_15727,N_15175,N_15483);
nand U15728 (N_15728,N_15437,N_15002);
and U15729 (N_15729,N_15327,N_15065);
and U15730 (N_15730,N_15480,N_15393);
xnor U15731 (N_15731,N_15384,N_15078);
nor U15732 (N_15732,N_15071,N_15496);
and U15733 (N_15733,N_15161,N_15067);
xnor U15734 (N_15734,N_15172,N_15051);
and U15735 (N_15735,N_15185,N_15255);
nand U15736 (N_15736,N_15154,N_15099);
and U15737 (N_15737,N_15292,N_15040);
xnor U15738 (N_15738,N_15039,N_15238);
and U15739 (N_15739,N_15391,N_15162);
or U15740 (N_15740,N_15484,N_15237);
xnor U15741 (N_15741,N_15056,N_15295);
nor U15742 (N_15742,N_15212,N_15479);
or U15743 (N_15743,N_15274,N_15317);
or U15744 (N_15744,N_15121,N_15299);
and U15745 (N_15745,N_15413,N_15253);
or U15746 (N_15746,N_15104,N_15320);
nand U15747 (N_15747,N_15443,N_15476);
or U15748 (N_15748,N_15349,N_15084);
xnor U15749 (N_15749,N_15241,N_15370);
nand U15750 (N_15750,N_15280,N_15122);
nor U15751 (N_15751,N_15296,N_15283);
or U15752 (N_15752,N_15351,N_15189);
and U15753 (N_15753,N_15370,N_15453);
nor U15754 (N_15754,N_15473,N_15488);
nand U15755 (N_15755,N_15459,N_15396);
nor U15756 (N_15756,N_15484,N_15416);
xor U15757 (N_15757,N_15463,N_15487);
or U15758 (N_15758,N_15186,N_15038);
or U15759 (N_15759,N_15403,N_15456);
and U15760 (N_15760,N_15178,N_15404);
nand U15761 (N_15761,N_15281,N_15360);
nand U15762 (N_15762,N_15157,N_15283);
nor U15763 (N_15763,N_15276,N_15342);
xor U15764 (N_15764,N_15347,N_15454);
nor U15765 (N_15765,N_15340,N_15465);
xor U15766 (N_15766,N_15477,N_15414);
and U15767 (N_15767,N_15082,N_15372);
nor U15768 (N_15768,N_15025,N_15032);
or U15769 (N_15769,N_15330,N_15482);
nand U15770 (N_15770,N_15395,N_15479);
and U15771 (N_15771,N_15202,N_15449);
nor U15772 (N_15772,N_15296,N_15172);
or U15773 (N_15773,N_15016,N_15211);
xor U15774 (N_15774,N_15127,N_15187);
nor U15775 (N_15775,N_15360,N_15143);
and U15776 (N_15776,N_15193,N_15139);
or U15777 (N_15777,N_15005,N_15324);
xor U15778 (N_15778,N_15307,N_15152);
nor U15779 (N_15779,N_15301,N_15077);
and U15780 (N_15780,N_15182,N_15154);
nor U15781 (N_15781,N_15234,N_15487);
or U15782 (N_15782,N_15476,N_15381);
xnor U15783 (N_15783,N_15242,N_15453);
xor U15784 (N_15784,N_15452,N_15404);
or U15785 (N_15785,N_15040,N_15350);
nand U15786 (N_15786,N_15187,N_15258);
or U15787 (N_15787,N_15219,N_15299);
nor U15788 (N_15788,N_15216,N_15228);
xnor U15789 (N_15789,N_15382,N_15188);
nand U15790 (N_15790,N_15090,N_15107);
and U15791 (N_15791,N_15362,N_15381);
nand U15792 (N_15792,N_15115,N_15047);
xnor U15793 (N_15793,N_15496,N_15338);
and U15794 (N_15794,N_15175,N_15289);
and U15795 (N_15795,N_15266,N_15059);
nor U15796 (N_15796,N_15274,N_15269);
nand U15797 (N_15797,N_15493,N_15266);
nand U15798 (N_15798,N_15233,N_15426);
and U15799 (N_15799,N_15479,N_15025);
xor U15800 (N_15800,N_15241,N_15349);
nor U15801 (N_15801,N_15449,N_15213);
nor U15802 (N_15802,N_15296,N_15490);
nor U15803 (N_15803,N_15158,N_15395);
nor U15804 (N_15804,N_15173,N_15493);
xnor U15805 (N_15805,N_15110,N_15368);
nand U15806 (N_15806,N_15319,N_15338);
nand U15807 (N_15807,N_15055,N_15029);
nor U15808 (N_15808,N_15145,N_15239);
nand U15809 (N_15809,N_15083,N_15146);
and U15810 (N_15810,N_15005,N_15063);
nor U15811 (N_15811,N_15182,N_15009);
nand U15812 (N_15812,N_15441,N_15290);
xor U15813 (N_15813,N_15146,N_15108);
or U15814 (N_15814,N_15345,N_15143);
and U15815 (N_15815,N_15390,N_15098);
or U15816 (N_15816,N_15317,N_15133);
xnor U15817 (N_15817,N_15412,N_15289);
xor U15818 (N_15818,N_15244,N_15451);
nor U15819 (N_15819,N_15218,N_15182);
nand U15820 (N_15820,N_15250,N_15378);
nand U15821 (N_15821,N_15125,N_15375);
nand U15822 (N_15822,N_15175,N_15104);
nand U15823 (N_15823,N_15252,N_15280);
or U15824 (N_15824,N_15288,N_15460);
nand U15825 (N_15825,N_15128,N_15455);
xor U15826 (N_15826,N_15433,N_15264);
or U15827 (N_15827,N_15185,N_15068);
and U15828 (N_15828,N_15235,N_15392);
xor U15829 (N_15829,N_15193,N_15175);
nand U15830 (N_15830,N_15360,N_15308);
nor U15831 (N_15831,N_15162,N_15120);
xnor U15832 (N_15832,N_15107,N_15325);
nand U15833 (N_15833,N_15171,N_15305);
or U15834 (N_15834,N_15097,N_15186);
xor U15835 (N_15835,N_15128,N_15042);
and U15836 (N_15836,N_15348,N_15030);
nor U15837 (N_15837,N_15260,N_15411);
or U15838 (N_15838,N_15290,N_15270);
nor U15839 (N_15839,N_15339,N_15465);
nor U15840 (N_15840,N_15065,N_15243);
nand U15841 (N_15841,N_15288,N_15154);
nor U15842 (N_15842,N_15492,N_15026);
nand U15843 (N_15843,N_15371,N_15208);
nand U15844 (N_15844,N_15035,N_15193);
nand U15845 (N_15845,N_15107,N_15147);
nand U15846 (N_15846,N_15313,N_15305);
and U15847 (N_15847,N_15188,N_15425);
nand U15848 (N_15848,N_15424,N_15203);
nor U15849 (N_15849,N_15003,N_15136);
and U15850 (N_15850,N_15306,N_15186);
xnor U15851 (N_15851,N_15481,N_15250);
and U15852 (N_15852,N_15403,N_15202);
xor U15853 (N_15853,N_15107,N_15088);
nand U15854 (N_15854,N_15069,N_15198);
and U15855 (N_15855,N_15269,N_15304);
and U15856 (N_15856,N_15072,N_15082);
or U15857 (N_15857,N_15105,N_15147);
nand U15858 (N_15858,N_15054,N_15479);
nand U15859 (N_15859,N_15307,N_15169);
or U15860 (N_15860,N_15389,N_15266);
and U15861 (N_15861,N_15050,N_15159);
nor U15862 (N_15862,N_15244,N_15254);
or U15863 (N_15863,N_15364,N_15250);
nand U15864 (N_15864,N_15457,N_15356);
and U15865 (N_15865,N_15444,N_15098);
xnor U15866 (N_15866,N_15135,N_15284);
nand U15867 (N_15867,N_15113,N_15213);
and U15868 (N_15868,N_15188,N_15047);
nand U15869 (N_15869,N_15450,N_15454);
nand U15870 (N_15870,N_15157,N_15331);
and U15871 (N_15871,N_15086,N_15021);
and U15872 (N_15872,N_15227,N_15197);
xor U15873 (N_15873,N_15418,N_15026);
and U15874 (N_15874,N_15282,N_15320);
and U15875 (N_15875,N_15307,N_15442);
nor U15876 (N_15876,N_15343,N_15295);
xor U15877 (N_15877,N_15078,N_15420);
nand U15878 (N_15878,N_15162,N_15381);
nor U15879 (N_15879,N_15394,N_15495);
or U15880 (N_15880,N_15197,N_15482);
nor U15881 (N_15881,N_15450,N_15464);
nor U15882 (N_15882,N_15334,N_15243);
nand U15883 (N_15883,N_15002,N_15450);
or U15884 (N_15884,N_15106,N_15197);
nand U15885 (N_15885,N_15291,N_15365);
nor U15886 (N_15886,N_15017,N_15360);
or U15887 (N_15887,N_15118,N_15234);
and U15888 (N_15888,N_15446,N_15174);
and U15889 (N_15889,N_15447,N_15084);
nand U15890 (N_15890,N_15359,N_15228);
and U15891 (N_15891,N_15311,N_15416);
nand U15892 (N_15892,N_15443,N_15219);
nor U15893 (N_15893,N_15405,N_15115);
nor U15894 (N_15894,N_15185,N_15475);
and U15895 (N_15895,N_15320,N_15175);
nand U15896 (N_15896,N_15358,N_15109);
and U15897 (N_15897,N_15078,N_15075);
nor U15898 (N_15898,N_15366,N_15293);
and U15899 (N_15899,N_15163,N_15475);
nor U15900 (N_15900,N_15458,N_15473);
xor U15901 (N_15901,N_15471,N_15064);
or U15902 (N_15902,N_15056,N_15344);
or U15903 (N_15903,N_15329,N_15209);
nand U15904 (N_15904,N_15175,N_15129);
or U15905 (N_15905,N_15059,N_15084);
xnor U15906 (N_15906,N_15243,N_15208);
nor U15907 (N_15907,N_15336,N_15441);
or U15908 (N_15908,N_15031,N_15346);
nand U15909 (N_15909,N_15273,N_15471);
xnor U15910 (N_15910,N_15061,N_15042);
or U15911 (N_15911,N_15189,N_15218);
nor U15912 (N_15912,N_15487,N_15153);
and U15913 (N_15913,N_15479,N_15278);
and U15914 (N_15914,N_15030,N_15021);
nand U15915 (N_15915,N_15113,N_15122);
nand U15916 (N_15916,N_15165,N_15220);
xnor U15917 (N_15917,N_15282,N_15389);
xor U15918 (N_15918,N_15469,N_15313);
xnor U15919 (N_15919,N_15218,N_15453);
nand U15920 (N_15920,N_15164,N_15248);
and U15921 (N_15921,N_15436,N_15049);
xnor U15922 (N_15922,N_15122,N_15441);
nand U15923 (N_15923,N_15143,N_15471);
and U15924 (N_15924,N_15022,N_15144);
nor U15925 (N_15925,N_15063,N_15062);
xor U15926 (N_15926,N_15424,N_15432);
and U15927 (N_15927,N_15012,N_15133);
or U15928 (N_15928,N_15317,N_15050);
nand U15929 (N_15929,N_15393,N_15213);
xnor U15930 (N_15930,N_15178,N_15043);
or U15931 (N_15931,N_15122,N_15382);
xor U15932 (N_15932,N_15193,N_15294);
nor U15933 (N_15933,N_15285,N_15406);
xor U15934 (N_15934,N_15076,N_15325);
nor U15935 (N_15935,N_15418,N_15221);
nor U15936 (N_15936,N_15192,N_15295);
or U15937 (N_15937,N_15123,N_15239);
or U15938 (N_15938,N_15145,N_15051);
nand U15939 (N_15939,N_15243,N_15108);
or U15940 (N_15940,N_15224,N_15457);
nor U15941 (N_15941,N_15282,N_15354);
or U15942 (N_15942,N_15015,N_15001);
nor U15943 (N_15943,N_15179,N_15398);
nand U15944 (N_15944,N_15258,N_15446);
nand U15945 (N_15945,N_15018,N_15243);
and U15946 (N_15946,N_15409,N_15332);
or U15947 (N_15947,N_15117,N_15213);
and U15948 (N_15948,N_15055,N_15113);
xor U15949 (N_15949,N_15313,N_15160);
and U15950 (N_15950,N_15075,N_15043);
nand U15951 (N_15951,N_15418,N_15314);
xnor U15952 (N_15952,N_15113,N_15400);
nand U15953 (N_15953,N_15426,N_15317);
and U15954 (N_15954,N_15128,N_15204);
and U15955 (N_15955,N_15330,N_15492);
or U15956 (N_15956,N_15372,N_15268);
xor U15957 (N_15957,N_15217,N_15455);
and U15958 (N_15958,N_15486,N_15293);
or U15959 (N_15959,N_15108,N_15010);
and U15960 (N_15960,N_15007,N_15464);
nand U15961 (N_15961,N_15487,N_15356);
nor U15962 (N_15962,N_15055,N_15122);
and U15963 (N_15963,N_15426,N_15154);
nand U15964 (N_15964,N_15306,N_15387);
and U15965 (N_15965,N_15348,N_15431);
nor U15966 (N_15966,N_15007,N_15043);
nor U15967 (N_15967,N_15042,N_15243);
nor U15968 (N_15968,N_15233,N_15456);
and U15969 (N_15969,N_15175,N_15453);
xnor U15970 (N_15970,N_15233,N_15152);
nor U15971 (N_15971,N_15383,N_15486);
and U15972 (N_15972,N_15408,N_15189);
nand U15973 (N_15973,N_15196,N_15471);
xnor U15974 (N_15974,N_15087,N_15330);
or U15975 (N_15975,N_15304,N_15352);
nor U15976 (N_15976,N_15076,N_15478);
or U15977 (N_15977,N_15193,N_15235);
nor U15978 (N_15978,N_15468,N_15053);
or U15979 (N_15979,N_15425,N_15306);
xnor U15980 (N_15980,N_15019,N_15198);
or U15981 (N_15981,N_15429,N_15494);
nand U15982 (N_15982,N_15274,N_15042);
xor U15983 (N_15983,N_15205,N_15307);
nor U15984 (N_15984,N_15104,N_15237);
and U15985 (N_15985,N_15410,N_15004);
nor U15986 (N_15986,N_15209,N_15236);
and U15987 (N_15987,N_15462,N_15195);
nand U15988 (N_15988,N_15170,N_15414);
nor U15989 (N_15989,N_15214,N_15264);
nor U15990 (N_15990,N_15279,N_15006);
nand U15991 (N_15991,N_15106,N_15254);
nor U15992 (N_15992,N_15098,N_15012);
and U15993 (N_15993,N_15444,N_15375);
or U15994 (N_15994,N_15371,N_15330);
and U15995 (N_15995,N_15110,N_15395);
and U15996 (N_15996,N_15029,N_15052);
or U15997 (N_15997,N_15033,N_15205);
and U15998 (N_15998,N_15368,N_15237);
nand U15999 (N_15999,N_15426,N_15031);
or U16000 (N_16000,N_15965,N_15789);
nor U16001 (N_16001,N_15980,N_15990);
or U16002 (N_16002,N_15732,N_15715);
nand U16003 (N_16003,N_15857,N_15870);
nor U16004 (N_16004,N_15853,N_15630);
nand U16005 (N_16005,N_15948,N_15929);
and U16006 (N_16006,N_15563,N_15879);
nor U16007 (N_16007,N_15687,N_15983);
nor U16008 (N_16008,N_15685,N_15609);
nand U16009 (N_16009,N_15916,N_15727);
or U16010 (N_16010,N_15644,N_15521);
and U16011 (N_16011,N_15860,N_15903);
and U16012 (N_16012,N_15695,N_15871);
and U16013 (N_16013,N_15790,N_15607);
xor U16014 (N_16014,N_15706,N_15925);
nand U16015 (N_16015,N_15680,N_15831);
xor U16016 (N_16016,N_15509,N_15873);
or U16017 (N_16017,N_15691,N_15745);
xor U16018 (N_16018,N_15812,N_15531);
nor U16019 (N_16019,N_15522,N_15885);
and U16020 (N_16020,N_15970,N_15798);
xnor U16021 (N_16021,N_15656,N_15985);
xor U16022 (N_16022,N_15973,N_15876);
nor U16023 (N_16023,N_15655,N_15517);
xor U16024 (N_16024,N_15843,N_15779);
xor U16025 (N_16025,N_15802,N_15746);
or U16026 (N_16026,N_15731,N_15847);
or U16027 (N_16027,N_15922,N_15835);
and U16028 (N_16028,N_15586,N_15780);
nand U16029 (N_16029,N_15976,N_15991);
nand U16030 (N_16030,N_15614,N_15765);
and U16031 (N_16031,N_15869,N_15744);
nor U16032 (N_16032,N_15776,N_15846);
nand U16033 (N_16033,N_15997,N_15712);
xor U16034 (N_16034,N_15883,N_15710);
and U16035 (N_16035,N_15815,N_15781);
nand U16036 (N_16036,N_15592,N_15625);
or U16037 (N_16037,N_15949,N_15877);
nor U16038 (N_16038,N_15714,N_15984);
xnor U16039 (N_16039,N_15761,N_15969);
nand U16040 (N_16040,N_15882,N_15955);
nor U16041 (N_16041,N_15633,N_15918);
or U16042 (N_16042,N_15737,N_15887);
nand U16043 (N_16043,N_15709,N_15844);
and U16044 (N_16044,N_15700,N_15594);
or U16045 (N_16045,N_15958,N_15551);
nand U16046 (N_16046,N_15937,N_15993);
or U16047 (N_16047,N_15787,N_15891);
and U16048 (N_16048,N_15747,N_15503);
and U16049 (N_16049,N_15565,N_15906);
xnor U16050 (N_16050,N_15632,N_15627);
xor U16051 (N_16051,N_15567,N_15834);
nand U16052 (N_16052,N_15688,N_15981);
or U16053 (N_16053,N_15571,N_15515);
nand U16054 (N_16054,N_15536,N_15880);
and U16055 (N_16055,N_15649,N_15783);
xor U16056 (N_16056,N_15543,N_15805);
nor U16057 (N_16057,N_15718,N_15865);
and U16058 (N_16058,N_15839,N_15568);
and U16059 (N_16059,N_15640,N_15862);
nor U16060 (N_16060,N_15824,N_15738);
nand U16061 (N_16061,N_15591,N_15678);
nor U16062 (N_16062,N_15754,N_15666);
nand U16063 (N_16063,N_15673,N_15942);
xor U16064 (N_16064,N_15537,N_15518);
xor U16065 (N_16065,N_15597,N_15777);
and U16066 (N_16066,N_15756,N_15613);
nand U16067 (N_16067,N_15966,N_15530);
nor U16068 (N_16068,N_15755,N_15811);
nand U16069 (N_16069,N_15622,N_15904);
nand U16070 (N_16070,N_15808,N_15936);
nand U16071 (N_16071,N_15897,N_15977);
and U16072 (N_16072,N_15672,N_15643);
nor U16073 (N_16073,N_15686,N_15516);
nor U16074 (N_16074,N_15513,N_15854);
nand U16075 (N_16075,N_15896,N_15730);
nor U16076 (N_16076,N_15758,N_15694);
nor U16077 (N_16077,N_15851,N_15769);
nor U16078 (N_16078,N_15574,N_15724);
and U16079 (N_16079,N_15674,N_15662);
or U16080 (N_16080,N_15697,N_15647);
xor U16081 (N_16081,N_15957,N_15905);
or U16082 (N_16082,N_15890,N_15593);
nor U16083 (N_16083,N_15935,N_15676);
xnor U16084 (N_16084,N_15863,N_15809);
nor U16085 (N_16085,N_15524,N_15610);
nor U16086 (N_16086,N_15941,N_15959);
nand U16087 (N_16087,N_15766,N_15519);
or U16088 (N_16088,N_15520,N_15864);
nor U16089 (N_16089,N_15919,N_15541);
xor U16090 (N_16090,N_15620,N_15884);
and U16091 (N_16091,N_15796,N_15719);
xnor U16092 (N_16092,N_15671,N_15585);
or U16093 (N_16093,N_15546,N_15911);
and U16094 (N_16094,N_15668,N_15635);
nand U16095 (N_16095,N_15927,N_15583);
and U16096 (N_16096,N_15791,N_15907);
nor U16097 (N_16097,N_15611,N_15713);
nor U16098 (N_16098,N_15921,N_15938);
xor U16099 (N_16099,N_15651,N_15703);
or U16100 (N_16100,N_15850,N_15828);
nor U16101 (N_16101,N_15657,N_15872);
nor U16102 (N_16102,N_15628,N_15721);
xor U16103 (N_16103,N_15582,N_15670);
and U16104 (N_16104,N_15764,N_15775);
or U16105 (N_16105,N_15733,N_15841);
nand U16106 (N_16106,N_15799,N_15636);
xor U16107 (N_16107,N_15848,N_15748);
and U16108 (N_16108,N_15621,N_15944);
nand U16109 (N_16109,N_15956,N_15501);
nand U16110 (N_16110,N_15605,N_15838);
and U16111 (N_16111,N_15507,N_15786);
and U16112 (N_16112,N_15974,N_15527);
and U16113 (N_16113,N_15868,N_15569);
and U16114 (N_16114,N_15542,N_15679);
xor U16115 (N_16115,N_15599,N_15665);
nor U16116 (N_16116,N_15639,N_15989);
nor U16117 (N_16117,N_15529,N_15742);
xnor U16118 (N_16118,N_15603,N_15951);
nor U16119 (N_16119,N_15578,N_15648);
xnor U16120 (N_16120,N_15999,N_15889);
and U16121 (N_16121,N_15823,N_15928);
or U16122 (N_16122,N_15506,N_15900);
or U16123 (N_16123,N_15945,N_15669);
or U16124 (N_16124,N_15555,N_15792);
nor U16125 (N_16125,N_15556,N_15553);
nand U16126 (N_16126,N_15508,N_15895);
and U16127 (N_16127,N_15913,N_15581);
xor U16128 (N_16128,N_15570,N_15892);
or U16129 (N_16129,N_15992,N_15881);
or U16130 (N_16130,N_15986,N_15740);
xnor U16131 (N_16131,N_15631,N_15914);
nand U16132 (N_16132,N_15500,N_15818);
xor U16133 (N_16133,N_15588,N_15767);
xnor U16134 (N_16134,N_15564,N_15893);
xor U16135 (N_16135,N_15601,N_15528);
nor U16136 (N_16136,N_15910,N_15988);
xor U16137 (N_16137,N_15600,N_15560);
and U16138 (N_16138,N_15624,N_15751);
xor U16139 (N_16139,N_15646,N_15902);
nand U16140 (N_16140,N_15573,N_15909);
and U16141 (N_16141,N_15923,N_15778);
xnor U16142 (N_16142,N_15874,N_15768);
xnor U16143 (N_16143,N_15523,N_15566);
xnor U16144 (N_16144,N_15736,N_15952);
xor U16145 (N_16145,N_15661,N_15511);
nand U16146 (N_16146,N_15595,N_15612);
nand U16147 (N_16147,N_15770,N_15899);
xnor U16148 (N_16148,N_15934,N_15699);
nand U16149 (N_16149,N_15852,N_15598);
nand U16150 (N_16150,N_15855,N_15596);
and U16151 (N_16151,N_15830,N_15728);
xnor U16152 (N_16152,N_15933,N_15637);
or U16153 (N_16153,N_15749,N_15978);
or U16154 (N_16154,N_15964,N_15616);
nand U16155 (N_16155,N_15832,N_15572);
or U16156 (N_16156,N_15998,N_15735);
nand U16157 (N_16157,N_15658,N_15793);
and U16158 (N_16158,N_15663,N_15619);
or U16159 (N_16159,N_15532,N_15510);
nor U16160 (N_16160,N_15842,N_15702);
or U16161 (N_16161,N_15734,N_15924);
xor U16162 (N_16162,N_15677,N_15514);
nand U16163 (N_16163,N_15642,N_15849);
or U16164 (N_16164,N_15693,N_15762);
and U16165 (N_16165,N_15682,N_15822);
or U16166 (N_16166,N_15757,N_15533);
or U16167 (N_16167,N_15804,N_15840);
nand U16168 (N_16168,N_15545,N_15926);
or U16169 (N_16169,N_15696,N_15547);
or U16170 (N_16170,N_15638,N_15615);
nor U16171 (N_16171,N_15602,N_15820);
or U16172 (N_16172,N_15716,N_15652);
nor U16173 (N_16173,N_15720,N_15741);
nor U16174 (N_16174,N_15554,N_15972);
and U16175 (N_16175,N_15813,N_15705);
nand U16176 (N_16176,N_15618,N_15759);
xnor U16177 (N_16177,N_15535,N_15894);
and U16178 (N_16178,N_15827,N_15801);
and U16179 (N_16179,N_15641,N_15502);
or U16180 (N_16180,N_15675,N_15794);
nor U16181 (N_16181,N_15587,N_15947);
and U16182 (N_16182,N_15689,N_15729);
nor U16183 (N_16183,N_15774,N_15539);
or U16184 (N_16184,N_15743,N_15845);
and U16185 (N_16185,N_15861,N_15963);
nand U16186 (N_16186,N_15698,N_15784);
or U16187 (N_16187,N_15722,N_15659);
nand U16188 (N_16188,N_15932,N_15653);
or U16189 (N_16189,N_15683,N_15617);
or U16190 (N_16190,N_15707,N_15577);
nand U16191 (N_16191,N_15561,N_15690);
xor U16192 (N_16192,N_15943,N_15623);
nand U16193 (N_16193,N_15858,N_15788);
or U16194 (N_16194,N_15821,N_15708);
and U16195 (N_16195,N_15975,N_15575);
nand U16196 (N_16196,N_15994,N_15711);
or U16197 (N_16197,N_15512,N_15557);
and U16198 (N_16198,N_15920,N_15684);
xnor U16199 (N_16199,N_15915,N_15559);
or U16200 (N_16200,N_15750,N_15886);
xor U16201 (N_16201,N_15837,N_15763);
or U16202 (N_16202,N_15540,N_15807);
or U16203 (N_16203,N_15645,N_15946);
or U16204 (N_16204,N_15650,N_15704);
nand U16205 (N_16205,N_15549,N_15829);
nand U16206 (N_16206,N_15795,N_15979);
xor U16207 (N_16207,N_15800,N_15898);
or U16208 (N_16208,N_15526,N_15917);
or U16209 (N_16209,N_15954,N_15908);
nand U16210 (N_16210,N_15717,N_15654);
xnor U16211 (N_16211,N_15785,N_15580);
xor U16212 (N_16212,N_15810,N_15552);
xnor U16213 (N_16213,N_15576,N_15548);
xnor U16214 (N_16214,N_15589,N_15558);
nor U16215 (N_16215,N_15782,N_15760);
nor U16216 (N_16216,N_15550,N_15982);
nand U16217 (N_16217,N_15803,N_15772);
or U16218 (N_16218,N_15836,N_15968);
and U16219 (N_16219,N_15953,N_15878);
or U16220 (N_16220,N_15701,N_15867);
nor U16221 (N_16221,N_15814,N_15660);
nand U16222 (N_16222,N_15826,N_15664);
or U16223 (N_16223,N_15995,N_15726);
xor U16224 (N_16224,N_15930,N_15875);
or U16225 (N_16225,N_15816,N_15856);
or U16226 (N_16226,N_15629,N_15725);
nor U16227 (N_16227,N_15866,N_15940);
xor U16228 (N_16228,N_15996,N_15971);
xnor U16229 (N_16229,N_15931,N_15634);
xor U16230 (N_16230,N_15544,N_15773);
or U16231 (N_16231,N_15590,N_15817);
xnor U16232 (N_16232,N_15505,N_15538);
nor U16233 (N_16233,N_15525,N_15833);
nand U16234 (N_16234,N_15753,N_15579);
xnor U16235 (N_16235,N_15771,N_15987);
xor U16236 (N_16236,N_15939,N_15606);
and U16237 (N_16237,N_15825,N_15608);
nand U16238 (N_16238,N_15723,N_15739);
or U16239 (N_16239,N_15819,N_15960);
nand U16240 (N_16240,N_15504,N_15584);
xnor U16241 (N_16241,N_15961,N_15562);
xor U16242 (N_16242,N_15534,N_15806);
nor U16243 (N_16243,N_15962,N_15797);
xor U16244 (N_16244,N_15626,N_15901);
and U16245 (N_16245,N_15692,N_15912);
nor U16246 (N_16246,N_15888,N_15950);
or U16247 (N_16247,N_15859,N_15667);
nor U16248 (N_16248,N_15604,N_15967);
nor U16249 (N_16249,N_15752,N_15681);
xnor U16250 (N_16250,N_15806,N_15796);
or U16251 (N_16251,N_15632,N_15966);
nand U16252 (N_16252,N_15641,N_15744);
nor U16253 (N_16253,N_15989,N_15665);
xor U16254 (N_16254,N_15977,N_15573);
xor U16255 (N_16255,N_15760,N_15650);
xor U16256 (N_16256,N_15570,N_15894);
nand U16257 (N_16257,N_15985,N_15955);
nand U16258 (N_16258,N_15847,N_15512);
nand U16259 (N_16259,N_15586,N_15847);
and U16260 (N_16260,N_15727,N_15924);
nand U16261 (N_16261,N_15820,N_15707);
nand U16262 (N_16262,N_15616,N_15829);
nand U16263 (N_16263,N_15728,N_15951);
and U16264 (N_16264,N_15837,N_15830);
nor U16265 (N_16265,N_15909,N_15554);
and U16266 (N_16266,N_15650,N_15872);
xnor U16267 (N_16267,N_15738,N_15702);
nor U16268 (N_16268,N_15885,N_15756);
or U16269 (N_16269,N_15605,N_15985);
and U16270 (N_16270,N_15688,N_15721);
nor U16271 (N_16271,N_15777,N_15974);
nand U16272 (N_16272,N_15802,N_15775);
or U16273 (N_16273,N_15763,N_15793);
xnor U16274 (N_16274,N_15917,N_15713);
or U16275 (N_16275,N_15790,N_15588);
nor U16276 (N_16276,N_15667,N_15564);
xor U16277 (N_16277,N_15811,N_15789);
and U16278 (N_16278,N_15682,N_15778);
nor U16279 (N_16279,N_15946,N_15632);
nor U16280 (N_16280,N_15668,N_15595);
nand U16281 (N_16281,N_15582,N_15545);
or U16282 (N_16282,N_15721,N_15637);
or U16283 (N_16283,N_15955,N_15800);
xor U16284 (N_16284,N_15827,N_15791);
nand U16285 (N_16285,N_15974,N_15966);
nand U16286 (N_16286,N_15936,N_15518);
or U16287 (N_16287,N_15788,N_15851);
and U16288 (N_16288,N_15989,N_15906);
nor U16289 (N_16289,N_15566,N_15618);
xor U16290 (N_16290,N_15836,N_15980);
xnor U16291 (N_16291,N_15804,N_15984);
nor U16292 (N_16292,N_15926,N_15585);
nor U16293 (N_16293,N_15649,N_15976);
or U16294 (N_16294,N_15907,N_15502);
nand U16295 (N_16295,N_15927,N_15920);
nand U16296 (N_16296,N_15506,N_15969);
xnor U16297 (N_16297,N_15874,N_15892);
or U16298 (N_16298,N_15542,N_15985);
xor U16299 (N_16299,N_15840,N_15602);
nand U16300 (N_16300,N_15565,N_15551);
and U16301 (N_16301,N_15564,N_15676);
xor U16302 (N_16302,N_15874,N_15715);
or U16303 (N_16303,N_15905,N_15590);
xor U16304 (N_16304,N_15846,N_15517);
xnor U16305 (N_16305,N_15711,N_15528);
nand U16306 (N_16306,N_15602,N_15633);
and U16307 (N_16307,N_15665,N_15628);
xnor U16308 (N_16308,N_15755,N_15715);
and U16309 (N_16309,N_15881,N_15977);
xnor U16310 (N_16310,N_15563,N_15954);
nand U16311 (N_16311,N_15642,N_15980);
xor U16312 (N_16312,N_15628,N_15991);
and U16313 (N_16313,N_15917,N_15576);
and U16314 (N_16314,N_15789,N_15648);
nor U16315 (N_16315,N_15570,N_15990);
or U16316 (N_16316,N_15782,N_15857);
and U16317 (N_16317,N_15991,N_15739);
or U16318 (N_16318,N_15601,N_15689);
nor U16319 (N_16319,N_15918,N_15745);
and U16320 (N_16320,N_15940,N_15981);
nand U16321 (N_16321,N_15787,N_15979);
nor U16322 (N_16322,N_15889,N_15544);
nor U16323 (N_16323,N_15880,N_15511);
nand U16324 (N_16324,N_15720,N_15893);
xor U16325 (N_16325,N_15675,N_15690);
xor U16326 (N_16326,N_15980,N_15942);
or U16327 (N_16327,N_15665,N_15847);
and U16328 (N_16328,N_15547,N_15887);
nand U16329 (N_16329,N_15967,N_15853);
or U16330 (N_16330,N_15787,N_15978);
xor U16331 (N_16331,N_15922,N_15589);
or U16332 (N_16332,N_15616,N_15614);
nand U16333 (N_16333,N_15985,N_15975);
nand U16334 (N_16334,N_15641,N_15662);
or U16335 (N_16335,N_15696,N_15942);
nand U16336 (N_16336,N_15999,N_15591);
nand U16337 (N_16337,N_15755,N_15897);
xor U16338 (N_16338,N_15926,N_15745);
or U16339 (N_16339,N_15552,N_15694);
and U16340 (N_16340,N_15794,N_15986);
nor U16341 (N_16341,N_15693,N_15936);
and U16342 (N_16342,N_15922,N_15692);
or U16343 (N_16343,N_15849,N_15621);
nor U16344 (N_16344,N_15788,N_15685);
and U16345 (N_16345,N_15560,N_15709);
xor U16346 (N_16346,N_15804,N_15519);
and U16347 (N_16347,N_15734,N_15629);
xor U16348 (N_16348,N_15566,N_15901);
and U16349 (N_16349,N_15799,N_15718);
and U16350 (N_16350,N_15734,N_15814);
nor U16351 (N_16351,N_15959,N_15884);
xor U16352 (N_16352,N_15977,N_15677);
nor U16353 (N_16353,N_15734,N_15893);
xnor U16354 (N_16354,N_15646,N_15864);
or U16355 (N_16355,N_15860,N_15898);
or U16356 (N_16356,N_15628,N_15911);
xnor U16357 (N_16357,N_15865,N_15703);
nand U16358 (N_16358,N_15941,N_15824);
xnor U16359 (N_16359,N_15850,N_15548);
nand U16360 (N_16360,N_15550,N_15825);
nor U16361 (N_16361,N_15951,N_15615);
xnor U16362 (N_16362,N_15932,N_15784);
and U16363 (N_16363,N_15802,N_15673);
nor U16364 (N_16364,N_15648,N_15636);
or U16365 (N_16365,N_15589,N_15730);
or U16366 (N_16366,N_15668,N_15976);
xor U16367 (N_16367,N_15746,N_15561);
nand U16368 (N_16368,N_15543,N_15777);
nand U16369 (N_16369,N_15512,N_15943);
and U16370 (N_16370,N_15916,N_15634);
nor U16371 (N_16371,N_15924,N_15790);
nand U16372 (N_16372,N_15537,N_15702);
and U16373 (N_16373,N_15598,N_15654);
xnor U16374 (N_16374,N_15988,N_15931);
nand U16375 (N_16375,N_15812,N_15895);
and U16376 (N_16376,N_15859,N_15568);
xnor U16377 (N_16377,N_15668,N_15784);
nor U16378 (N_16378,N_15795,N_15774);
and U16379 (N_16379,N_15873,N_15645);
xor U16380 (N_16380,N_15599,N_15626);
or U16381 (N_16381,N_15933,N_15980);
or U16382 (N_16382,N_15985,N_15766);
xor U16383 (N_16383,N_15933,N_15939);
nor U16384 (N_16384,N_15564,N_15697);
nand U16385 (N_16385,N_15624,N_15819);
or U16386 (N_16386,N_15739,N_15561);
and U16387 (N_16387,N_15687,N_15822);
nor U16388 (N_16388,N_15726,N_15840);
nor U16389 (N_16389,N_15567,N_15912);
nor U16390 (N_16390,N_15780,N_15750);
nor U16391 (N_16391,N_15876,N_15715);
xor U16392 (N_16392,N_15717,N_15903);
and U16393 (N_16393,N_15603,N_15590);
xor U16394 (N_16394,N_15867,N_15517);
and U16395 (N_16395,N_15588,N_15895);
nand U16396 (N_16396,N_15751,N_15913);
nand U16397 (N_16397,N_15690,N_15691);
and U16398 (N_16398,N_15735,N_15700);
nand U16399 (N_16399,N_15945,N_15633);
and U16400 (N_16400,N_15682,N_15836);
nand U16401 (N_16401,N_15726,N_15819);
or U16402 (N_16402,N_15818,N_15681);
nor U16403 (N_16403,N_15663,N_15880);
nor U16404 (N_16404,N_15896,N_15655);
xnor U16405 (N_16405,N_15996,N_15715);
xor U16406 (N_16406,N_15657,N_15785);
nand U16407 (N_16407,N_15952,N_15988);
nor U16408 (N_16408,N_15870,N_15523);
or U16409 (N_16409,N_15555,N_15663);
nor U16410 (N_16410,N_15579,N_15720);
nor U16411 (N_16411,N_15570,N_15508);
nand U16412 (N_16412,N_15984,N_15829);
nand U16413 (N_16413,N_15961,N_15722);
nor U16414 (N_16414,N_15996,N_15525);
nor U16415 (N_16415,N_15527,N_15648);
or U16416 (N_16416,N_15848,N_15695);
nand U16417 (N_16417,N_15642,N_15928);
nor U16418 (N_16418,N_15639,N_15752);
xnor U16419 (N_16419,N_15969,N_15972);
nand U16420 (N_16420,N_15771,N_15952);
xnor U16421 (N_16421,N_15576,N_15697);
or U16422 (N_16422,N_15502,N_15615);
xnor U16423 (N_16423,N_15609,N_15727);
or U16424 (N_16424,N_15818,N_15637);
nor U16425 (N_16425,N_15857,N_15970);
and U16426 (N_16426,N_15840,N_15868);
or U16427 (N_16427,N_15572,N_15506);
nor U16428 (N_16428,N_15560,N_15943);
nor U16429 (N_16429,N_15985,N_15771);
nor U16430 (N_16430,N_15543,N_15844);
xnor U16431 (N_16431,N_15993,N_15883);
and U16432 (N_16432,N_15730,N_15638);
xnor U16433 (N_16433,N_15762,N_15806);
nor U16434 (N_16434,N_15793,N_15709);
nor U16435 (N_16435,N_15618,N_15906);
xnor U16436 (N_16436,N_15605,N_15818);
nand U16437 (N_16437,N_15915,N_15707);
xor U16438 (N_16438,N_15607,N_15660);
or U16439 (N_16439,N_15656,N_15931);
nand U16440 (N_16440,N_15799,N_15791);
nand U16441 (N_16441,N_15709,N_15551);
or U16442 (N_16442,N_15623,N_15557);
and U16443 (N_16443,N_15567,N_15703);
nand U16444 (N_16444,N_15760,N_15959);
xor U16445 (N_16445,N_15782,N_15564);
or U16446 (N_16446,N_15992,N_15731);
xnor U16447 (N_16447,N_15500,N_15540);
nand U16448 (N_16448,N_15895,N_15505);
xnor U16449 (N_16449,N_15836,N_15856);
xor U16450 (N_16450,N_15640,N_15501);
nand U16451 (N_16451,N_15727,N_15555);
nor U16452 (N_16452,N_15502,N_15714);
xor U16453 (N_16453,N_15800,N_15697);
nand U16454 (N_16454,N_15623,N_15585);
nor U16455 (N_16455,N_15961,N_15719);
nor U16456 (N_16456,N_15676,N_15969);
nand U16457 (N_16457,N_15742,N_15908);
nand U16458 (N_16458,N_15996,N_15687);
xor U16459 (N_16459,N_15807,N_15878);
nor U16460 (N_16460,N_15566,N_15703);
or U16461 (N_16461,N_15661,N_15873);
nand U16462 (N_16462,N_15527,N_15697);
or U16463 (N_16463,N_15695,N_15829);
nand U16464 (N_16464,N_15884,N_15677);
and U16465 (N_16465,N_15591,N_15553);
nand U16466 (N_16466,N_15997,N_15870);
and U16467 (N_16467,N_15543,N_15930);
or U16468 (N_16468,N_15645,N_15505);
nor U16469 (N_16469,N_15504,N_15690);
xnor U16470 (N_16470,N_15817,N_15919);
and U16471 (N_16471,N_15500,N_15875);
nor U16472 (N_16472,N_15803,N_15559);
or U16473 (N_16473,N_15581,N_15797);
xor U16474 (N_16474,N_15747,N_15782);
nor U16475 (N_16475,N_15990,N_15985);
nor U16476 (N_16476,N_15623,N_15939);
or U16477 (N_16477,N_15544,N_15852);
or U16478 (N_16478,N_15622,N_15965);
and U16479 (N_16479,N_15568,N_15521);
nand U16480 (N_16480,N_15966,N_15883);
xnor U16481 (N_16481,N_15977,N_15714);
nor U16482 (N_16482,N_15747,N_15728);
nand U16483 (N_16483,N_15562,N_15660);
xor U16484 (N_16484,N_15541,N_15899);
and U16485 (N_16485,N_15656,N_15686);
and U16486 (N_16486,N_15521,N_15923);
nor U16487 (N_16487,N_15927,N_15644);
or U16488 (N_16488,N_15547,N_15851);
or U16489 (N_16489,N_15993,N_15840);
nand U16490 (N_16490,N_15707,N_15639);
nor U16491 (N_16491,N_15532,N_15892);
and U16492 (N_16492,N_15551,N_15639);
nand U16493 (N_16493,N_15590,N_15751);
nor U16494 (N_16494,N_15528,N_15737);
or U16495 (N_16495,N_15912,N_15600);
and U16496 (N_16496,N_15915,N_15923);
or U16497 (N_16497,N_15526,N_15814);
nand U16498 (N_16498,N_15692,N_15565);
and U16499 (N_16499,N_15758,N_15757);
nand U16500 (N_16500,N_16429,N_16204);
nand U16501 (N_16501,N_16348,N_16147);
nor U16502 (N_16502,N_16279,N_16412);
or U16503 (N_16503,N_16100,N_16109);
nand U16504 (N_16504,N_16413,N_16395);
nor U16505 (N_16505,N_16058,N_16067);
nand U16506 (N_16506,N_16486,N_16146);
nor U16507 (N_16507,N_16021,N_16115);
nand U16508 (N_16508,N_16207,N_16469);
and U16509 (N_16509,N_16209,N_16051);
nor U16510 (N_16510,N_16497,N_16337);
or U16511 (N_16511,N_16231,N_16088);
nor U16512 (N_16512,N_16199,N_16305);
xnor U16513 (N_16513,N_16011,N_16349);
or U16514 (N_16514,N_16483,N_16151);
xnor U16515 (N_16515,N_16158,N_16030);
and U16516 (N_16516,N_16422,N_16185);
nand U16517 (N_16517,N_16291,N_16217);
and U16518 (N_16518,N_16474,N_16317);
or U16519 (N_16519,N_16376,N_16138);
nor U16520 (N_16520,N_16351,N_16297);
and U16521 (N_16521,N_16073,N_16491);
or U16522 (N_16522,N_16382,N_16066);
or U16523 (N_16523,N_16284,N_16262);
and U16524 (N_16524,N_16300,N_16442);
xnor U16525 (N_16525,N_16356,N_16290);
and U16526 (N_16526,N_16293,N_16229);
xnor U16527 (N_16527,N_16467,N_16246);
or U16528 (N_16528,N_16411,N_16294);
and U16529 (N_16529,N_16244,N_16122);
or U16530 (N_16530,N_16312,N_16225);
nand U16531 (N_16531,N_16424,N_16368);
and U16532 (N_16532,N_16272,N_16227);
nor U16533 (N_16533,N_16091,N_16380);
and U16534 (N_16534,N_16438,N_16040);
and U16535 (N_16535,N_16069,N_16439);
or U16536 (N_16536,N_16488,N_16035);
nor U16537 (N_16537,N_16453,N_16235);
or U16538 (N_16538,N_16492,N_16403);
nand U16539 (N_16539,N_16302,N_16077);
nand U16540 (N_16540,N_16134,N_16277);
nand U16541 (N_16541,N_16287,N_16344);
nor U16542 (N_16542,N_16331,N_16318);
xor U16543 (N_16543,N_16308,N_16280);
nor U16544 (N_16544,N_16118,N_16081);
nand U16545 (N_16545,N_16187,N_16445);
nand U16546 (N_16546,N_16420,N_16216);
nand U16547 (N_16547,N_16096,N_16360);
nor U16548 (N_16548,N_16477,N_16201);
nor U16549 (N_16549,N_16464,N_16027);
and U16550 (N_16550,N_16196,N_16385);
and U16551 (N_16551,N_16044,N_16084);
and U16552 (N_16552,N_16493,N_16458);
nand U16553 (N_16553,N_16093,N_16128);
nand U16554 (N_16554,N_16316,N_16325);
or U16555 (N_16555,N_16019,N_16400);
nand U16556 (N_16556,N_16462,N_16392);
or U16557 (N_16557,N_16228,N_16259);
or U16558 (N_16558,N_16358,N_16215);
xor U16559 (N_16559,N_16264,N_16029);
xnor U16560 (N_16560,N_16393,N_16127);
nand U16561 (N_16561,N_16188,N_16136);
and U16562 (N_16562,N_16328,N_16074);
nor U16563 (N_16563,N_16242,N_16489);
xor U16564 (N_16564,N_16025,N_16444);
xnor U16565 (N_16565,N_16432,N_16056);
or U16566 (N_16566,N_16310,N_16042);
nand U16567 (N_16567,N_16336,N_16140);
nand U16568 (N_16568,N_16105,N_16343);
xnor U16569 (N_16569,N_16386,N_16252);
and U16570 (N_16570,N_16065,N_16114);
xor U16571 (N_16571,N_16379,N_16017);
nor U16572 (N_16572,N_16320,N_16145);
xnor U16573 (N_16573,N_16452,N_16388);
xor U16574 (N_16574,N_16164,N_16237);
and U16575 (N_16575,N_16226,N_16457);
or U16576 (N_16576,N_16223,N_16407);
and U16577 (N_16577,N_16428,N_16311);
or U16578 (N_16578,N_16482,N_16046);
and U16579 (N_16579,N_16039,N_16345);
nor U16580 (N_16580,N_16406,N_16057);
nand U16581 (N_16581,N_16346,N_16431);
or U16582 (N_16582,N_16273,N_16433);
nand U16583 (N_16583,N_16110,N_16381);
nor U16584 (N_16584,N_16068,N_16212);
or U16585 (N_16585,N_16255,N_16000);
nand U16586 (N_16586,N_16248,N_16132);
and U16587 (N_16587,N_16022,N_16135);
nand U16588 (N_16588,N_16269,N_16236);
nor U16589 (N_16589,N_16072,N_16218);
and U16590 (N_16590,N_16309,N_16090);
or U16591 (N_16591,N_16026,N_16409);
nor U16592 (N_16592,N_16028,N_16276);
xor U16593 (N_16593,N_16113,N_16166);
nor U16594 (N_16594,N_16327,N_16447);
or U16595 (N_16595,N_16408,N_16001);
nor U16596 (N_16596,N_16338,N_16366);
and U16597 (N_16597,N_16171,N_16283);
nand U16598 (N_16598,N_16373,N_16275);
nor U16599 (N_16599,N_16485,N_16377);
nor U16600 (N_16600,N_16410,N_16415);
nand U16601 (N_16601,N_16052,N_16043);
nor U16602 (N_16602,N_16150,N_16210);
nand U16603 (N_16603,N_16154,N_16459);
and U16604 (N_16604,N_16195,N_16045);
or U16605 (N_16605,N_16258,N_16031);
xor U16606 (N_16606,N_16002,N_16103);
nor U16607 (N_16607,N_16354,N_16288);
nand U16608 (N_16608,N_16323,N_16430);
xor U16609 (N_16609,N_16086,N_16170);
and U16610 (N_16610,N_16121,N_16004);
nor U16611 (N_16611,N_16374,N_16123);
or U16612 (N_16612,N_16340,N_16324);
nand U16613 (N_16613,N_16174,N_16125);
or U16614 (N_16614,N_16361,N_16448);
nand U16615 (N_16615,N_16167,N_16142);
or U16616 (N_16616,N_16478,N_16451);
nor U16617 (N_16617,N_16414,N_16062);
and U16618 (N_16618,N_16268,N_16071);
and U16619 (N_16619,N_16461,N_16394);
nand U16620 (N_16620,N_16137,N_16080);
and U16621 (N_16621,N_16243,N_16033);
nand U16622 (N_16622,N_16494,N_16261);
nor U16623 (N_16623,N_16397,N_16296);
nor U16624 (N_16624,N_16423,N_16247);
nand U16625 (N_16625,N_16334,N_16363);
xor U16626 (N_16626,N_16401,N_16214);
and U16627 (N_16627,N_16260,N_16139);
nor U16628 (N_16628,N_16176,N_16319);
xor U16629 (N_16629,N_16342,N_16326);
nor U16630 (N_16630,N_16463,N_16211);
and U16631 (N_16631,N_16330,N_16203);
or U16632 (N_16632,N_16208,N_16435);
nor U16633 (N_16633,N_16239,N_16119);
nor U16634 (N_16634,N_16107,N_16177);
xor U16635 (N_16635,N_16092,N_16498);
xnor U16636 (N_16636,N_16220,N_16322);
or U16637 (N_16637,N_16153,N_16369);
and U16638 (N_16638,N_16362,N_16111);
and U16639 (N_16639,N_16253,N_16126);
nor U16640 (N_16640,N_16129,N_16499);
or U16641 (N_16641,N_16353,N_16417);
xnor U16642 (N_16642,N_16321,N_16249);
or U16643 (N_16643,N_16180,N_16120);
nor U16644 (N_16644,N_16152,N_16335);
and U16645 (N_16645,N_16426,N_16131);
and U16646 (N_16646,N_16257,N_16101);
xor U16647 (N_16647,N_16018,N_16263);
or U16648 (N_16648,N_16076,N_16198);
nor U16649 (N_16649,N_16173,N_16367);
nor U16650 (N_16650,N_16020,N_16148);
xor U16651 (N_16651,N_16289,N_16405);
or U16652 (N_16652,N_16479,N_16099);
xor U16653 (N_16653,N_16161,N_16292);
nor U16654 (N_16654,N_16496,N_16034);
nand U16655 (N_16655,N_16265,N_16443);
and U16656 (N_16656,N_16314,N_16238);
xor U16657 (N_16657,N_16281,N_16476);
or U16658 (N_16658,N_16475,N_16450);
nor U16659 (N_16659,N_16172,N_16008);
or U16660 (N_16660,N_16102,N_16495);
or U16661 (N_16661,N_16456,N_16285);
and U16662 (N_16662,N_16425,N_16094);
nand U16663 (N_16663,N_16159,N_16224);
nor U16664 (N_16664,N_16160,N_16181);
nand U16665 (N_16665,N_16014,N_16041);
nor U16666 (N_16666,N_16064,N_16012);
or U16667 (N_16667,N_16480,N_16295);
xnor U16668 (N_16668,N_16434,N_16047);
xor U16669 (N_16669,N_16192,N_16390);
and U16670 (N_16670,N_16075,N_16191);
and U16671 (N_16671,N_16329,N_16481);
and U16672 (N_16672,N_16149,N_16465);
nor U16673 (N_16673,N_16083,N_16350);
xnor U16674 (N_16674,N_16383,N_16054);
and U16675 (N_16675,N_16355,N_16155);
or U16676 (N_16676,N_16274,N_16055);
xnor U16677 (N_16677,N_16095,N_16440);
nor U16678 (N_16678,N_16182,N_16230);
xnor U16679 (N_16679,N_16124,N_16163);
nor U16680 (N_16680,N_16162,N_16384);
nor U16681 (N_16681,N_16063,N_16112);
and U16682 (N_16682,N_16468,N_16282);
xnor U16683 (N_16683,N_16206,N_16190);
or U16684 (N_16684,N_16036,N_16251);
and U16685 (N_16685,N_16396,N_16009);
nor U16686 (N_16686,N_16427,N_16306);
or U16687 (N_16687,N_16378,N_16232);
nor U16688 (N_16688,N_16003,N_16298);
nand U16689 (N_16689,N_16446,N_16179);
nand U16690 (N_16690,N_16490,N_16472);
and U16691 (N_16691,N_16078,N_16133);
nand U16692 (N_16692,N_16303,N_16389);
nand U16693 (N_16693,N_16471,N_16089);
xnor U16694 (N_16694,N_16024,N_16202);
xnor U16695 (N_16695,N_16304,N_16183);
nand U16696 (N_16696,N_16193,N_16240);
nand U16697 (N_16697,N_16016,N_16184);
xnor U16698 (N_16698,N_16038,N_16416);
xor U16699 (N_16699,N_16418,N_16359);
xnor U16700 (N_16700,N_16387,N_16347);
or U16701 (N_16701,N_16286,N_16254);
and U16702 (N_16702,N_16157,N_16398);
xor U16703 (N_16703,N_16484,N_16301);
nand U16704 (N_16704,N_16333,N_16130);
or U16705 (N_16705,N_16194,N_16156);
xor U16706 (N_16706,N_16106,N_16189);
or U16707 (N_16707,N_16050,N_16460);
and U16708 (N_16708,N_16233,N_16267);
and U16709 (N_16709,N_16271,N_16175);
or U16710 (N_16710,N_16085,N_16010);
xor U16711 (N_16711,N_16487,N_16013);
or U16712 (N_16712,N_16169,N_16200);
nor U16713 (N_16713,N_16313,N_16372);
and U16714 (N_16714,N_16339,N_16473);
nor U16715 (N_16715,N_16007,N_16219);
and U16716 (N_16716,N_16245,N_16061);
nand U16717 (N_16717,N_16168,N_16186);
xnor U16718 (N_16718,N_16421,N_16278);
and U16719 (N_16719,N_16116,N_16234);
xor U16720 (N_16720,N_16441,N_16332);
nand U16721 (N_16721,N_16087,N_16023);
xnor U16722 (N_16722,N_16391,N_16419);
or U16723 (N_16723,N_16082,N_16352);
nand U16724 (N_16724,N_16375,N_16037);
and U16725 (N_16725,N_16222,N_16365);
nor U16726 (N_16726,N_16032,N_16404);
nand U16727 (N_16727,N_16466,N_16307);
or U16728 (N_16728,N_16049,N_16048);
or U16729 (N_16729,N_16470,N_16165);
and U16730 (N_16730,N_16006,N_16144);
and U16731 (N_16731,N_16059,N_16449);
nand U16732 (N_16732,N_16436,N_16437);
xnor U16733 (N_16733,N_16060,N_16299);
nor U16734 (N_16734,N_16221,N_16399);
or U16735 (N_16735,N_16108,N_16371);
xor U16736 (N_16736,N_16213,N_16370);
and U16737 (N_16737,N_16005,N_16250);
nand U16738 (N_16738,N_16256,N_16141);
nor U16739 (N_16739,N_16315,N_16117);
nor U16740 (N_16740,N_16454,N_16053);
xnor U16741 (N_16741,N_16079,N_16015);
nand U16742 (N_16742,N_16178,N_16270);
xor U16743 (N_16743,N_16143,N_16197);
nand U16744 (N_16744,N_16364,N_16357);
or U16745 (N_16745,N_16341,N_16097);
nand U16746 (N_16746,N_16070,N_16455);
nand U16747 (N_16747,N_16241,N_16402);
and U16748 (N_16748,N_16098,N_16205);
or U16749 (N_16749,N_16266,N_16104);
nor U16750 (N_16750,N_16436,N_16190);
and U16751 (N_16751,N_16265,N_16108);
xnor U16752 (N_16752,N_16226,N_16277);
or U16753 (N_16753,N_16020,N_16309);
and U16754 (N_16754,N_16099,N_16469);
or U16755 (N_16755,N_16151,N_16262);
nor U16756 (N_16756,N_16361,N_16216);
xnor U16757 (N_16757,N_16391,N_16055);
nor U16758 (N_16758,N_16025,N_16282);
nor U16759 (N_16759,N_16368,N_16413);
and U16760 (N_16760,N_16188,N_16322);
xnor U16761 (N_16761,N_16255,N_16191);
or U16762 (N_16762,N_16318,N_16270);
or U16763 (N_16763,N_16419,N_16013);
or U16764 (N_16764,N_16098,N_16252);
or U16765 (N_16765,N_16234,N_16123);
nor U16766 (N_16766,N_16415,N_16307);
and U16767 (N_16767,N_16266,N_16445);
nor U16768 (N_16768,N_16183,N_16387);
and U16769 (N_16769,N_16478,N_16115);
nand U16770 (N_16770,N_16412,N_16483);
and U16771 (N_16771,N_16069,N_16109);
nor U16772 (N_16772,N_16024,N_16395);
and U16773 (N_16773,N_16169,N_16129);
xnor U16774 (N_16774,N_16023,N_16085);
nand U16775 (N_16775,N_16416,N_16121);
and U16776 (N_16776,N_16063,N_16430);
and U16777 (N_16777,N_16241,N_16465);
xnor U16778 (N_16778,N_16186,N_16094);
xnor U16779 (N_16779,N_16289,N_16473);
nor U16780 (N_16780,N_16073,N_16107);
nor U16781 (N_16781,N_16303,N_16160);
xor U16782 (N_16782,N_16078,N_16307);
or U16783 (N_16783,N_16196,N_16383);
nand U16784 (N_16784,N_16240,N_16369);
xnor U16785 (N_16785,N_16057,N_16096);
or U16786 (N_16786,N_16242,N_16182);
xor U16787 (N_16787,N_16338,N_16178);
nand U16788 (N_16788,N_16409,N_16121);
nand U16789 (N_16789,N_16345,N_16464);
or U16790 (N_16790,N_16378,N_16436);
nor U16791 (N_16791,N_16009,N_16270);
nand U16792 (N_16792,N_16216,N_16329);
nor U16793 (N_16793,N_16463,N_16215);
or U16794 (N_16794,N_16463,N_16147);
and U16795 (N_16795,N_16192,N_16269);
xor U16796 (N_16796,N_16292,N_16173);
xor U16797 (N_16797,N_16089,N_16403);
xnor U16798 (N_16798,N_16387,N_16118);
or U16799 (N_16799,N_16077,N_16191);
nor U16800 (N_16800,N_16343,N_16115);
nand U16801 (N_16801,N_16064,N_16346);
nor U16802 (N_16802,N_16283,N_16480);
xor U16803 (N_16803,N_16442,N_16269);
nand U16804 (N_16804,N_16290,N_16382);
and U16805 (N_16805,N_16293,N_16228);
and U16806 (N_16806,N_16236,N_16127);
nor U16807 (N_16807,N_16260,N_16351);
xnor U16808 (N_16808,N_16089,N_16133);
nor U16809 (N_16809,N_16445,N_16175);
or U16810 (N_16810,N_16100,N_16388);
nor U16811 (N_16811,N_16420,N_16277);
xor U16812 (N_16812,N_16127,N_16026);
nor U16813 (N_16813,N_16039,N_16037);
and U16814 (N_16814,N_16149,N_16213);
or U16815 (N_16815,N_16136,N_16050);
nor U16816 (N_16816,N_16308,N_16055);
nor U16817 (N_16817,N_16129,N_16073);
and U16818 (N_16818,N_16102,N_16237);
xnor U16819 (N_16819,N_16389,N_16159);
nor U16820 (N_16820,N_16157,N_16426);
and U16821 (N_16821,N_16134,N_16488);
nor U16822 (N_16822,N_16359,N_16111);
nand U16823 (N_16823,N_16298,N_16011);
xnor U16824 (N_16824,N_16073,N_16056);
nand U16825 (N_16825,N_16217,N_16298);
and U16826 (N_16826,N_16022,N_16371);
or U16827 (N_16827,N_16450,N_16200);
or U16828 (N_16828,N_16017,N_16197);
nor U16829 (N_16829,N_16044,N_16188);
and U16830 (N_16830,N_16231,N_16009);
nand U16831 (N_16831,N_16397,N_16328);
nand U16832 (N_16832,N_16432,N_16487);
and U16833 (N_16833,N_16461,N_16095);
nor U16834 (N_16834,N_16026,N_16398);
nand U16835 (N_16835,N_16237,N_16498);
nand U16836 (N_16836,N_16218,N_16019);
and U16837 (N_16837,N_16056,N_16209);
and U16838 (N_16838,N_16338,N_16121);
nand U16839 (N_16839,N_16199,N_16396);
nor U16840 (N_16840,N_16379,N_16277);
nand U16841 (N_16841,N_16259,N_16433);
nand U16842 (N_16842,N_16253,N_16089);
nor U16843 (N_16843,N_16034,N_16392);
xor U16844 (N_16844,N_16052,N_16346);
xnor U16845 (N_16845,N_16207,N_16354);
nor U16846 (N_16846,N_16195,N_16492);
or U16847 (N_16847,N_16340,N_16297);
and U16848 (N_16848,N_16292,N_16132);
and U16849 (N_16849,N_16264,N_16364);
nand U16850 (N_16850,N_16336,N_16348);
nand U16851 (N_16851,N_16474,N_16173);
nor U16852 (N_16852,N_16287,N_16460);
nor U16853 (N_16853,N_16087,N_16414);
or U16854 (N_16854,N_16068,N_16176);
nand U16855 (N_16855,N_16265,N_16163);
nor U16856 (N_16856,N_16415,N_16271);
nand U16857 (N_16857,N_16175,N_16412);
nand U16858 (N_16858,N_16285,N_16108);
nand U16859 (N_16859,N_16016,N_16077);
and U16860 (N_16860,N_16207,N_16189);
and U16861 (N_16861,N_16218,N_16144);
and U16862 (N_16862,N_16231,N_16115);
nor U16863 (N_16863,N_16325,N_16025);
nor U16864 (N_16864,N_16359,N_16014);
and U16865 (N_16865,N_16200,N_16167);
or U16866 (N_16866,N_16282,N_16392);
nand U16867 (N_16867,N_16154,N_16402);
xor U16868 (N_16868,N_16435,N_16206);
nand U16869 (N_16869,N_16063,N_16176);
and U16870 (N_16870,N_16356,N_16173);
and U16871 (N_16871,N_16106,N_16386);
nand U16872 (N_16872,N_16073,N_16271);
and U16873 (N_16873,N_16345,N_16143);
and U16874 (N_16874,N_16323,N_16046);
nand U16875 (N_16875,N_16125,N_16178);
xnor U16876 (N_16876,N_16415,N_16405);
and U16877 (N_16877,N_16330,N_16120);
nand U16878 (N_16878,N_16147,N_16014);
and U16879 (N_16879,N_16422,N_16137);
nand U16880 (N_16880,N_16034,N_16029);
or U16881 (N_16881,N_16422,N_16144);
xor U16882 (N_16882,N_16121,N_16472);
nand U16883 (N_16883,N_16147,N_16315);
and U16884 (N_16884,N_16131,N_16452);
and U16885 (N_16885,N_16146,N_16131);
nand U16886 (N_16886,N_16079,N_16061);
or U16887 (N_16887,N_16196,N_16063);
xnor U16888 (N_16888,N_16191,N_16347);
nor U16889 (N_16889,N_16343,N_16308);
nand U16890 (N_16890,N_16191,N_16267);
xnor U16891 (N_16891,N_16315,N_16482);
nor U16892 (N_16892,N_16108,N_16302);
nor U16893 (N_16893,N_16100,N_16081);
xnor U16894 (N_16894,N_16273,N_16197);
and U16895 (N_16895,N_16108,N_16391);
and U16896 (N_16896,N_16088,N_16488);
nand U16897 (N_16897,N_16294,N_16275);
and U16898 (N_16898,N_16030,N_16155);
and U16899 (N_16899,N_16155,N_16275);
and U16900 (N_16900,N_16422,N_16386);
nor U16901 (N_16901,N_16218,N_16058);
nand U16902 (N_16902,N_16029,N_16162);
nor U16903 (N_16903,N_16275,N_16240);
or U16904 (N_16904,N_16276,N_16045);
or U16905 (N_16905,N_16241,N_16369);
xnor U16906 (N_16906,N_16260,N_16246);
xor U16907 (N_16907,N_16394,N_16330);
xor U16908 (N_16908,N_16328,N_16140);
and U16909 (N_16909,N_16327,N_16332);
or U16910 (N_16910,N_16054,N_16120);
or U16911 (N_16911,N_16196,N_16118);
and U16912 (N_16912,N_16029,N_16105);
xnor U16913 (N_16913,N_16255,N_16032);
xnor U16914 (N_16914,N_16116,N_16484);
or U16915 (N_16915,N_16149,N_16273);
or U16916 (N_16916,N_16322,N_16405);
or U16917 (N_16917,N_16491,N_16467);
xnor U16918 (N_16918,N_16071,N_16270);
nor U16919 (N_16919,N_16354,N_16186);
nor U16920 (N_16920,N_16140,N_16201);
nand U16921 (N_16921,N_16164,N_16042);
nor U16922 (N_16922,N_16120,N_16023);
nor U16923 (N_16923,N_16443,N_16354);
or U16924 (N_16924,N_16355,N_16315);
xor U16925 (N_16925,N_16176,N_16128);
and U16926 (N_16926,N_16163,N_16015);
xnor U16927 (N_16927,N_16323,N_16367);
and U16928 (N_16928,N_16021,N_16440);
or U16929 (N_16929,N_16452,N_16001);
and U16930 (N_16930,N_16384,N_16294);
xor U16931 (N_16931,N_16080,N_16302);
or U16932 (N_16932,N_16357,N_16235);
and U16933 (N_16933,N_16438,N_16042);
xnor U16934 (N_16934,N_16449,N_16472);
nand U16935 (N_16935,N_16099,N_16482);
or U16936 (N_16936,N_16155,N_16130);
nor U16937 (N_16937,N_16177,N_16001);
and U16938 (N_16938,N_16248,N_16215);
nand U16939 (N_16939,N_16026,N_16317);
or U16940 (N_16940,N_16481,N_16293);
and U16941 (N_16941,N_16048,N_16229);
nand U16942 (N_16942,N_16410,N_16360);
nand U16943 (N_16943,N_16089,N_16395);
xor U16944 (N_16944,N_16063,N_16497);
nor U16945 (N_16945,N_16087,N_16491);
xor U16946 (N_16946,N_16209,N_16080);
xnor U16947 (N_16947,N_16401,N_16024);
or U16948 (N_16948,N_16334,N_16001);
xor U16949 (N_16949,N_16470,N_16125);
xor U16950 (N_16950,N_16366,N_16459);
nor U16951 (N_16951,N_16271,N_16385);
nand U16952 (N_16952,N_16294,N_16041);
and U16953 (N_16953,N_16257,N_16046);
and U16954 (N_16954,N_16218,N_16289);
and U16955 (N_16955,N_16369,N_16198);
nand U16956 (N_16956,N_16175,N_16275);
or U16957 (N_16957,N_16469,N_16070);
nand U16958 (N_16958,N_16173,N_16428);
or U16959 (N_16959,N_16094,N_16312);
and U16960 (N_16960,N_16162,N_16172);
nor U16961 (N_16961,N_16034,N_16306);
or U16962 (N_16962,N_16497,N_16085);
nor U16963 (N_16963,N_16256,N_16333);
and U16964 (N_16964,N_16000,N_16345);
nor U16965 (N_16965,N_16466,N_16360);
xor U16966 (N_16966,N_16487,N_16193);
nor U16967 (N_16967,N_16203,N_16301);
nand U16968 (N_16968,N_16351,N_16061);
xnor U16969 (N_16969,N_16324,N_16143);
nand U16970 (N_16970,N_16073,N_16401);
and U16971 (N_16971,N_16153,N_16079);
nand U16972 (N_16972,N_16041,N_16023);
nor U16973 (N_16973,N_16443,N_16278);
xnor U16974 (N_16974,N_16456,N_16095);
nor U16975 (N_16975,N_16067,N_16414);
nor U16976 (N_16976,N_16462,N_16430);
nand U16977 (N_16977,N_16006,N_16021);
or U16978 (N_16978,N_16071,N_16008);
nand U16979 (N_16979,N_16066,N_16158);
and U16980 (N_16980,N_16002,N_16482);
nand U16981 (N_16981,N_16134,N_16153);
and U16982 (N_16982,N_16203,N_16194);
xnor U16983 (N_16983,N_16232,N_16379);
nand U16984 (N_16984,N_16292,N_16414);
nor U16985 (N_16985,N_16338,N_16439);
or U16986 (N_16986,N_16490,N_16437);
and U16987 (N_16987,N_16396,N_16383);
nor U16988 (N_16988,N_16286,N_16152);
nand U16989 (N_16989,N_16248,N_16079);
nand U16990 (N_16990,N_16332,N_16178);
nor U16991 (N_16991,N_16486,N_16481);
nand U16992 (N_16992,N_16116,N_16486);
xnor U16993 (N_16993,N_16097,N_16406);
or U16994 (N_16994,N_16493,N_16326);
nor U16995 (N_16995,N_16113,N_16176);
nand U16996 (N_16996,N_16330,N_16168);
nand U16997 (N_16997,N_16444,N_16036);
nor U16998 (N_16998,N_16269,N_16239);
xnor U16999 (N_16999,N_16484,N_16079);
or U17000 (N_17000,N_16829,N_16690);
nand U17001 (N_17001,N_16992,N_16824);
or U17002 (N_17002,N_16589,N_16865);
xor U17003 (N_17003,N_16750,N_16915);
xnor U17004 (N_17004,N_16518,N_16601);
and U17005 (N_17005,N_16925,N_16657);
nand U17006 (N_17006,N_16924,N_16831);
and U17007 (N_17007,N_16728,N_16999);
and U17008 (N_17008,N_16904,N_16959);
nor U17009 (N_17009,N_16563,N_16774);
nor U17010 (N_17010,N_16797,N_16997);
nand U17011 (N_17011,N_16842,N_16650);
nand U17012 (N_17012,N_16662,N_16964);
and U17013 (N_17013,N_16530,N_16920);
nor U17014 (N_17014,N_16562,N_16729);
nand U17015 (N_17015,N_16653,N_16916);
or U17016 (N_17016,N_16626,N_16863);
xor U17017 (N_17017,N_16605,N_16591);
and U17018 (N_17018,N_16879,N_16509);
nor U17019 (N_17019,N_16955,N_16980);
and U17020 (N_17020,N_16620,N_16779);
nor U17021 (N_17021,N_16917,N_16841);
nand U17022 (N_17022,N_16953,N_16641);
or U17023 (N_17023,N_16813,N_16952);
xnor U17024 (N_17024,N_16806,N_16903);
nand U17025 (N_17025,N_16547,N_16584);
or U17026 (N_17026,N_16968,N_16646);
nand U17027 (N_17027,N_16988,N_16642);
and U17028 (N_17028,N_16840,N_16960);
xor U17029 (N_17029,N_16738,N_16748);
nor U17030 (N_17030,N_16501,N_16633);
xor U17031 (N_17031,N_16719,N_16782);
nand U17032 (N_17032,N_16614,N_16781);
or U17033 (N_17033,N_16585,N_16943);
nor U17034 (N_17034,N_16812,N_16613);
and U17035 (N_17035,N_16640,N_16730);
and U17036 (N_17036,N_16686,N_16818);
and U17037 (N_17037,N_16921,N_16820);
or U17038 (N_17038,N_16939,N_16993);
or U17039 (N_17039,N_16823,N_16805);
xnor U17040 (N_17040,N_16891,N_16977);
nor U17041 (N_17041,N_16809,N_16656);
or U17042 (N_17042,N_16691,N_16886);
xor U17043 (N_17043,N_16660,N_16994);
nor U17044 (N_17044,N_16654,N_16767);
or U17045 (N_17045,N_16757,N_16510);
nor U17046 (N_17046,N_16529,N_16937);
or U17047 (N_17047,N_16864,N_16958);
xor U17048 (N_17048,N_16696,N_16976);
nand U17049 (N_17049,N_16735,N_16555);
nand U17050 (N_17050,N_16918,N_16670);
or U17051 (N_17051,N_16740,N_16768);
and U17052 (N_17052,N_16710,N_16896);
and U17053 (N_17053,N_16931,N_16972);
or U17054 (N_17054,N_16847,N_16693);
nor U17055 (N_17055,N_16618,N_16973);
xor U17056 (N_17056,N_16553,N_16786);
and U17057 (N_17057,N_16857,N_16926);
and U17058 (N_17058,N_16877,N_16844);
and U17059 (N_17059,N_16705,N_16861);
nor U17060 (N_17060,N_16900,N_16734);
or U17061 (N_17061,N_16628,N_16834);
nand U17062 (N_17062,N_16808,N_16636);
xnor U17063 (N_17063,N_16989,N_16739);
or U17064 (N_17064,N_16957,N_16694);
or U17065 (N_17065,N_16575,N_16982);
or U17066 (N_17066,N_16978,N_16720);
nand U17067 (N_17067,N_16607,N_16707);
nor U17068 (N_17068,N_16761,N_16559);
and U17069 (N_17069,N_16769,N_16528);
xor U17070 (N_17070,N_16838,N_16600);
nand U17071 (N_17071,N_16552,N_16764);
or U17072 (N_17072,N_16661,N_16651);
nor U17073 (N_17073,N_16744,N_16872);
nand U17074 (N_17074,N_16731,N_16550);
nand U17075 (N_17075,N_16860,N_16602);
or U17076 (N_17076,N_16914,N_16579);
nor U17077 (N_17077,N_16790,N_16793);
and U17078 (N_17078,N_16679,N_16548);
and U17079 (N_17079,N_16996,N_16565);
nand U17080 (N_17080,N_16827,N_16783);
nor U17081 (N_17081,N_16839,N_16540);
or U17082 (N_17082,N_16658,N_16810);
or U17083 (N_17083,N_16507,N_16789);
or U17084 (N_17084,N_16909,N_16560);
and U17085 (N_17085,N_16544,N_16723);
nand U17086 (N_17086,N_16913,N_16668);
nor U17087 (N_17087,N_16522,N_16755);
or U17088 (N_17088,N_16527,N_16950);
or U17089 (N_17089,N_16692,N_16675);
xor U17090 (N_17090,N_16711,N_16749);
or U17091 (N_17091,N_16811,N_16845);
nor U17092 (N_17092,N_16951,N_16816);
xor U17093 (N_17093,N_16590,N_16532);
and U17094 (N_17094,N_16667,N_16780);
nand U17095 (N_17095,N_16569,N_16718);
nor U17096 (N_17096,N_16502,N_16644);
and U17097 (N_17097,N_16849,N_16724);
and U17098 (N_17098,N_16526,N_16936);
xor U17099 (N_17099,N_16851,N_16508);
nand U17100 (N_17100,N_16583,N_16715);
and U17101 (N_17101,N_16500,N_16520);
nand U17102 (N_17102,N_16868,N_16700);
or U17103 (N_17103,N_16677,N_16762);
xor U17104 (N_17104,N_16716,N_16514);
nand U17105 (N_17105,N_16615,N_16745);
xor U17106 (N_17106,N_16776,N_16676);
nand U17107 (N_17107,N_16948,N_16524);
xnor U17108 (N_17108,N_16846,N_16963);
or U17109 (N_17109,N_16717,N_16746);
and U17110 (N_17110,N_16558,N_16604);
and U17111 (N_17111,N_16645,N_16611);
xor U17112 (N_17112,N_16892,N_16938);
or U17113 (N_17113,N_16732,N_16832);
and U17114 (N_17114,N_16855,N_16525);
nor U17115 (N_17115,N_16850,N_16534);
nand U17116 (N_17116,N_16619,N_16798);
and U17117 (N_17117,N_16856,N_16754);
nand U17118 (N_17118,N_16687,N_16815);
and U17119 (N_17119,N_16801,N_16582);
nor U17120 (N_17120,N_16505,N_16616);
nand U17121 (N_17121,N_16617,N_16803);
and U17122 (N_17122,N_16947,N_16802);
xnor U17123 (N_17123,N_16567,N_16852);
xor U17124 (N_17124,N_16987,N_16946);
and U17125 (N_17125,N_16698,N_16597);
or U17126 (N_17126,N_16871,N_16737);
and U17127 (N_17127,N_16566,N_16956);
nand U17128 (N_17128,N_16873,N_16685);
and U17129 (N_17129,N_16772,N_16709);
nor U17130 (N_17130,N_16941,N_16674);
nand U17131 (N_17131,N_16659,N_16577);
nor U17132 (N_17132,N_16893,N_16919);
nor U17133 (N_17133,N_16539,N_16778);
xor U17134 (N_17134,N_16609,N_16983);
nand U17135 (N_17135,N_16549,N_16874);
nor U17136 (N_17136,N_16859,N_16817);
nand U17137 (N_17137,N_16837,N_16875);
nor U17138 (N_17138,N_16683,N_16912);
xnor U17139 (N_17139,N_16537,N_16635);
nor U17140 (N_17140,N_16869,N_16760);
nor U17141 (N_17141,N_16966,N_16985);
or U17142 (N_17142,N_16504,N_16631);
nand U17143 (N_17143,N_16519,N_16800);
nor U17144 (N_17144,N_16627,N_16954);
or U17145 (N_17145,N_16536,N_16557);
and U17146 (N_17146,N_16703,N_16799);
nand U17147 (N_17147,N_16721,N_16521);
or U17148 (N_17148,N_16588,N_16680);
xor U17149 (N_17149,N_16511,N_16922);
nand U17150 (N_17150,N_16796,N_16682);
nor U17151 (N_17151,N_16830,N_16759);
or U17152 (N_17152,N_16777,N_16571);
and U17153 (N_17153,N_16974,N_16541);
xor U17154 (N_17154,N_16971,N_16833);
or U17155 (N_17155,N_16699,N_16940);
and U17156 (N_17156,N_16867,N_16901);
or U17157 (N_17157,N_16906,N_16836);
or U17158 (N_17158,N_16995,N_16902);
and U17159 (N_17159,N_16932,N_16928);
or U17160 (N_17160,N_16881,N_16681);
xnor U17161 (N_17161,N_16763,N_16606);
or U17162 (N_17162,N_16515,N_16714);
nor U17163 (N_17163,N_16701,N_16625);
nor U17164 (N_17164,N_16791,N_16770);
xor U17165 (N_17165,N_16758,N_16581);
nand U17166 (N_17166,N_16910,N_16826);
or U17167 (N_17167,N_16942,N_16969);
and U17168 (N_17168,N_16962,N_16652);
or U17169 (N_17169,N_16596,N_16773);
xor U17170 (N_17170,N_16848,N_16853);
nand U17171 (N_17171,N_16890,N_16599);
nand U17172 (N_17172,N_16538,N_16570);
nor U17173 (N_17173,N_16756,N_16885);
nand U17174 (N_17174,N_16897,N_16608);
nand U17175 (N_17175,N_16592,N_16632);
xnor U17176 (N_17176,N_16513,N_16543);
xor U17177 (N_17177,N_16672,N_16648);
nand U17178 (N_17178,N_16967,N_16878);
nor U17179 (N_17179,N_16965,N_16533);
xor U17180 (N_17180,N_16678,N_16568);
xor U17181 (N_17181,N_16512,N_16899);
or U17182 (N_17182,N_16843,N_16908);
nand U17183 (N_17183,N_16586,N_16564);
and U17184 (N_17184,N_16784,N_16727);
nand U17185 (N_17185,N_16561,N_16930);
and U17186 (N_17186,N_16907,N_16753);
xor U17187 (N_17187,N_16695,N_16663);
xor U17188 (N_17188,N_16647,N_16911);
and U17189 (N_17189,N_16828,N_16979);
and U17190 (N_17190,N_16580,N_16517);
nor U17191 (N_17191,N_16629,N_16503);
nand U17192 (N_17192,N_16598,N_16637);
or U17193 (N_17193,N_16933,N_16551);
nand U17194 (N_17194,N_16638,N_16702);
or U17195 (N_17195,N_16506,N_16794);
nor U17196 (N_17196,N_16572,N_16889);
or U17197 (N_17197,N_16593,N_16944);
xor U17198 (N_17198,N_16991,N_16788);
or U17199 (N_17199,N_16535,N_16821);
xor U17200 (N_17200,N_16825,N_16895);
nor U17201 (N_17201,N_16523,N_16587);
nor U17202 (N_17202,N_16929,N_16949);
and U17203 (N_17203,N_16733,N_16649);
and U17204 (N_17204,N_16595,N_16574);
or U17205 (N_17205,N_16765,N_16655);
xor U17206 (N_17206,N_16643,N_16634);
xor U17207 (N_17207,N_16858,N_16725);
and U17208 (N_17208,N_16712,N_16981);
or U17209 (N_17209,N_16854,N_16822);
and U17210 (N_17210,N_16751,N_16545);
or U17211 (N_17211,N_16708,N_16706);
xnor U17212 (N_17212,N_16623,N_16819);
nand U17213 (N_17213,N_16887,N_16766);
or U17214 (N_17214,N_16612,N_16870);
or U17215 (N_17215,N_16961,N_16713);
and U17216 (N_17216,N_16945,N_16894);
or U17217 (N_17217,N_16882,N_16923);
nand U17218 (N_17218,N_16876,N_16927);
nor U17219 (N_17219,N_16554,N_16556);
nand U17220 (N_17220,N_16835,N_16984);
and U17221 (N_17221,N_16576,N_16741);
nand U17222 (N_17222,N_16624,N_16630);
xnor U17223 (N_17223,N_16666,N_16747);
nand U17224 (N_17224,N_16888,N_16787);
and U17225 (N_17225,N_16622,N_16664);
and U17226 (N_17226,N_16807,N_16880);
xor U17227 (N_17227,N_16603,N_16722);
xnor U17228 (N_17228,N_16516,N_16986);
xor U17229 (N_17229,N_16688,N_16704);
nor U17230 (N_17230,N_16814,N_16792);
nor U17231 (N_17231,N_16573,N_16785);
nand U17232 (N_17232,N_16742,N_16898);
and U17233 (N_17233,N_16884,N_16697);
and U17234 (N_17234,N_16671,N_16736);
nand U17235 (N_17235,N_16998,N_16970);
xnor U17236 (N_17236,N_16905,N_16684);
or U17237 (N_17237,N_16669,N_16752);
nor U17238 (N_17238,N_16804,N_16990);
or U17239 (N_17239,N_16531,N_16934);
nand U17240 (N_17240,N_16542,N_16883);
and U17241 (N_17241,N_16639,N_16975);
or U17242 (N_17242,N_16621,N_16726);
nor U17243 (N_17243,N_16689,N_16610);
and U17244 (N_17244,N_16673,N_16795);
or U17245 (N_17245,N_16546,N_16594);
xnor U17246 (N_17246,N_16775,N_16862);
and U17247 (N_17247,N_16866,N_16578);
and U17248 (N_17248,N_16743,N_16771);
nand U17249 (N_17249,N_16935,N_16665);
xor U17250 (N_17250,N_16774,N_16760);
xnor U17251 (N_17251,N_16970,N_16529);
nand U17252 (N_17252,N_16979,N_16592);
nand U17253 (N_17253,N_16852,N_16748);
nand U17254 (N_17254,N_16689,N_16845);
xnor U17255 (N_17255,N_16950,N_16863);
xnor U17256 (N_17256,N_16820,N_16702);
and U17257 (N_17257,N_16679,N_16875);
or U17258 (N_17258,N_16729,N_16764);
or U17259 (N_17259,N_16829,N_16976);
xor U17260 (N_17260,N_16964,N_16619);
or U17261 (N_17261,N_16564,N_16515);
or U17262 (N_17262,N_16813,N_16715);
nor U17263 (N_17263,N_16804,N_16699);
nor U17264 (N_17264,N_16513,N_16629);
nor U17265 (N_17265,N_16584,N_16898);
and U17266 (N_17266,N_16953,N_16997);
xnor U17267 (N_17267,N_16851,N_16929);
nand U17268 (N_17268,N_16677,N_16658);
nor U17269 (N_17269,N_16952,N_16662);
and U17270 (N_17270,N_16769,N_16843);
or U17271 (N_17271,N_16897,N_16610);
and U17272 (N_17272,N_16874,N_16665);
and U17273 (N_17273,N_16525,N_16597);
nor U17274 (N_17274,N_16572,N_16588);
nor U17275 (N_17275,N_16553,N_16620);
xnor U17276 (N_17276,N_16986,N_16597);
nor U17277 (N_17277,N_16848,N_16814);
nand U17278 (N_17278,N_16787,N_16866);
xor U17279 (N_17279,N_16815,N_16517);
nor U17280 (N_17280,N_16718,N_16754);
xnor U17281 (N_17281,N_16742,N_16722);
nor U17282 (N_17282,N_16884,N_16721);
nand U17283 (N_17283,N_16863,N_16788);
and U17284 (N_17284,N_16600,N_16612);
or U17285 (N_17285,N_16752,N_16609);
nand U17286 (N_17286,N_16598,N_16870);
or U17287 (N_17287,N_16610,N_16994);
xor U17288 (N_17288,N_16509,N_16613);
or U17289 (N_17289,N_16929,N_16778);
nand U17290 (N_17290,N_16986,N_16696);
nand U17291 (N_17291,N_16671,N_16755);
and U17292 (N_17292,N_16609,N_16734);
xor U17293 (N_17293,N_16931,N_16748);
xnor U17294 (N_17294,N_16866,N_16614);
xnor U17295 (N_17295,N_16648,N_16828);
nand U17296 (N_17296,N_16985,N_16761);
xnor U17297 (N_17297,N_16632,N_16739);
or U17298 (N_17298,N_16856,N_16595);
or U17299 (N_17299,N_16824,N_16853);
xnor U17300 (N_17300,N_16864,N_16912);
nor U17301 (N_17301,N_16584,N_16593);
or U17302 (N_17302,N_16898,N_16992);
nand U17303 (N_17303,N_16511,N_16919);
or U17304 (N_17304,N_16736,N_16917);
nand U17305 (N_17305,N_16574,N_16880);
and U17306 (N_17306,N_16624,N_16620);
xor U17307 (N_17307,N_16690,N_16979);
nor U17308 (N_17308,N_16526,N_16925);
nand U17309 (N_17309,N_16633,N_16622);
or U17310 (N_17310,N_16832,N_16725);
or U17311 (N_17311,N_16696,N_16542);
nor U17312 (N_17312,N_16658,N_16829);
nand U17313 (N_17313,N_16839,N_16643);
or U17314 (N_17314,N_16548,N_16806);
nor U17315 (N_17315,N_16583,N_16828);
nand U17316 (N_17316,N_16949,N_16549);
or U17317 (N_17317,N_16917,N_16892);
xor U17318 (N_17318,N_16895,N_16872);
or U17319 (N_17319,N_16781,N_16678);
and U17320 (N_17320,N_16751,N_16643);
and U17321 (N_17321,N_16522,N_16862);
xnor U17322 (N_17322,N_16725,N_16743);
xor U17323 (N_17323,N_16770,N_16544);
and U17324 (N_17324,N_16524,N_16705);
nand U17325 (N_17325,N_16730,N_16544);
xnor U17326 (N_17326,N_16664,N_16747);
nor U17327 (N_17327,N_16674,N_16517);
and U17328 (N_17328,N_16609,N_16616);
nand U17329 (N_17329,N_16595,N_16874);
nand U17330 (N_17330,N_16719,N_16600);
xor U17331 (N_17331,N_16730,N_16961);
or U17332 (N_17332,N_16800,N_16877);
xnor U17333 (N_17333,N_16759,N_16519);
xor U17334 (N_17334,N_16775,N_16818);
nand U17335 (N_17335,N_16728,N_16866);
xnor U17336 (N_17336,N_16876,N_16775);
nand U17337 (N_17337,N_16780,N_16500);
nand U17338 (N_17338,N_16831,N_16556);
xor U17339 (N_17339,N_16502,N_16733);
nand U17340 (N_17340,N_16719,N_16696);
and U17341 (N_17341,N_16941,N_16526);
or U17342 (N_17342,N_16751,N_16936);
or U17343 (N_17343,N_16806,N_16859);
xor U17344 (N_17344,N_16872,N_16816);
or U17345 (N_17345,N_16562,N_16649);
or U17346 (N_17346,N_16801,N_16605);
and U17347 (N_17347,N_16915,N_16701);
and U17348 (N_17348,N_16953,N_16642);
nor U17349 (N_17349,N_16671,N_16648);
or U17350 (N_17350,N_16823,N_16917);
xor U17351 (N_17351,N_16643,N_16833);
xor U17352 (N_17352,N_16938,N_16934);
nand U17353 (N_17353,N_16886,N_16851);
nor U17354 (N_17354,N_16707,N_16703);
xor U17355 (N_17355,N_16860,N_16685);
nand U17356 (N_17356,N_16621,N_16795);
and U17357 (N_17357,N_16569,N_16738);
or U17358 (N_17358,N_16549,N_16524);
xnor U17359 (N_17359,N_16607,N_16826);
nand U17360 (N_17360,N_16632,N_16926);
or U17361 (N_17361,N_16991,N_16544);
nor U17362 (N_17362,N_16953,N_16512);
xor U17363 (N_17363,N_16866,N_16948);
nor U17364 (N_17364,N_16867,N_16804);
nand U17365 (N_17365,N_16829,N_16564);
nor U17366 (N_17366,N_16577,N_16602);
nor U17367 (N_17367,N_16703,N_16885);
nand U17368 (N_17368,N_16571,N_16809);
and U17369 (N_17369,N_16588,N_16515);
or U17370 (N_17370,N_16965,N_16992);
or U17371 (N_17371,N_16686,N_16965);
nor U17372 (N_17372,N_16725,N_16703);
xor U17373 (N_17373,N_16952,N_16968);
and U17374 (N_17374,N_16571,N_16957);
xor U17375 (N_17375,N_16786,N_16510);
xor U17376 (N_17376,N_16975,N_16509);
nand U17377 (N_17377,N_16660,N_16690);
and U17378 (N_17378,N_16627,N_16922);
or U17379 (N_17379,N_16837,N_16834);
nor U17380 (N_17380,N_16605,N_16841);
and U17381 (N_17381,N_16713,N_16810);
nor U17382 (N_17382,N_16854,N_16871);
and U17383 (N_17383,N_16960,N_16616);
nand U17384 (N_17384,N_16543,N_16879);
or U17385 (N_17385,N_16664,N_16857);
and U17386 (N_17386,N_16515,N_16911);
nand U17387 (N_17387,N_16759,N_16695);
nand U17388 (N_17388,N_16653,N_16767);
nor U17389 (N_17389,N_16843,N_16796);
xor U17390 (N_17390,N_16905,N_16978);
and U17391 (N_17391,N_16822,N_16916);
or U17392 (N_17392,N_16571,N_16902);
nor U17393 (N_17393,N_16503,N_16908);
nand U17394 (N_17394,N_16661,N_16867);
nand U17395 (N_17395,N_16685,N_16581);
and U17396 (N_17396,N_16836,N_16710);
nand U17397 (N_17397,N_16551,N_16648);
or U17398 (N_17398,N_16625,N_16780);
nor U17399 (N_17399,N_16887,N_16576);
xor U17400 (N_17400,N_16510,N_16958);
nor U17401 (N_17401,N_16867,N_16645);
nor U17402 (N_17402,N_16947,N_16811);
and U17403 (N_17403,N_16590,N_16548);
or U17404 (N_17404,N_16665,N_16963);
nor U17405 (N_17405,N_16692,N_16805);
nor U17406 (N_17406,N_16988,N_16790);
or U17407 (N_17407,N_16580,N_16585);
nor U17408 (N_17408,N_16801,N_16916);
or U17409 (N_17409,N_16999,N_16784);
xnor U17410 (N_17410,N_16759,N_16644);
nand U17411 (N_17411,N_16896,N_16767);
or U17412 (N_17412,N_16762,N_16980);
nor U17413 (N_17413,N_16575,N_16788);
and U17414 (N_17414,N_16510,N_16691);
nand U17415 (N_17415,N_16777,N_16833);
or U17416 (N_17416,N_16540,N_16781);
nor U17417 (N_17417,N_16842,N_16710);
nand U17418 (N_17418,N_16622,N_16707);
nand U17419 (N_17419,N_16706,N_16526);
nor U17420 (N_17420,N_16983,N_16958);
nand U17421 (N_17421,N_16995,N_16629);
xnor U17422 (N_17422,N_16553,N_16556);
nor U17423 (N_17423,N_16705,N_16678);
xor U17424 (N_17424,N_16737,N_16558);
xnor U17425 (N_17425,N_16784,N_16862);
xnor U17426 (N_17426,N_16702,N_16999);
or U17427 (N_17427,N_16619,N_16772);
xor U17428 (N_17428,N_16533,N_16960);
xor U17429 (N_17429,N_16644,N_16760);
nor U17430 (N_17430,N_16590,N_16588);
nand U17431 (N_17431,N_16866,N_16670);
nand U17432 (N_17432,N_16505,N_16894);
or U17433 (N_17433,N_16855,N_16606);
nand U17434 (N_17434,N_16968,N_16698);
or U17435 (N_17435,N_16765,N_16662);
and U17436 (N_17436,N_16550,N_16735);
xor U17437 (N_17437,N_16890,N_16833);
and U17438 (N_17438,N_16568,N_16664);
nor U17439 (N_17439,N_16855,N_16545);
xor U17440 (N_17440,N_16999,N_16507);
or U17441 (N_17441,N_16792,N_16862);
and U17442 (N_17442,N_16744,N_16657);
xor U17443 (N_17443,N_16747,N_16661);
nor U17444 (N_17444,N_16722,N_16926);
xnor U17445 (N_17445,N_16881,N_16525);
and U17446 (N_17446,N_16973,N_16923);
nor U17447 (N_17447,N_16685,N_16925);
xor U17448 (N_17448,N_16933,N_16791);
nand U17449 (N_17449,N_16900,N_16690);
nand U17450 (N_17450,N_16641,N_16732);
nor U17451 (N_17451,N_16647,N_16802);
xor U17452 (N_17452,N_16903,N_16582);
nor U17453 (N_17453,N_16884,N_16637);
nand U17454 (N_17454,N_16605,N_16599);
nand U17455 (N_17455,N_16558,N_16972);
nand U17456 (N_17456,N_16650,N_16733);
xor U17457 (N_17457,N_16683,N_16915);
nor U17458 (N_17458,N_16976,N_16859);
and U17459 (N_17459,N_16764,N_16854);
or U17460 (N_17460,N_16895,N_16918);
nor U17461 (N_17461,N_16517,N_16558);
nand U17462 (N_17462,N_16726,N_16729);
and U17463 (N_17463,N_16774,N_16978);
nor U17464 (N_17464,N_16972,N_16550);
or U17465 (N_17465,N_16579,N_16926);
nand U17466 (N_17466,N_16987,N_16510);
and U17467 (N_17467,N_16914,N_16985);
nor U17468 (N_17468,N_16538,N_16971);
and U17469 (N_17469,N_16685,N_16732);
nand U17470 (N_17470,N_16653,N_16781);
xnor U17471 (N_17471,N_16704,N_16838);
xnor U17472 (N_17472,N_16507,N_16951);
or U17473 (N_17473,N_16676,N_16759);
nand U17474 (N_17474,N_16729,N_16620);
xnor U17475 (N_17475,N_16643,N_16983);
nor U17476 (N_17476,N_16883,N_16914);
xor U17477 (N_17477,N_16945,N_16734);
nand U17478 (N_17478,N_16695,N_16728);
nor U17479 (N_17479,N_16642,N_16688);
nand U17480 (N_17480,N_16980,N_16726);
and U17481 (N_17481,N_16816,N_16577);
or U17482 (N_17482,N_16923,N_16591);
xor U17483 (N_17483,N_16649,N_16876);
nor U17484 (N_17484,N_16548,N_16551);
xnor U17485 (N_17485,N_16761,N_16756);
and U17486 (N_17486,N_16654,N_16900);
xor U17487 (N_17487,N_16542,N_16794);
and U17488 (N_17488,N_16977,N_16561);
nor U17489 (N_17489,N_16923,N_16991);
and U17490 (N_17490,N_16926,N_16600);
nor U17491 (N_17491,N_16802,N_16905);
or U17492 (N_17492,N_16871,N_16773);
nor U17493 (N_17493,N_16591,N_16834);
nor U17494 (N_17494,N_16511,N_16767);
and U17495 (N_17495,N_16603,N_16655);
and U17496 (N_17496,N_16980,N_16731);
xnor U17497 (N_17497,N_16657,N_16535);
nand U17498 (N_17498,N_16843,N_16699);
xnor U17499 (N_17499,N_16777,N_16647);
or U17500 (N_17500,N_17135,N_17233);
xor U17501 (N_17501,N_17075,N_17450);
nand U17502 (N_17502,N_17032,N_17193);
nor U17503 (N_17503,N_17222,N_17069);
xnor U17504 (N_17504,N_17191,N_17317);
or U17505 (N_17505,N_17371,N_17001);
and U17506 (N_17506,N_17441,N_17307);
xnor U17507 (N_17507,N_17171,N_17038);
and U17508 (N_17508,N_17043,N_17202);
nor U17509 (N_17509,N_17091,N_17260);
or U17510 (N_17510,N_17452,N_17010);
xnor U17511 (N_17511,N_17068,N_17026);
and U17512 (N_17512,N_17420,N_17086);
nand U17513 (N_17513,N_17146,N_17312);
and U17514 (N_17514,N_17466,N_17006);
or U17515 (N_17515,N_17361,N_17300);
xor U17516 (N_17516,N_17322,N_17347);
xor U17517 (N_17517,N_17412,N_17031);
or U17518 (N_17518,N_17495,N_17132);
nand U17519 (N_17519,N_17157,N_17351);
nand U17520 (N_17520,N_17207,N_17363);
nor U17521 (N_17521,N_17235,N_17267);
or U17522 (N_17522,N_17030,N_17172);
nor U17523 (N_17523,N_17044,N_17040);
xor U17524 (N_17524,N_17138,N_17360);
nor U17525 (N_17525,N_17074,N_17173);
nand U17526 (N_17526,N_17185,N_17309);
nand U17527 (N_17527,N_17170,N_17252);
nand U17528 (N_17528,N_17458,N_17011);
nand U17529 (N_17529,N_17117,N_17061);
xnor U17530 (N_17530,N_17045,N_17463);
and U17531 (N_17531,N_17291,N_17262);
xnor U17532 (N_17532,N_17413,N_17257);
nand U17533 (N_17533,N_17015,N_17096);
nor U17534 (N_17534,N_17399,N_17389);
and U17535 (N_17535,N_17147,N_17244);
or U17536 (N_17536,N_17439,N_17438);
nand U17537 (N_17537,N_17085,N_17034);
nor U17538 (N_17538,N_17018,N_17167);
and U17539 (N_17539,N_17239,N_17002);
and U17540 (N_17540,N_17268,N_17430);
xor U17541 (N_17541,N_17014,N_17070);
xnor U17542 (N_17542,N_17111,N_17421);
and U17543 (N_17543,N_17273,N_17393);
or U17544 (N_17544,N_17052,N_17459);
nor U17545 (N_17545,N_17050,N_17008);
or U17546 (N_17546,N_17081,N_17119);
nand U17547 (N_17547,N_17094,N_17051);
nor U17548 (N_17548,N_17246,N_17118);
nand U17549 (N_17549,N_17021,N_17457);
nand U17550 (N_17550,N_17107,N_17293);
nand U17551 (N_17551,N_17376,N_17342);
nor U17552 (N_17552,N_17472,N_17180);
xnor U17553 (N_17553,N_17100,N_17469);
and U17554 (N_17554,N_17326,N_17440);
nor U17555 (N_17555,N_17210,N_17255);
xnor U17556 (N_17556,N_17057,N_17302);
xor U17557 (N_17557,N_17323,N_17264);
xnor U17558 (N_17558,N_17324,N_17343);
and U17559 (N_17559,N_17033,N_17159);
or U17560 (N_17560,N_17238,N_17189);
and U17561 (N_17561,N_17158,N_17102);
nor U17562 (N_17562,N_17053,N_17071);
or U17563 (N_17563,N_17039,N_17179);
nand U17564 (N_17564,N_17137,N_17063);
and U17565 (N_17565,N_17289,N_17296);
and U17566 (N_17566,N_17298,N_17041);
or U17567 (N_17567,N_17073,N_17403);
or U17568 (N_17568,N_17271,N_17320);
and U17569 (N_17569,N_17223,N_17446);
xor U17570 (N_17570,N_17279,N_17388);
nand U17571 (N_17571,N_17082,N_17286);
or U17572 (N_17572,N_17473,N_17407);
nor U17573 (N_17573,N_17048,N_17319);
or U17574 (N_17574,N_17359,N_17381);
nand U17575 (N_17575,N_17192,N_17400);
nand U17576 (N_17576,N_17449,N_17288);
nor U17577 (N_17577,N_17250,N_17416);
or U17578 (N_17578,N_17247,N_17303);
nand U17579 (N_17579,N_17292,N_17136);
and U17580 (N_17580,N_17467,N_17164);
nor U17581 (N_17581,N_17425,N_17422);
nor U17582 (N_17582,N_17224,N_17313);
xnor U17583 (N_17583,N_17127,N_17434);
and U17584 (N_17584,N_17465,N_17261);
nor U17585 (N_17585,N_17116,N_17499);
and U17586 (N_17586,N_17204,N_17398);
nor U17587 (N_17587,N_17301,N_17232);
or U17588 (N_17588,N_17408,N_17148);
or U17589 (N_17589,N_17195,N_17060);
xnor U17590 (N_17590,N_17089,N_17215);
or U17591 (N_17591,N_17236,N_17329);
xnor U17592 (N_17592,N_17353,N_17378);
or U17593 (N_17593,N_17188,N_17419);
nor U17594 (N_17594,N_17212,N_17256);
and U17595 (N_17595,N_17428,N_17203);
xnor U17596 (N_17596,N_17155,N_17476);
and U17597 (N_17597,N_17377,N_17427);
xnor U17598 (N_17598,N_17345,N_17078);
nand U17599 (N_17599,N_17237,N_17042);
nand U17600 (N_17600,N_17186,N_17474);
nor U17601 (N_17601,N_17219,N_17477);
or U17602 (N_17602,N_17093,N_17498);
xnor U17603 (N_17603,N_17409,N_17218);
xor U17604 (N_17604,N_17201,N_17475);
and U17605 (N_17605,N_17415,N_17028);
xnor U17606 (N_17606,N_17274,N_17337);
nor U17607 (N_17607,N_17493,N_17490);
nand U17608 (N_17608,N_17013,N_17206);
nand U17609 (N_17609,N_17375,N_17278);
nand U17610 (N_17610,N_17331,N_17327);
nand U17611 (N_17611,N_17036,N_17373);
nor U17612 (N_17612,N_17007,N_17484);
xnor U17613 (N_17613,N_17338,N_17437);
and U17614 (N_17614,N_17027,N_17384);
nand U17615 (N_17615,N_17395,N_17494);
nor U17616 (N_17616,N_17083,N_17456);
nor U17617 (N_17617,N_17272,N_17295);
xor U17618 (N_17618,N_17374,N_17339);
xor U17619 (N_17619,N_17284,N_17299);
nor U17620 (N_17620,N_17460,N_17294);
nor U17621 (N_17621,N_17162,N_17253);
nand U17622 (N_17622,N_17165,N_17401);
or U17623 (N_17623,N_17280,N_17304);
and U17624 (N_17624,N_17357,N_17243);
xnor U17625 (N_17625,N_17056,N_17417);
xor U17626 (N_17626,N_17000,N_17480);
or U17627 (N_17627,N_17208,N_17121);
nor U17628 (N_17628,N_17453,N_17491);
nand U17629 (N_17629,N_17194,N_17470);
nor U17630 (N_17630,N_17362,N_17391);
xor U17631 (N_17631,N_17321,N_17168);
nor U17632 (N_17632,N_17198,N_17305);
xor U17633 (N_17633,N_17332,N_17226);
and U17634 (N_17634,N_17064,N_17025);
or U17635 (N_17635,N_17405,N_17190);
and U17636 (N_17636,N_17108,N_17023);
nand U17637 (N_17637,N_17140,N_17481);
or U17638 (N_17638,N_17390,N_17153);
nand U17639 (N_17639,N_17095,N_17080);
nor U17640 (N_17640,N_17176,N_17315);
nand U17641 (N_17641,N_17468,N_17330);
and U17642 (N_17642,N_17358,N_17414);
nor U17643 (N_17643,N_17240,N_17266);
nor U17644 (N_17644,N_17325,N_17258);
xnor U17645 (N_17645,N_17003,N_17187);
xor U17646 (N_17646,N_17058,N_17386);
and U17647 (N_17647,N_17249,N_17139);
xnor U17648 (N_17648,N_17103,N_17149);
and U17649 (N_17649,N_17120,N_17334);
or U17650 (N_17650,N_17145,N_17211);
nor U17651 (N_17651,N_17005,N_17088);
xnor U17652 (N_17652,N_17055,N_17230);
or U17653 (N_17653,N_17114,N_17163);
nor U17654 (N_17654,N_17483,N_17352);
or U17655 (N_17655,N_17369,N_17380);
nand U17656 (N_17656,N_17287,N_17461);
xor U17657 (N_17657,N_17115,N_17076);
and U17658 (N_17658,N_17444,N_17426);
and U17659 (N_17659,N_17471,N_17451);
and U17660 (N_17660,N_17183,N_17382);
or U17661 (N_17661,N_17442,N_17123);
or U17662 (N_17662,N_17150,N_17418);
or U17663 (N_17663,N_17336,N_17281);
nand U17664 (N_17664,N_17049,N_17454);
xor U17665 (N_17665,N_17314,N_17318);
nand U17666 (N_17666,N_17367,N_17310);
nor U17667 (N_17667,N_17035,N_17077);
nand U17668 (N_17668,N_17356,N_17277);
nand U17669 (N_17669,N_17184,N_17365);
or U17670 (N_17670,N_17346,N_17199);
and U17671 (N_17671,N_17406,N_17251);
or U17672 (N_17672,N_17479,N_17349);
and U17673 (N_17673,N_17112,N_17282);
and U17674 (N_17674,N_17104,N_17269);
xnor U17675 (N_17675,N_17228,N_17105);
and U17676 (N_17676,N_17205,N_17079);
xnor U17677 (N_17677,N_17241,N_17344);
or U17678 (N_17678,N_17128,N_17254);
xnor U17679 (N_17679,N_17029,N_17098);
nor U17680 (N_17680,N_17177,N_17259);
nand U17681 (N_17681,N_17020,N_17364);
and U17682 (N_17682,N_17169,N_17379);
xnor U17683 (N_17683,N_17265,N_17174);
nor U17684 (N_17684,N_17178,N_17248);
nor U17685 (N_17685,N_17004,N_17024);
and U17686 (N_17686,N_17209,N_17221);
nor U17687 (N_17687,N_17429,N_17047);
nor U17688 (N_17688,N_17097,N_17276);
or U17689 (N_17689,N_17012,N_17046);
xor U17690 (N_17690,N_17113,N_17016);
or U17691 (N_17691,N_17066,N_17059);
and U17692 (N_17692,N_17090,N_17348);
nor U17693 (N_17693,N_17435,N_17072);
or U17694 (N_17694,N_17160,N_17242);
and U17695 (N_17695,N_17355,N_17485);
or U17696 (N_17696,N_17270,N_17133);
and U17697 (N_17697,N_17106,N_17433);
or U17698 (N_17698,N_17328,N_17445);
xnor U17699 (N_17699,N_17350,N_17341);
nor U17700 (N_17700,N_17436,N_17297);
or U17701 (N_17701,N_17492,N_17464);
xor U17702 (N_17702,N_17496,N_17488);
nand U17703 (N_17703,N_17216,N_17110);
or U17704 (N_17704,N_17037,N_17129);
or U17705 (N_17705,N_17290,N_17275);
or U17706 (N_17706,N_17154,N_17234);
and U17707 (N_17707,N_17394,N_17144);
xnor U17708 (N_17708,N_17431,N_17245);
or U17709 (N_17709,N_17125,N_17443);
and U17710 (N_17710,N_17387,N_17231);
and U17711 (N_17711,N_17368,N_17308);
nor U17712 (N_17712,N_17447,N_17383);
nor U17713 (N_17713,N_17099,N_17152);
xnor U17714 (N_17714,N_17166,N_17196);
xor U17715 (N_17715,N_17062,N_17065);
or U17716 (N_17716,N_17109,N_17067);
and U17717 (N_17717,N_17311,N_17462);
or U17718 (N_17718,N_17432,N_17370);
nor U17719 (N_17719,N_17283,N_17130);
and U17720 (N_17720,N_17423,N_17092);
nand U17721 (N_17721,N_17126,N_17486);
or U17722 (N_17722,N_17333,N_17217);
and U17723 (N_17723,N_17009,N_17410);
xor U17724 (N_17724,N_17087,N_17017);
nor U17725 (N_17725,N_17131,N_17151);
nor U17726 (N_17726,N_17455,N_17022);
or U17727 (N_17727,N_17392,N_17487);
xor U17728 (N_17728,N_17225,N_17124);
nand U17729 (N_17729,N_17213,N_17424);
and U17730 (N_17730,N_17220,N_17084);
xor U17731 (N_17731,N_17134,N_17316);
nor U17732 (N_17732,N_17229,N_17497);
nand U17733 (N_17733,N_17200,N_17402);
xor U17734 (N_17734,N_17197,N_17122);
xor U17735 (N_17735,N_17448,N_17482);
nand U17736 (N_17736,N_17181,N_17404);
nor U17737 (N_17737,N_17227,N_17411);
xor U17738 (N_17738,N_17143,N_17054);
nor U17739 (N_17739,N_17019,N_17478);
nor U17740 (N_17740,N_17285,N_17372);
xnor U17741 (N_17741,N_17306,N_17156);
xnor U17742 (N_17742,N_17263,N_17340);
xor U17743 (N_17743,N_17175,N_17141);
xor U17744 (N_17744,N_17489,N_17397);
nand U17745 (N_17745,N_17385,N_17354);
nor U17746 (N_17746,N_17366,N_17335);
or U17747 (N_17747,N_17142,N_17101);
nand U17748 (N_17748,N_17214,N_17396);
xnor U17749 (N_17749,N_17161,N_17182);
nand U17750 (N_17750,N_17413,N_17018);
nor U17751 (N_17751,N_17493,N_17058);
nand U17752 (N_17752,N_17214,N_17170);
xnor U17753 (N_17753,N_17095,N_17034);
nor U17754 (N_17754,N_17297,N_17131);
and U17755 (N_17755,N_17185,N_17110);
and U17756 (N_17756,N_17238,N_17311);
nor U17757 (N_17757,N_17210,N_17406);
xor U17758 (N_17758,N_17304,N_17217);
or U17759 (N_17759,N_17207,N_17275);
or U17760 (N_17760,N_17095,N_17146);
nand U17761 (N_17761,N_17476,N_17138);
xnor U17762 (N_17762,N_17421,N_17021);
nand U17763 (N_17763,N_17252,N_17197);
xor U17764 (N_17764,N_17353,N_17447);
xor U17765 (N_17765,N_17013,N_17409);
nand U17766 (N_17766,N_17173,N_17295);
xor U17767 (N_17767,N_17198,N_17269);
xnor U17768 (N_17768,N_17180,N_17413);
nor U17769 (N_17769,N_17277,N_17029);
xor U17770 (N_17770,N_17076,N_17066);
and U17771 (N_17771,N_17015,N_17410);
xor U17772 (N_17772,N_17332,N_17449);
or U17773 (N_17773,N_17042,N_17232);
nor U17774 (N_17774,N_17023,N_17124);
and U17775 (N_17775,N_17156,N_17147);
and U17776 (N_17776,N_17213,N_17294);
and U17777 (N_17777,N_17395,N_17116);
nand U17778 (N_17778,N_17471,N_17115);
nor U17779 (N_17779,N_17288,N_17322);
nor U17780 (N_17780,N_17329,N_17116);
xnor U17781 (N_17781,N_17471,N_17333);
and U17782 (N_17782,N_17429,N_17360);
xor U17783 (N_17783,N_17117,N_17450);
nand U17784 (N_17784,N_17289,N_17000);
xnor U17785 (N_17785,N_17451,N_17413);
nor U17786 (N_17786,N_17488,N_17135);
and U17787 (N_17787,N_17115,N_17024);
nor U17788 (N_17788,N_17304,N_17404);
xor U17789 (N_17789,N_17123,N_17203);
and U17790 (N_17790,N_17464,N_17495);
and U17791 (N_17791,N_17466,N_17245);
nor U17792 (N_17792,N_17249,N_17077);
or U17793 (N_17793,N_17400,N_17279);
nor U17794 (N_17794,N_17100,N_17212);
and U17795 (N_17795,N_17495,N_17383);
xnor U17796 (N_17796,N_17498,N_17082);
nand U17797 (N_17797,N_17372,N_17172);
or U17798 (N_17798,N_17367,N_17268);
nand U17799 (N_17799,N_17012,N_17351);
nor U17800 (N_17800,N_17019,N_17223);
or U17801 (N_17801,N_17094,N_17430);
xnor U17802 (N_17802,N_17252,N_17171);
nand U17803 (N_17803,N_17137,N_17132);
and U17804 (N_17804,N_17455,N_17484);
nand U17805 (N_17805,N_17331,N_17407);
xnor U17806 (N_17806,N_17203,N_17219);
nand U17807 (N_17807,N_17380,N_17010);
or U17808 (N_17808,N_17275,N_17395);
and U17809 (N_17809,N_17104,N_17370);
or U17810 (N_17810,N_17074,N_17419);
or U17811 (N_17811,N_17462,N_17176);
nand U17812 (N_17812,N_17109,N_17456);
xor U17813 (N_17813,N_17122,N_17258);
xnor U17814 (N_17814,N_17049,N_17326);
and U17815 (N_17815,N_17425,N_17358);
nand U17816 (N_17816,N_17187,N_17328);
xor U17817 (N_17817,N_17237,N_17324);
nand U17818 (N_17818,N_17004,N_17180);
xnor U17819 (N_17819,N_17429,N_17463);
xnor U17820 (N_17820,N_17499,N_17095);
nor U17821 (N_17821,N_17451,N_17456);
nor U17822 (N_17822,N_17364,N_17101);
xnor U17823 (N_17823,N_17340,N_17296);
or U17824 (N_17824,N_17419,N_17494);
xnor U17825 (N_17825,N_17234,N_17342);
nor U17826 (N_17826,N_17405,N_17385);
xor U17827 (N_17827,N_17151,N_17362);
or U17828 (N_17828,N_17328,N_17078);
nor U17829 (N_17829,N_17098,N_17060);
xor U17830 (N_17830,N_17341,N_17436);
and U17831 (N_17831,N_17404,N_17484);
and U17832 (N_17832,N_17218,N_17302);
or U17833 (N_17833,N_17337,N_17449);
nor U17834 (N_17834,N_17415,N_17494);
nor U17835 (N_17835,N_17242,N_17195);
nor U17836 (N_17836,N_17222,N_17313);
or U17837 (N_17837,N_17183,N_17466);
nor U17838 (N_17838,N_17130,N_17338);
nand U17839 (N_17839,N_17463,N_17069);
nand U17840 (N_17840,N_17058,N_17293);
or U17841 (N_17841,N_17051,N_17134);
nand U17842 (N_17842,N_17274,N_17363);
and U17843 (N_17843,N_17054,N_17466);
and U17844 (N_17844,N_17346,N_17021);
nor U17845 (N_17845,N_17017,N_17493);
and U17846 (N_17846,N_17143,N_17262);
xor U17847 (N_17847,N_17296,N_17294);
nor U17848 (N_17848,N_17422,N_17351);
nand U17849 (N_17849,N_17050,N_17369);
or U17850 (N_17850,N_17381,N_17046);
nor U17851 (N_17851,N_17142,N_17090);
or U17852 (N_17852,N_17070,N_17382);
or U17853 (N_17853,N_17381,N_17456);
or U17854 (N_17854,N_17169,N_17088);
xnor U17855 (N_17855,N_17234,N_17395);
nor U17856 (N_17856,N_17206,N_17175);
nor U17857 (N_17857,N_17310,N_17104);
nor U17858 (N_17858,N_17158,N_17209);
nand U17859 (N_17859,N_17020,N_17055);
and U17860 (N_17860,N_17261,N_17478);
and U17861 (N_17861,N_17150,N_17435);
xnor U17862 (N_17862,N_17189,N_17453);
and U17863 (N_17863,N_17267,N_17170);
or U17864 (N_17864,N_17434,N_17456);
nand U17865 (N_17865,N_17486,N_17482);
nand U17866 (N_17866,N_17268,N_17364);
and U17867 (N_17867,N_17229,N_17068);
nand U17868 (N_17868,N_17437,N_17282);
or U17869 (N_17869,N_17384,N_17464);
or U17870 (N_17870,N_17076,N_17042);
nor U17871 (N_17871,N_17337,N_17261);
xnor U17872 (N_17872,N_17409,N_17321);
nor U17873 (N_17873,N_17216,N_17090);
xor U17874 (N_17874,N_17368,N_17276);
nor U17875 (N_17875,N_17305,N_17307);
xnor U17876 (N_17876,N_17366,N_17395);
nor U17877 (N_17877,N_17015,N_17052);
nor U17878 (N_17878,N_17160,N_17101);
xnor U17879 (N_17879,N_17153,N_17197);
nor U17880 (N_17880,N_17405,N_17439);
nand U17881 (N_17881,N_17300,N_17043);
or U17882 (N_17882,N_17273,N_17091);
xor U17883 (N_17883,N_17199,N_17393);
nand U17884 (N_17884,N_17131,N_17451);
nand U17885 (N_17885,N_17225,N_17236);
nor U17886 (N_17886,N_17364,N_17357);
nand U17887 (N_17887,N_17062,N_17229);
nor U17888 (N_17888,N_17320,N_17098);
and U17889 (N_17889,N_17266,N_17047);
and U17890 (N_17890,N_17231,N_17021);
and U17891 (N_17891,N_17075,N_17000);
xnor U17892 (N_17892,N_17489,N_17325);
and U17893 (N_17893,N_17253,N_17470);
or U17894 (N_17894,N_17016,N_17442);
or U17895 (N_17895,N_17487,N_17424);
or U17896 (N_17896,N_17068,N_17366);
nand U17897 (N_17897,N_17369,N_17467);
nor U17898 (N_17898,N_17206,N_17464);
nand U17899 (N_17899,N_17421,N_17494);
xnor U17900 (N_17900,N_17326,N_17313);
xor U17901 (N_17901,N_17250,N_17307);
xnor U17902 (N_17902,N_17338,N_17085);
or U17903 (N_17903,N_17085,N_17493);
nand U17904 (N_17904,N_17113,N_17317);
and U17905 (N_17905,N_17029,N_17436);
nand U17906 (N_17906,N_17412,N_17494);
and U17907 (N_17907,N_17274,N_17373);
and U17908 (N_17908,N_17166,N_17459);
or U17909 (N_17909,N_17070,N_17388);
and U17910 (N_17910,N_17492,N_17252);
or U17911 (N_17911,N_17295,N_17347);
nor U17912 (N_17912,N_17448,N_17307);
and U17913 (N_17913,N_17297,N_17279);
nand U17914 (N_17914,N_17274,N_17468);
and U17915 (N_17915,N_17023,N_17487);
xnor U17916 (N_17916,N_17191,N_17283);
or U17917 (N_17917,N_17203,N_17448);
nand U17918 (N_17918,N_17254,N_17100);
xor U17919 (N_17919,N_17111,N_17171);
or U17920 (N_17920,N_17170,N_17120);
or U17921 (N_17921,N_17245,N_17240);
and U17922 (N_17922,N_17050,N_17142);
and U17923 (N_17923,N_17233,N_17250);
and U17924 (N_17924,N_17236,N_17193);
and U17925 (N_17925,N_17131,N_17216);
or U17926 (N_17926,N_17221,N_17359);
nor U17927 (N_17927,N_17239,N_17422);
and U17928 (N_17928,N_17317,N_17090);
and U17929 (N_17929,N_17476,N_17177);
xor U17930 (N_17930,N_17175,N_17188);
nor U17931 (N_17931,N_17257,N_17207);
nand U17932 (N_17932,N_17168,N_17326);
nor U17933 (N_17933,N_17437,N_17216);
nor U17934 (N_17934,N_17016,N_17282);
or U17935 (N_17935,N_17096,N_17499);
and U17936 (N_17936,N_17163,N_17023);
and U17937 (N_17937,N_17208,N_17151);
nor U17938 (N_17938,N_17388,N_17396);
nor U17939 (N_17939,N_17390,N_17498);
and U17940 (N_17940,N_17419,N_17395);
xnor U17941 (N_17941,N_17177,N_17214);
nand U17942 (N_17942,N_17433,N_17429);
nor U17943 (N_17943,N_17051,N_17036);
or U17944 (N_17944,N_17400,N_17322);
and U17945 (N_17945,N_17203,N_17253);
and U17946 (N_17946,N_17226,N_17285);
nand U17947 (N_17947,N_17272,N_17008);
xor U17948 (N_17948,N_17085,N_17351);
xnor U17949 (N_17949,N_17454,N_17446);
nand U17950 (N_17950,N_17113,N_17290);
nand U17951 (N_17951,N_17146,N_17426);
or U17952 (N_17952,N_17114,N_17018);
xnor U17953 (N_17953,N_17090,N_17281);
xor U17954 (N_17954,N_17204,N_17491);
nor U17955 (N_17955,N_17046,N_17040);
nor U17956 (N_17956,N_17367,N_17012);
or U17957 (N_17957,N_17304,N_17187);
or U17958 (N_17958,N_17243,N_17297);
or U17959 (N_17959,N_17126,N_17134);
xnor U17960 (N_17960,N_17464,N_17397);
nand U17961 (N_17961,N_17492,N_17401);
xnor U17962 (N_17962,N_17179,N_17439);
nor U17963 (N_17963,N_17276,N_17443);
nor U17964 (N_17964,N_17210,N_17101);
nor U17965 (N_17965,N_17062,N_17464);
nand U17966 (N_17966,N_17386,N_17478);
nand U17967 (N_17967,N_17308,N_17494);
or U17968 (N_17968,N_17419,N_17370);
nor U17969 (N_17969,N_17266,N_17032);
and U17970 (N_17970,N_17020,N_17163);
xor U17971 (N_17971,N_17389,N_17137);
or U17972 (N_17972,N_17277,N_17137);
and U17973 (N_17973,N_17245,N_17486);
xnor U17974 (N_17974,N_17050,N_17386);
or U17975 (N_17975,N_17499,N_17377);
nor U17976 (N_17976,N_17362,N_17174);
nand U17977 (N_17977,N_17453,N_17035);
xor U17978 (N_17978,N_17238,N_17452);
or U17979 (N_17979,N_17054,N_17058);
or U17980 (N_17980,N_17215,N_17430);
and U17981 (N_17981,N_17416,N_17081);
nor U17982 (N_17982,N_17107,N_17019);
xnor U17983 (N_17983,N_17233,N_17083);
and U17984 (N_17984,N_17469,N_17190);
nor U17985 (N_17985,N_17249,N_17006);
or U17986 (N_17986,N_17198,N_17439);
and U17987 (N_17987,N_17279,N_17103);
or U17988 (N_17988,N_17162,N_17343);
and U17989 (N_17989,N_17135,N_17484);
nand U17990 (N_17990,N_17192,N_17398);
nor U17991 (N_17991,N_17051,N_17207);
and U17992 (N_17992,N_17461,N_17312);
nand U17993 (N_17993,N_17340,N_17473);
nor U17994 (N_17994,N_17158,N_17350);
xor U17995 (N_17995,N_17299,N_17438);
and U17996 (N_17996,N_17256,N_17396);
or U17997 (N_17997,N_17017,N_17281);
nand U17998 (N_17998,N_17336,N_17092);
or U17999 (N_17999,N_17112,N_17433);
and U18000 (N_18000,N_17716,N_17919);
nor U18001 (N_18001,N_17545,N_17900);
nor U18002 (N_18002,N_17557,N_17760);
or U18003 (N_18003,N_17834,N_17932);
xnor U18004 (N_18004,N_17500,N_17647);
and U18005 (N_18005,N_17561,N_17794);
nand U18006 (N_18006,N_17526,N_17844);
nand U18007 (N_18007,N_17995,N_17720);
xnor U18008 (N_18008,N_17642,N_17683);
xor U18009 (N_18009,N_17841,N_17584);
or U18010 (N_18010,N_17539,N_17676);
and U18011 (N_18011,N_17871,N_17908);
or U18012 (N_18012,N_17651,N_17795);
nand U18013 (N_18013,N_17961,N_17641);
nor U18014 (N_18014,N_17743,N_17784);
nand U18015 (N_18015,N_17680,N_17935);
or U18016 (N_18016,N_17772,N_17733);
or U18017 (N_18017,N_17863,N_17707);
nor U18018 (N_18018,N_17629,N_17549);
or U18019 (N_18019,N_17677,N_17832);
xnor U18020 (N_18020,N_17839,N_17816);
xnor U18021 (N_18021,N_17893,N_17659);
nand U18022 (N_18022,N_17594,N_17997);
and U18023 (N_18023,N_17735,N_17656);
or U18024 (N_18024,N_17525,N_17737);
or U18025 (N_18025,N_17521,N_17886);
or U18026 (N_18026,N_17681,N_17567);
xor U18027 (N_18027,N_17591,N_17955);
nand U18028 (N_18028,N_17652,N_17954);
nor U18029 (N_18029,N_17933,N_17714);
xor U18030 (N_18030,N_17805,N_17732);
nor U18031 (N_18031,N_17501,N_17729);
and U18032 (N_18032,N_17630,N_17906);
nand U18033 (N_18033,N_17688,N_17994);
xor U18034 (N_18034,N_17595,N_17851);
nand U18035 (N_18035,N_17813,N_17943);
nand U18036 (N_18036,N_17510,N_17940);
xor U18037 (N_18037,N_17699,N_17705);
and U18038 (N_18038,N_17614,N_17740);
or U18039 (N_18039,N_17667,N_17782);
and U18040 (N_18040,N_17827,N_17708);
xor U18041 (N_18041,N_17867,N_17610);
or U18042 (N_18042,N_17559,N_17694);
or U18043 (N_18043,N_17796,N_17921);
nand U18044 (N_18044,N_17996,N_17789);
nand U18045 (N_18045,N_17853,N_17605);
nor U18046 (N_18046,N_17530,N_17578);
and U18047 (N_18047,N_17535,N_17777);
or U18048 (N_18048,N_17976,N_17689);
xor U18049 (N_18049,N_17527,N_17768);
nor U18050 (N_18050,N_17883,N_17751);
nor U18051 (N_18051,N_17670,N_17956);
nor U18052 (N_18052,N_17581,N_17508);
and U18053 (N_18053,N_17988,N_17985);
xnor U18054 (N_18054,N_17929,N_17661);
nor U18055 (N_18055,N_17907,N_17672);
nor U18056 (N_18056,N_17738,N_17809);
or U18057 (N_18057,N_17514,N_17815);
and U18058 (N_18058,N_17939,N_17653);
and U18059 (N_18059,N_17566,N_17627);
xor U18060 (N_18060,N_17766,N_17990);
nand U18061 (N_18061,N_17711,N_17519);
and U18062 (N_18062,N_17606,N_17828);
and U18063 (N_18063,N_17818,N_17978);
nand U18064 (N_18064,N_17646,N_17687);
nand U18065 (N_18065,N_17846,N_17590);
nor U18066 (N_18066,N_17531,N_17986);
or U18067 (N_18067,N_17973,N_17702);
nand U18068 (N_18068,N_17821,N_17660);
and U18069 (N_18069,N_17979,N_17645);
and U18070 (N_18070,N_17504,N_17838);
xnor U18071 (N_18071,N_17896,N_17833);
nand U18072 (N_18072,N_17502,N_17779);
xor U18073 (N_18073,N_17989,N_17593);
xor U18074 (N_18074,N_17690,N_17715);
nand U18075 (N_18075,N_17901,N_17542);
nor U18076 (N_18076,N_17761,N_17587);
nand U18077 (N_18077,N_17904,N_17505);
xor U18078 (N_18078,N_17764,N_17773);
or U18079 (N_18079,N_17727,N_17635);
or U18080 (N_18080,N_17543,N_17685);
and U18081 (N_18081,N_17836,N_17599);
or U18082 (N_18082,N_17897,N_17889);
nand U18083 (N_18083,N_17586,N_17754);
and U18084 (N_18084,N_17970,N_17802);
xnor U18085 (N_18085,N_17930,N_17856);
or U18086 (N_18086,N_17806,N_17657);
or U18087 (N_18087,N_17537,N_17516);
xnor U18088 (N_18088,N_17544,N_17880);
and U18089 (N_18089,N_17726,N_17905);
or U18090 (N_18090,N_17790,N_17756);
or U18091 (N_18091,N_17673,N_17810);
and U18092 (N_18092,N_17850,N_17881);
nand U18093 (N_18093,N_17574,N_17875);
and U18094 (N_18094,N_17892,N_17983);
nor U18095 (N_18095,N_17520,N_17580);
nand U18096 (N_18096,N_17511,N_17858);
and U18097 (N_18097,N_17588,N_17603);
xor U18098 (N_18098,N_17987,N_17826);
nand U18099 (N_18099,N_17678,N_17728);
or U18100 (N_18100,N_17895,N_17854);
nand U18101 (N_18101,N_17665,N_17925);
and U18102 (N_18102,N_17982,N_17874);
or U18103 (N_18103,N_17757,N_17697);
nand U18104 (N_18104,N_17840,N_17877);
and U18105 (N_18105,N_17931,N_17554);
or U18106 (N_18106,N_17734,N_17541);
xnor U18107 (N_18107,N_17755,N_17664);
or U18108 (N_18108,N_17583,N_17902);
xnor U18109 (N_18109,N_17991,N_17859);
nand U18110 (N_18110,N_17601,N_17555);
nand U18111 (N_18111,N_17631,N_17825);
nor U18112 (N_18112,N_17914,N_17577);
or U18113 (N_18113,N_17695,N_17948);
and U18114 (N_18114,N_17634,N_17941);
nand U18115 (N_18115,N_17831,N_17636);
or U18116 (N_18116,N_17524,N_17960);
and U18117 (N_18117,N_17920,N_17959);
and U18118 (N_18118,N_17602,N_17675);
or U18119 (N_18119,N_17934,N_17648);
nor U18120 (N_18120,N_17776,N_17649);
nor U18121 (N_18121,N_17517,N_17589);
xnor U18122 (N_18122,N_17951,N_17563);
xor U18123 (N_18123,N_17927,N_17797);
xnor U18124 (N_18124,N_17758,N_17829);
and U18125 (N_18125,N_17891,N_17512);
and U18126 (N_18126,N_17570,N_17503);
nor U18127 (N_18127,N_17977,N_17770);
and U18128 (N_18128,N_17894,N_17852);
and U18129 (N_18129,N_17903,N_17696);
xnor U18130 (N_18130,N_17736,N_17966);
and U18131 (N_18131,N_17866,N_17981);
or U18132 (N_18132,N_17556,N_17739);
or U18133 (N_18133,N_17864,N_17868);
xor U18134 (N_18134,N_17682,N_17597);
nand U18135 (N_18135,N_17767,N_17741);
xor U18136 (N_18136,N_17565,N_17620);
or U18137 (N_18137,N_17742,N_17807);
or U18138 (N_18138,N_17873,N_17536);
or U18139 (N_18139,N_17862,N_17624);
xnor U18140 (N_18140,N_17532,N_17638);
xnor U18141 (N_18141,N_17747,N_17618);
xor U18142 (N_18142,N_17709,N_17604);
nor U18143 (N_18143,N_17529,N_17533);
xor U18144 (N_18144,N_17662,N_17560);
xor U18145 (N_18145,N_17621,N_17655);
nor U18146 (N_18146,N_17969,N_17749);
and U18147 (N_18147,N_17980,N_17644);
and U18148 (N_18148,N_17824,N_17540);
and U18149 (N_18149,N_17633,N_17804);
and U18150 (N_18150,N_17684,N_17534);
xnor U18151 (N_18151,N_17548,N_17949);
nand U18152 (N_18152,N_17700,N_17942);
xor U18153 (N_18153,N_17759,N_17924);
nand U18154 (N_18154,N_17632,N_17912);
and U18155 (N_18155,N_17884,N_17855);
and U18156 (N_18156,N_17974,N_17928);
nand U18157 (N_18157,N_17745,N_17781);
or U18158 (N_18158,N_17706,N_17639);
and U18159 (N_18159,N_17569,N_17946);
nor U18160 (N_18160,N_17619,N_17817);
and U18161 (N_18161,N_17944,N_17686);
and U18162 (N_18162,N_17801,N_17936);
nor U18163 (N_18163,N_17722,N_17710);
or U18164 (N_18164,N_17808,N_17958);
xnor U18165 (N_18165,N_17669,N_17547);
xnor U18166 (N_18166,N_17962,N_17721);
and U18167 (N_18167,N_17528,N_17857);
nand U18168 (N_18168,N_17837,N_17507);
and U18169 (N_18169,N_17800,N_17622);
or U18170 (N_18170,N_17992,N_17788);
nor U18171 (N_18171,N_17953,N_17885);
and U18172 (N_18172,N_17693,N_17568);
and U18173 (N_18173,N_17765,N_17842);
nand U18174 (N_18174,N_17803,N_17812);
nor U18175 (N_18175,N_17799,N_17957);
or U18176 (N_18176,N_17872,N_17998);
and U18177 (N_18177,N_17650,N_17964);
or U18178 (N_18178,N_17876,N_17783);
nand U18179 (N_18179,N_17774,N_17820);
and U18180 (N_18180,N_17848,N_17637);
or U18181 (N_18181,N_17778,N_17769);
nand U18182 (N_18182,N_17792,N_17691);
nand U18183 (N_18183,N_17909,N_17922);
nor U18184 (N_18184,N_17882,N_17518);
xnor U18185 (N_18185,N_17615,N_17698);
xor U18186 (N_18186,N_17625,N_17692);
and U18187 (N_18187,N_17551,N_17550);
xnor U18188 (N_18188,N_17582,N_17911);
or U18189 (N_18189,N_17823,N_17609);
or U18190 (N_18190,N_17787,N_17849);
xnor U18191 (N_18191,N_17965,N_17835);
xor U18192 (N_18192,N_17916,N_17972);
and U18193 (N_18193,N_17878,N_17666);
nor U18194 (N_18194,N_17717,N_17592);
nand U18195 (N_18195,N_17918,N_17861);
xnor U18196 (N_18196,N_17975,N_17626);
nand U18197 (N_18197,N_17730,N_17719);
and U18198 (N_18198,N_17963,N_17811);
and U18199 (N_18199,N_17617,N_17763);
or U18200 (N_18200,N_17562,N_17843);
nor U18201 (N_18201,N_17658,N_17564);
nor U18202 (N_18202,N_17579,N_17993);
nand U18203 (N_18203,N_17845,N_17654);
xnor U18204 (N_18204,N_17913,N_17786);
and U18205 (N_18205,N_17546,N_17725);
and U18206 (N_18206,N_17600,N_17643);
nor U18207 (N_18207,N_17628,N_17744);
nand U18208 (N_18208,N_17679,N_17890);
and U18209 (N_18209,N_17713,N_17746);
xor U18210 (N_18210,N_17814,N_17952);
or U18211 (N_18211,N_17509,N_17750);
xnor U18212 (N_18212,N_17984,N_17910);
nor U18213 (N_18213,N_17847,N_17723);
xor U18214 (N_18214,N_17771,N_17576);
and U18215 (N_18215,N_17879,N_17611);
xor U18216 (N_18216,N_17785,N_17869);
nand U18217 (N_18217,N_17572,N_17608);
xnor U18218 (N_18218,N_17674,N_17596);
or U18219 (N_18219,N_17506,N_17967);
nand U18220 (N_18220,N_17513,N_17780);
and U18221 (N_18221,N_17748,N_17860);
and U18222 (N_18222,N_17950,N_17671);
and U18223 (N_18223,N_17623,N_17898);
nand U18224 (N_18224,N_17752,N_17515);
or U18225 (N_18225,N_17870,N_17753);
and U18226 (N_18226,N_17917,N_17703);
nor U18227 (N_18227,N_17724,N_17937);
and U18228 (N_18228,N_17668,N_17573);
and U18229 (N_18229,N_17915,N_17762);
xor U18230 (N_18230,N_17865,N_17968);
nand U18231 (N_18231,N_17616,N_17775);
xnor U18232 (N_18232,N_17971,N_17523);
nand U18233 (N_18233,N_17798,N_17791);
and U18234 (N_18234,N_17819,N_17887);
nand U18235 (N_18235,N_17712,N_17899);
and U18236 (N_18236,N_17613,N_17598);
xor U18237 (N_18237,N_17926,N_17522);
xor U18238 (N_18238,N_17663,N_17553);
and U18239 (N_18239,N_17552,N_17607);
and U18240 (N_18240,N_17945,N_17701);
or U18241 (N_18241,N_17612,N_17947);
and U18242 (N_18242,N_17704,N_17938);
nor U18243 (N_18243,N_17999,N_17793);
nor U18244 (N_18244,N_17640,N_17538);
nand U18245 (N_18245,N_17731,N_17575);
nor U18246 (N_18246,N_17923,N_17830);
nor U18247 (N_18247,N_17558,N_17571);
xnor U18248 (N_18248,N_17822,N_17718);
nor U18249 (N_18249,N_17585,N_17888);
nand U18250 (N_18250,N_17760,N_17512);
or U18251 (N_18251,N_17830,N_17888);
nor U18252 (N_18252,N_17713,N_17788);
or U18253 (N_18253,N_17810,N_17978);
or U18254 (N_18254,N_17711,N_17762);
and U18255 (N_18255,N_17545,N_17847);
and U18256 (N_18256,N_17771,N_17568);
and U18257 (N_18257,N_17756,N_17506);
nand U18258 (N_18258,N_17581,N_17831);
xor U18259 (N_18259,N_17503,N_17837);
nand U18260 (N_18260,N_17861,N_17986);
nor U18261 (N_18261,N_17878,N_17738);
and U18262 (N_18262,N_17995,N_17568);
nor U18263 (N_18263,N_17868,N_17991);
or U18264 (N_18264,N_17829,N_17822);
nand U18265 (N_18265,N_17971,N_17527);
nor U18266 (N_18266,N_17562,N_17641);
nand U18267 (N_18267,N_17875,N_17843);
nor U18268 (N_18268,N_17933,N_17659);
and U18269 (N_18269,N_17536,N_17800);
nor U18270 (N_18270,N_17522,N_17679);
nor U18271 (N_18271,N_17566,N_17660);
and U18272 (N_18272,N_17829,N_17685);
and U18273 (N_18273,N_17765,N_17668);
or U18274 (N_18274,N_17820,N_17671);
xor U18275 (N_18275,N_17743,N_17641);
nor U18276 (N_18276,N_17607,N_17617);
or U18277 (N_18277,N_17938,N_17906);
nand U18278 (N_18278,N_17965,N_17843);
and U18279 (N_18279,N_17840,N_17971);
nand U18280 (N_18280,N_17714,N_17904);
nand U18281 (N_18281,N_17875,N_17593);
xnor U18282 (N_18282,N_17905,N_17744);
or U18283 (N_18283,N_17728,N_17569);
nand U18284 (N_18284,N_17920,N_17744);
or U18285 (N_18285,N_17981,N_17790);
nand U18286 (N_18286,N_17549,N_17837);
and U18287 (N_18287,N_17524,N_17947);
or U18288 (N_18288,N_17823,N_17935);
xnor U18289 (N_18289,N_17629,N_17852);
or U18290 (N_18290,N_17645,N_17777);
and U18291 (N_18291,N_17776,N_17769);
and U18292 (N_18292,N_17758,N_17820);
and U18293 (N_18293,N_17664,N_17641);
and U18294 (N_18294,N_17948,N_17784);
or U18295 (N_18295,N_17946,N_17501);
xor U18296 (N_18296,N_17655,N_17770);
xnor U18297 (N_18297,N_17622,N_17560);
or U18298 (N_18298,N_17846,N_17994);
or U18299 (N_18299,N_17822,N_17863);
or U18300 (N_18300,N_17725,N_17649);
xor U18301 (N_18301,N_17781,N_17737);
or U18302 (N_18302,N_17532,N_17868);
and U18303 (N_18303,N_17792,N_17748);
and U18304 (N_18304,N_17683,N_17948);
xnor U18305 (N_18305,N_17938,N_17703);
xnor U18306 (N_18306,N_17950,N_17839);
and U18307 (N_18307,N_17908,N_17707);
nand U18308 (N_18308,N_17549,N_17600);
nand U18309 (N_18309,N_17757,N_17532);
nor U18310 (N_18310,N_17653,N_17740);
or U18311 (N_18311,N_17582,N_17607);
xor U18312 (N_18312,N_17646,N_17934);
nor U18313 (N_18313,N_17746,N_17901);
nand U18314 (N_18314,N_17814,N_17606);
or U18315 (N_18315,N_17705,N_17857);
nor U18316 (N_18316,N_17710,N_17899);
and U18317 (N_18317,N_17558,N_17927);
nor U18318 (N_18318,N_17926,N_17524);
or U18319 (N_18319,N_17853,N_17502);
or U18320 (N_18320,N_17719,N_17883);
or U18321 (N_18321,N_17548,N_17844);
nor U18322 (N_18322,N_17963,N_17952);
nor U18323 (N_18323,N_17799,N_17604);
nor U18324 (N_18324,N_17533,N_17931);
xnor U18325 (N_18325,N_17660,N_17548);
or U18326 (N_18326,N_17922,N_17520);
nor U18327 (N_18327,N_17805,N_17776);
xnor U18328 (N_18328,N_17906,N_17574);
or U18329 (N_18329,N_17796,N_17899);
xor U18330 (N_18330,N_17822,N_17577);
nor U18331 (N_18331,N_17951,N_17769);
nor U18332 (N_18332,N_17544,N_17509);
nand U18333 (N_18333,N_17517,N_17803);
xnor U18334 (N_18334,N_17525,N_17662);
nand U18335 (N_18335,N_17521,N_17792);
nor U18336 (N_18336,N_17675,N_17932);
or U18337 (N_18337,N_17699,N_17882);
nand U18338 (N_18338,N_17848,N_17834);
or U18339 (N_18339,N_17885,N_17513);
nand U18340 (N_18340,N_17594,N_17750);
or U18341 (N_18341,N_17735,N_17819);
nand U18342 (N_18342,N_17823,N_17840);
and U18343 (N_18343,N_17543,N_17887);
or U18344 (N_18344,N_17994,N_17925);
or U18345 (N_18345,N_17803,N_17811);
nor U18346 (N_18346,N_17589,N_17899);
and U18347 (N_18347,N_17899,N_17609);
xnor U18348 (N_18348,N_17963,N_17903);
nor U18349 (N_18349,N_17957,N_17866);
nor U18350 (N_18350,N_17657,N_17925);
nand U18351 (N_18351,N_17894,N_17569);
xor U18352 (N_18352,N_17887,N_17782);
xnor U18353 (N_18353,N_17702,N_17911);
and U18354 (N_18354,N_17528,N_17840);
nand U18355 (N_18355,N_17709,N_17722);
nor U18356 (N_18356,N_17770,N_17798);
xor U18357 (N_18357,N_17934,N_17820);
and U18358 (N_18358,N_17667,N_17718);
xnor U18359 (N_18359,N_17621,N_17617);
nand U18360 (N_18360,N_17613,N_17890);
nor U18361 (N_18361,N_17507,N_17722);
or U18362 (N_18362,N_17791,N_17920);
nand U18363 (N_18363,N_17810,N_17812);
or U18364 (N_18364,N_17863,N_17930);
and U18365 (N_18365,N_17526,N_17748);
nor U18366 (N_18366,N_17642,N_17959);
or U18367 (N_18367,N_17815,N_17641);
or U18368 (N_18368,N_17957,N_17541);
nand U18369 (N_18369,N_17510,N_17764);
and U18370 (N_18370,N_17821,N_17826);
and U18371 (N_18371,N_17906,N_17817);
or U18372 (N_18372,N_17623,N_17635);
and U18373 (N_18373,N_17753,N_17633);
xor U18374 (N_18374,N_17527,N_17545);
and U18375 (N_18375,N_17972,N_17631);
nor U18376 (N_18376,N_17967,N_17973);
nand U18377 (N_18377,N_17961,N_17694);
nand U18378 (N_18378,N_17882,N_17735);
nand U18379 (N_18379,N_17631,N_17838);
and U18380 (N_18380,N_17676,N_17975);
and U18381 (N_18381,N_17612,N_17974);
or U18382 (N_18382,N_17990,N_17747);
and U18383 (N_18383,N_17741,N_17967);
or U18384 (N_18384,N_17797,N_17794);
xor U18385 (N_18385,N_17851,N_17853);
or U18386 (N_18386,N_17612,N_17642);
nand U18387 (N_18387,N_17824,N_17935);
nor U18388 (N_18388,N_17715,N_17883);
and U18389 (N_18389,N_17660,N_17567);
xor U18390 (N_18390,N_17960,N_17935);
xnor U18391 (N_18391,N_17737,N_17897);
or U18392 (N_18392,N_17556,N_17934);
or U18393 (N_18393,N_17791,N_17995);
and U18394 (N_18394,N_17960,N_17878);
or U18395 (N_18395,N_17520,N_17578);
xor U18396 (N_18396,N_17611,N_17853);
or U18397 (N_18397,N_17854,N_17824);
and U18398 (N_18398,N_17675,N_17956);
or U18399 (N_18399,N_17985,N_17937);
xor U18400 (N_18400,N_17616,N_17523);
or U18401 (N_18401,N_17838,N_17648);
nand U18402 (N_18402,N_17985,N_17796);
and U18403 (N_18403,N_17640,N_17861);
and U18404 (N_18404,N_17965,N_17712);
nand U18405 (N_18405,N_17690,N_17536);
nand U18406 (N_18406,N_17662,N_17621);
and U18407 (N_18407,N_17639,N_17965);
or U18408 (N_18408,N_17913,N_17945);
xor U18409 (N_18409,N_17998,N_17849);
nor U18410 (N_18410,N_17538,N_17614);
and U18411 (N_18411,N_17668,N_17888);
nor U18412 (N_18412,N_17858,N_17979);
nor U18413 (N_18413,N_17566,N_17541);
or U18414 (N_18414,N_17748,N_17841);
and U18415 (N_18415,N_17740,N_17902);
xnor U18416 (N_18416,N_17835,N_17946);
and U18417 (N_18417,N_17842,N_17810);
xnor U18418 (N_18418,N_17748,N_17788);
nor U18419 (N_18419,N_17891,N_17727);
or U18420 (N_18420,N_17785,N_17965);
nor U18421 (N_18421,N_17962,N_17567);
or U18422 (N_18422,N_17907,N_17978);
or U18423 (N_18423,N_17667,N_17813);
xor U18424 (N_18424,N_17783,N_17909);
xnor U18425 (N_18425,N_17974,N_17601);
and U18426 (N_18426,N_17505,N_17553);
nand U18427 (N_18427,N_17933,N_17894);
nand U18428 (N_18428,N_17540,N_17935);
nand U18429 (N_18429,N_17948,N_17987);
xor U18430 (N_18430,N_17644,N_17529);
nor U18431 (N_18431,N_17721,N_17809);
nand U18432 (N_18432,N_17588,N_17685);
or U18433 (N_18433,N_17802,N_17554);
nand U18434 (N_18434,N_17929,N_17657);
and U18435 (N_18435,N_17910,N_17947);
nor U18436 (N_18436,N_17749,N_17610);
nor U18437 (N_18437,N_17911,N_17759);
and U18438 (N_18438,N_17856,N_17752);
and U18439 (N_18439,N_17503,N_17690);
xnor U18440 (N_18440,N_17832,N_17874);
or U18441 (N_18441,N_17504,N_17584);
nand U18442 (N_18442,N_17774,N_17957);
or U18443 (N_18443,N_17971,N_17917);
or U18444 (N_18444,N_17746,N_17814);
xor U18445 (N_18445,N_17547,N_17693);
xor U18446 (N_18446,N_17501,N_17704);
or U18447 (N_18447,N_17701,N_17517);
and U18448 (N_18448,N_17533,N_17943);
nand U18449 (N_18449,N_17919,N_17542);
or U18450 (N_18450,N_17751,N_17757);
nor U18451 (N_18451,N_17680,N_17712);
and U18452 (N_18452,N_17980,N_17828);
or U18453 (N_18453,N_17780,N_17824);
xor U18454 (N_18454,N_17927,N_17501);
or U18455 (N_18455,N_17600,N_17938);
or U18456 (N_18456,N_17850,N_17972);
xnor U18457 (N_18457,N_17838,N_17914);
nand U18458 (N_18458,N_17750,N_17913);
and U18459 (N_18459,N_17950,N_17840);
nor U18460 (N_18460,N_17582,N_17790);
or U18461 (N_18461,N_17713,N_17702);
nor U18462 (N_18462,N_17952,N_17727);
and U18463 (N_18463,N_17613,N_17778);
xnor U18464 (N_18464,N_17710,N_17795);
or U18465 (N_18465,N_17589,N_17706);
nand U18466 (N_18466,N_17781,N_17893);
and U18467 (N_18467,N_17763,N_17707);
and U18468 (N_18468,N_17978,N_17980);
or U18469 (N_18469,N_17739,N_17638);
and U18470 (N_18470,N_17944,N_17997);
or U18471 (N_18471,N_17577,N_17531);
and U18472 (N_18472,N_17658,N_17964);
and U18473 (N_18473,N_17935,N_17983);
or U18474 (N_18474,N_17545,N_17733);
xor U18475 (N_18475,N_17711,N_17705);
nand U18476 (N_18476,N_17997,N_17753);
nor U18477 (N_18477,N_17818,N_17918);
and U18478 (N_18478,N_17986,N_17660);
nand U18479 (N_18479,N_17748,N_17897);
xor U18480 (N_18480,N_17645,N_17724);
nor U18481 (N_18481,N_17672,N_17760);
or U18482 (N_18482,N_17734,N_17903);
or U18483 (N_18483,N_17930,N_17834);
nand U18484 (N_18484,N_17768,N_17686);
nor U18485 (N_18485,N_17861,N_17679);
xnor U18486 (N_18486,N_17753,N_17899);
or U18487 (N_18487,N_17832,N_17611);
nor U18488 (N_18488,N_17773,N_17797);
or U18489 (N_18489,N_17718,N_17757);
nor U18490 (N_18490,N_17559,N_17616);
nand U18491 (N_18491,N_17538,N_17660);
or U18492 (N_18492,N_17824,N_17939);
nor U18493 (N_18493,N_17703,N_17981);
nor U18494 (N_18494,N_17762,N_17824);
xor U18495 (N_18495,N_17930,N_17841);
or U18496 (N_18496,N_17816,N_17929);
nand U18497 (N_18497,N_17788,N_17687);
and U18498 (N_18498,N_17700,N_17883);
nand U18499 (N_18499,N_17661,N_17980);
nand U18500 (N_18500,N_18235,N_18294);
or U18501 (N_18501,N_18431,N_18257);
nand U18502 (N_18502,N_18231,N_18360);
nand U18503 (N_18503,N_18044,N_18003);
nor U18504 (N_18504,N_18107,N_18036);
and U18505 (N_18505,N_18207,N_18081);
and U18506 (N_18506,N_18262,N_18027);
or U18507 (N_18507,N_18308,N_18042);
and U18508 (N_18508,N_18296,N_18392);
nor U18509 (N_18509,N_18472,N_18031);
nor U18510 (N_18510,N_18118,N_18218);
nand U18511 (N_18511,N_18212,N_18088);
xnor U18512 (N_18512,N_18171,N_18223);
nor U18513 (N_18513,N_18409,N_18421);
xor U18514 (N_18514,N_18200,N_18237);
nor U18515 (N_18515,N_18238,N_18375);
nand U18516 (N_18516,N_18195,N_18180);
nor U18517 (N_18517,N_18252,N_18468);
and U18518 (N_18518,N_18402,N_18350);
or U18519 (N_18519,N_18112,N_18080);
or U18520 (N_18520,N_18256,N_18436);
nand U18521 (N_18521,N_18249,N_18199);
and U18522 (N_18522,N_18444,N_18440);
xor U18523 (N_18523,N_18220,N_18029);
xnor U18524 (N_18524,N_18267,N_18158);
xor U18525 (N_18525,N_18263,N_18279);
xnor U18526 (N_18526,N_18014,N_18146);
nand U18527 (N_18527,N_18433,N_18202);
nand U18528 (N_18528,N_18108,N_18119);
or U18529 (N_18529,N_18287,N_18345);
and U18530 (N_18530,N_18365,N_18101);
or U18531 (N_18531,N_18289,N_18227);
xor U18532 (N_18532,N_18273,N_18366);
xnor U18533 (N_18533,N_18483,N_18233);
and U18534 (N_18534,N_18145,N_18232);
xor U18535 (N_18535,N_18429,N_18214);
nor U18536 (N_18536,N_18068,N_18412);
nor U18537 (N_18537,N_18466,N_18122);
nand U18538 (N_18538,N_18166,N_18435);
nand U18539 (N_18539,N_18033,N_18248);
xor U18540 (N_18540,N_18061,N_18425);
nor U18541 (N_18541,N_18246,N_18497);
and U18542 (N_18542,N_18177,N_18082);
and U18543 (N_18543,N_18313,N_18096);
nand U18544 (N_18544,N_18405,N_18292);
nand U18545 (N_18545,N_18376,N_18150);
nand U18546 (N_18546,N_18113,N_18131);
nor U18547 (N_18547,N_18488,N_18278);
nand U18548 (N_18548,N_18115,N_18407);
and U18549 (N_18549,N_18028,N_18323);
xnor U18550 (N_18550,N_18187,N_18021);
or U18551 (N_18551,N_18379,N_18138);
and U18552 (N_18552,N_18346,N_18065);
nand U18553 (N_18553,N_18439,N_18271);
nor U18554 (N_18554,N_18190,N_18169);
or U18555 (N_18555,N_18456,N_18192);
or U18556 (N_18556,N_18000,N_18393);
nand U18557 (N_18557,N_18400,N_18210);
xnor U18558 (N_18558,N_18089,N_18451);
nor U18559 (N_18559,N_18418,N_18134);
xnor U18560 (N_18560,N_18243,N_18165);
and U18561 (N_18561,N_18139,N_18458);
nor U18562 (N_18562,N_18160,N_18354);
or U18563 (N_18563,N_18475,N_18416);
nand U18564 (N_18564,N_18266,N_18136);
xor U18565 (N_18565,N_18219,N_18198);
nor U18566 (N_18566,N_18361,N_18176);
and U18567 (N_18567,N_18070,N_18413);
or U18568 (N_18568,N_18324,N_18058);
nor U18569 (N_18569,N_18364,N_18447);
nand U18570 (N_18570,N_18295,N_18063);
nor U18571 (N_18571,N_18201,N_18423);
and U18572 (N_18572,N_18084,N_18445);
or U18573 (N_18573,N_18216,N_18245);
xor U18574 (N_18574,N_18135,N_18124);
and U18575 (N_18575,N_18410,N_18196);
nand U18576 (N_18576,N_18398,N_18155);
and U18577 (N_18577,N_18277,N_18471);
xnor U18578 (N_18578,N_18325,N_18351);
nand U18579 (N_18579,N_18406,N_18330);
nor U18580 (N_18580,N_18002,N_18012);
nor U18581 (N_18581,N_18013,N_18420);
or U18582 (N_18582,N_18380,N_18174);
nand U18583 (N_18583,N_18034,N_18419);
nand U18584 (N_18584,N_18011,N_18017);
xnor U18585 (N_18585,N_18205,N_18025);
xor U18586 (N_18586,N_18432,N_18301);
nand U18587 (N_18587,N_18041,N_18496);
nand U18588 (N_18588,N_18396,N_18322);
nand U18589 (N_18589,N_18315,N_18016);
xor U18590 (N_18590,N_18372,N_18007);
and U18591 (N_18591,N_18282,N_18338);
or U18592 (N_18592,N_18052,N_18043);
and U18593 (N_18593,N_18355,N_18302);
and U18594 (N_18594,N_18085,N_18023);
and U18595 (N_18595,N_18288,N_18339);
nand U18596 (N_18596,N_18224,N_18247);
nand U18597 (N_18597,N_18069,N_18344);
and U18598 (N_18598,N_18242,N_18334);
nor U18599 (N_18599,N_18141,N_18056);
and U18600 (N_18600,N_18464,N_18481);
and U18601 (N_18601,N_18328,N_18213);
nor U18602 (N_18602,N_18221,N_18388);
nand U18603 (N_18603,N_18280,N_18422);
nand U18604 (N_18604,N_18083,N_18179);
nand U18605 (N_18605,N_18383,N_18127);
xnor U18606 (N_18606,N_18045,N_18222);
nor U18607 (N_18607,N_18309,N_18125);
nand U18608 (N_18608,N_18241,N_18097);
or U18609 (N_18609,N_18321,N_18186);
nor U18610 (N_18610,N_18395,N_18384);
xor U18611 (N_18611,N_18251,N_18206);
xor U18612 (N_18612,N_18073,N_18164);
xor U18613 (N_18613,N_18306,N_18106);
or U18614 (N_18614,N_18123,N_18074);
and U18615 (N_18615,N_18281,N_18168);
nand U18616 (N_18616,N_18269,N_18454);
or U18617 (N_18617,N_18417,N_18408);
nor U18618 (N_18618,N_18092,N_18250);
and U18619 (N_18619,N_18030,N_18414);
or U18620 (N_18620,N_18485,N_18318);
nand U18621 (N_18621,N_18194,N_18154);
nor U18622 (N_18622,N_18078,N_18102);
xnor U18623 (N_18623,N_18491,N_18381);
xnor U18624 (N_18624,N_18461,N_18236);
xnor U18625 (N_18625,N_18182,N_18293);
and U18626 (N_18626,N_18310,N_18151);
or U18627 (N_18627,N_18153,N_18071);
xor U18628 (N_18628,N_18333,N_18480);
xnor U18629 (N_18629,N_18215,N_18457);
nand U18630 (N_18630,N_18140,N_18050);
and U18631 (N_18631,N_18387,N_18019);
and U18632 (N_18632,N_18047,N_18455);
xnor U18633 (N_18633,N_18428,N_18109);
nor U18634 (N_18634,N_18188,N_18357);
nor U18635 (N_18635,N_18048,N_18037);
or U18636 (N_18636,N_18314,N_18087);
xnor U18637 (N_18637,N_18356,N_18385);
xnor U18638 (N_18638,N_18265,N_18172);
and U18639 (N_18639,N_18446,N_18072);
nor U18640 (N_18640,N_18337,N_18253);
nand U18641 (N_18641,N_18430,N_18374);
nand U18642 (N_18642,N_18272,N_18264);
and U18643 (N_18643,N_18448,N_18476);
xnor U18644 (N_18644,N_18283,N_18258);
and U18645 (N_18645,N_18185,N_18130);
nor U18646 (N_18646,N_18303,N_18067);
or U18647 (N_18647,N_18137,N_18059);
nor U18648 (N_18648,N_18291,N_18299);
nor U18649 (N_18649,N_18259,N_18053);
and U18650 (N_18650,N_18449,N_18015);
xnor U18651 (N_18651,N_18347,N_18204);
and U18652 (N_18652,N_18352,N_18482);
and U18653 (N_18653,N_18434,N_18394);
nand U18654 (N_18654,N_18142,N_18152);
xnor U18655 (N_18655,N_18285,N_18450);
xor U18656 (N_18656,N_18270,N_18427);
and U18657 (N_18657,N_18358,N_18051);
xnor U18658 (N_18658,N_18239,N_18319);
nand U18659 (N_18659,N_18305,N_18184);
xor U18660 (N_18660,N_18062,N_18167);
and U18661 (N_18661,N_18484,N_18170);
or U18662 (N_18662,N_18441,N_18369);
and U18663 (N_18663,N_18230,N_18143);
nand U18664 (N_18664,N_18474,N_18329);
nor U18665 (N_18665,N_18103,N_18286);
nor U18666 (N_18666,N_18075,N_18367);
nor U18667 (N_18667,N_18126,N_18090);
nand U18668 (N_18668,N_18401,N_18371);
and U18669 (N_18669,N_18320,N_18426);
and U18670 (N_18670,N_18095,N_18332);
xor U18671 (N_18671,N_18175,N_18260);
and U18672 (N_18672,N_18348,N_18462);
or U18673 (N_18673,N_18024,N_18159);
and U18674 (N_18674,N_18039,N_18349);
or U18675 (N_18675,N_18261,N_18006);
and U18676 (N_18676,N_18133,N_18276);
nor U18677 (N_18677,N_18386,N_18226);
or U18678 (N_18678,N_18486,N_18442);
nand U18679 (N_18679,N_18121,N_18370);
or U18680 (N_18680,N_18217,N_18336);
xnor U18681 (N_18681,N_18162,N_18004);
and U18682 (N_18682,N_18255,N_18064);
xor U18683 (N_18683,N_18490,N_18335);
xnor U18684 (N_18684,N_18390,N_18066);
xnor U18685 (N_18685,N_18353,N_18437);
xor U18686 (N_18686,N_18001,N_18403);
and U18687 (N_18687,N_18443,N_18300);
xnor U18688 (N_18688,N_18312,N_18094);
and U18689 (N_18689,N_18228,N_18368);
nor U18690 (N_18690,N_18391,N_18341);
or U18691 (N_18691,N_18010,N_18077);
nor U18692 (N_18692,N_18467,N_18378);
and U18693 (N_18693,N_18163,N_18203);
nand U18694 (N_18694,N_18463,N_18492);
nand U18695 (N_18695,N_18415,N_18040);
or U18696 (N_18696,N_18307,N_18178);
and U18697 (N_18697,N_18284,N_18487);
xor U18698 (N_18698,N_18197,N_18477);
nand U18699 (N_18699,N_18297,N_18149);
and U18700 (N_18700,N_18499,N_18093);
nor U18701 (N_18701,N_18193,N_18018);
nand U18702 (N_18702,N_18128,N_18234);
and U18703 (N_18703,N_18469,N_18331);
and U18704 (N_18704,N_18020,N_18493);
nor U18705 (N_18705,N_18452,N_18240);
xnor U18706 (N_18706,N_18110,N_18022);
xor U18707 (N_18707,N_18032,N_18129);
and U18708 (N_18708,N_18116,N_18148);
xnor U18709 (N_18709,N_18343,N_18111);
or U18710 (N_18710,N_18120,N_18498);
or U18711 (N_18711,N_18459,N_18317);
or U18712 (N_18712,N_18495,N_18114);
nand U18713 (N_18713,N_18311,N_18225);
xnor U18714 (N_18714,N_18091,N_18086);
nor U18715 (N_18715,N_18161,N_18183);
nor U18716 (N_18716,N_18211,N_18340);
and U18717 (N_18717,N_18274,N_18399);
xnor U18718 (N_18718,N_18099,N_18460);
nor U18719 (N_18719,N_18104,N_18147);
and U18720 (N_18720,N_18009,N_18229);
nand U18721 (N_18721,N_18005,N_18290);
nand U18722 (N_18722,N_18268,N_18060);
xnor U18723 (N_18723,N_18411,N_18173);
or U18724 (N_18724,N_18181,N_18494);
and U18725 (N_18725,N_18342,N_18326);
nand U18726 (N_18726,N_18362,N_18054);
or U18727 (N_18727,N_18156,N_18035);
xor U18728 (N_18728,N_18098,N_18100);
xnor U18729 (N_18729,N_18438,N_18046);
and U18730 (N_18730,N_18208,N_18244);
nand U18731 (N_18731,N_18008,N_18453);
or U18732 (N_18732,N_18327,N_18038);
or U18733 (N_18733,N_18465,N_18117);
xor U18734 (N_18734,N_18209,N_18389);
nand U18735 (N_18735,N_18304,N_18479);
nor U18736 (N_18736,N_18105,N_18026);
nand U18737 (N_18737,N_18359,N_18382);
xnor U18738 (N_18738,N_18316,N_18473);
nor U18739 (N_18739,N_18144,N_18404);
xor U18740 (N_18740,N_18470,N_18076);
and U18741 (N_18741,N_18055,N_18057);
or U18742 (N_18742,N_18049,N_18157);
nand U18743 (N_18743,N_18189,N_18254);
or U18744 (N_18744,N_18489,N_18424);
or U18745 (N_18745,N_18079,N_18298);
xnor U18746 (N_18746,N_18191,N_18373);
nand U18747 (N_18747,N_18132,N_18478);
nor U18748 (N_18748,N_18275,N_18377);
xor U18749 (N_18749,N_18397,N_18363);
xor U18750 (N_18750,N_18141,N_18413);
nor U18751 (N_18751,N_18284,N_18007);
nor U18752 (N_18752,N_18084,N_18486);
xnor U18753 (N_18753,N_18091,N_18088);
nand U18754 (N_18754,N_18149,N_18390);
nor U18755 (N_18755,N_18117,N_18008);
and U18756 (N_18756,N_18302,N_18000);
or U18757 (N_18757,N_18156,N_18257);
xnor U18758 (N_18758,N_18015,N_18026);
nor U18759 (N_18759,N_18383,N_18349);
xor U18760 (N_18760,N_18179,N_18178);
or U18761 (N_18761,N_18385,N_18408);
nand U18762 (N_18762,N_18111,N_18348);
and U18763 (N_18763,N_18382,N_18017);
and U18764 (N_18764,N_18242,N_18498);
xnor U18765 (N_18765,N_18483,N_18013);
xor U18766 (N_18766,N_18325,N_18192);
nand U18767 (N_18767,N_18381,N_18395);
xor U18768 (N_18768,N_18394,N_18244);
and U18769 (N_18769,N_18366,N_18142);
nor U18770 (N_18770,N_18415,N_18414);
xor U18771 (N_18771,N_18199,N_18021);
nand U18772 (N_18772,N_18334,N_18368);
xor U18773 (N_18773,N_18003,N_18339);
nor U18774 (N_18774,N_18402,N_18050);
nand U18775 (N_18775,N_18470,N_18336);
or U18776 (N_18776,N_18298,N_18426);
nor U18777 (N_18777,N_18071,N_18174);
xnor U18778 (N_18778,N_18210,N_18124);
or U18779 (N_18779,N_18086,N_18251);
xnor U18780 (N_18780,N_18199,N_18246);
and U18781 (N_18781,N_18251,N_18218);
nor U18782 (N_18782,N_18366,N_18111);
xor U18783 (N_18783,N_18146,N_18350);
or U18784 (N_18784,N_18304,N_18307);
xnor U18785 (N_18785,N_18263,N_18475);
nand U18786 (N_18786,N_18446,N_18241);
nor U18787 (N_18787,N_18297,N_18231);
and U18788 (N_18788,N_18255,N_18202);
nor U18789 (N_18789,N_18444,N_18145);
nand U18790 (N_18790,N_18001,N_18290);
xor U18791 (N_18791,N_18102,N_18399);
nor U18792 (N_18792,N_18295,N_18463);
nand U18793 (N_18793,N_18457,N_18052);
nor U18794 (N_18794,N_18016,N_18397);
nor U18795 (N_18795,N_18362,N_18125);
or U18796 (N_18796,N_18412,N_18353);
or U18797 (N_18797,N_18481,N_18074);
nor U18798 (N_18798,N_18292,N_18431);
or U18799 (N_18799,N_18496,N_18150);
nor U18800 (N_18800,N_18378,N_18478);
and U18801 (N_18801,N_18081,N_18088);
nand U18802 (N_18802,N_18126,N_18318);
and U18803 (N_18803,N_18109,N_18404);
and U18804 (N_18804,N_18099,N_18348);
xnor U18805 (N_18805,N_18135,N_18334);
nor U18806 (N_18806,N_18371,N_18201);
nor U18807 (N_18807,N_18135,N_18458);
or U18808 (N_18808,N_18029,N_18476);
xnor U18809 (N_18809,N_18252,N_18475);
and U18810 (N_18810,N_18064,N_18338);
or U18811 (N_18811,N_18019,N_18102);
or U18812 (N_18812,N_18464,N_18143);
nand U18813 (N_18813,N_18111,N_18282);
or U18814 (N_18814,N_18128,N_18424);
nand U18815 (N_18815,N_18427,N_18436);
xor U18816 (N_18816,N_18207,N_18349);
nor U18817 (N_18817,N_18433,N_18247);
nor U18818 (N_18818,N_18453,N_18057);
nor U18819 (N_18819,N_18280,N_18302);
and U18820 (N_18820,N_18236,N_18391);
nand U18821 (N_18821,N_18320,N_18342);
or U18822 (N_18822,N_18205,N_18478);
nor U18823 (N_18823,N_18075,N_18387);
and U18824 (N_18824,N_18035,N_18346);
xor U18825 (N_18825,N_18369,N_18475);
nand U18826 (N_18826,N_18133,N_18064);
or U18827 (N_18827,N_18220,N_18207);
nor U18828 (N_18828,N_18192,N_18096);
or U18829 (N_18829,N_18461,N_18023);
xor U18830 (N_18830,N_18237,N_18471);
or U18831 (N_18831,N_18276,N_18271);
or U18832 (N_18832,N_18346,N_18429);
or U18833 (N_18833,N_18037,N_18417);
nor U18834 (N_18834,N_18436,N_18134);
nor U18835 (N_18835,N_18250,N_18439);
xnor U18836 (N_18836,N_18481,N_18425);
nand U18837 (N_18837,N_18375,N_18131);
nand U18838 (N_18838,N_18064,N_18053);
or U18839 (N_18839,N_18091,N_18215);
and U18840 (N_18840,N_18268,N_18266);
or U18841 (N_18841,N_18389,N_18207);
and U18842 (N_18842,N_18291,N_18020);
and U18843 (N_18843,N_18324,N_18301);
and U18844 (N_18844,N_18329,N_18495);
and U18845 (N_18845,N_18137,N_18142);
or U18846 (N_18846,N_18469,N_18302);
and U18847 (N_18847,N_18025,N_18482);
nand U18848 (N_18848,N_18115,N_18490);
and U18849 (N_18849,N_18305,N_18398);
xor U18850 (N_18850,N_18290,N_18033);
nand U18851 (N_18851,N_18452,N_18199);
nand U18852 (N_18852,N_18317,N_18399);
xnor U18853 (N_18853,N_18107,N_18098);
or U18854 (N_18854,N_18387,N_18446);
and U18855 (N_18855,N_18127,N_18156);
and U18856 (N_18856,N_18015,N_18365);
xor U18857 (N_18857,N_18351,N_18131);
xor U18858 (N_18858,N_18132,N_18262);
and U18859 (N_18859,N_18397,N_18086);
nor U18860 (N_18860,N_18274,N_18443);
and U18861 (N_18861,N_18038,N_18176);
nand U18862 (N_18862,N_18123,N_18065);
nor U18863 (N_18863,N_18428,N_18007);
nand U18864 (N_18864,N_18426,N_18493);
nor U18865 (N_18865,N_18247,N_18199);
xnor U18866 (N_18866,N_18280,N_18174);
nor U18867 (N_18867,N_18278,N_18482);
xnor U18868 (N_18868,N_18073,N_18395);
nand U18869 (N_18869,N_18168,N_18079);
or U18870 (N_18870,N_18229,N_18460);
nand U18871 (N_18871,N_18010,N_18261);
nor U18872 (N_18872,N_18170,N_18193);
nand U18873 (N_18873,N_18208,N_18402);
or U18874 (N_18874,N_18340,N_18039);
xnor U18875 (N_18875,N_18302,N_18142);
xor U18876 (N_18876,N_18245,N_18110);
xnor U18877 (N_18877,N_18457,N_18219);
nor U18878 (N_18878,N_18054,N_18192);
nand U18879 (N_18879,N_18102,N_18229);
nand U18880 (N_18880,N_18302,N_18022);
nand U18881 (N_18881,N_18488,N_18241);
or U18882 (N_18882,N_18390,N_18410);
or U18883 (N_18883,N_18497,N_18057);
or U18884 (N_18884,N_18450,N_18454);
and U18885 (N_18885,N_18349,N_18367);
xor U18886 (N_18886,N_18050,N_18058);
or U18887 (N_18887,N_18181,N_18050);
nand U18888 (N_18888,N_18145,N_18300);
nor U18889 (N_18889,N_18272,N_18436);
xnor U18890 (N_18890,N_18407,N_18277);
and U18891 (N_18891,N_18381,N_18422);
or U18892 (N_18892,N_18057,N_18257);
xor U18893 (N_18893,N_18252,N_18005);
or U18894 (N_18894,N_18096,N_18115);
nor U18895 (N_18895,N_18463,N_18001);
xnor U18896 (N_18896,N_18252,N_18358);
nand U18897 (N_18897,N_18487,N_18148);
xnor U18898 (N_18898,N_18321,N_18029);
nor U18899 (N_18899,N_18034,N_18346);
nor U18900 (N_18900,N_18070,N_18310);
and U18901 (N_18901,N_18075,N_18199);
and U18902 (N_18902,N_18481,N_18168);
and U18903 (N_18903,N_18457,N_18417);
nand U18904 (N_18904,N_18220,N_18090);
and U18905 (N_18905,N_18326,N_18128);
nand U18906 (N_18906,N_18228,N_18343);
xor U18907 (N_18907,N_18396,N_18221);
nor U18908 (N_18908,N_18222,N_18444);
and U18909 (N_18909,N_18089,N_18108);
nor U18910 (N_18910,N_18166,N_18248);
xor U18911 (N_18911,N_18375,N_18253);
or U18912 (N_18912,N_18144,N_18174);
nor U18913 (N_18913,N_18181,N_18464);
xor U18914 (N_18914,N_18113,N_18149);
nor U18915 (N_18915,N_18063,N_18071);
nand U18916 (N_18916,N_18249,N_18376);
nor U18917 (N_18917,N_18051,N_18085);
xor U18918 (N_18918,N_18277,N_18302);
nor U18919 (N_18919,N_18248,N_18160);
nor U18920 (N_18920,N_18103,N_18041);
xnor U18921 (N_18921,N_18372,N_18316);
and U18922 (N_18922,N_18462,N_18483);
or U18923 (N_18923,N_18313,N_18273);
nor U18924 (N_18924,N_18474,N_18355);
or U18925 (N_18925,N_18086,N_18335);
and U18926 (N_18926,N_18137,N_18109);
or U18927 (N_18927,N_18059,N_18158);
or U18928 (N_18928,N_18446,N_18158);
xor U18929 (N_18929,N_18025,N_18020);
or U18930 (N_18930,N_18018,N_18208);
nand U18931 (N_18931,N_18073,N_18497);
or U18932 (N_18932,N_18343,N_18281);
nor U18933 (N_18933,N_18407,N_18166);
nand U18934 (N_18934,N_18460,N_18081);
and U18935 (N_18935,N_18257,N_18412);
and U18936 (N_18936,N_18313,N_18136);
or U18937 (N_18937,N_18016,N_18454);
and U18938 (N_18938,N_18436,N_18408);
or U18939 (N_18939,N_18108,N_18060);
nor U18940 (N_18940,N_18054,N_18136);
nor U18941 (N_18941,N_18318,N_18423);
xnor U18942 (N_18942,N_18339,N_18178);
nand U18943 (N_18943,N_18266,N_18488);
xnor U18944 (N_18944,N_18044,N_18269);
nand U18945 (N_18945,N_18156,N_18280);
or U18946 (N_18946,N_18126,N_18426);
xnor U18947 (N_18947,N_18432,N_18398);
and U18948 (N_18948,N_18010,N_18030);
nor U18949 (N_18949,N_18382,N_18050);
or U18950 (N_18950,N_18362,N_18453);
nand U18951 (N_18951,N_18241,N_18377);
or U18952 (N_18952,N_18365,N_18098);
or U18953 (N_18953,N_18033,N_18420);
or U18954 (N_18954,N_18287,N_18376);
or U18955 (N_18955,N_18215,N_18090);
nand U18956 (N_18956,N_18266,N_18048);
nand U18957 (N_18957,N_18169,N_18269);
or U18958 (N_18958,N_18445,N_18054);
nand U18959 (N_18959,N_18135,N_18002);
nand U18960 (N_18960,N_18026,N_18102);
xnor U18961 (N_18961,N_18296,N_18467);
xnor U18962 (N_18962,N_18328,N_18443);
and U18963 (N_18963,N_18160,N_18093);
and U18964 (N_18964,N_18325,N_18426);
and U18965 (N_18965,N_18081,N_18213);
nor U18966 (N_18966,N_18326,N_18041);
or U18967 (N_18967,N_18199,N_18019);
nor U18968 (N_18968,N_18397,N_18227);
nor U18969 (N_18969,N_18086,N_18184);
nor U18970 (N_18970,N_18279,N_18337);
xor U18971 (N_18971,N_18266,N_18322);
or U18972 (N_18972,N_18113,N_18465);
xor U18973 (N_18973,N_18340,N_18320);
nand U18974 (N_18974,N_18494,N_18307);
and U18975 (N_18975,N_18417,N_18169);
nand U18976 (N_18976,N_18231,N_18072);
nand U18977 (N_18977,N_18389,N_18077);
nor U18978 (N_18978,N_18255,N_18275);
nor U18979 (N_18979,N_18358,N_18065);
nand U18980 (N_18980,N_18127,N_18288);
and U18981 (N_18981,N_18272,N_18302);
and U18982 (N_18982,N_18203,N_18294);
xor U18983 (N_18983,N_18160,N_18176);
nor U18984 (N_18984,N_18401,N_18122);
or U18985 (N_18985,N_18370,N_18131);
or U18986 (N_18986,N_18301,N_18103);
and U18987 (N_18987,N_18259,N_18376);
nor U18988 (N_18988,N_18064,N_18342);
nand U18989 (N_18989,N_18176,N_18447);
or U18990 (N_18990,N_18451,N_18432);
xor U18991 (N_18991,N_18459,N_18140);
nand U18992 (N_18992,N_18333,N_18275);
nor U18993 (N_18993,N_18395,N_18003);
nor U18994 (N_18994,N_18129,N_18366);
nor U18995 (N_18995,N_18196,N_18093);
nor U18996 (N_18996,N_18247,N_18293);
nand U18997 (N_18997,N_18379,N_18268);
and U18998 (N_18998,N_18423,N_18450);
or U18999 (N_18999,N_18115,N_18308);
xor U19000 (N_19000,N_18516,N_18648);
xnor U19001 (N_19001,N_18582,N_18927);
nand U19002 (N_19002,N_18738,N_18896);
and U19003 (N_19003,N_18803,N_18628);
xor U19004 (N_19004,N_18814,N_18613);
xor U19005 (N_19005,N_18694,N_18609);
or U19006 (N_19006,N_18710,N_18602);
xor U19007 (N_19007,N_18600,N_18715);
nor U19008 (N_19008,N_18765,N_18953);
or U19009 (N_19009,N_18566,N_18721);
or U19010 (N_19010,N_18698,N_18911);
nand U19011 (N_19011,N_18697,N_18769);
or U19012 (N_19012,N_18887,N_18846);
nor U19013 (N_19013,N_18825,N_18674);
nand U19014 (N_19014,N_18834,N_18699);
xor U19015 (N_19015,N_18794,N_18914);
or U19016 (N_19016,N_18865,N_18513);
nor U19017 (N_19017,N_18923,N_18898);
nand U19018 (N_19018,N_18536,N_18977);
nor U19019 (N_19019,N_18922,N_18562);
nor U19020 (N_19020,N_18855,N_18670);
nand U19021 (N_19021,N_18622,N_18596);
xor U19022 (N_19022,N_18877,N_18618);
xor U19023 (N_19023,N_18610,N_18564);
nand U19024 (N_19024,N_18666,N_18965);
xor U19025 (N_19025,N_18508,N_18505);
nor U19026 (N_19026,N_18815,N_18942);
xor U19027 (N_19027,N_18801,N_18890);
or U19028 (N_19028,N_18547,N_18879);
nand U19029 (N_19029,N_18621,N_18617);
or U19030 (N_19030,N_18510,N_18591);
nand U19031 (N_19031,N_18875,N_18827);
and U19032 (N_19032,N_18806,N_18581);
or U19033 (N_19033,N_18974,N_18878);
or U19034 (N_19034,N_18804,N_18713);
nand U19035 (N_19035,N_18862,N_18893);
nand U19036 (N_19036,N_18656,N_18573);
or U19037 (N_19037,N_18538,N_18945);
and U19038 (N_19038,N_18662,N_18722);
nor U19039 (N_19039,N_18627,N_18657);
and U19040 (N_19040,N_18521,N_18874);
or U19041 (N_19041,N_18841,N_18908);
xor U19042 (N_19042,N_18671,N_18660);
or U19043 (N_19043,N_18557,N_18859);
nand U19044 (N_19044,N_18623,N_18525);
xnor U19045 (N_19045,N_18812,N_18523);
and U19046 (N_19046,N_18730,N_18552);
xnor U19047 (N_19047,N_18732,N_18717);
nand U19048 (N_19048,N_18941,N_18588);
nor U19049 (N_19049,N_18541,N_18635);
and U19050 (N_19050,N_18807,N_18767);
and U19051 (N_19051,N_18861,N_18586);
or U19052 (N_19052,N_18719,N_18615);
and U19053 (N_19053,N_18864,N_18823);
xnor U19054 (N_19054,N_18759,N_18956);
nand U19055 (N_19055,N_18842,N_18917);
and U19056 (N_19056,N_18770,N_18563);
nand U19057 (N_19057,N_18661,N_18796);
nor U19058 (N_19058,N_18940,N_18681);
xor U19059 (N_19059,N_18958,N_18675);
nor U19060 (N_19060,N_18542,N_18649);
and U19061 (N_19061,N_18873,N_18976);
xor U19062 (N_19062,N_18659,N_18998);
xor U19063 (N_19063,N_18668,N_18575);
nand U19064 (N_19064,N_18565,N_18546);
nor U19065 (N_19065,N_18848,N_18718);
xor U19066 (N_19066,N_18789,N_18757);
xnor U19067 (N_19067,N_18943,N_18933);
nand U19068 (N_19068,N_18693,N_18678);
or U19069 (N_19069,N_18733,N_18947);
nor U19070 (N_19070,N_18828,N_18840);
and U19071 (N_19071,N_18534,N_18500);
xor U19072 (N_19072,N_18626,N_18743);
nor U19073 (N_19073,N_18737,N_18851);
nand U19074 (N_19074,N_18589,N_18816);
nor U19075 (N_19075,N_18689,N_18640);
or U19076 (N_19076,N_18792,N_18558);
and U19077 (N_19077,N_18939,N_18909);
or U19078 (N_19078,N_18752,N_18625);
or U19079 (N_19079,N_18768,N_18745);
xnor U19080 (N_19080,N_18696,N_18643);
and U19081 (N_19081,N_18756,N_18912);
and U19082 (N_19082,N_18795,N_18820);
xnor U19083 (N_19083,N_18830,N_18747);
and U19084 (N_19084,N_18599,N_18568);
nand U19085 (N_19085,N_18906,N_18734);
nand U19086 (N_19086,N_18835,N_18569);
and U19087 (N_19087,N_18603,N_18714);
nand U19088 (N_19088,N_18856,N_18637);
nor U19089 (N_19089,N_18687,N_18780);
or U19090 (N_19090,N_18870,N_18549);
nor U19091 (N_19091,N_18785,N_18584);
nor U19092 (N_19092,N_18818,N_18900);
xor U19093 (N_19093,N_18918,N_18969);
nand U19094 (N_19094,N_18968,N_18984);
or U19095 (N_19095,N_18781,N_18983);
nor U19096 (N_19096,N_18527,N_18624);
nor U19097 (N_19097,N_18892,N_18629);
and U19098 (N_19098,N_18799,N_18838);
xnor U19099 (N_19099,N_18729,N_18886);
and U19100 (N_19100,N_18520,N_18614);
nand U19101 (N_19101,N_18979,N_18533);
nor U19102 (N_19102,N_18994,N_18949);
or U19103 (N_19103,N_18790,N_18559);
xor U19104 (N_19104,N_18779,N_18585);
and U19105 (N_19105,N_18880,N_18881);
xor U19106 (N_19106,N_18630,N_18951);
and U19107 (N_19107,N_18761,N_18511);
nor U19108 (N_19108,N_18579,N_18889);
xor U19109 (N_19109,N_18946,N_18805);
xnor U19110 (N_19110,N_18636,N_18616);
nor U19111 (N_19111,N_18858,N_18695);
or U19112 (N_19112,N_18903,N_18854);
nand U19113 (N_19113,N_18791,N_18829);
and U19114 (N_19114,N_18691,N_18680);
xor U19115 (N_19115,N_18905,N_18529);
xnor U19116 (N_19116,N_18611,N_18959);
and U19117 (N_19117,N_18888,N_18783);
nor U19118 (N_19118,N_18831,N_18571);
nor U19119 (N_19119,N_18995,N_18703);
xnor U19120 (N_19120,N_18782,N_18576);
and U19121 (N_19121,N_18619,N_18587);
and U19122 (N_19122,N_18607,N_18988);
nand U19123 (N_19123,N_18742,N_18836);
or U19124 (N_19124,N_18952,N_18999);
or U19125 (N_19125,N_18981,N_18773);
nand U19126 (N_19126,N_18899,N_18819);
nor U19127 (N_19127,N_18705,N_18539);
and U19128 (N_19128,N_18650,N_18750);
or U19129 (N_19129,N_18688,N_18669);
nand U19130 (N_19130,N_18551,N_18679);
nor U19131 (N_19131,N_18894,N_18583);
or U19132 (N_19132,N_18633,N_18727);
nand U19133 (N_19133,N_18808,N_18639);
nand U19134 (N_19134,N_18777,N_18548);
nor U19135 (N_19135,N_18537,N_18793);
or U19136 (N_19136,N_18686,N_18904);
nand U19137 (N_19137,N_18802,N_18753);
nor U19138 (N_19138,N_18967,N_18866);
or U19139 (N_19139,N_18936,N_18833);
xnor U19140 (N_19140,N_18692,N_18701);
or U19141 (N_19141,N_18944,N_18519);
nand U19142 (N_19142,N_18535,N_18708);
or U19143 (N_19143,N_18684,N_18755);
or U19144 (N_19144,N_18762,N_18658);
and U19145 (N_19145,N_18707,N_18677);
xor U19146 (N_19146,N_18740,N_18863);
nor U19147 (N_19147,N_18673,N_18950);
nor U19148 (N_19148,N_18506,N_18891);
xor U19149 (N_19149,N_18665,N_18849);
or U19150 (N_19150,N_18934,N_18763);
xor U19151 (N_19151,N_18960,N_18731);
nand U19152 (N_19152,N_18991,N_18797);
or U19153 (N_19153,N_18578,N_18935);
nand U19154 (N_19154,N_18663,N_18593);
nor U19155 (N_19155,N_18570,N_18809);
nor U19156 (N_19156,N_18826,N_18970);
and U19157 (N_19157,N_18672,N_18915);
nor U19158 (N_19158,N_18822,N_18509);
or U19159 (N_19159,N_18852,N_18726);
nand U19160 (N_19160,N_18544,N_18774);
or U19161 (N_19161,N_18844,N_18594);
or U19162 (N_19162,N_18992,N_18735);
and U19163 (N_19163,N_18772,N_18642);
and U19164 (N_19164,N_18524,N_18530);
nand U19165 (N_19165,N_18932,N_18518);
or U19166 (N_19166,N_18653,N_18634);
nor U19167 (N_19167,N_18645,N_18954);
xnor U19168 (N_19168,N_18916,N_18595);
and U19169 (N_19169,N_18728,N_18925);
nand U19170 (N_19170,N_18667,N_18771);
nand U19171 (N_19171,N_18741,N_18545);
and U19172 (N_19172,N_18647,N_18683);
or U19173 (N_19173,N_18567,N_18857);
nor U19174 (N_19174,N_18504,N_18522);
and U19175 (N_19175,N_18937,N_18920);
and U19176 (N_19176,N_18971,N_18832);
xnor U19177 (N_19177,N_18641,N_18929);
and U19178 (N_19178,N_18989,N_18902);
nor U19179 (N_19179,N_18601,N_18948);
and U19180 (N_19180,N_18690,N_18612);
and U19181 (N_19181,N_18543,N_18860);
and U19182 (N_19182,N_18501,N_18554);
nor U19183 (N_19183,N_18926,N_18850);
nor U19184 (N_19184,N_18608,N_18644);
xnor U19185 (N_19185,N_18638,N_18990);
nand U19186 (N_19186,N_18813,N_18606);
nand U19187 (N_19187,N_18532,N_18632);
and U19188 (N_19188,N_18955,N_18821);
nor U19189 (N_19189,N_18883,N_18555);
xnor U19190 (N_19190,N_18716,N_18869);
or U19191 (N_19191,N_18775,N_18884);
nor U19192 (N_19192,N_18872,N_18682);
or U19193 (N_19193,N_18592,N_18928);
nand U19194 (N_19194,N_18963,N_18997);
or U19195 (N_19195,N_18924,N_18910);
and U19196 (N_19196,N_18938,N_18655);
and U19197 (N_19197,N_18982,N_18531);
and U19198 (N_19198,N_18597,N_18764);
nor U19199 (N_19199,N_18986,N_18550);
nor U19200 (N_19200,N_18574,N_18885);
xor U19201 (N_19201,N_18975,N_18631);
nand U19202 (N_19202,N_18503,N_18811);
xnor U19203 (N_19203,N_18706,N_18972);
xnor U19204 (N_19204,N_18867,N_18786);
nor U19205 (N_19205,N_18652,N_18810);
and U19206 (N_19206,N_18853,N_18528);
or U19207 (N_19207,N_18847,N_18572);
xor U19208 (N_19208,N_18739,N_18664);
xor U19209 (N_19209,N_18973,N_18845);
nor U19210 (N_19210,N_18798,N_18766);
xor U19211 (N_19211,N_18711,N_18676);
xnor U19212 (N_19212,N_18560,N_18839);
nor U19213 (N_19213,N_18784,N_18748);
nand U19214 (N_19214,N_18871,N_18709);
or U19215 (N_19215,N_18685,N_18540);
nor U19216 (N_19216,N_18744,N_18978);
and U19217 (N_19217,N_18980,N_18749);
or U19218 (N_19218,N_18646,N_18843);
nor U19219 (N_19219,N_18580,N_18913);
nand U19220 (N_19220,N_18651,N_18895);
or U19221 (N_19221,N_18962,N_18526);
nand U19222 (N_19222,N_18907,N_18987);
nor U19223 (N_19223,N_18620,N_18961);
nor U19224 (N_19224,N_18901,N_18882);
or U19225 (N_19225,N_18760,N_18800);
nand U19226 (N_19226,N_18868,N_18778);
or U19227 (N_19227,N_18702,N_18515);
and U19228 (N_19228,N_18930,N_18931);
and U19229 (N_19229,N_18512,N_18712);
xor U19230 (N_19230,N_18577,N_18897);
and U19231 (N_19231,N_18704,N_18725);
nor U19232 (N_19232,N_18590,N_18921);
and U19233 (N_19233,N_18754,N_18966);
nor U19234 (N_19234,N_18957,N_18556);
nand U19235 (N_19235,N_18605,N_18758);
nor U19236 (N_19236,N_18985,N_18788);
or U19237 (N_19237,N_18787,N_18824);
and U19238 (N_19238,N_18751,N_18817);
nand U19239 (N_19239,N_18723,N_18700);
nor U19240 (N_19240,N_18507,N_18837);
and U19241 (N_19241,N_18876,N_18553);
xor U19242 (N_19242,N_18746,N_18517);
xnor U19243 (N_19243,N_18720,N_18502);
nand U19244 (N_19244,N_18919,N_18776);
and U19245 (N_19245,N_18654,N_18724);
nand U19246 (N_19246,N_18993,N_18964);
or U19247 (N_19247,N_18561,N_18604);
nand U19248 (N_19248,N_18598,N_18736);
xnor U19249 (N_19249,N_18514,N_18996);
nand U19250 (N_19250,N_18683,N_18924);
nand U19251 (N_19251,N_18888,N_18983);
or U19252 (N_19252,N_18743,N_18985);
nand U19253 (N_19253,N_18770,N_18645);
or U19254 (N_19254,N_18704,N_18876);
and U19255 (N_19255,N_18702,N_18610);
or U19256 (N_19256,N_18628,N_18815);
nand U19257 (N_19257,N_18637,N_18525);
or U19258 (N_19258,N_18966,N_18749);
xor U19259 (N_19259,N_18649,N_18798);
or U19260 (N_19260,N_18632,N_18597);
or U19261 (N_19261,N_18523,N_18653);
nor U19262 (N_19262,N_18731,N_18940);
nand U19263 (N_19263,N_18912,N_18544);
or U19264 (N_19264,N_18543,N_18537);
nor U19265 (N_19265,N_18664,N_18926);
xnor U19266 (N_19266,N_18620,N_18746);
nand U19267 (N_19267,N_18610,N_18538);
nor U19268 (N_19268,N_18834,N_18744);
and U19269 (N_19269,N_18557,N_18972);
nor U19270 (N_19270,N_18824,N_18585);
or U19271 (N_19271,N_18686,N_18666);
and U19272 (N_19272,N_18584,N_18669);
nor U19273 (N_19273,N_18620,N_18733);
nand U19274 (N_19274,N_18643,N_18718);
nand U19275 (N_19275,N_18654,N_18845);
nand U19276 (N_19276,N_18805,N_18867);
nand U19277 (N_19277,N_18839,N_18769);
nand U19278 (N_19278,N_18727,N_18867);
nand U19279 (N_19279,N_18938,N_18926);
xnor U19280 (N_19280,N_18944,N_18824);
or U19281 (N_19281,N_18693,N_18845);
and U19282 (N_19282,N_18743,N_18845);
and U19283 (N_19283,N_18746,N_18573);
xnor U19284 (N_19284,N_18618,N_18689);
or U19285 (N_19285,N_18777,N_18931);
nor U19286 (N_19286,N_18755,N_18610);
xnor U19287 (N_19287,N_18988,N_18826);
and U19288 (N_19288,N_18858,N_18907);
and U19289 (N_19289,N_18662,N_18502);
xor U19290 (N_19290,N_18729,N_18764);
xor U19291 (N_19291,N_18611,N_18637);
nand U19292 (N_19292,N_18951,N_18654);
and U19293 (N_19293,N_18595,N_18981);
nand U19294 (N_19294,N_18892,N_18595);
nor U19295 (N_19295,N_18766,N_18787);
xor U19296 (N_19296,N_18633,N_18808);
and U19297 (N_19297,N_18584,N_18544);
and U19298 (N_19298,N_18730,N_18692);
or U19299 (N_19299,N_18746,N_18603);
nor U19300 (N_19300,N_18875,N_18617);
and U19301 (N_19301,N_18773,N_18657);
and U19302 (N_19302,N_18580,N_18625);
xor U19303 (N_19303,N_18962,N_18886);
or U19304 (N_19304,N_18605,N_18558);
nor U19305 (N_19305,N_18663,N_18921);
and U19306 (N_19306,N_18725,N_18524);
nor U19307 (N_19307,N_18547,N_18632);
nand U19308 (N_19308,N_18501,N_18582);
or U19309 (N_19309,N_18873,N_18827);
nand U19310 (N_19310,N_18829,N_18931);
nand U19311 (N_19311,N_18732,N_18744);
nand U19312 (N_19312,N_18636,N_18663);
and U19313 (N_19313,N_18599,N_18794);
and U19314 (N_19314,N_18799,N_18860);
or U19315 (N_19315,N_18780,N_18881);
nor U19316 (N_19316,N_18870,N_18993);
and U19317 (N_19317,N_18772,N_18747);
nor U19318 (N_19318,N_18659,N_18599);
nand U19319 (N_19319,N_18603,N_18840);
nor U19320 (N_19320,N_18806,N_18848);
and U19321 (N_19321,N_18843,N_18522);
and U19322 (N_19322,N_18774,N_18763);
xor U19323 (N_19323,N_18803,N_18835);
nand U19324 (N_19324,N_18717,N_18787);
or U19325 (N_19325,N_18753,N_18643);
or U19326 (N_19326,N_18815,N_18827);
nand U19327 (N_19327,N_18711,N_18675);
nand U19328 (N_19328,N_18833,N_18582);
or U19329 (N_19329,N_18859,N_18684);
nand U19330 (N_19330,N_18575,N_18885);
xnor U19331 (N_19331,N_18886,N_18781);
xnor U19332 (N_19332,N_18789,N_18665);
nand U19333 (N_19333,N_18659,N_18686);
nand U19334 (N_19334,N_18993,N_18673);
nand U19335 (N_19335,N_18847,N_18511);
xnor U19336 (N_19336,N_18986,N_18643);
or U19337 (N_19337,N_18888,N_18622);
nor U19338 (N_19338,N_18670,N_18939);
xnor U19339 (N_19339,N_18947,N_18877);
xnor U19340 (N_19340,N_18982,N_18766);
and U19341 (N_19341,N_18749,N_18627);
nand U19342 (N_19342,N_18515,N_18838);
nand U19343 (N_19343,N_18961,N_18539);
xnor U19344 (N_19344,N_18805,N_18568);
xnor U19345 (N_19345,N_18757,N_18754);
nand U19346 (N_19346,N_18741,N_18929);
and U19347 (N_19347,N_18986,N_18696);
and U19348 (N_19348,N_18584,N_18680);
and U19349 (N_19349,N_18926,N_18637);
or U19350 (N_19350,N_18947,N_18556);
and U19351 (N_19351,N_18985,N_18752);
xnor U19352 (N_19352,N_18663,N_18689);
xor U19353 (N_19353,N_18615,N_18864);
and U19354 (N_19354,N_18772,N_18537);
and U19355 (N_19355,N_18787,N_18987);
or U19356 (N_19356,N_18502,N_18903);
nand U19357 (N_19357,N_18636,N_18915);
or U19358 (N_19358,N_18905,N_18915);
nor U19359 (N_19359,N_18665,N_18991);
nor U19360 (N_19360,N_18584,N_18781);
xor U19361 (N_19361,N_18989,N_18740);
and U19362 (N_19362,N_18963,N_18613);
and U19363 (N_19363,N_18749,N_18800);
nor U19364 (N_19364,N_18719,N_18986);
nand U19365 (N_19365,N_18857,N_18959);
nand U19366 (N_19366,N_18522,N_18823);
nand U19367 (N_19367,N_18688,N_18522);
and U19368 (N_19368,N_18963,N_18885);
or U19369 (N_19369,N_18997,N_18567);
nor U19370 (N_19370,N_18947,N_18832);
nor U19371 (N_19371,N_18737,N_18560);
xor U19372 (N_19372,N_18571,N_18689);
nor U19373 (N_19373,N_18888,N_18878);
and U19374 (N_19374,N_18712,N_18944);
nor U19375 (N_19375,N_18842,N_18535);
nor U19376 (N_19376,N_18755,N_18515);
nor U19377 (N_19377,N_18619,N_18794);
or U19378 (N_19378,N_18852,N_18597);
xnor U19379 (N_19379,N_18658,N_18724);
nor U19380 (N_19380,N_18746,N_18783);
nand U19381 (N_19381,N_18758,N_18570);
nor U19382 (N_19382,N_18784,N_18759);
or U19383 (N_19383,N_18692,N_18541);
and U19384 (N_19384,N_18569,N_18944);
or U19385 (N_19385,N_18815,N_18609);
nand U19386 (N_19386,N_18672,N_18945);
nor U19387 (N_19387,N_18818,N_18959);
or U19388 (N_19388,N_18707,N_18878);
and U19389 (N_19389,N_18854,N_18802);
nor U19390 (N_19390,N_18746,N_18979);
xor U19391 (N_19391,N_18783,N_18937);
nor U19392 (N_19392,N_18504,N_18512);
nor U19393 (N_19393,N_18918,N_18625);
nor U19394 (N_19394,N_18991,N_18664);
xor U19395 (N_19395,N_18841,N_18513);
nand U19396 (N_19396,N_18896,N_18515);
or U19397 (N_19397,N_18606,N_18514);
xnor U19398 (N_19398,N_18801,N_18724);
xnor U19399 (N_19399,N_18861,N_18869);
and U19400 (N_19400,N_18914,N_18541);
xnor U19401 (N_19401,N_18584,N_18909);
nand U19402 (N_19402,N_18792,N_18544);
or U19403 (N_19403,N_18690,N_18744);
xor U19404 (N_19404,N_18676,N_18555);
or U19405 (N_19405,N_18845,N_18688);
nand U19406 (N_19406,N_18881,N_18964);
and U19407 (N_19407,N_18780,N_18684);
nand U19408 (N_19408,N_18577,N_18783);
and U19409 (N_19409,N_18922,N_18890);
nand U19410 (N_19410,N_18768,N_18782);
and U19411 (N_19411,N_18504,N_18641);
xnor U19412 (N_19412,N_18748,N_18815);
nand U19413 (N_19413,N_18596,N_18922);
xnor U19414 (N_19414,N_18574,N_18795);
or U19415 (N_19415,N_18764,N_18780);
and U19416 (N_19416,N_18832,N_18872);
and U19417 (N_19417,N_18987,N_18877);
nand U19418 (N_19418,N_18955,N_18820);
and U19419 (N_19419,N_18652,N_18654);
nor U19420 (N_19420,N_18733,N_18595);
nor U19421 (N_19421,N_18842,N_18952);
and U19422 (N_19422,N_18949,N_18913);
nor U19423 (N_19423,N_18545,N_18781);
nand U19424 (N_19424,N_18570,N_18939);
and U19425 (N_19425,N_18773,N_18633);
or U19426 (N_19426,N_18921,N_18870);
xor U19427 (N_19427,N_18684,N_18644);
and U19428 (N_19428,N_18844,N_18654);
nor U19429 (N_19429,N_18578,N_18714);
nor U19430 (N_19430,N_18819,N_18697);
nor U19431 (N_19431,N_18889,N_18650);
nand U19432 (N_19432,N_18669,N_18683);
nand U19433 (N_19433,N_18781,N_18951);
and U19434 (N_19434,N_18621,N_18828);
or U19435 (N_19435,N_18748,N_18871);
or U19436 (N_19436,N_18543,N_18748);
or U19437 (N_19437,N_18579,N_18777);
xnor U19438 (N_19438,N_18843,N_18688);
nand U19439 (N_19439,N_18764,N_18749);
xnor U19440 (N_19440,N_18861,N_18739);
or U19441 (N_19441,N_18650,N_18538);
and U19442 (N_19442,N_18918,N_18764);
xor U19443 (N_19443,N_18670,N_18841);
nor U19444 (N_19444,N_18851,N_18557);
xor U19445 (N_19445,N_18529,N_18964);
and U19446 (N_19446,N_18869,N_18778);
nand U19447 (N_19447,N_18960,N_18686);
nand U19448 (N_19448,N_18974,N_18704);
nand U19449 (N_19449,N_18919,N_18678);
xnor U19450 (N_19450,N_18662,N_18638);
nand U19451 (N_19451,N_18574,N_18945);
nand U19452 (N_19452,N_18621,N_18894);
and U19453 (N_19453,N_18866,N_18885);
or U19454 (N_19454,N_18608,N_18748);
xor U19455 (N_19455,N_18908,N_18692);
and U19456 (N_19456,N_18852,N_18948);
and U19457 (N_19457,N_18630,N_18667);
or U19458 (N_19458,N_18611,N_18572);
or U19459 (N_19459,N_18819,N_18894);
and U19460 (N_19460,N_18741,N_18677);
and U19461 (N_19461,N_18554,N_18914);
xor U19462 (N_19462,N_18537,N_18588);
nor U19463 (N_19463,N_18579,N_18605);
and U19464 (N_19464,N_18871,N_18923);
xnor U19465 (N_19465,N_18547,N_18945);
nor U19466 (N_19466,N_18879,N_18599);
xnor U19467 (N_19467,N_18679,N_18881);
and U19468 (N_19468,N_18839,N_18638);
nand U19469 (N_19469,N_18543,N_18753);
nor U19470 (N_19470,N_18516,N_18616);
nor U19471 (N_19471,N_18568,N_18597);
and U19472 (N_19472,N_18883,N_18510);
nand U19473 (N_19473,N_18885,N_18879);
or U19474 (N_19474,N_18803,N_18758);
and U19475 (N_19475,N_18793,N_18918);
and U19476 (N_19476,N_18869,N_18528);
or U19477 (N_19477,N_18978,N_18910);
xor U19478 (N_19478,N_18868,N_18703);
nand U19479 (N_19479,N_18589,N_18740);
nor U19480 (N_19480,N_18854,N_18889);
nand U19481 (N_19481,N_18504,N_18721);
nand U19482 (N_19482,N_18537,N_18875);
nor U19483 (N_19483,N_18667,N_18573);
or U19484 (N_19484,N_18616,N_18621);
nand U19485 (N_19485,N_18984,N_18985);
nand U19486 (N_19486,N_18626,N_18836);
and U19487 (N_19487,N_18881,N_18713);
nand U19488 (N_19488,N_18672,N_18713);
nand U19489 (N_19489,N_18667,N_18856);
and U19490 (N_19490,N_18766,N_18730);
nand U19491 (N_19491,N_18858,N_18856);
nand U19492 (N_19492,N_18967,N_18964);
nand U19493 (N_19493,N_18542,N_18986);
and U19494 (N_19494,N_18619,N_18902);
and U19495 (N_19495,N_18560,N_18768);
or U19496 (N_19496,N_18744,N_18997);
and U19497 (N_19497,N_18783,N_18657);
or U19498 (N_19498,N_18563,N_18900);
nor U19499 (N_19499,N_18941,N_18944);
or U19500 (N_19500,N_19041,N_19390);
nor U19501 (N_19501,N_19208,N_19031);
nor U19502 (N_19502,N_19488,N_19355);
xor U19503 (N_19503,N_19048,N_19085);
nand U19504 (N_19504,N_19172,N_19144);
nor U19505 (N_19505,N_19203,N_19409);
nor U19506 (N_19506,N_19387,N_19275);
nor U19507 (N_19507,N_19450,N_19246);
and U19508 (N_19508,N_19110,N_19054);
nor U19509 (N_19509,N_19474,N_19078);
or U19510 (N_19510,N_19029,N_19370);
nand U19511 (N_19511,N_19030,N_19118);
and U19512 (N_19512,N_19006,N_19353);
nor U19513 (N_19513,N_19490,N_19362);
or U19514 (N_19514,N_19478,N_19371);
nand U19515 (N_19515,N_19004,N_19157);
xor U19516 (N_19516,N_19057,N_19485);
nor U19517 (N_19517,N_19161,N_19454);
nor U19518 (N_19518,N_19201,N_19402);
and U19519 (N_19519,N_19050,N_19411);
or U19520 (N_19520,N_19467,N_19090);
and U19521 (N_19521,N_19284,N_19372);
and U19522 (N_19522,N_19245,N_19329);
nor U19523 (N_19523,N_19391,N_19218);
xor U19524 (N_19524,N_19084,N_19468);
and U19525 (N_19525,N_19385,N_19496);
xor U19526 (N_19526,N_19212,N_19102);
nand U19527 (N_19527,N_19347,N_19170);
nand U19528 (N_19528,N_19338,N_19486);
nor U19529 (N_19529,N_19357,N_19290);
xnor U19530 (N_19530,N_19247,N_19120);
and U19531 (N_19531,N_19470,N_19099);
nand U19532 (N_19532,N_19452,N_19018);
and U19533 (N_19533,N_19475,N_19015);
or U19534 (N_19534,N_19428,N_19294);
xnor U19535 (N_19535,N_19077,N_19440);
nand U19536 (N_19536,N_19130,N_19379);
or U19537 (N_19537,N_19472,N_19262);
xnor U19538 (N_19538,N_19274,N_19152);
and U19539 (N_19539,N_19021,N_19455);
xor U19540 (N_19540,N_19369,N_19378);
xor U19541 (N_19541,N_19185,N_19192);
and U19542 (N_19542,N_19451,N_19066);
or U19543 (N_19543,N_19356,N_19125);
or U19544 (N_19544,N_19222,N_19105);
or U19545 (N_19545,N_19361,N_19182);
xor U19546 (N_19546,N_19477,N_19173);
nor U19547 (N_19547,N_19424,N_19331);
or U19548 (N_19548,N_19304,N_19292);
or U19549 (N_19549,N_19232,N_19237);
xnor U19550 (N_19550,N_19079,N_19163);
or U19551 (N_19551,N_19059,N_19098);
nor U19552 (N_19552,N_19473,N_19028);
nor U19553 (N_19553,N_19335,N_19121);
nor U19554 (N_19554,N_19134,N_19049);
nand U19555 (N_19555,N_19180,N_19449);
or U19556 (N_19556,N_19136,N_19492);
nor U19557 (N_19557,N_19311,N_19219);
and U19558 (N_19558,N_19147,N_19471);
nand U19559 (N_19559,N_19312,N_19149);
nor U19560 (N_19560,N_19154,N_19322);
or U19561 (N_19561,N_19314,N_19352);
nand U19562 (N_19562,N_19268,N_19253);
xor U19563 (N_19563,N_19422,N_19122);
nor U19564 (N_19564,N_19297,N_19325);
nor U19565 (N_19565,N_19377,N_19350);
nand U19566 (N_19566,N_19256,N_19324);
nand U19567 (N_19567,N_19403,N_19309);
or U19568 (N_19568,N_19106,N_19288);
nor U19569 (N_19569,N_19072,N_19466);
and U19570 (N_19570,N_19263,N_19448);
xnor U19571 (N_19571,N_19407,N_19260);
nor U19572 (N_19572,N_19364,N_19044);
nor U19573 (N_19573,N_19367,N_19039);
nor U19574 (N_19574,N_19053,N_19373);
or U19575 (N_19575,N_19123,N_19483);
or U19576 (N_19576,N_19231,N_19287);
nand U19577 (N_19577,N_19129,N_19255);
xor U19578 (N_19578,N_19220,N_19051);
nand U19579 (N_19579,N_19209,N_19417);
nor U19580 (N_19580,N_19458,N_19023);
and U19581 (N_19581,N_19183,N_19086);
and U19582 (N_19582,N_19376,N_19103);
nor U19583 (N_19583,N_19150,N_19139);
xor U19584 (N_19584,N_19360,N_19349);
xnor U19585 (N_19585,N_19251,N_19065);
or U19586 (N_19586,N_19404,N_19459);
and U19587 (N_19587,N_19092,N_19064);
and U19588 (N_19588,N_19261,N_19199);
or U19589 (N_19589,N_19258,N_19341);
nor U19590 (N_19590,N_19318,N_19439);
nor U19591 (N_19591,N_19188,N_19215);
or U19592 (N_19592,N_19076,N_19233);
xor U19593 (N_19593,N_19224,N_19271);
and U19594 (N_19594,N_19043,N_19151);
xor U19595 (N_19595,N_19040,N_19011);
nor U19596 (N_19596,N_19302,N_19249);
or U19597 (N_19597,N_19229,N_19205);
nor U19598 (N_19598,N_19116,N_19239);
or U19599 (N_19599,N_19425,N_19264);
xor U19600 (N_19600,N_19259,N_19083);
nor U19601 (N_19601,N_19197,N_19286);
xor U19602 (N_19602,N_19137,N_19115);
or U19603 (N_19603,N_19438,N_19382);
or U19604 (N_19604,N_19421,N_19346);
or U19605 (N_19605,N_19034,N_19181);
nor U19606 (N_19606,N_19025,N_19305);
xor U19607 (N_19607,N_19445,N_19423);
xor U19608 (N_19608,N_19000,N_19447);
or U19609 (N_19609,N_19081,N_19014);
nand U19610 (N_19610,N_19374,N_19111);
nand U19611 (N_19611,N_19155,N_19291);
xnor U19612 (N_19612,N_19293,N_19345);
nand U19613 (N_19613,N_19190,N_19316);
nor U19614 (N_19614,N_19026,N_19446);
xnor U19615 (N_19615,N_19127,N_19300);
nand U19616 (N_19616,N_19009,N_19141);
xor U19617 (N_19617,N_19340,N_19088);
or U19618 (N_19618,N_19126,N_19204);
or U19619 (N_19619,N_19265,N_19442);
nand U19620 (N_19620,N_19375,N_19207);
xor U19621 (N_19621,N_19179,N_19279);
nand U19622 (N_19622,N_19413,N_19463);
xor U19623 (N_19623,N_19153,N_19412);
and U19624 (N_19624,N_19384,N_19461);
and U19625 (N_19625,N_19113,N_19241);
nand U19626 (N_19626,N_19061,N_19317);
and U19627 (N_19627,N_19401,N_19348);
xnor U19628 (N_19628,N_19499,N_19080);
xnor U19629 (N_19629,N_19491,N_19476);
nor U19630 (N_19630,N_19295,N_19187);
or U19631 (N_19631,N_19368,N_19269);
and U19632 (N_19632,N_19160,N_19315);
nand U19633 (N_19633,N_19069,N_19097);
nor U19634 (N_19634,N_19132,N_19138);
nand U19635 (N_19635,N_19252,N_19464);
xnor U19636 (N_19636,N_19244,N_19414);
and U19637 (N_19637,N_19223,N_19082);
xnor U19638 (N_19638,N_19013,N_19298);
or U19639 (N_19639,N_19142,N_19308);
xnor U19640 (N_19640,N_19381,N_19321);
xor U19641 (N_19641,N_19481,N_19266);
nor U19642 (N_19642,N_19363,N_19052);
nand U19643 (N_19643,N_19482,N_19008);
or U19644 (N_19644,N_19426,N_19395);
and U19645 (N_19645,N_19332,N_19389);
or U19646 (N_19646,N_19135,N_19174);
nand U19647 (N_19647,N_19193,N_19035);
xor U19648 (N_19648,N_19437,N_19457);
xnor U19649 (N_19649,N_19243,N_19480);
nand U19650 (N_19650,N_19068,N_19393);
xnor U19651 (N_19651,N_19012,N_19280);
or U19652 (N_19652,N_19211,N_19055);
nand U19653 (N_19653,N_19184,N_19328);
or U19654 (N_19654,N_19435,N_19186);
and U19655 (N_19655,N_19443,N_19177);
and U19656 (N_19656,N_19162,N_19380);
nor U19657 (N_19657,N_19001,N_19165);
nand U19658 (N_19658,N_19326,N_19104);
or U19659 (N_19659,N_19276,N_19176);
or U19660 (N_19660,N_19415,N_19418);
or U19661 (N_19661,N_19221,N_19063);
xnor U19662 (N_19662,N_19416,N_19303);
and U19663 (N_19663,N_19198,N_19108);
nand U19664 (N_19664,N_19285,N_19432);
and U19665 (N_19665,N_19479,N_19330);
nand U19666 (N_19666,N_19107,N_19214);
nor U19667 (N_19667,N_19436,N_19230);
nand U19668 (N_19668,N_19433,N_19250);
xnor U19669 (N_19669,N_19489,N_19272);
and U19670 (N_19670,N_19046,N_19128);
nor U19671 (N_19671,N_19366,N_19327);
nor U19672 (N_19672,N_19140,N_19234);
nand U19673 (N_19673,N_19019,N_19278);
or U19674 (N_19674,N_19020,N_19202);
or U19675 (N_19675,N_19277,N_19156);
nor U19676 (N_19676,N_19047,N_19392);
nand U19677 (N_19677,N_19112,N_19343);
xnor U19678 (N_19678,N_19096,N_19216);
and U19679 (N_19679,N_19313,N_19166);
or U19680 (N_19680,N_19117,N_19164);
and U19681 (N_19681,N_19095,N_19281);
nor U19682 (N_19682,N_19310,N_19073);
and U19683 (N_19683,N_19235,N_19124);
or U19684 (N_19684,N_19351,N_19217);
nor U19685 (N_19685,N_19242,N_19060);
and U19686 (N_19686,N_19408,N_19419);
or U19687 (N_19687,N_19024,N_19226);
and U19688 (N_19688,N_19365,N_19400);
and U19689 (N_19689,N_19087,N_19159);
xnor U19690 (N_19690,N_19194,N_19210);
xnor U19691 (N_19691,N_19067,N_19131);
and U19692 (N_19692,N_19460,N_19089);
nor U19693 (N_19693,N_19213,N_19167);
nand U19694 (N_19694,N_19075,N_19236);
xnor U19695 (N_19695,N_19036,N_19495);
nand U19696 (N_19696,N_19420,N_19484);
xnor U19697 (N_19697,N_19133,N_19058);
xnor U19698 (N_19698,N_19022,N_19070);
and U19699 (N_19699,N_19100,N_19228);
nand U19700 (N_19700,N_19359,N_19227);
nand U19701 (N_19701,N_19248,N_19431);
nor U19702 (N_19702,N_19168,N_19270);
and U19703 (N_19703,N_19320,N_19358);
nand U19704 (N_19704,N_19319,N_19143);
nor U19705 (N_19705,N_19429,N_19394);
xor U19706 (N_19706,N_19169,N_19101);
or U19707 (N_19707,N_19396,N_19042);
or U19708 (N_19708,N_19397,N_19033);
and U19709 (N_19709,N_19487,N_19427);
nor U19710 (N_19710,N_19497,N_19091);
nor U19711 (N_19711,N_19002,N_19453);
nor U19712 (N_19712,N_19037,N_19145);
nand U19713 (N_19713,N_19109,N_19225);
or U19714 (N_19714,N_19257,N_19462);
nor U19715 (N_19715,N_19189,N_19158);
nand U19716 (N_19716,N_19398,N_19175);
nor U19717 (N_19717,N_19191,N_19196);
xnor U19718 (N_19718,N_19405,N_19032);
nor U19719 (N_19719,N_19456,N_19074);
xnor U19720 (N_19720,N_19114,N_19017);
nor U19721 (N_19721,N_19289,N_19296);
and U19722 (N_19722,N_19056,N_19465);
or U19723 (N_19723,N_19273,N_19494);
and U19724 (N_19724,N_19430,N_19469);
and U19725 (N_19725,N_19386,N_19045);
xnor U19726 (N_19726,N_19383,N_19240);
nor U19727 (N_19727,N_19333,N_19007);
and U19728 (N_19728,N_19301,N_19342);
xnor U19729 (N_19729,N_19306,N_19119);
xor U19730 (N_19730,N_19282,N_19038);
nor U19731 (N_19731,N_19094,N_19254);
xor U19732 (N_19732,N_19399,N_19005);
nor U19733 (N_19733,N_19406,N_19323);
xor U19734 (N_19734,N_19334,N_19238);
nand U19735 (N_19735,N_19434,N_19010);
xnor U19736 (N_19736,N_19093,N_19206);
and U19737 (N_19737,N_19354,N_19003);
xor U19738 (N_19738,N_19062,N_19200);
and U19739 (N_19739,N_19171,N_19146);
nand U19740 (N_19740,N_19337,N_19444);
nor U19741 (N_19741,N_19283,N_19336);
nand U19742 (N_19742,N_19498,N_19071);
and U19743 (N_19743,N_19148,N_19307);
or U19744 (N_19744,N_19267,N_19178);
or U19745 (N_19745,N_19410,N_19195);
nor U19746 (N_19746,N_19299,N_19441);
nor U19747 (N_19747,N_19027,N_19339);
xnor U19748 (N_19748,N_19388,N_19016);
nor U19749 (N_19749,N_19344,N_19493);
nor U19750 (N_19750,N_19423,N_19400);
nand U19751 (N_19751,N_19239,N_19393);
or U19752 (N_19752,N_19499,N_19497);
or U19753 (N_19753,N_19158,N_19092);
nand U19754 (N_19754,N_19457,N_19166);
nor U19755 (N_19755,N_19234,N_19253);
or U19756 (N_19756,N_19026,N_19321);
nand U19757 (N_19757,N_19051,N_19486);
or U19758 (N_19758,N_19316,N_19416);
or U19759 (N_19759,N_19267,N_19207);
nand U19760 (N_19760,N_19418,N_19444);
and U19761 (N_19761,N_19076,N_19199);
xnor U19762 (N_19762,N_19091,N_19324);
xor U19763 (N_19763,N_19385,N_19280);
xor U19764 (N_19764,N_19325,N_19428);
nand U19765 (N_19765,N_19384,N_19322);
or U19766 (N_19766,N_19167,N_19217);
nand U19767 (N_19767,N_19075,N_19290);
nor U19768 (N_19768,N_19302,N_19420);
nor U19769 (N_19769,N_19201,N_19213);
xnor U19770 (N_19770,N_19244,N_19365);
and U19771 (N_19771,N_19102,N_19431);
xor U19772 (N_19772,N_19110,N_19394);
nor U19773 (N_19773,N_19252,N_19001);
xor U19774 (N_19774,N_19331,N_19366);
xor U19775 (N_19775,N_19028,N_19411);
or U19776 (N_19776,N_19061,N_19338);
nor U19777 (N_19777,N_19281,N_19370);
or U19778 (N_19778,N_19055,N_19422);
nor U19779 (N_19779,N_19065,N_19302);
xor U19780 (N_19780,N_19470,N_19272);
nand U19781 (N_19781,N_19205,N_19476);
and U19782 (N_19782,N_19085,N_19126);
and U19783 (N_19783,N_19444,N_19199);
nand U19784 (N_19784,N_19481,N_19066);
xor U19785 (N_19785,N_19172,N_19412);
nor U19786 (N_19786,N_19424,N_19443);
nand U19787 (N_19787,N_19237,N_19396);
and U19788 (N_19788,N_19146,N_19310);
nor U19789 (N_19789,N_19433,N_19016);
xor U19790 (N_19790,N_19196,N_19062);
and U19791 (N_19791,N_19035,N_19381);
xnor U19792 (N_19792,N_19162,N_19465);
nand U19793 (N_19793,N_19057,N_19479);
or U19794 (N_19794,N_19353,N_19072);
xnor U19795 (N_19795,N_19306,N_19261);
or U19796 (N_19796,N_19331,N_19170);
xor U19797 (N_19797,N_19393,N_19210);
xor U19798 (N_19798,N_19118,N_19296);
nand U19799 (N_19799,N_19248,N_19163);
and U19800 (N_19800,N_19197,N_19159);
xnor U19801 (N_19801,N_19333,N_19252);
and U19802 (N_19802,N_19083,N_19466);
nand U19803 (N_19803,N_19172,N_19394);
or U19804 (N_19804,N_19389,N_19168);
or U19805 (N_19805,N_19145,N_19286);
xnor U19806 (N_19806,N_19089,N_19358);
xnor U19807 (N_19807,N_19186,N_19383);
and U19808 (N_19808,N_19032,N_19230);
or U19809 (N_19809,N_19185,N_19382);
nor U19810 (N_19810,N_19399,N_19136);
nor U19811 (N_19811,N_19472,N_19352);
nand U19812 (N_19812,N_19156,N_19493);
nand U19813 (N_19813,N_19081,N_19349);
xor U19814 (N_19814,N_19327,N_19140);
xor U19815 (N_19815,N_19386,N_19154);
nor U19816 (N_19816,N_19396,N_19239);
xor U19817 (N_19817,N_19012,N_19018);
xnor U19818 (N_19818,N_19169,N_19032);
nor U19819 (N_19819,N_19043,N_19352);
or U19820 (N_19820,N_19133,N_19310);
xor U19821 (N_19821,N_19003,N_19402);
and U19822 (N_19822,N_19109,N_19179);
nand U19823 (N_19823,N_19016,N_19202);
nor U19824 (N_19824,N_19310,N_19170);
and U19825 (N_19825,N_19051,N_19353);
xor U19826 (N_19826,N_19107,N_19441);
or U19827 (N_19827,N_19257,N_19464);
and U19828 (N_19828,N_19101,N_19025);
and U19829 (N_19829,N_19198,N_19012);
and U19830 (N_19830,N_19144,N_19432);
nor U19831 (N_19831,N_19298,N_19315);
and U19832 (N_19832,N_19104,N_19236);
or U19833 (N_19833,N_19314,N_19455);
nor U19834 (N_19834,N_19457,N_19176);
or U19835 (N_19835,N_19298,N_19245);
xnor U19836 (N_19836,N_19026,N_19372);
or U19837 (N_19837,N_19071,N_19092);
nor U19838 (N_19838,N_19475,N_19140);
nor U19839 (N_19839,N_19423,N_19073);
and U19840 (N_19840,N_19333,N_19445);
xor U19841 (N_19841,N_19321,N_19406);
and U19842 (N_19842,N_19091,N_19137);
nor U19843 (N_19843,N_19044,N_19219);
or U19844 (N_19844,N_19383,N_19488);
and U19845 (N_19845,N_19301,N_19295);
xor U19846 (N_19846,N_19485,N_19390);
nand U19847 (N_19847,N_19382,N_19316);
nand U19848 (N_19848,N_19035,N_19461);
nor U19849 (N_19849,N_19088,N_19392);
xor U19850 (N_19850,N_19406,N_19175);
nand U19851 (N_19851,N_19105,N_19089);
nand U19852 (N_19852,N_19083,N_19058);
xor U19853 (N_19853,N_19047,N_19369);
nand U19854 (N_19854,N_19293,N_19474);
xor U19855 (N_19855,N_19226,N_19082);
nand U19856 (N_19856,N_19240,N_19093);
xnor U19857 (N_19857,N_19224,N_19396);
xor U19858 (N_19858,N_19354,N_19147);
or U19859 (N_19859,N_19449,N_19027);
nand U19860 (N_19860,N_19297,N_19387);
or U19861 (N_19861,N_19139,N_19213);
nor U19862 (N_19862,N_19000,N_19418);
xnor U19863 (N_19863,N_19012,N_19347);
and U19864 (N_19864,N_19168,N_19152);
nor U19865 (N_19865,N_19158,N_19098);
nand U19866 (N_19866,N_19454,N_19170);
nor U19867 (N_19867,N_19306,N_19404);
nor U19868 (N_19868,N_19364,N_19293);
or U19869 (N_19869,N_19444,N_19014);
nor U19870 (N_19870,N_19004,N_19294);
nor U19871 (N_19871,N_19421,N_19475);
xor U19872 (N_19872,N_19213,N_19056);
nand U19873 (N_19873,N_19393,N_19423);
or U19874 (N_19874,N_19115,N_19367);
nand U19875 (N_19875,N_19472,N_19451);
and U19876 (N_19876,N_19278,N_19217);
or U19877 (N_19877,N_19373,N_19485);
and U19878 (N_19878,N_19041,N_19043);
and U19879 (N_19879,N_19277,N_19173);
nand U19880 (N_19880,N_19484,N_19072);
and U19881 (N_19881,N_19261,N_19397);
and U19882 (N_19882,N_19156,N_19475);
nand U19883 (N_19883,N_19475,N_19294);
nand U19884 (N_19884,N_19391,N_19193);
nand U19885 (N_19885,N_19206,N_19215);
or U19886 (N_19886,N_19279,N_19441);
nor U19887 (N_19887,N_19459,N_19243);
nand U19888 (N_19888,N_19477,N_19163);
nor U19889 (N_19889,N_19006,N_19214);
nor U19890 (N_19890,N_19034,N_19321);
nor U19891 (N_19891,N_19388,N_19183);
nand U19892 (N_19892,N_19000,N_19098);
nor U19893 (N_19893,N_19420,N_19405);
nand U19894 (N_19894,N_19007,N_19039);
nand U19895 (N_19895,N_19304,N_19414);
and U19896 (N_19896,N_19048,N_19137);
xnor U19897 (N_19897,N_19390,N_19384);
or U19898 (N_19898,N_19125,N_19013);
nand U19899 (N_19899,N_19032,N_19261);
nor U19900 (N_19900,N_19247,N_19472);
xor U19901 (N_19901,N_19345,N_19489);
nand U19902 (N_19902,N_19251,N_19019);
or U19903 (N_19903,N_19480,N_19054);
and U19904 (N_19904,N_19137,N_19398);
or U19905 (N_19905,N_19034,N_19380);
or U19906 (N_19906,N_19043,N_19204);
or U19907 (N_19907,N_19113,N_19445);
xor U19908 (N_19908,N_19375,N_19393);
nand U19909 (N_19909,N_19215,N_19373);
xor U19910 (N_19910,N_19141,N_19284);
nand U19911 (N_19911,N_19279,N_19296);
nor U19912 (N_19912,N_19181,N_19491);
or U19913 (N_19913,N_19338,N_19258);
or U19914 (N_19914,N_19316,N_19099);
or U19915 (N_19915,N_19229,N_19253);
nor U19916 (N_19916,N_19489,N_19387);
nand U19917 (N_19917,N_19131,N_19226);
nand U19918 (N_19918,N_19195,N_19238);
and U19919 (N_19919,N_19155,N_19170);
xor U19920 (N_19920,N_19065,N_19217);
nand U19921 (N_19921,N_19013,N_19264);
or U19922 (N_19922,N_19331,N_19041);
nand U19923 (N_19923,N_19040,N_19053);
nor U19924 (N_19924,N_19267,N_19285);
nor U19925 (N_19925,N_19101,N_19273);
or U19926 (N_19926,N_19464,N_19125);
xnor U19927 (N_19927,N_19211,N_19489);
and U19928 (N_19928,N_19152,N_19313);
nand U19929 (N_19929,N_19407,N_19303);
or U19930 (N_19930,N_19480,N_19321);
or U19931 (N_19931,N_19189,N_19279);
xnor U19932 (N_19932,N_19484,N_19461);
nand U19933 (N_19933,N_19050,N_19314);
nor U19934 (N_19934,N_19497,N_19272);
and U19935 (N_19935,N_19298,N_19080);
or U19936 (N_19936,N_19319,N_19346);
xor U19937 (N_19937,N_19263,N_19226);
nor U19938 (N_19938,N_19367,N_19393);
nand U19939 (N_19939,N_19377,N_19462);
and U19940 (N_19940,N_19032,N_19147);
nand U19941 (N_19941,N_19497,N_19356);
nor U19942 (N_19942,N_19258,N_19159);
xor U19943 (N_19943,N_19454,N_19480);
or U19944 (N_19944,N_19169,N_19281);
xnor U19945 (N_19945,N_19492,N_19395);
nand U19946 (N_19946,N_19311,N_19210);
or U19947 (N_19947,N_19275,N_19173);
and U19948 (N_19948,N_19344,N_19006);
or U19949 (N_19949,N_19148,N_19273);
and U19950 (N_19950,N_19224,N_19244);
or U19951 (N_19951,N_19219,N_19383);
nand U19952 (N_19952,N_19254,N_19294);
xor U19953 (N_19953,N_19260,N_19138);
nand U19954 (N_19954,N_19307,N_19044);
nor U19955 (N_19955,N_19478,N_19130);
and U19956 (N_19956,N_19494,N_19465);
nor U19957 (N_19957,N_19144,N_19000);
and U19958 (N_19958,N_19241,N_19345);
xnor U19959 (N_19959,N_19352,N_19213);
and U19960 (N_19960,N_19373,N_19495);
nand U19961 (N_19961,N_19008,N_19144);
and U19962 (N_19962,N_19349,N_19094);
or U19963 (N_19963,N_19219,N_19341);
nor U19964 (N_19964,N_19329,N_19244);
xnor U19965 (N_19965,N_19489,N_19349);
and U19966 (N_19966,N_19216,N_19393);
and U19967 (N_19967,N_19069,N_19410);
and U19968 (N_19968,N_19216,N_19429);
xnor U19969 (N_19969,N_19462,N_19466);
nand U19970 (N_19970,N_19160,N_19464);
and U19971 (N_19971,N_19251,N_19240);
nand U19972 (N_19972,N_19000,N_19161);
nand U19973 (N_19973,N_19411,N_19314);
nand U19974 (N_19974,N_19185,N_19062);
and U19975 (N_19975,N_19243,N_19112);
and U19976 (N_19976,N_19369,N_19226);
nand U19977 (N_19977,N_19272,N_19132);
nand U19978 (N_19978,N_19082,N_19047);
nor U19979 (N_19979,N_19485,N_19446);
nand U19980 (N_19980,N_19171,N_19246);
nand U19981 (N_19981,N_19276,N_19005);
nor U19982 (N_19982,N_19092,N_19475);
and U19983 (N_19983,N_19197,N_19470);
nand U19984 (N_19984,N_19418,N_19023);
nor U19985 (N_19985,N_19330,N_19260);
xor U19986 (N_19986,N_19470,N_19004);
nand U19987 (N_19987,N_19059,N_19021);
or U19988 (N_19988,N_19474,N_19276);
nand U19989 (N_19989,N_19314,N_19253);
or U19990 (N_19990,N_19309,N_19393);
or U19991 (N_19991,N_19478,N_19172);
nand U19992 (N_19992,N_19267,N_19433);
xnor U19993 (N_19993,N_19072,N_19240);
and U19994 (N_19994,N_19370,N_19380);
nand U19995 (N_19995,N_19484,N_19404);
and U19996 (N_19996,N_19327,N_19386);
xnor U19997 (N_19997,N_19109,N_19449);
or U19998 (N_19998,N_19388,N_19417);
xor U19999 (N_19999,N_19042,N_19426);
and U20000 (N_20000,N_19938,N_19501);
nor U20001 (N_20001,N_19572,N_19964);
nand U20002 (N_20002,N_19549,N_19635);
nand U20003 (N_20003,N_19646,N_19943);
xor U20004 (N_20004,N_19510,N_19776);
nand U20005 (N_20005,N_19534,N_19750);
or U20006 (N_20006,N_19911,N_19888);
nor U20007 (N_20007,N_19773,N_19584);
or U20008 (N_20008,N_19931,N_19759);
xor U20009 (N_20009,N_19642,N_19804);
xnor U20010 (N_20010,N_19553,N_19955);
and U20011 (N_20011,N_19603,N_19959);
nor U20012 (N_20012,N_19504,N_19652);
xor U20013 (N_20013,N_19641,N_19640);
nand U20014 (N_20014,N_19707,N_19538);
nor U20015 (N_20015,N_19799,N_19928);
nor U20016 (N_20016,N_19583,N_19841);
or U20017 (N_20017,N_19587,N_19594);
nand U20018 (N_20018,N_19827,N_19850);
xnor U20019 (N_20019,N_19973,N_19612);
and U20020 (N_20020,N_19919,N_19765);
or U20021 (N_20021,N_19671,N_19621);
and U20022 (N_20022,N_19548,N_19654);
xnor U20023 (N_20023,N_19902,N_19697);
and U20024 (N_20024,N_19744,N_19520);
nor U20025 (N_20025,N_19904,N_19905);
nor U20026 (N_20026,N_19505,N_19556);
nand U20027 (N_20027,N_19801,N_19714);
nand U20028 (N_20028,N_19561,N_19960);
or U20029 (N_20029,N_19713,N_19916);
nor U20030 (N_20030,N_19982,N_19562);
nand U20031 (N_20031,N_19715,N_19996);
nor U20032 (N_20032,N_19558,N_19547);
or U20033 (N_20033,N_19808,N_19829);
nor U20034 (N_20034,N_19567,N_19734);
or U20035 (N_20035,N_19786,N_19596);
or U20036 (N_20036,N_19760,N_19889);
and U20037 (N_20037,N_19580,N_19880);
and U20038 (N_20038,N_19639,N_19855);
xnor U20039 (N_20039,N_19585,N_19545);
and U20040 (N_20040,N_19803,N_19978);
or U20041 (N_20041,N_19766,N_19686);
or U20042 (N_20042,N_19975,N_19897);
and U20043 (N_20043,N_19814,N_19944);
nand U20044 (N_20044,N_19624,N_19593);
nor U20045 (N_20045,N_19840,N_19632);
or U20046 (N_20046,N_19576,N_19798);
or U20047 (N_20047,N_19950,N_19650);
nand U20048 (N_20048,N_19992,N_19859);
xor U20049 (N_20049,N_19660,N_19991);
and U20050 (N_20050,N_19569,N_19873);
xnor U20051 (N_20051,N_19695,N_19664);
nand U20052 (N_20052,N_19941,N_19949);
xnor U20053 (N_20053,N_19772,N_19761);
xor U20054 (N_20054,N_19541,N_19856);
or U20055 (N_20055,N_19817,N_19825);
xnor U20056 (N_20056,N_19729,N_19974);
xor U20057 (N_20057,N_19833,N_19939);
nor U20058 (N_20058,N_19655,N_19672);
xor U20059 (N_20059,N_19812,N_19636);
or U20060 (N_20060,N_19935,N_19564);
nand U20061 (N_20061,N_19756,N_19649);
nand U20062 (N_20062,N_19927,N_19770);
and U20063 (N_20063,N_19622,N_19809);
or U20064 (N_20064,N_19507,N_19990);
xnor U20065 (N_20065,N_19847,N_19518);
and U20066 (N_20066,N_19945,N_19717);
nand U20067 (N_20067,N_19539,N_19733);
or U20068 (N_20068,N_19876,N_19883);
xnor U20069 (N_20069,N_19846,N_19780);
xor U20070 (N_20070,N_19669,N_19531);
or U20071 (N_20071,N_19681,N_19957);
or U20072 (N_20072,N_19623,N_19871);
or U20073 (N_20073,N_19923,N_19896);
nand U20074 (N_20074,N_19647,N_19824);
nand U20075 (N_20075,N_19618,N_19511);
nand U20076 (N_20076,N_19685,N_19542);
xnor U20077 (N_20077,N_19674,N_19638);
and U20078 (N_20078,N_19626,N_19863);
or U20079 (N_20079,N_19735,N_19702);
or U20080 (N_20080,N_19987,N_19683);
and U20081 (N_20081,N_19673,N_19696);
or U20082 (N_20082,N_19559,N_19966);
xor U20083 (N_20083,N_19630,N_19512);
and U20084 (N_20084,N_19728,N_19557);
xnor U20085 (N_20085,N_19693,N_19778);
nor U20086 (N_20086,N_19680,N_19924);
nand U20087 (N_20087,N_19595,N_19692);
nand U20088 (N_20088,N_19738,N_19627);
nor U20089 (N_20089,N_19901,N_19956);
or U20090 (N_20090,N_19740,N_19936);
and U20091 (N_20091,N_19907,N_19918);
nor U20092 (N_20092,N_19732,N_19894);
and U20093 (N_20093,N_19563,N_19749);
and U20094 (N_20094,N_19581,N_19684);
and U20095 (N_20095,N_19881,N_19795);
nor U20096 (N_20096,N_19926,N_19645);
and U20097 (N_20097,N_19570,N_19958);
and U20098 (N_20098,N_19983,N_19860);
and U20099 (N_20099,N_19678,N_19842);
nor U20100 (N_20100,N_19723,N_19857);
or U20101 (N_20101,N_19599,N_19746);
nand U20102 (N_20102,N_19797,N_19884);
and U20103 (N_20103,N_19724,N_19699);
and U20104 (N_20104,N_19834,N_19914);
nor U20105 (N_20105,N_19946,N_19609);
xnor U20106 (N_20106,N_19980,N_19818);
xor U20107 (N_20107,N_19767,N_19870);
xor U20108 (N_20108,N_19589,N_19568);
nand U20109 (N_20109,N_19885,N_19947);
nand U20110 (N_20110,N_19970,N_19700);
nor U20111 (N_20111,N_19868,N_19689);
nor U20112 (N_20112,N_19648,N_19525);
xnor U20113 (N_20113,N_19940,N_19743);
and U20114 (N_20114,N_19910,N_19832);
or U20115 (N_20115,N_19509,N_19688);
or U20116 (N_20116,N_19872,N_19782);
nor U20117 (N_20117,N_19785,N_19800);
and U20118 (N_20118,N_19816,N_19995);
nor U20119 (N_20119,N_19573,N_19844);
nand U20120 (N_20120,N_19830,N_19516);
nand U20121 (N_20121,N_19535,N_19532);
and U20122 (N_20122,N_19577,N_19591);
xnor U20123 (N_20123,N_19691,N_19615);
and U20124 (N_20124,N_19722,N_19537);
and U20125 (N_20125,N_19755,N_19579);
or U20126 (N_20126,N_19985,N_19783);
nand U20127 (N_20127,N_19920,N_19790);
nor U20128 (N_20128,N_19574,N_19758);
nor U20129 (N_20129,N_19874,N_19513);
and U20130 (N_20130,N_19932,N_19745);
nand U20131 (N_20131,N_19858,N_19961);
and U20132 (N_20132,N_19762,N_19952);
and U20133 (N_20133,N_19588,N_19708);
or U20134 (N_20134,N_19706,N_19592);
nand U20135 (N_20135,N_19741,N_19682);
or U20136 (N_20136,N_19566,N_19900);
xnor U20137 (N_20137,N_19668,N_19677);
nor U20138 (N_20138,N_19586,N_19796);
xnor U20139 (N_20139,N_19552,N_19862);
nor U20140 (N_20140,N_19820,N_19815);
nand U20141 (N_20141,N_19962,N_19779);
and U20142 (N_20142,N_19752,N_19698);
xnor U20143 (N_20143,N_19794,N_19965);
nand U20144 (N_20144,N_19667,N_19554);
and U20145 (N_20145,N_19725,N_19726);
and U20146 (N_20146,N_19831,N_19748);
or U20147 (N_20147,N_19533,N_19502);
nor U20148 (N_20148,N_19625,N_19967);
nor U20149 (N_20149,N_19663,N_19720);
xor U20150 (N_20150,N_19527,N_19988);
nand U20151 (N_20151,N_19895,N_19736);
nor U20152 (N_20152,N_19969,N_19613);
and U20153 (N_20153,N_19540,N_19709);
xor U20154 (N_20154,N_19948,N_19757);
nand U20155 (N_20155,N_19807,N_19875);
nor U20156 (N_20156,N_19629,N_19546);
and U20157 (N_20157,N_19751,N_19930);
and U20158 (N_20158,N_19519,N_19915);
and U20159 (N_20159,N_19971,N_19887);
xor U20160 (N_20160,N_19933,N_19620);
xor U20161 (N_20161,N_19838,N_19739);
xor U20162 (N_20162,N_19628,N_19777);
xnor U20163 (N_20163,N_19784,N_19703);
or U20164 (N_20164,N_19616,N_19694);
nor U20165 (N_20165,N_19602,N_19651);
xor U20166 (N_20166,N_19747,N_19854);
xor U20167 (N_20167,N_19524,N_19523);
xor U20168 (N_20168,N_19822,N_19659);
nand U20169 (N_20169,N_19789,N_19575);
nand U20170 (N_20170,N_19921,N_19662);
or U20171 (N_20171,N_19802,N_19909);
nor U20172 (N_20172,N_19879,N_19528);
and U20173 (N_20173,N_19690,N_19601);
or U20174 (N_20174,N_19536,N_19611);
nor U20175 (N_20175,N_19771,N_19637);
or U20176 (N_20176,N_19890,N_19643);
xor U20177 (N_20177,N_19836,N_19845);
and U20178 (N_20178,N_19631,N_19604);
and U20179 (N_20179,N_19806,N_19508);
and U20180 (N_20180,N_19837,N_19633);
nor U20181 (N_20181,N_19993,N_19763);
nor U20182 (N_20182,N_19793,N_19805);
and U20183 (N_20183,N_19644,N_19737);
or U20184 (N_20184,N_19898,N_19530);
and U20185 (N_20185,N_19658,N_19653);
and U20186 (N_20186,N_19582,N_19781);
nor U20187 (N_20187,N_19503,N_19819);
nor U20188 (N_20188,N_19989,N_19634);
xor U20189 (N_20189,N_19598,N_19984);
nor U20190 (N_20190,N_19705,N_19500);
xor U20191 (N_20191,N_19753,N_19711);
xor U20192 (N_20192,N_19867,N_19712);
xor U20193 (N_20193,N_19614,N_19986);
xor U20194 (N_20194,N_19590,N_19953);
and U20195 (N_20195,N_19605,N_19828);
nand U20196 (N_20196,N_19981,N_19864);
and U20197 (N_20197,N_19517,N_19908);
and U20198 (N_20198,N_19687,N_19768);
xnor U20199 (N_20199,N_19925,N_19994);
nor U20200 (N_20200,N_19544,N_19791);
nand U20201 (N_20201,N_19730,N_19977);
and U20202 (N_20202,N_19891,N_19515);
xnor U20203 (N_20203,N_19954,N_19656);
or U20204 (N_20204,N_19719,N_19821);
nor U20205 (N_20205,N_19787,N_19619);
nor U20206 (N_20206,N_19522,N_19917);
nand U20207 (N_20207,N_19848,N_19839);
xor U20208 (N_20208,N_19843,N_19666);
xnor U20209 (N_20209,N_19865,N_19972);
and U20210 (N_20210,N_19882,N_19861);
xor U20211 (N_20211,N_19937,N_19657);
xor U20212 (N_20212,N_19979,N_19929);
nand U20213 (N_20213,N_19661,N_19716);
nand U20214 (N_20214,N_19792,N_19529);
nand U20215 (N_20215,N_19769,N_19710);
or U20216 (N_20216,N_19823,N_19997);
xor U20217 (N_20217,N_19665,N_19565);
nor U20218 (N_20218,N_19718,N_19835);
and U20219 (N_20219,N_19721,N_19934);
xnor U20220 (N_20220,N_19886,N_19893);
and U20221 (N_20221,N_19810,N_19550);
nor U20222 (N_20222,N_19906,N_19899);
and U20223 (N_20223,N_19774,N_19788);
nor U20224 (N_20224,N_19764,N_19560);
or U20225 (N_20225,N_19968,N_19878);
or U20226 (N_20226,N_19892,N_19963);
and U20227 (N_20227,N_19727,N_19754);
xor U20228 (N_20228,N_19852,N_19670);
nor U20229 (N_20229,N_19851,N_19869);
nand U20230 (N_20230,N_19675,N_19555);
and U20231 (N_20231,N_19976,N_19600);
nor U20232 (N_20232,N_19826,N_19922);
nor U20233 (N_20233,N_19704,N_19617);
nor U20234 (N_20234,N_19942,N_19526);
and U20235 (N_20235,N_19877,N_19912);
xnor U20236 (N_20236,N_19571,N_19731);
xnor U20237 (N_20237,N_19775,N_19607);
xnor U20238 (N_20238,N_19951,N_19813);
nand U20239 (N_20239,N_19543,N_19903);
nand U20240 (N_20240,N_19849,N_19742);
and U20241 (N_20241,N_19521,N_19551);
nand U20242 (N_20242,N_19679,N_19676);
or U20243 (N_20243,N_19913,N_19606);
nor U20244 (N_20244,N_19998,N_19811);
and U20245 (N_20245,N_19999,N_19866);
or U20246 (N_20246,N_19853,N_19597);
and U20247 (N_20247,N_19701,N_19608);
and U20248 (N_20248,N_19514,N_19610);
or U20249 (N_20249,N_19578,N_19506);
and U20250 (N_20250,N_19780,N_19525);
and U20251 (N_20251,N_19703,N_19686);
nand U20252 (N_20252,N_19582,N_19720);
or U20253 (N_20253,N_19907,N_19668);
xor U20254 (N_20254,N_19681,N_19867);
and U20255 (N_20255,N_19778,N_19937);
nor U20256 (N_20256,N_19671,N_19634);
xor U20257 (N_20257,N_19734,N_19874);
nor U20258 (N_20258,N_19779,N_19785);
nand U20259 (N_20259,N_19514,N_19718);
nand U20260 (N_20260,N_19936,N_19922);
and U20261 (N_20261,N_19909,N_19789);
or U20262 (N_20262,N_19822,N_19836);
nand U20263 (N_20263,N_19857,N_19782);
xnor U20264 (N_20264,N_19713,N_19897);
and U20265 (N_20265,N_19656,N_19707);
xnor U20266 (N_20266,N_19964,N_19619);
nor U20267 (N_20267,N_19927,N_19835);
xor U20268 (N_20268,N_19724,N_19739);
or U20269 (N_20269,N_19695,N_19828);
xnor U20270 (N_20270,N_19897,N_19517);
xnor U20271 (N_20271,N_19997,N_19904);
and U20272 (N_20272,N_19953,N_19966);
xnor U20273 (N_20273,N_19998,N_19551);
xor U20274 (N_20274,N_19575,N_19815);
nor U20275 (N_20275,N_19827,N_19911);
xor U20276 (N_20276,N_19684,N_19681);
and U20277 (N_20277,N_19742,N_19708);
xor U20278 (N_20278,N_19947,N_19955);
and U20279 (N_20279,N_19717,N_19725);
xnor U20280 (N_20280,N_19610,N_19743);
and U20281 (N_20281,N_19848,N_19799);
xor U20282 (N_20282,N_19954,N_19741);
nand U20283 (N_20283,N_19637,N_19559);
nand U20284 (N_20284,N_19627,N_19932);
or U20285 (N_20285,N_19833,N_19838);
xor U20286 (N_20286,N_19535,N_19593);
nor U20287 (N_20287,N_19772,N_19783);
or U20288 (N_20288,N_19665,N_19812);
xor U20289 (N_20289,N_19763,N_19912);
nand U20290 (N_20290,N_19910,N_19786);
nand U20291 (N_20291,N_19685,N_19883);
or U20292 (N_20292,N_19924,N_19928);
xnor U20293 (N_20293,N_19746,N_19704);
xor U20294 (N_20294,N_19606,N_19922);
nor U20295 (N_20295,N_19630,N_19962);
nor U20296 (N_20296,N_19841,N_19920);
or U20297 (N_20297,N_19872,N_19905);
nand U20298 (N_20298,N_19684,N_19558);
and U20299 (N_20299,N_19521,N_19893);
nand U20300 (N_20300,N_19534,N_19749);
or U20301 (N_20301,N_19974,N_19990);
and U20302 (N_20302,N_19636,N_19566);
or U20303 (N_20303,N_19757,N_19925);
nand U20304 (N_20304,N_19527,N_19811);
xor U20305 (N_20305,N_19977,N_19954);
xnor U20306 (N_20306,N_19984,N_19972);
or U20307 (N_20307,N_19551,N_19528);
nand U20308 (N_20308,N_19671,N_19850);
nand U20309 (N_20309,N_19679,N_19568);
nor U20310 (N_20310,N_19899,N_19923);
nor U20311 (N_20311,N_19931,N_19987);
nor U20312 (N_20312,N_19576,N_19848);
and U20313 (N_20313,N_19794,N_19694);
nor U20314 (N_20314,N_19835,N_19833);
xor U20315 (N_20315,N_19597,N_19750);
and U20316 (N_20316,N_19978,N_19561);
or U20317 (N_20317,N_19769,N_19751);
nand U20318 (N_20318,N_19635,N_19986);
nand U20319 (N_20319,N_19712,N_19767);
nand U20320 (N_20320,N_19541,N_19973);
nor U20321 (N_20321,N_19566,N_19632);
and U20322 (N_20322,N_19528,N_19661);
and U20323 (N_20323,N_19816,N_19552);
xnor U20324 (N_20324,N_19859,N_19850);
nor U20325 (N_20325,N_19739,N_19719);
nand U20326 (N_20326,N_19752,N_19712);
and U20327 (N_20327,N_19614,N_19633);
nand U20328 (N_20328,N_19596,N_19816);
or U20329 (N_20329,N_19694,N_19506);
and U20330 (N_20330,N_19863,N_19572);
nor U20331 (N_20331,N_19598,N_19912);
nand U20332 (N_20332,N_19749,N_19922);
nor U20333 (N_20333,N_19552,N_19678);
xor U20334 (N_20334,N_19525,N_19806);
and U20335 (N_20335,N_19751,N_19646);
or U20336 (N_20336,N_19663,N_19660);
nand U20337 (N_20337,N_19713,N_19517);
and U20338 (N_20338,N_19874,N_19621);
nor U20339 (N_20339,N_19993,N_19658);
or U20340 (N_20340,N_19997,N_19890);
or U20341 (N_20341,N_19648,N_19818);
or U20342 (N_20342,N_19651,N_19517);
and U20343 (N_20343,N_19852,N_19573);
nor U20344 (N_20344,N_19728,N_19724);
nor U20345 (N_20345,N_19726,N_19599);
nand U20346 (N_20346,N_19766,N_19950);
and U20347 (N_20347,N_19785,N_19601);
nor U20348 (N_20348,N_19863,N_19813);
nor U20349 (N_20349,N_19817,N_19782);
or U20350 (N_20350,N_19863,N_19596);
and U20351 (N_20351,N_19835,N_19545);
and U20352 (N_20352,N_19845,N_19694);
and U20353 (N_20353,N_19564,N_19823);
and U20354 (N_20354,N_19859,N_19714);
and U20355 (N_20355,N_19837,N_19849);
and U20356 (N_20356,N_19504,N_19908);
or U20357 (N_20357,N_19538,N_19985);
nand U20358 (N_20358,N_19617,N_19966);
xor U20359 (N_20359,N_19766,N_19516);
nand U20360 (N_20360,N_19849,N_19860);
nor U20361 (N_20361,N_19819,N_19629);
or U20362 (N_20362,N_19830,N_19613);
or U20363 (N_20363,N_19651,N_19505);
nor U20364 (N_20364,N_19682,N_19977);
or U20365 (N_20365,N_19933,N_19694);
and U20366 (N_20366,N_19741,N_19715);
and U20367 (N_20367,N_19706,N_19690);
and U20368 (N_20368,N_19685,N_19644);
xnor U20369 (N_20369,N_19554,N_19551);
and U20370 (N_20370,N_19659,N_19764);
nor U20371 (N_20371,N_19673,N_19742);
or U20372 (N_20372,N_19817,N_19785);
and U20373 (N_20373,N_19843,N_19805);
and U20374 (N_20374,N_19788,N_19604);
nor U20375 (N_20375,N_19549,N_19604);
nor U20376 (N_20376,N_19939,N_19572);
xor U20377 (N_20377,N_19503,N_19821);
nor U20378 (N_20378,N_19939,N_19851);
or U20379 (N_20379,N_19805,N_19865);
nor U20380 (N_20380,N_19767,N_19884);
xor U20381 (N_20381,N_19776,N_19603);
and U20382 (N_20382,N_19629,N_19550);
or U20383 (N_20383,N_19788,N_19889);
and U20384 (N_20384,N_19701,N_19556);
or U20385 (N_20385,N_19967,N_19894);
or U20386 (N_20386,N_19661,N_19691);
nand U20387 (N_20387,N_19662,N_19538);
and U20388 (N_20388,N_19990,N_19948);
nand U20389 (N_20389,N_19611,N_19712);
nand U20390 (N_20390,N_19648,N_19635);
xnor U20391 (N_20391,N_19598,N_19907);
and U20392 (N_20392,N_19814,N_19645);
or U20393 (N_20393,N_19765,N_19501);
nand U20394 (N_20394,N_19574,N_19982);
nand U20395 (N_20395,N_19503,N_19540);
and U20396 (N_20396,N_19634,N_19765);
xor U20397 (N_20397,N_19999,N_19608);
and U20398 (N_20398,N_19919,N_19767);
nand U20399 (N_20399,N_19533,N_19568);
nand U20400 (N_20400,N_19645,N_19745);
nor U20401 (N_20401,N_19961,N_19855);
and U20402 (N_20402,N_19749,N_19832);
xnor U20403 (N_20403,N_19547,N_19696);
nor U20404 (N_20404,N_19988,N_19931);
nor U20405 (N_20405,N_19671,N_19847);
xnor U20406 (N_20406,N_19573,N_19716);
nand U20407 (N_20407,N_19978,N_19971);
nor U20408 (N_20408,N_19543,N_19862);
nand U20409 (N_20409,N_19867,N_19548);
and U20410 (N_20410,N_19905,N_19703);
or U20411 (N_20411,N_19522,N_19788);
xor U20412 (N_20412,N_19849,N_19596);
or U20413 (N_20413,N_19555,N_19805);
and U20414 (N_20414,N_19920,N_19636);
nand U20415 (N_20415,N_19776,N_19952);
and U20416 (N_20416,N_19627,N_19914);
nand U20417 (N_20417,N_19885,N_19929);
and U20418 (N_20418,N_19944,N_19671);
or U20419 (N_20419,N_19724,N_19848);
nand U20420 (N_20420,N_19800,N_19968);
or U20421 (N_20421,N_19805,N_19985);
nor U20422 (N_20422,N_19939,N_19694);
and U20423 (N_20423,N_19562,N_19808);
or U20424 (N_20424,N_19898,N_19981);
and U20425 (N_20425,N_19967,N_19532);
and U20426 (N_20426,N_19898,N_19605);
nand U20427 (N_20427,N_19512,N_19820);
nor U20428 (N_20428,N_19767,N_19954);
or U20429 (N_20429,N_19898,N_19956);
nand U20430 (N_20430,N_19622,N_19946);
nand U20431 (N_20431,N_19725,N_19748);
xnor U20432 (N_20432,N_19618,N_19848);
nand U20433 (N_20433,N_19728,N_19685);
or U20434 (N_20434,N_19674,N_19866);
nor U20435 (N_20435,N_19719,N_19922);
nor U20436 (N_20436,N_19722,N_19732);
and U20437 (N_20437,N_19593,N_19995);
nand U20438 (N_20438,N_19787,N_19796);
nand U20439 (N_20439,N_19737,N_19540);
nor U20440 (N_20440,N_19632,N_19647);
nand U20441 (N_20441,N_19763,N_19680);
nor U20442 (N_20442,N_19760,N_19507);
nand U20443 (N_20443,N_19768,N_19742);
or U20444 (N_20444,N_19704,N_19647);
and U20445 (N_20445,N_19987,N_19558);
and U20446 (N_20446,N_19942,N_19920);
and U20447 (N_20447,N_19915,N_19664);
nor U20448 (N_20448,N_19896,N_19638);
or U20449 (N_20449,N_19723,N_19825);
nor U20450 (N_20450,N_19862,N_19536);
nor U20451 (N_20451,N_19806,N_19542);
nand U20452 (N_20452,N_19761,N_19998);
or U20453 (N_20453,N_19953,N_19844);
xor U20454 (N_20454,N_19906,N_19992);
or U20455 (N_20455,N_19952,N_19985);
or U20456 (N_20456,N_19861,N_19982);
or U20457 (N_20457,N_19717,N_19793);
nor U20458 (N_20458,N_19527,N_19969);
and U20459 (N_20459,N_19970,N_19856);
and U20460 (N_20460,N_19759,N_19691);
nand U20461 (N_20461,N_19756,N_19843);
nand U20462 (N_20462,N_19662,N_19987);
xor U20463 (N_20463,N_19600,N_19532);
and U20464 (N_20464,N_19801,N_19630);
or U20465 (N_20465,N_19839,N_19897);
nand U20466 (N_20466,N_19616,N_19841);
xnor U20467 (N_20467,N_19912,N_19786);
xor U20468 (N_20468,N_19758,N_19683);
nand U20469 (N_20469,N_19787,N_19772);
and U20470 (N_20470,N_19725,N_19700);
xor U20471 (N_20471,N_19893,N_19722);
nor U20472 (N_20472,N_19579,N_19904);
xnor U20473 (N_20473,N_19688,N_19895);
and U20474 (N_20474,N_19600,N_19940);
or U20475 (N_20475,N_19945,N_19827);
nor U20476 (N_20476,N_19861,N_19626);
nor U20477 (N_20477,N_19836,N_19625);
nor U20478 (N_20478,N_19848,N_19609);
or U20479 (N_20479,N_19998,N_19665);
and U20480 (N_20480,N_19659,N_19635);
nor U20481 (N_20481,N_19952,N_19745);
and U20482 (N_20482,N_19688,N_19664);
and U20483 (N_20483,N_19838,N_19642);
nand U20484 (N_20484,N_19638,N_19783);
or U20485 (N_20485,N_19898,N_19752);
nor U20486 (N_20486,N_19824,N_19550);
nand U20487 (N_20487,N_19513,N_19740);
and U20488 (N_20488,N_19610,N_19637);
xnor U20489 (N_20489,N_19580,N_19804);
nand U20490 (N_20490,N_19813,N_19718);
xor U20491 (N_20491,N_19659,N_19692);
and U20492 (N_20492,N_19928,N_19506);
xor U20493 (N_20493,N_19734,N_19792);
or U20494 (N_20494,N_19990,N_19664);
xor U20495 (N_20495,N_19643,N_19778);
nand U20496 (N_20496,N_19703,N_19963);
and U20497 (N_20497,N_19593,N_19924);
nor U20498 (N_20498,N_19845,N_19973);
or U20499 (N_20499,N_19936,N_19920);
xnor U20500 (N_20500,N_20199,N_20149);
or U20501 (N_20501,N_20073,N_20295);
and U20502 (N_20502,N_20190,N_20092);
nand U20503 (N_20503,N_20291,N_20211);
nor U20504 (N_20504,N_20287,N_20377);
and U20505 (N_20505,N_20054,N_20138);
nand U20506 (N_20506,N_20242,N_20479);
xor U20507 (N_20507,N_20449,N_20387);
and U20508 (N_20508,N_20484,N_20297);
or U20509 (N_20509,N_20298,N_20410);
nand U20510 (N_20510,N_20011,N_20186);
or U20511 (N_20511,N_20458,N_20396);
nand U20512 (N_20512,N_20355,N_20338);
xor U20513 (N_20513,N_20215,N_20266);
nor U20514 (N_20514,N_20476,N_20084);
nand U20515 (N_20515,N_20263,N_20280);
and U20516 (N_20516,N_20093,N_20462);
xnor U20517 (N_20517,N_20113,N_20038);
xor U20518 (N_20518,N_20028,N_20294);
xor U20519 (N_20519,N_20078,N_20408);
nor U20520 (N_20520,N_20130,N_20374);
nor U20521 (N_20521,N_20002,N_20053);
xor U20522 (N_20522,N_20492,N_20421);
and U20523 (N_20523,N_20496,N_20499);
nand U20524 (N_20524,N_20075,N_20279);
xnor U20525 (N_20525,N_20224,N_20193);
or U20526 (N_20526,N_20292,N_20276);
or U20527 (N_20527,N_20386,N_20069);
nand U20528 (N_20528,N_20248,N_20413);
and U20529 (N_20529,N_20445,N_20335);
and U20530 (N_20530,N_20465,N_20346);
and U20531 (N_20531,N_20194,N_20083);
nand U20532 (N_20532,N_20375,N_20045);
or U20533 (N_20533,N_20226,N_20336);
xnor U20534 (N_20534,N_20475,N_20156);
xor U20535 (N_20535,N_20343,N_20316);
nand U20536 (N_20536,N_20022,N_20174);
xor U20537 (N_20537,N_20409,N_20125);
nand U20538 (N_20538,N_20042,N_20129);
xor U20539 (N_20539,N_20000,N_20383);
or U20540 (N_20540,N_20014,N_20171);
or U20541 (N_20541,N_20235,N_20183);
nor U20542 (N_20542,N_20210,N_20371);
xor U20543 (N_20543,N_20332,N_20036);
and U20544 (N_20544,N_20273,N_20357);
or U20545 (N_20545,N_20139,N_20019);
xnor U20546 (N_20546,N_20488,N_20257);
nor U20547 (N_20547,N_20310,N_20351);
nand U20548 (N_20548,N_20182,N_20450);
nor U20549 (N_20549,N_20474,N_20286);
nor U20550 (N_20550,N_20430,N_20392);
xor U20551 (N_20551,N_20487,N_20285);
nand U20552 (N_20552,N_20344,N_20153);
and U20553 (N_20553,N_20065,N_20158);
or U20554 (N_20554,N_20018,N_20366);
nor U20555 (N_20555,N_20068,N_20032);
and U20556 (N_20556,N_20233,N_20031);
nor U20557 (N_20557,N_20241,N_20380);
and U20558 (N_20558,N_20472,N_20363);
nor U20559 (N_20559,N_20200,N_20132);
xor U20560 (N_20560,N_20320,N_20070);
xor U20561 (N_20561,N_20391,N_20003);
nor U20562 (N_20562,N_20309,N_20164);
nand U20563 (N_20563,N_20091,N_20090);
and U20564 (N_20564,N_20117,N_20107);
and U20565 (N_20565,N_20096,N_20470);
and U20566 (N_20566,N_20037,N_20122);
nand U20567 (N_20567,N_20061,N_20317);
and U20568 (N_20568,N_20364,N_20238);
xnor U20569 (N_20569,N_20469,N_20035);
xor U20570 (N_20570,N_20218,N_20356);
nor U20571 (N_20571,N_20467,N_20017);
or U20572 (N_20572,N_20397,N_20486);
nand U20573 (N_20573,N_20063,N_20362);
and U20574 (N_20574,N_20024,N_20209);
xnor U20575 (N_20575,N_20227,N_20460);
nand U20576 (N_20576,N_20468,N_20105);
xor U20577 (N_20577,N_20439,N_20051);
and U20578 (N_20578,N_20121,N_20142);
or U20579 (N_20579,N_20172,N_20013);
nor U20580 (N_20580,N_20119,N_20217);
and U20581 (N_20581,N_20106,N_20365);
and U20582 (N_20582,N_20389,N_20066);
nand U20583 (N_20583,N_20097,N_20133);
nor U20584 (N_20584,N_20278,N_20456);
nand U20585 (N_20585,N_20021,N_20373);
nor U20586 (N_20586,N_20085,N_20252);
nor U20587 (N_20587,N_20060,N_20195);
or U20588 (N_20588,N_20128,N_20020);
nor U20589 (N_20589,N_20342,N_20434);
xnor U20590 (N_20590,N_20322,N_20141);
and U20591 (N_20591,N_20176,N_20481);
or U20592 (N_20592,N_20400,N_20345);
or U20593 (N_20593,N_20290,N_20206);
xnor U20594 (N_20594,N_20111,N_20094);
and U20595 (N_20595,N_20010,N_20333);
and U20596 (N_20596,N_20426,N_20379);
nand U20597 (N_20597,N_20267,N_20131);
xnor U20598 (N_20598,N_20464,N_20431);
and U20599 (N_20599,N_20260,N_20315);
and U20600 (N_20600,N_20359,N_20148);
or U20601 (N_20601,N_20382,N_20079);
xor U20602 (N_20602,N_20304,N_20212);
or U20603 (N_20603,N_20247,N_20098);
nor U20604 (N_20604,N_20104,N_20127);
or U20605 (N_20605,N_20436,N_20058);
xor U20606 (N_20606,N_20205,N_20432);
nand U20607 (N_20607,N_20394,N_20015);
nand U20608 (N_20608,N_20480,N_20393);
nor U20609 (N_20609,N_20422,N_20180);
nor U20610 (N_20610,N_20477,N_20440);
nand U20611 (N_20611,N_20323,N_20214);
nand U20612 (N_20612,N_20006,N_20026);
or U20613 (N_20613,N_20497,N_20428);
nor U20614 (N_20614,N_20225,N_20262);
xnor U20615 (N_20615,N_20245,N_20367);
and U20616 (N_20616,N_20419,N_20289);
or U20617 (N_20617,N_20123,N_20049);
nand U20618 (N_20618,N_20108,N_20404);
and U20619 (N_20619,N_20187,N_20348);
xor U20620 (N_20620,N_20059,N_20326);
nor U20621 (N_20621,N_20376,N_20237);
or U20622 (N_20622,N_20269,N_20112);
nand U20623 (N_20623,N_20466,N_20258);
and U20624 (N_20624,N_20378,N_20438);
nor U20625 (N_20625,N_20372,N_20160);
nor U20626 (N_20626,N_20064,N_20314);
nand U20627 (N_20627,N_20411,N_20330);
xnor U20628 (N_20628,N_20056,N_20213);
xnor U20629 (N_20629,N_20340,N_20169);
xor U20630 (N_20630,N_20143,N_20243);
or U20631 (N_20631,N_20159,N_20162);
nor U20632 (N_20632,N_20087,N_20151);
xnor U20633 (N_20633,N_20170,N_20116);
nor U20634 (N_20634,N_20435,N_20145);
nand U20635 (N_20635,N_20339,N_20412);
or U20636 (N_20636,N_20095,N_20255);
nor U20637 (N_20637,N_20253,N_20249);
and U20638 (N_20638,N_20007,N_20202);
nor U20639 (N_20639,N_20448,N_20334);
and U20640 (N_20640,N_20204,N_20030);
nand U20641 (N_20641,N_20076,N_20441);
nor U20642 (N_20642,N_20306,N_20381);
nand U20643 (N_20643,N_20126,N_20039);
xnor U20644 (N_20644,N_20178,N_20311);
and U20645 (N_20645,N_20259,N_20296);
nand U20646 (N_20646,N_20181,N_20246);
nand U20647 (N_20647,N_20443,N_20293);
nor U20648 (N_20648,N_20319,N_20067);
nand U20649 (N_20649,N_20461,N_20114);
or U20650 (N_20650,N_20220,N_20155);
nand U20651 (N_20651,N_20184,N_20407);
nor U20652 (N_20652,N_20228,N_20299);
xnor U20653 (N_20653,N_20175,N_20350);
nand U20654 (N_20654,N_20166,N_20025);
and U20655 (N_20655,N_20109,N_20425);
nor U20656 (N_20656,N_20074,N_20288);
or U20657 (N_20657,N_20082,N_20254);
nor U20658 (N_20658,N_20232,N_20444);
xnor U20659 (N_20659,N_20327,N_20268);
nand U20660 (N_20660,N_20361,N_20427);
xnor U20661 (N_20661,N_20052,N_20009);
and U20662 (N_20662,N_20437,N_20004);
nor U20663 (N_20663,N_20473,N_20385);
or U20664 (N_20664,N_20349,N_20368);
xnor U20665 (N_20665,N_20399,N_20231);
or U20666 (N_20666,N_20494,N_20086);
nor U20667 (N_20667,N_20207,N_20453);
and U20668 (N_20668,N_20077,N_20150);
or U20669 (N_20669,N_20047,N_20489);
or U20670 (N_20670,N_20390,N_20457);
xor U20671 (N_20671,N_20167,N_20491);
xor U20672 (N_20672,N_20040,N_20118);
or U20673 (N_20673,N_20274,N_20302);
and U20674 (N_20674,N_20272,N_20081);
nor U20675 (N_20675,N_20454,N_20188);
xor U20676 (N_20676,N_20250,N_20418);
or U20677 (N_20677,N_20301,N_20201);
nor U20678 (N_20678,N_20482,N_20023);
nor U20679 (N_20679,N_20307,N_20414);
nand U20680 (N_20680,N_20451,N_20203);
xnor U20681 (N_20681,N_20275,N_20029);
nand U20682 (N_20682,N_20134,N_20221);
nand U20683 (N_20683,N_20463,N_20271);
or U20684 (N_20684,N_20189,N_20395);
and U20685 (N_20685,N_20354,N_20165);
and U20686 (N_20686,N_20337,N_20027);
xor U20687 (N_20687,N_20384,N_20401);
nand U20688 (N_20688,N_20452,N_20196);
xor U20689 (N_20689,N_20177,N_20041);
xnor U20690 (N_20690,N_20168,N_20099);
nor U20691 (N_20691,N_20230,N_20048);
nor U20692 (N_20692,N_20495,N_20137);
nor U20693 (N_20693,N_20352,N_20417);
nor U20694 (N_20694,N_20423,N_20324);
nand U20695 (N_20695,N_20146,N_20191);
and U20696 (N_20696,N_20234,N_20163);
xor U20697 (N_20697,N_20341,N_20208);
and U20698 (N_20698,N_20223,N_20012);
or U20699 (N_20699,N_20001,N_20455);
xnor U20700 (N_20700,N_20147,N_20144);
nand U20701 (N_20701,N_20135,N_20016);
nor U20702 (N_20702,N_20173,N_20062);
nand U20703 (N_20703,N_20124,N_20033);
nor U20704 (N_20704,N_20120,N_20136);
nand U20705 (N_20705,N_20157,N_20369);
and U20706 (N_20706,N_20005,N_20222);
or U20707 (N_20707,N_20325,N_20043);
or U20708 (N_20708,N_20328,N_20313);
or U20709 (N_20709,N_20198,N_20265);
nor U20710 (N_20710,N_20321,N_20072);
or U20711 (N_20711,N_20402,N_20442);
xor U20712 (N_20712,N_20034,N_20197);
nor U20713 (N_20713,N_20420,N_20088);
nand U20714 (N_20714,N_20493,N_20300);
xor U20715 (N_20715,N_20050,N_20219);
nand U20716 (N_20716,N_20485,N_20115);
and U20717 (N_20717,N_20008,N_20490);
nor U20718 (N_20718,N_20110,N_20406);
nand U20719 (N_20719,N_20284,N_20471);
or U20720 (N_20720,N_20353,N_20370);
nor U20721 (N_20721,N_20282,N_20152);
nor U20722 (N_20722,N_20283,N_20192);
xnor U20723 (N_20723,N_20046,N_20478);
nand U20724 (N_20724,N_20303,N_20483);
nor U20725 (N_20725,N_20447,N_20261);
nor U20726 (N_20726,N_20429,N_20229);
and U20727 (N_20727,N_20102,N_20398);
and U20728 (N_20728,N_20305,N_20277);
nand U20729 (N_20729,N_20459,N_20071);
and U20730 (N_20730,N_20358,N_20100);
xnor U20731 (N_20731,N_20415,N_20433);
nand U20732 (N_20732,N_20236,N_20154);
or U20733 (N_20733,N_20264,N_20360);
nand U20734 (N_20734,N_20179,N_20057);
or U20735 (N_20735,N_20101,N_20244);
xor U20736 (N_20736,N_20140,N_20329);
nor U20737 (N_20737,N_20331,N_20388);
and U20738 (N_20738,N_20312,N_20251);
and U20739 (N_20739,N_20239,N_20405);
xor U20740 (N_20740,N_20256,N_20403);
nand U20741 (N_20741,N_20416,N_20498);
or U20742 (N_20742,N_20103,N_20318);
nor U20743 (N_20743,N_20270,N_20044);
nand U20744 (N_20744,N_20161,N_20446);
nand U20745 (N_20745,N_20424,N_20240);
nor U20746 (N_20746,N_20216,N_20347);
or U20747 (N_20747,N_20308,N_20089);
nor U20748 (N_20748,N_20281,N_20080);
nand U20749 (N_20749,N_20185,N_20055);
or U20750 (N_20750,N_20276,N_20203);
and U20751 (N_20751,N_20175,N_20317);
and U20752 (N_20752,N_20448,N_20298);
xor U20753 (N_20753,N_20409,N_20199);
or U20754 (N_20754,N_20366,N_20147);
nand U20755 (N_20755,N_20142,N_20083);
or U20756 (N_20756,N_20386,N_20071);
and U20757 (N_20757,N_20443,N_20201);
nand U20758 (N_20758,N_20480,N_20227);
nand U20759 (N_20759,N_20058,N_20071);
or U20760 (N_20760,N_20257,N_20311);
xor U20761 (N_20761,N_20310,N_20331);
and U20762 (N_20762,N_20227,N_20442);
nand U20763 (N_20763,N_20172,N_20278);
nand U20764 (N_20764,N_20281,N_20246);
nand U20765 (N_20765,N_20420,N_20042);
nand U20766 (N_20766,N_20307,N_20493);
xnor U20767 (N_20767,N_20158,N_20421);
and U20768 (N_20768,N_20092,N_20165);
xnor U20769 (N_20769,N_20005,N_20130);
and U20770 (N_20770,N_20090,N_20098);
or U20771 (N_20771,N_20071,N_20227);
nor U20772 (N_20772,N_20173,N_20003);
xnor U20773 (N_20773,N_20234,N_20463);
or U20774 (N_20774,N_20240,N_20046);
nor U20775 (N_20775,N_20436,N_20162);
or U20776 (N_20776,N_20041,N_20328);
and U20777 (N_20777,N_20459,N_20417);
xor U20778 (N_20778,N_20206,N_20317);
nor U20779 (N_20779,N_20275,N_20494);
xnor U20780 (N_20780,N_20371,N_20452);
xnor U20781 (N_20781,N_20347,N_20147);
nor U20782 (N_20782,N_20147,N_20358);
nor U20783 (N_20783,N_20176,N_20049);
nand U20784 (N_20784,N_20272,N_20309);
nor U20785 (N_20785,N_20095,N_20233);
or U20786 (N_20786,N_20496,N_20102);
xor U20787 (N_20787,N_20474,N_20128);
nand U20788 (N_20788,N_20140,N_20069);
xnor U20789 (N_20789,N_20366,N_20365);
and U20790 (N_20790,N_20441,N_20077);
nand U20791 (N_20791,N_20347,N_20356);
and U20792 (N_20792,N_20068,N_20088);
or U20793 (N_20793,N_20428,N_20142);
or U20794 (N_20794,N_20266,N_20330);
nor U20795 (N_20795,N_20231,N_20261);
nor U20796 (N_20796,N_20164,N_20186);
and U20797 (N_20797,N_20218,N_20457);
nand U20798 (N_20798,N_20344,N_20295);
or U20799 (N_20799,N_20429,N_20481);
nor U20800 (N_20800,N_20293,N_20252);
nor U20801 (N_20801,N_20092,N_20063);
nor U20802 (N_20802,N_20074,N_20197);
nor U20803 (N_20803,N_20346,N_20460);
or U20804 (N_20804,N_20122,N_20446);
nor U20805 (N_20805,N_20147,N_20268);
or U20806 (N_20806,N_20215,N_20150);
nand U20807 (N_20807,N_20491,N_20247);
or U20808 (N_20808,N_20486,N_20293);
and U20809 (N_20809,N_20119,N_20218);
nand U20810 (N_20810,N_20242,N_20203);
nor U20811 (N_20811,N_20397,N_20306);
nor U20812 (N_20812,N_20492,N_20473);
nand U20813 (N_20813,N_20205,N_20165);
and U20814 (N_20814,N_20297,N_20089);
or U20815 (N_20815,N_20194,N_20170);
nor U20816 (N_20816,N_20158,N_20118);
and U20817 (N_20817,N_20021,N_20357);
xor U20818 (N_20818,N_20277,N_20301);
nand U20819 (N_20819,N_20040,N_20434);
nand U20820 (N_20820,N_20101,N_20085);
and U20821 (N_20821,N_20076,N_20461);
nand U20822 (N_20822,N_20115,N_20250);
nand U20823 (N_20823,N_20369,N_20463);
or U20824 (N_20824,N_20071,N_20442);
nand U20825 (N_20825,N_20019,N_20438);
nor U20826 (N_20826,N_20120,N_20474);
xor U20827 (N_20827,N_20306,N_20067);
nand U20828 (N_20828,N_20022,N_20478);
or U20829 (N_20829,N_20114,N_20060);
nor U20830 (N_20830,N_20178,N_20264);
nand U20831 (N_20831,N_20452,N_20495);
xor U20832 (N_20832,N_20403,N_20387);
nor U20833 (N_20833,N_20099,N_20317);
nor U20834 (N_20834,N_20391,N_20396);
xor U20835 (N_20835,N_20124,N_20101);
or U20836 (N_20836,N_20391,N_20373);
xnor U20837 (N_20837,N_20362,N_20243);
and U20838 (N_20838,N_20482,N_20111);
or U20839 (N_20839,N_20366,N_20156);
and U20840 (N_20840,N_20163,N_20155);
nor U20841 (N_20841,N_20334,N_20422);
nor U20842 (N_20842,N_20047,N_20117);
nor U20843 (N_20843,N_20027,N_20311);
and U20844 (N_20844,N_20415,N_20332);
and U20845 (N_20845,N_20021,N_20019);
or U20846 (N_20846,N_20035,N_20099);
and U20847 (N_20847,N_20445,N_20485);
nand U20848 (N_20848,N_20460,N_20359);
or U20849 (N_20849,N_20187,N_20166);
and U20850 (N_20850,N_20334,N_20364);
and U20851 (N_20851,N_20230,N_20120);
nand U20852 (N_20852,N_20107,N_20079);
nand U20853 (N_20853,N_20194,N_20291);
xnor U20854 (N_20854,N_20155,N_20125);
nor U20855 (N_20855,N_20149,N_20494);
and U20856 (N_20856,N_20160,N_20305);
nand U20857 (N_20857,N_20114,N_20293);
and U20858 (N_20858,N_20452,N_20210);
xnor U20859 (N_20859,N_20361,N_20189);
nor U20860 (N_20860,N_20438,N_20181);
and U20861 (N_20861,N_20361,N_20352);
xnor U20862 (N_20862,N_20388,N_20024);
nor U20863 (N_20863,N_20073,N_20165);
nor U20864 (N_20864,N_20120,N_20064);
nor U20865 (N_20865,N_20111,N_20330);
or U20866 (N_20866,N_20368,N_20237);
or U20867 (N_20867,N_20208,N_20365);
or U20868 (N_20868,N_20238,N_20309);
xor U20869 (N_20869,N_20061,N_20459);
nor U20870 (N_20870,N_20471,N_20356);
xnor U20871 (N_20871,N_20008,N_20042);
or U20872 (N_20872,N_20398,N_20273);
nand U20873 (N_20873,N_20456,N_20411);
nor U20874 (N_20874,N_20369,N_20160);
nand U20875 (N_20875,N_20019,N_20159);
nand U20876 (N_20876,N_20130,N_20174);
nor U20877 (N_20877,N_20210,N_20030);
nor U20878 (N_20878,N_20319,N_20216);
nor U20879 (N_20879,N_20080,N_20111);
or U20880 (N_20880,N_20214,N_20434);
and U20881 (N_20881,N_20201,N_20400);
nor U20882 (N_20882,N_20309,N_20303);
nand U20883 (N_20883,N_20054,N_20077);
and U20884 (N_20884,N_20436,N_20490);
nor U20885 (N_20885,N_20364,N_20321);
and U20886 (N_20886,N_20301,N_20467);
nand U20887 (N_20887,N_20358,N_20437);
or U20888 (N_20888,N_20001,N_20315);
xnor U20889 (N_20889,N_20260,N_20378);
nand U20890 (N_20890,N_20497,N_20335);
nor U20891 (N_20891,N_20397,N_20269);
nor U20892 (N_20892,N_20382,N_20499);
xor U20893 (N_20893,N_20294,N_20361);
and U20894 (N_20894,N_20200,N_20285);
nand U20895 (N_20895,N_20345,N_20201);
xor U20896 (N_20896,N_20130,N_20373);
or U20897 (N_20897,N_20462,N_20136);
or U20898 (N_20898,N_20009,N_20390);
nand U20899 (N_20899,N_20462,N_20089);
or U20900 (N_20900,N_20361,N_20041);
or U20901 (N_20901,N_20491,N_20451);
and U20902 (N_20902,N_20358,N_20062);
and U20903 (N_20903,N_20013,N_20049);
nor U20904 (N_20904,N_20385,N_20380);
and U20905 (N_20905,N_20262,N_20273);
xor U20906 (N_20906,N_20281,N_20215);
xnor U20907 (N_20907,N_20248,N_20244);
nand U20908 (N_20908,N_20149,N_20173);
and U20909 (N_20909,N_20418,N_20219);
nand U20910 (N_20910,N_20134,N_20012);
and U20911 (N_20911,N_20059,N_20284);
and U20912 (N_20912,N_20206,N_20367);
or U20913 (N_20913,N_20328,N_20048);
nand U20914 (N_20914,N_20010,N_20098);
nor U20915 (N_20915,N_20106,N_20044);
nor U20916 (N_20916,N_20053,N_20184);
xor U20917 (N_20917,N_20130,N_20054);
nor U20918 (N_20918,N_20218,N_20323);
xnor U20919 (N_20919,N_20321,N_20342);
nand U20920 (N_20920,N_20076,N_20106);
and U20921 (N_20921,N_20434,N_20186);
xnor U20922 (N_20922,N_20352,N_20455);
or U20923 (N_20923,N_20198,N_20068);
xnor U20924 (N_20924,N_20438,N_20235);
nand U20925 (N_20925,N_20115,N_20431);
or U20926 (N_20926,N_20186,N_20240);
xor U20927 (N_20927,N_20328,N_20277);
and U20928 (N_20928,N_20283,N_20078);
or U20929 (N_20929,N_20033,N_20138);
nand U20930 (N_20930,N_20172,N_20441);
and U20931 (N_20931,N_20024,N_20065);
nand U20932 (N_20932,N_20387,N_20239);
and U20933 (N_20933,N_20080,N_20380);
nor U20934 (N_20934,N_20092,N_20273);
and U20935 (N_20935,N_20033,N_20067);
or U20936 (N_20936,N_20318,N_20280);
or U20937 (N_20937,N_20178,N_20128);
and U20938 (N_20938,N_20010,N_20485);
xnor U20939 (N_20939,N_20265,N_20099);
nand U20940 (N_20940,N_20287,N_20183);
xnor U20941 (N_20941,N_20160,N_20210);
nand U20942 (N_20942,N_20476,N_20108);
and U20943 (N_20943,N_20085,N_20330);
and U20944 (N_20944,N_20256,N_20428);
and U20945 (N_20945,N_20046,N_20122);
nor U20946 (N_20946,N_20383,N_20316);
or U20947 (N_20947,N_20411,N_20347);
nand U20948 (N_20948,N_20455,N_20475);
and U20949 (N_20949,N_20348,N_20317);
and U20950 (N_20950,N_20200,N_20230);
nand U20951 (N_20951,N_20063,N_20112);
nor U20952 (N_20952,N_20085,N_20454);
xnor U20953 (N_20953,N_20313,N_20342);
xor U20954 (N_20954,N_20002,N_20068);
or U20955 (N_20955,N_20187,N_20414);
nand U20956 (N_20956,N_20113,N_20246);
and U20957 (N_20957,N_20330,N_20472);
nand U20958 (N_20958,N_20488,N_20135);
nand U20959 (N_20959,N_20371,N_20039);
xor U20960 (N_20960,N_20219,N_20252);
nor U20961 (N_20961,N_20311,N_20410);
xnor U20962 (N_20962,N_20483,N_20338);
and U20963 (N_20963,N_20014,N_20016);
xnor U20964 (N_20964,N_20425,N_20085);
nand U20965 (N_20965,N_20011,N_20010);
xor U20966 (N_20966,N_20225,N_20358);
or U20967 (N_20967,N_20100,N_20391);
nor U20968 (N_20968,N_20479,N_20354);
nor U20969 (N_20969,N_20119,N_20233);
nand U20970 (N_20970,N_20252,N_20390);
and U20971 (N_20971,N_20194,N_20001);
nand U20972 (N_20972,N_20083,N_20121);
nand U20973 (N_20973,N_20198,N_20276);
nand U20974 (N_20974,N_20098,N_20069);
nand U20975 (N_20975,N_20410,N_20440);
and U20976 (N_20976,N_20049,N_20209);
xnor U20977 (N_20977,N_20141,N_20476);
nand U20978 (N_20978,N_20132,N_20201);
xnor U20979 (N_20979,N_20075,N_20490);
and U20980 (N_20980,N_20235,N_20247);
nor U20981 (N_20981,N_20189,N_20343);
and U20982 (N_20982,N_20000,N_20225);
or U20983 (N_20983,N_20167,N_20108);
or U20984 (N_20984,N_20127,N_20409);
xnor U20985 (N_20985,N_20176,N_20392);
nor U20986 (N_20986,N_20159,N_20333);
nand U20987 (N_20987,N_20178,N_20171);
or U20988 (N_20988,N_20315,N_20353);
and U20989 (N_20989,N_20135,N_20402);
or U20990 (N_20990,N_20052,N_20271);
xor U20991 (N_20991,N_20418,N_20066);
nand U20992 (N_20992,N_20275,N_20007);
xnor U20993 (N_20993,N_20343,N_20207);
nand U20994 (N_20994,N_20486,N_20097);
or U20995 (N_20995,N_20414,N_20484);
nor U20996 (N_20996,N_20476,N_20338);
nor U20997 (N_20997,N_20018,N_20498);
or U20998 (N_20998,N_20395,N_20237);
or U20999 (N_20999,N_20467,N_20223);
nor U21000 (N_21000,N_20686,N_20935);
and U21001 (N_21001,N_20577,N_20851);
or U21002 (N_21002,N_20683,N_20729);
nand U21003 (N_21003,N_20775,N_20873);
or U21004 (N_21004,N_20774,N_20987);
nor U21005 (N_21005,N_20556,N_20739);
or U21006 (N_21006,N_20822,N_20823);
and U21007 (N_21007,N_20595,N_20842);
nor U21008 (N_21008,N_20985,N_20995);
and U21009 (N_21009,N_20876,N_20703);
xor U21010 (N_21010,N_20788,N_20634);
nand U21011 (N_21011,N_20535,N_20777);
xnor U21012 (N_21012,N_20562,N_20812);
nor U21013 (N_21013,N_20815,N_20802);
nand U21014 (N_21014,N_20897,N_20648);
xnor U21015 (N_21015,N_20704,N_20807);
nand U21016 (N_21016,N_20869,N_20701);
and U21017 (N_21017,N_20772,N_20982);
and U21018 (N_21018,N_20708,N_20500);
nor U21019 (N_21019,N_20575,N_20814);
nand U21020 (N_21020,N_20790,N_20916);
nand U21021 (N_21021,N_20921,N_20994);
xor U21022 (N_21022,N_20793,N_20977);
nand U21023 (N_21023,N_20817,N_20714);
or U21024 (N_21024,N_20555,N_20620);
and U21025 (N_21025,N_20863,N_20549);
nor U21026 (N_21026,N_20796,N_20617);
or U21027 (N_21027,N_20780,N_20972);
and U21028 (N_21028,N_20637,N_20606);
nand U21029 (N_21029,N_20582,N_20888);
nand U21030 (N_21030,N_20861,N_20874);
or U21031 (N_21031,N_20760,N_20502);
and U21032 (N_21032,N_20964,N_20924);
or U21033 (N_21033,N_20587,N_20979);
and U21034 (N_21034,N_20510,N_20532);
xor U21035 (N_21035,N_20955,N_20651);
or U21036 (N_21036,N_20682,N_20635);
nor U21037 (N_21037,N_20693,N_20768);
nand U21038 (N_21038,N_20834,N_20759);
and U21039 (N_21039,N_20737,N_20613);
nor U21040 (N_21040,N_20854,N_20791);
nor U21041 (N_21041,N_20557,N_20969);
xor U21042 (N_21042,N_20545,N_20699);
or U21043 (N_21043,N_20709,N_20917);
and U21044 (N_21044,N_20561,N_20801);
nor U21045 (N_21045,N_20860,N_20521);
xor U21046 (N_21046,N_20622,N_20731);
xnor U21047 (N_21047,N_20586,N_20734);
nand U21048 (N_21048,N_20886,N_20929);
xor U21049 (N_21049,N_20570,N_20804);
xor U21050 (N_21050,N_20836,N_20880);
nand U21051 (N_21051,N_20903,N_20781);
nand U21052 (N_21052,N_20654,N_20517);
and U21053 (N_21053,N_20677,N_20710);
nor U21054 (N_21054,N_20787,N_20938);
xnor U21055 (N_21055,N_20658,N_20685);
and U21056 (N_21056,N_20958,N_20576);
xor U21057 (N_21057,N_20928,N_20741);
nor U21058 (N_21058,N_20516,N_20852);
nand U21059 (N_21059,N_20689,N_20945);
and U21060 (N_21060,N_20946,N_20883);
or U21061 (N_21061,N_20809,N_20800);
xor U21062 (N_21062,N_20831,N_20980);
nand U21063 (N_21063,N_20891,N_20999);
xnor U21064 (N_21064,N_20871,N_20530);
nand U21065 (N_21065,N_20782,N_20757);
nand U21066 (N_21066,N_20910,N_20642);
nor U21067 (N_21067,N_20653,N_20966);
xnor U21068 (N_21068,N_20518,N_20858);
and U21069 (N_21069,N_20813,N_20771);
and U21070 (N_21070,N_20625,N_20738);
nor U21071 (N_21071,N_20748,N_20660);
nor U21072 (N_21072,N_20553,N_20845);
and U21073 (N_21073,N_20566,N_20519);
xor U21074 (N_21074,N_20743,N_20909);
nand U21075 (N_21075,N_20522,N_20536);
xnor U21076 (N_21076,N_20592,N_20616);
and U21077 (N_21077,N_20922,N_20583);
xor U21078 (N_21078,N_20900,N_20511);
and U21079 (N_21079,N_20914,N_20661);
xor U21080 (N_21080,N_20630,N_20712);
nor U21081 (N_21081,N_20786,N_20546);
nand U21082 (N_21082,N_20855,N_20572);
xnor U21083 (N_21083,N_20636,N_20803);
and U21084 (N_21084,N_20565,N_20941);
nor U21085 (N_21085,N_20974,N_20758);
or U21086 (N_21086,N_20794,N_20749);
nand U21087 (N_21087,N_20767,N_20605);
nand U21088 (N_21088,N_20618,N_20829);
and U21089 (N_21089,N_20779,N_20621);
nand U21090 (N_21090,N_20598,N_20992);
nand U21091 (N_21091,N_20745,N_20652);
xor U21092 (N_21092,N_20765,N_20944);
and U21093 (N_21093,N_20655,N_20720);
nor U21094 (N_21094,N_20906,N_20997);
nand U21095 (N_21095,N_20911,N_20872);
or U21096 (N_21096,N_20590,N_20918);
and U21097 (N_21097,N_20523,N_20819);
nor U21098 (N_21098,N_20976,N_20559);
xnor U21099 (N_21099,N_20789,N_20931);
or U21100 (N_21100,N_20600,N_20956);
or U21101 (N_21101,N_20848,N_20747);
xor U21102 (N_21102,N_20970,N_20730);
nor U21103 (N_21103,N_20627,N_20604);
xor U21104 (N_21104,N_20593,N_20965);
xor U21105 (N_21105,N_20534,N_20681);
or U21106 (N_21106,N_20769,N_20713);
or U21107 (N_21107,N_20707,N_20609);
nand U21108 (N_21108,N_20671,N_20948);
nor U21109 (N_21109,N_20614,N_20908);
xor U21110 (N_21110,N_20702,N_20742);
or U21111 (N_21111,N_20950,N_20665);
xnor U21112 (N_21112,N_20889,N_20875);
or U21113 (N_21113,N_20723,N_20878);
and U21114 (N_21114,N_20961,N_20727);
xor U21115 (N_21115,N_20988,N_20859);
nor U21116 (N_21116,N_20744,N_20513);
nor U21117 (N_21117,N_20694,N_20962);
and U21118 (N_21118,N_20646,N_20560);
nand U21119 (N_21119,N_20773,N_20752);
or U21120 (N_21120,N_20993,N_20514);
or U21121 (N_21121,N_20700,N_20501);
or U21122 (N_21122,N_20567,N_20968);
or U21123 (N_21123,N_20507,N_20971);
and U21124 (N_21124,N_20776,N_20608);
xor U21125 (N_21125,N_20890,N_20839);
nor U21126 (N_21126,N_20877,N_20750);
xnor U21127 (N_21127,N_20597,N_20864);
nand U21128 (N_21128,N_20862,N_20715);
nand U21129 (N_21129,N_20571,N_20824);
nor U21130 (N_21130,N_20520,N_20659);
or U21131 (N_21131,N_20975,N_20939);
and U21132 (N_21132,N_20850,N_20662);
xor U21133 (N_21133,N_20695,N_20755);
xor U21134 (N_21134,N_20996,N_20509);
nand U21135 (N_21135,N_20797,N_20675);
or U21136 (N_21136,N_20547,N_20647);
nor U21137 (N_21137,N_20746,N_20936);
nand U21138 (N_21138,N_20603,N_20952);
xor U21139 (N_21139,N_20882,N_20820);
xor U21140 (N_21140,N_20633,N_20933);
nand U21141 (N_21141,N_20692,N_20830);
nor U21142 (N_21142,N_20960,N_20624);
and U21143 (N_21143,N_20816,N_20940);
xor U21144 (N_21144,N_20973,N_20825);
nand U21145 (N_21145,N_20806,N_20934);
or U21146 (N_21146,N_20528,N_20919);
or U21147 (N_21147,N_20687,N_20649);
and U21148 (N_21148,N_20684,N_20574);
xnor U21149 (N_21149,N_20601,N_20548);
and U21150 (N_21150,N_20542,N_20515);
xnor U21151 (N_21151,N_20539,N_20896);
nand U21152 (N_21152,N_20953,N_20835);
or U21153 (N_21153,N_20963,N_20912);
and U21154 (N_21154,N_20725,N_20990);
or U21155 (N_21155,N_20833,N_20674);
nor U21156 (N_21156,N_20766,N_20881);
xnor U21157 (N_21157,N_20778,N_20599);
and U21158 (N_21158,N_20923,N_20808);
nand U21159 (N_21159,N_20657,N_20696);
xor U21160 (N_21160,N_20641,N_20672);
nor U21161 (N_21161,N_20615,N_20705);
nand U21162 (N_21162,N_20623,N_20638);
or U21163 (N_21163,N_20679,N_20949);
or U21164 (N_21164,N_20650,N_20524);
xor U21165 (N_21165,N_20721,N_20552);
or U21166 (N_21166,N_20763,N_20884);
or U21167 (N_21167,N_20591,N_20895);
or U21168 (N_21168,N_20792,N_20733);
xor U21169 (N_21169,N_20840,N_20538);
nor U21170 (N_21170,N_20826,N_20865);
nand U21171 (N_21171,N_20740,N_20664);
nor U21172 (N_21172,N_20920,N_20680);
or U21173 (N_21173,N_20558,N_20785);
nand U21174 (N_21174,N_20578,N_20942);
or U21175 (N_21175,N_20619,N_20991);
xor U21176 (N_21176,N_20540,N_20887);
nand U21177 (N_21177,N_20588,N_20580);
xor U21178 (N_21178,N_20818,N_20579);
and U21179 (N_21179,N_20899,N_20879);
or U21180 (N_21180,N_20525,N_20736);
xnor U21181 (N_21181,N_20596,N_20563);
or U21182 (N_21182,N_20554,N_20568);
nor U21183 (N_21183,N_20584,N_20867);
nor U21184 (N_21184,N_20629,N_20989);
xnor U21185 (N_21185,N_20676,N_20645);
nand U21186 (N_21186,N_20898,N_20986);
and U21187 (N_21187,N_20810,N_20569);
and U21188 (N_21188,N_20951,N_20508);
nor U21189 (N_21189,N_20644,N_20663);
and U21190 (N_21190,N_20668,N_20849);
xor U21191 (N_21191,N_20504,N_20706);
xor U21192 (N_21192,N_20550,N_20904);
nor U21193 (N_21193,N_20902,N_20581);
nand U21194 (N_21194,N_20711,N_20954);
or U21195 (N_21195,N_20784,N_20512);
nor U21196 (N_21196,N_20602,N_20631);
nor U21197 (N_21197,N_20527,N_20957);
or U21198 (N_21198,N_20719,N_20856);
xor U21199 (N_21199,N_20640,N_20594);
nand U21200 (N_21200,N_20844,N_20998);
or U21201 (N_21201,N_20892,N_20959);
xor U21202 (N_21202,N_20698,N_20901);
or U21203 (N_21203,N_20632,N_20841);
nor U21204 (N_21204,N_20503,N_20761);
xor U21205 (N_21205,N_20506,N_20837);
nand U21206 (N_21206,N_20827,N_20915);
nand U21207 (N_21207,N_20905,N_20610);
nor U21208 (N_21208,N_20543,N_20930);
or U21209 (N_21209,N_20564,N_20531);
nor U21210 (N_21210,N_20691,N_20770);
and U21211 (N_21211,N_20756,N_20795);
xor U21212 (N_21212,N_20893,N_20639);
nand U21213 (N_21213,N_20868,N_20667);
nand U21214 (N_21214,N_20754,N_20870);
nand U21215 (N_21215,N_20724,N_20533);
nand U21216 (N_21216,N_20716,N_20798);
or U21217 (N_21217,N_20811,N_20983);
nor U21218 (N_21218,N_20669,N_20753);
nand U21219 (N_21219,N_20947,N_20678);
nor U21220 (N_21220,N_20762,N_20937);
or U21221 (N_21221,N_20732,N_20894);
nor U21222 (N_21222,N_20828,N_20673);
or U21223 (N_21223,N_20666,N_20735);
xnor U21224 (N_21224,N_20670,N_20541);
xnor U21225 (N_21225,N_20907,N_20529);
or U21226 (N_21226,N_20611,N_20926);
or U21227 (N_21227,N_20656,N_20726);
nor U21228 (N_21228,N_20607,N_20751);
or U21229 (N_21229,N_20967,N_20626);
nand U21230 (N_21230,N_20857,N_20913);
nor U21231 (N_21231,N_20832,N_20526);
xnor U21232 (N_21232,N_20589,N_20612);
or U21233 (N_21233,N_20838,N_20925);
or U21234 (N_21234,N_20847,N_20573);
xnor U21235 (N_21235,N_20764,N_20551);
nor U21236 (N_21236,N_20843,N_20805);
nand U21237 (N_21237,N_20783,N_20537);
nand U21238 (N_21238,N_20697,N_20505);
nand U21239 (N_21239,N_20688,N_20690);
or U21240 (N_21240,N_20718,N_20628);
nor U21241 (N_21241,N_20585,N_20981);
nand U21242 (N_21242,N_20866,N_20932);
nor U21243 (N_21243,N_20728,N_20722);
and U21244 (N_21244,N_20885,N_20821);
nand U21245 (N_21245,N_20846,N_20978);
and U21246 (N_21246,N_20984,N_20927);
nor U21247 (N_21247,N_20643,N_20799);
and U21248 (N_21248,N_20717,N_20943);
or U21249 (N_21249,N_20544,N_20853);
nor U21250 (N_21250,N_20965,N_20940);
or U21251 (N_21251,N_20874,N_20872);
nand U21252 (N_21252,N_20902,N_20593);
nor U21253 (N_21253,N_20946,N_20942);
xor U21254 (N_21254,N_20591,N_20568);
nor U21255 (N_21255,N_20844,N_20552);
nand U21256 (N_21256,N_20651,N_20999);
nand U21257 (N_21257,N_20512,N_20780);
or U21258 (N_21258,N_20706,N_20983);
xor U21259 (N_21259,N_20932,N_20721);
and U21260 (N_21260,N_20676,N_20565);
and U21261 (N_21261,N_20687,N_20603);
nand U21262 (N_21262,N_20628,N_20567);
and U21263 (N_21263,N_20856,N_20635);
or U21264 (N_21264,N_20829,N_20776);
and U21265 (N_21265,N_20788,N_20770);
nor U21266 (N_21266,N_20763,N_20553);
xnor U21267 (N_21267,N_20510,N_20737);
or U21268 (N_21268,N_20550,N_20526);
nor U21269 (N_21269,N_20651,N_20831);
nor U21270 (N_21270,N_20701,N_20690);
xnor U21271 (N_21271,N_20697,N_20729);
xnor U21272 (N_21272,N_20837,N_20905);
or U21273 (N_21273,N_20558,N_20896);
nor U21274 (N_21274,N_20577,N_20894);
and U21275 (N_21275,N_20953,N_20910);
and U21276 (N_21276,N_20559,N_20852);
or U21277 (N_21277,N_20609,N_20899);
nand U21278 (N_21278,N_20694,N_20558);
xor U21279 (N_21279,N_20733,N_20974);
or U21280 (N_21280,N_20804,N_20977);
xnor U21281 (N_21281,N_20856,N_20731);
nor U21282 (N_21282,N_20852,N_20647);
and U21283 (N_21283,N_20839,N_20994);
nor U21284 (N_21284,N_20797,N_20968);
and U21285 (N_21285,N_20774,N_20519);
and U21286 (N_21286,N_20700,N_20511);
nor U21287 (N_21287,N_20698,N_20729);
xor U21288 (N_21288,N_20935,N_20732);
xor U21289 (N_21289,N_20703,N_20761);
and U21290 (N_21290,N_20653,N_20576);
xor U21291 (N_21291,N_20781,N_20841);
nor U21292 (N_21292,N_20792,N_20611);
nor U21293 (N_21293,N_20909,N_20581);
and U21294 (N_21294,N_20525,N_20808);
nand U21295 (N_21295,N_20560,N_20576);
xor U21296 (N_21296,N_20751,N_20513);
or U21297 (N_21297,N_20923,N_20914);
or U21298 (N_21298,N_20694,N_20647);
and U21299 (N_21299,N_20990,N_20910);
nand U21300 (N_21300,N_20988,N_20743);
nor U21301 (N_21301,N_20546,N_20886);
or U21302 (N_21302,N_20547,N_20827);
nand U21303 (N_21303,N_20620,N_20992);
or U21304 (N_21304,N_20501,N_20636);
and U21305 (N_21305,N_20899,N_20682);
or U21306 (N_21306,N_20606,N_20946);
or U21307 (N_21307,N_20984,N_20582);
and U21308 (N_21308,N_20804,N_20611);
xnor U21309 (N_21309,N_20943,N_20904);
or U21310 (N_21310,N_20753,N_20860);
nor U21311 (N_21311,N_20874,N_20783);
and U21312 (N_21312,N_20650,N_20734);
and U21313 (N_21313,N_20752,N_20860);
nand U21314 (N_21314,N_20988,N_20787);
nor U21315 (N_21315,N_20960,N_20843);
nand U21316 (N_21316,N_20578,N_20790);
xnor U21317 (N_21317,N_20852,N_20864);
xor U21318 (N_21318,N_20728,N_20996);
nand U21319 (N_21319,N_20932,N_20642);
nand U21320 (N_21320,N_20791,N_20664);
or U21321 (N_21321,N_20958,N_20654);
nand U21322 (N_21322,N_20772,N_20541);
and U21323 (N_21323,N_20975,N_20960);
nor U21324 (N_21324,N_20670,N_20932);
or U21325 (N_21325,N_20565,N_20973);
nor U21326 (N_21326,N_20774,N_20602);
or U21327 (N_21327,N_20990,N_20956);
nor U21328 (N_21328,N_20752,N_20642);
nand U21329 (N_21329,N_20920,N_20509);
xor U21330 (N_21330,N_20793,N_20581);
xnor U21331 (N_21331,N_20684,N_20757);
xor U21332 (N_21332,N_20613,N_20933);
and U21333 (N_21333,N_20662,N_20867);
xnor U21334 (N_21334,N_20614,N_20667);
nand U21335 (N_21335,N_20941,N_20647);
or U21336 (N_21336,N_20903,N_20820);
or U21337 (N_21337,N_20703,N_20962);
and U21338 (N_21338,N_20663,N_20650);
xor U21339 (N_21339,N_20871,N_20843);
nor U21340 (N_21340,N_20940,N_20764);
and U21341 (N_21341,N_20931,N_20956);
nor U21342 (N_21342,N_20710,N_20748);
xnor U21343 (N_21343,N_20625,N_20578);
nor U21344 (N_21344,N_20988,N_20881);
xor U21345 (N_21345,N_20741,N_20836);
nand U21346 (N_21346,N_20787,N_20756);
nand U21347 (N_21347,N_20965,N_20885);
or U21348 (N_21348,N_20941,N_20963);
xor U21349 (N_21349,N_20874,N_20752);
nand U21350 (N_21350,N_20926,N_20861);
nand U21351 (N_21351,N_20550,N_20838);
or U21352 (N_21352,N_20870,N_20769);
and U21353 (N_21353,N_20954,N_20975);
or U21354 (N_21354,N_20619,N_20974);
and U21355 (N_21355,N_20835,N_20803);
xnor U21356 (N_21356,N_20728,N_20531);
xnor U21357 (N_21357,N_20630,N_20639);
nor U21358 (N_21358,N_20669,N_20852);
nor U21359 (N_21359,N_20978,N_20506);
and U21360 (N_21360,N_20858,N_20614);
and U21361 (N_21361,N_20823,N_20601);
xnor U21362 (N_21362,N_20698,N_20970);
xor U21363 (N_21363,N_20549,N_20980);
nand U21364 (N_21364,N_20854,N_20530);
nand U21365 (N_21365,N_20926,N_20901);
and U21366 (N_21366,N_20943,N_20888);
and U21367 (N_21367,N_20881,N_20791);
nor U21368 (N_21368,N_20559,N_20784);
xnor U21369 (N_21369,N_20582,N_20708);
nand U21370 (N_21370,N_20804,N_20871);
nor U21371 (N_21371,N_20776,N_20710);
and U21372 (N_21372,N_20740,N_20507);
xnor U21373 (N_21373,N_20962,N_20827);
and U21374 (N_21374,N_20842,N_20711);
and U21375 (N_21375,N_20897,N_20761);
nor U21376 (N_21376,N_20680,N_20942);
and U21377 (N_21377,N_20509,N_20814);
nor U21378 (N_21378,N_20517,N_20648);
xnor U21379 (N_21379,N_20922,N_20752);
and U21380 (N_21380,N_20882,N_20909);
and U21381 (N_21381,N_20906,N_20739);
nor U21382 (N_21382,N_20944,N_20911);
nor U21383 (N_21383,N_20677,N_20621);
xor U21384 (N_21384,N_20688,N_20524);
nor U21385 (N_21385,N_20813,N_20632);
and U21386 (N_21386,N_20679,N_20981);
xnor U21387 (N_21387,N_20838,N_20776);
xnor U21388 (N_21388,N_20997,N_20656);
or U21389 (N_21389,N_20855,N_20994);
xor U21390 (N_21390,N_20949,N_20894);
nor U21391 (N_21391,N_20521,N_20558);
and U21392 (N_21392,N_20989,N_20700);
and U21393 (N_21393,N_20884,N_20809);
or U21394 (N_21394,N_20957,N_20562);
nand U21395 (N_21395,N_20630,N_20802);
or U21396 (N_21396,N_20618,N_20603);
nor U21397 (N_21397,N_20579,N_20919);
nand U21398 (N_21398,N_20689,N_20661);
nand U21399 (N_21399,N_20566,N_20717);
and U21400 (N_21400,N_20845,N_20737);
and U21401 (N_21401,N_20523,N_20959);
xor U21402 (N_21402,N_20602,N_20809);
and U21403 (N_21403,N_20757,N_20645);
or U21404 (N_21404,N_20737,N_20935);
or U21405 (N_21405,N_20853,N_20736);
or U21406 (N_21406,N_20538,N_20803);
nor U21407 (N_21407,N_20510,N_20719);
and U21408 (N_21408,N_20530,N_20535);
xor U21409 (N_21409,N_20853,N_20979);
or U21410 (N_21410,N_20567,N_20542);
nand U21411 (N_21411,N_20639,N_20866);
nor U21412 (N_21412,N_20519,N_20908);
or U21413 (N_21413,N_20531,N_20856);
and U21414 (N_21414,N_20621,N_20737);
or U21415 (N_21415,N_20737,N_20819);
nand U21416 (N_21416,N_20858,N_20812);
nand U21417 (N_21417,N_20651,N_20847);
or U21418 (N_21418,N_20862,N_20719);
nor U21419 (N_21419,N_20775,N_20966);
xnor U21420 (N_21420,N_20797,N_20507);
nand U21421 (N_21421,N_20638,N_20504);
nand U21422 (N_21422,N_20601,N_20912);
nor U21423 (N_21423,N_20588,N_20974);
or U21424 (N_21424,N_20858,N_20674);
and U21425 (N_21425,N_20992,N_20875);
and U21426 (N_21426,N_20870,N_20920);
nand U21427 (N_21427,N_20911,N_20884);
or U21428 (N_21428,N_20792,N_20956);
xnor U21429 (N_21429,N_20537,N_20837);
nand U21430 (N_21430,N_20958,N_20704);
and U21431 (N_21431,N_20805,N_20504);
nor U21432 (N_21432,N_20743,N_20891);
xor U21433 (N_21433,N_20668,N_20569);
nor U21434 (N_21434,N_20714,N_20602);
xor U21435 (N_21435,N_20600,N_20889);
or U21436 (N_21436,N_20658,N_20841);
and U21437 (N_21437,N_20800,N_20689);
or U21438 (N_21438,N_20750,N_20932);
nor U21439 (N_21439,N_20755,N_20592);
or U21440 (N_21440,N_20836,N_20528);
xor U21441 (N_21441,N_20937,N_20983);
xnor U21442 (N_21442,N_20991,N_20696);
nor U21443 (N_21443,N_20930,N_20672);
and U21444 (N_21444,N_20535,N_20585);
and U21445 (N_21445,N_20839,N_20621);
xnor U21446 (N_21446,N_20876,N_20603);
and U21447 (N_21447,N_20639,N_20602);
and U21448 (N_21448,N_20629,N_20912);
xnor U21449 (N_21449,N_20506,N_20975);
nor U21450 (N_21450,N_20873,N_20721);
and U21451 (N_21451,N_20857,N_20527);
xor U21452 (N_21452,N_20945,N_20619);
and U21453 (N_21453,N_20694,N_20873);
or U21454 (N_21454,N_20957,N_20809);
nor U21455 (N_21455,N_20665,N_20501);
and U21456 (N_21456,N_20684,N_20619);
or U21457 (N_21457,N_20934,N_20607);
xnor U21458 (N_21458,N_20762,N_20688);
nand U21459 (N_21459,N_20670,N_20793);
or U21460 (N_21460,N_20960,N_20503);
xor U21461 (N_21461,N_20587,N_20618);
or U21462 (N_21462,N_20988,N_20765);
nor U21463 (N_21463,N_20937,N_20651);
nor U21464 (N_21464,N_20547,N_20900);
nor U21465 (N_21465,N_20633,N_20543);
or U21466 (N_21466,N_20509,N_20955);
and U21467 (N_21467,N_20726,N_20568);
xnor U21468 (N_21468,N_20588,N_20968);
nand U21469 (N_21469,N_20551,N_20745);
xnor U21470 (N_21470,N_20561,N_20730);
nand U21471 (N_21471,N_20829,N_20750);
nand U21472 (N_21472,N_20986,N_20526);
nor U21473 (N_21473,N_20741,N_20777);
nor U21474 (N_21474,N_20943,N_20500);
and U21475 (N_21475,N_20809,N_20720);
and U21476 (N_21476,N_20669,N_20706);
nor U21477 (N_21477,N_20952,N_20589);
nor U21478 (N_21478,N_20862,N_20759);
xor U21479 (N_21479,N_20719,N_20953);
nand U21480 (N_21480,N_20611,N_20551);
or U21481 (N_21481,N_20517,N_20813);
nand U21482 (N_21482,N_20779,N_20515);
and U21483 (N_21483,N_20548,N_20527);
nand U21484 (N_21484,N_20776,N_20933);
nand U21485 (N_21485,N_20885,N_20765);
nor U21486 (N_21486,N_20732,N_20790);
nor U21487 (N_21487,N_20907,N_20676);
or U21488 (N_21488,N_20640,N_20510);
xnor U21489 (N_21489,N_20584,N_20585);
or U21490 (N_21490,N_20582,N_20742);
or U21491 (N_21491,N_20997,N_20994);
or U21492 (N_21492,N_20709,N_20614);
and U21493 (N_21493,N_20982,N_20580);
or U21494 (N_21494,N_20529,N_20762);
or U21495 (N_21495,N_20590,N_20722);
nor U21496 (N_21496,N_20839,N_20730);
xnor U21497 (N_21497,N_20855,N_20675);
or U21498 (N_21498,N_20895,N_20638);
nor U21499 (N_21499,N_20738,N_20886);
or U21500 (N_21500,N_21050,N_21000);
nor U21501 (N_21501,N_21248,N_21081);
or U21502 (N_21502,N_21013,N_21322);
and U21503 (N_21503,N_21175,N_21225);
xor U21504 (N_21504,N_21121,N_21386);
nor U21505 (N_21505,N_21069,N_21339);
xnor U21506 (N_21506,N_21015,N_21398);
and U21507 (N_21507,N_21369,N_21291);
or U21508 (N_21508,N_21349,N_21469);
and U21509 (N_21509,N_21003,N_21061);
and U21510 (N_21510,N_21303,N_21265);
nor U21511 (N_21511,N_21337,N_21222);
xor U21512 (N_21512,N_21362,N_21219);
and U21513 (N_21513,N_21004,N_21371);
xor U21514 (N_21514,N_21320,N_21016);
nor U21515 (N_21515,N_21131,N_21007);
nand U21516 (N_21516,N_21193,N_21101);
xnor U21517 (N_21517,N_21278,N_21289);
or U21518 (N_21518,N_21318,N_21251);
or U21519 (N_21519,N_21275,N_21042);
nor U21520 (N_21520,N_21233,N_21305);
and U21521 (N_21521,N_21370,N_21238);
or U21522 (N_21522,N_21394,N_21208);
xor U21523 (N_21523,N_21221,N_21209);
nand U21524 (N_21524,N_21354,N_21380);
and U21525 (N_21525,N_21206,N_21237);
nor U21526 (N_21526,N_21105,N_21342);
and U21527 (N_21527,N_21256,N_21145);
or U21528 (N_21528,N_21249,N_21134);
and U21529 (N_21529,N_21123,N_21387);
nand U21530 (N_21530,N_21276,N_21325);
or U21531 (N_21531,N_21491,N_21189);
or U21532 (N_21532,N_21271,N_21070);
nand U21533 (N_21533,N_21396,N_21176);
nand U21534 (N_21534,N_21058,N_21299);
nand U21535 (N_21535,N_21037,N_21292);
or U21536 (N_21536,N_21444,N_21281);
nor U21537 (N_21537,N_21467,N_21104);
and U21538 (N_21538,N_21122,N_21077);
or U21539 (N_21539,N_21462,N_21019);
or U21540 (N_21540,N_21112,N_21253);
and U21541 (N_21541,N_21190,N_21470);
xor U21542 (N_21542,N_21002,N_21096);
nand U21543 (N_21543,N_21451,N_21199);
nand U21544 (N_21544,N_21423,N_21492);
xnor U21545 (N_21545,N_21267,N_21164);
nor U21546 (N_21546,N_21018,N_21067);
nor U21547 (N_21547,N_21390,N_21376);
nand U21548 (N_21548,N_21202,N_21167);
xnor U21549 (N_21549,N_21383,N_21316);
nand U21550 (N_21550,N_21433,N_21029);
nand U21551 (N_21551,N_21187,N_21283);
and U21552 (N_21552,N_21153,N_21051);
nor U21553 (N_21553,N_21488,N_21047);
or U21554 (N_21554,N_21389,N_21413);
nor U21555 (N_21555,N_21140,N_21288);
or U21556 (N_21556,N_21091,N_21473);
nand U21557 (N_21557,N_21118,N_21446);
or U21558 (N_21558,N_21100,N_21461);
nand U21559 (N_21559,N_21268,N_21310);
xor U21560 (N_21560,N_21366,N_21098);
or U21561 (N_21561,N_21132,N_21054);
nor U21562 (N_21562,N_21409,N_21165);
and U21563 (N_21563,N_21186,N_21447);
nand U21564 (N_21564,N_21484,N_21162);
xor U21565 (N_21565,N_21106,N_21391);
nor U21566 (N_21566,N_21232,N_21368);
xnor U21567 (N_21567,N_21177,N_21143);
or U21568 (N_21568,N_21308,N_21043);
nand U21569 (N_21569,N_21490,N_21057);
nor U21570 (N_21570,N_21319,N_21372);
nand U21571 (N_21571,N_21163,N_21374);
nand U21572 (N_21572,N_21393,N_21453);
or U21573 (N_21573,N_21068,N_21183);
nand U21574 (N_21574,N_21297,N_21378);
nor U21575 (N_21575,N_21156,N_21420);
nor U21576 (N_21576,N_21180,N_21464);
nand U21577 (N_21577,N_21139,N_21185);
and U21578 (N_21578,N_21345,N_21152);
nand U21579 (N_21579,N_21330,N_21290);
xor U21580 (N_21580,N_21487,N_21463);
nor U21581 (N_21581,N_21023,N_21410);
nor U21582 (N_21582,N_21381,N_21363);
xnor U21583 (N_21583,N_21338,N_21294);
nand U21584 (N_21584,N_21382,N_21074);
or U21585 (N_21585,N_21497,N_21472);
or U21586 (N_21586,N_21264,N_21195);
nor U21587 (N_21587,N_21111,N_21135);
nand U21588 (N_21588,N_21073,N_21173);
and U21589 (N_21589,N_21129,N_21483);
nand U21590 (N_21590,N_21244,N_21486);
nor U21591 (N_21591,N_21107,N_21441);
xnor U21592 (N_21592,N_21285,N_21109);
and U21593 (N_21593,N_21346,N_21242);
xnor U21594 (N_21594,N_21332,N_21422);
nor U21595 (N_21595,N_21060,N_21343);
nand U21596 (N_21596,N_21494,N_21384);
and U21597 (N_21597,N_21099,N_21204);
nor U21598 (N_21598,N_21009,N_21127);
xor U21599 (N_21599,N_21026,N_21427);
xor U21600 (N_21600,N_21076,N_21336);
and U21601 (N_21601,N_21226,N_21030);
nand U21602 (N_21602,N_21352,N_21149);
nor U21603 (N_21603,N_21179,N_21459);
nor U21604 (N_21604,N_21207,N_21457);
nor U21605 (N_21605,N_21412,N_21033);
or U21606 (N_21606,N_21090,N_21010);
and U21607 (N_21607,N_21089,N_21216);
and U21608 (N_21608,N_21421,N_21194);
xnor U21609 (N_21609,N_21182,N_21357);
or U21610 (N_21610,N_21114,N_21071);
or U21611 (N_21611,N_21450,N_21388);
nor U21612 (N_21612,N_21128,N_21085);
xor U21613 (N_21613,N_21148,N_21498);
nor U21614 (N_21614,N_21306,N_21418);
nor U21615 (N_21615,N_21046,N_21031);
nand U21616 (N_21616,N_21400,N_21203);
nor U21617 (N_21617,N_21240,N_21417);
xnor U21618 (N_21618,N_21373,N_21274);
or U21619 (N_21619,N_21367,N_21228);
or U21620 (N_21620,N_21062,N_21477);
or U21621 (N_21621,N_21399,N_21028);
xor U21622 (N_21622,N_21205,N_21301);
and U21623 (N_21623,N_21088,N_21334);
and U21624 (N_21624,N_21379,N_21136);
and U21625 (N_21625,N_21331,N_21084);
nor U21626 (N_21626,N_21001,N_21231);
xor U21627 (N_21627,N_21113,N_21279);
or U21628 (N_21628,N_21227,N_21375);
or U21629 (N_21629,N_21284,N_21311);
xor U21630 (N_21630,N_21347,N_21474);
nor U21631 (N_21631,N_21430,N_21086);
xor U21632 (N_21632,N_21220,N_21295);
nor U21633 (N_21633,N_21293,N_21055);
nand U21634 (N_21634,N_21272,N_21201);
xor U21635 (N_21635,N_21236,N_21468);
nor U21636 (N_21636,N_21082,N_21150);
nand U21637 (N_21637,N_21261,N_21116);
nor U21638 (N_21638,N_21258,N_21364);
xor U21639 (N_21639,N_21286,N_21321);
nand U21640 (N_21640,N_21198,N_21213);
and U21641 (N_21641,N_21215,N_21138);
nor U21642 (N_21642,N_21260,N_21212);
and U21643 (N_21643,N_21239,N_21166);
nand U21644 (N_21644,N_21020,N_21419);
and U21645 (N_21645,N_21263,N_21200);
nand U21646 (N_21646,N_21171,N_21095);
nor U21647 (N_21647,N_21103,N_21429);
xor U21648 (N_21648,N_21436,N_21063);
nor U21649 (N_21649,N_21155,N_21437);
nand U21650 (N_21650,N_21035,N_21078);
nand U21651 (N_21651,N_21392,N_21426);
and U21652 (N_21652,N_21326,N_21435);
nand U21653 (N_21653,N_21197,N_21277);
or U21654 (N_21654,N_21348,N_21401);
and U21655 (N_21655,N_21097,N_21022);
xnor U21656 (N_21656,N_21353,N_21178);
and U21657 (N_21657,N_21324,N_21270);
nor U21658 (N_21658,N_21328,N_21036);
and U21659 (N_21659,N_21262,N_21048);
and U21660 (N_21660,N_21038,N_21172);
or U21661 (N_21661,N_21287,N_21312);
xor U21662 (N_21662,N_21188,N_21094);
or U21663 (N_21663,N_21146,N_21092);
and U21664 (N_21664,N_21317,N_21191);
nor U21665 (N_21665,N_21025,N_21234);
xor U21666 (N_21666,N_21259,N_21449);
xor U21667 (N_21667,N_21455,N_21170);
and U21668 (N_21668,N_21224,N_21014);
xnor U21669 (N_21669,N_21385,N_21458);
nor U21670 (N_21670,N_21083,N_21255);
xor U21671 (N_21671,N_21159,N_21452);
and U21672 (N_21672,N_21425,N_21323);
nor U21673 (N_21673,N_21137,N_21117);
xnor U21674 (N_21674,N_21245,N_21438);
xor U21675 (N_21675,N_21456,N_21360);
or U21676 (N_21676,N_21006,N_21125);
xor U21677 (N_21677,N_21196,N_21169);
and U21678 (N_21678,N_21223,N_21499);
xnor U21679 (N_21679,N_21493,N_21160);
or U21680 (N_21680,N_21482,N_21039);
or U21681 (N_21681,N_21307,N_21478);
nor U21682 (N_21682,N_21314,N_21102);
or U21683 (N_21683,N_21126,N_21230);
xnor U21684 (N_21684,N_21056,N_21415);
nor U21685 (N_21685,N_21243,N_21174);
xnor U21686 (N_21686,N_21403,N_21327);
nor U21687 (N_21687,N_21049,N_21355);
nor U21688 (N_21688,N_21075,N_21108);
or U21689 (N_21689,N_21133,N_21481);
nand U21690 (N_21690,N_21034,N_21309);
nand U21691 (N_21691,N_21157,N_21066);
xor U21692 (N_21692,N_21405,N_21141);
nor U21693 (N_21693,N_21021,N_21431);
and U21694 (N_21694,N_21032,N_21445);
xnor U21695 (N_21695,N_21466,N_21080);
nor U21696 (N_21696,N_21124,N_21340);
and U21697 (N_21697,N_21341,N_21252);
xor U21698 (N_21698,N_21211,N_21300);
nor U21699 (N_21699,N_21052,N_21011);
and U21700 (N_21700,N_21130,N_21296);
or U21701 (N_21701,N_21072,N_21079);
xnor U21702 (N_21702,N_21407,N_21087);
and U21703 (N_21703,N_21440,N_21344);
xnor U21704 (N_21704,N_21465,N_21428);
nor U21705 (N_21705,N_21257,N_21192);
and U21706 (N_21706,N_21110,N_21161);
or U21707 (N_21707,N_21147,N_21280);
nor U21708 (N_21708,N_21335,N_21432);
nand U21709 (N_21709,N_21093,N_21443);
nor U21710 (N_21710,N_21184,N_21214);
nand U21711 (N_21711,N_21005,N_21210);
nor U21712 (N_21712,N_21476,N_21024);
and U21713 (N_21713,N_21304,N_21475);
and U21714 (N_21714,N_21115,N_21246);
or U21715 (N_21715,N_21471,N_21496);
or U21716 (N_21716,N_21142,N_21358);
xor U21717 (N_21717,N_21151,N_21416);
and U21718 (N_21718,N_21064,N_21485);
and U21719 (N_21719,N_21329,N_21424);
xnor U21720 (N_21720,N_21377,N_21313);
nand U21721 (N_21721,N_21008,N_21247);
and U21722 (N_21722,N_21158,N_21442);
and U21723 (N_21723,N_21250,N_21315);
or U21724 (N_21724,N_21448,N_21404);
nand U21725 (N_21725,N_21439,N_21241);
nor U21726 (N_21726,N_21351,N_21012);
nor U21727 (N_21727,N_21411,N_21144);
nor U21728 (N_21728,N_21402,N_21395);
and U21729 (N_21729,N_21269,N_21053);
xnor U21730 (N_21730,N_21480,N_21406);
and U21731 (N_21731,N_21495,N_21365);
nand U21732 (N_21732,N_21040,N_21460);
xor U21733 (N_21733,N_21065,N_21119);
xor U21734 (N_21734,N_21414,N_21059);
and U21735 (N_21735,N_21027,N_21489);
or U21736 (N_21736,N_21408,N_21041);
xor U21737 (N_21737,N_21218,N_21282);
nor U21738 (N_21738,N_21217,N_21479);
or U21739 (N_21739,N_21181,N_21235);
or U21740 (N_21740,N_21229,N_21302);
nor U21741 (N_21741,N_21333,N_21154);
xnor U21742 (N_21742,N_21397,N_21359);
nor U21743 (N_21743,N_21361,N_21044);
nor U21744 (N_21744,N_21350,N_21045);
nand U21745 (N_21745,N_21356,N_21168);
xnor U21746 (N_21746,N_21434,N_21017);
nor U21747 (N_21747,N_21254,N_21454);
and U21748 (N_21748,N_21266,N_21298);
nor U21749 (N_21749,N_21120,N_21273);
xor U21750 (N_21750,N_21206,N_21494);
nor U21751 (N_21751,N_21251,N_21325);
nand U21752 (N_21752,N_21025,N_21080);
nand U21753 (N_21753,N_21045,N_21474);
xnor U21754 (N_21754,N_21114,N_21116);
or U21755 (N_21755,N_21285,N_21090);
or U21756 (N_21756,N_21255,N_21298);
xnor U21757 (N_21757,N_21143,N_21449);
nand U21758 (N_21758,N_21287,N_21425);
xor U21759 (N_21759,N_21493,N_21326);
xnor U21760 (N_21760,N_21293,N_21241);
or U21761 (N_21761,N_21317,N_21166);
xnor U21762 (N_21762,N_21218,N_21060);
nor U21763 (N_21763,N_21118,N_21084);
nand U21764 (N_21764,N_21019,N_21394);
or U21765 (N_21765,N_21241,N_21156);
nand U21766 (N_21766,N_21140,N_21109);
xor U21767 (N_21767,N_21073,N_21316);
nand U21768 (N_21768,N_21258,N_21076);
xor U21769 (N_21769,N_21205,N_21068);
or U21770 (N_21770,N_21397,N_21081);
nor U21771 (N_21771,N_21054,N_21163);
nor U21772 (N_21772,N_21289,N_21480);
and U21773 (N_21773,N_21492,N_21193);
nand U21774 (N_21774,N_21000,N_21119);
and U21775 (N_21775,N_21245,N_21108);
xnor U21776 (N_21776,N_21124,N_21222);
nand U21777 (N_21777,N_21136,N_21257);
or U21778 (N_21778,N_21435,N_21141);
xnor U21779 (N_21779,N_21408,N_21238);
or U21780 (N_21780,N_21261,N_21105);
nand U21781 (N_21781,N_21062,N_21016);
and U21782 (N_21782,N_21092,N_21304);
nand U21783 (N_21783,N_21230,N_21233);
nor U21784 (N_21784,N_21035,N_21010);
nand U21785 (N_21785,N_21285,N_21326);
xnor U21786 (N_21786,N_21378,N_21475);
xor U21787 (N_21787,N_21399,N_21054);
or U21788 (N_21788,N_21135,N_21427);
and U21789 (N_21789,N_21423,N_21201);
nor U21790 (N_21790,N_21003,N_21317);
nand U21791 (N_21791,N_21068,N_21319);
nand U21792 (N_21792,N_21435,N_21101);
nand U21793 (N_21793,N_21234,N_21417);
and U21794 (N_21794,N_21493,N_21203);
nor U21795 (N_21795,N_21111,N_21398);
and U21796 (N_21796,N_21415,N_21123);
nand U21797 (N_21797,N_21388,N_21421);
nand U21798 (N_21798,N_21378,N_21066);
nand U21799 (N_21799,N_21361,N_21422);
xnor U21800 (N_21800,N_21323,N_21043);
nand U21801 (N_21801,N_21386,N_21002);
nor U21802 (N_21802,N_21160,N_21107);
nand U21803 (N_21803,N_21033,N_21030);
nor U21804 (N_21804,N_21033,N_21178);
nand U21805 (N_21805,N_21138,N_21404);
and U21806 (N_21806,N_21188,N_21021);
or U21807 (N_21807,N_21342,N_21421);
nand U21808 (N_21808,N_21040,N_21242);
or U21809 (N_21809,N_21336,N_21131);
nor U21810 (N_21810,N_21219,N_21471);
nor U21811 (N_21811,N_21455,N_21317);
xnor U21812 (N_21812,N_21435,N_21404);
xnor U21813 (N_21813,N_21223,N_21074);
and U21814 (N_21814,N_21075,N_21359);
nand U21815 (N_21815,N_21180,N_21111);
nand U21816 (N_21816,N_21078,N_21294);
xor U21817 (N_21817,N_21401,N_21116);
and U21818 (N_21818,N_21181,N_21152);
or U21819 (N_21819,N_21408,N_21025);
or U21820 (N_21820,N_21488,N_21313);
or U21821 (N_21821,N_21086,N_21255);
nor U21822 (N_21822,N_21243,N_21425);
and U21823 (N_21823,N_21069,N_21189);
nor U21824 (N_21824,N_21300,N_21297);
xor U21825 (N_21825,N_21252,N_21134);
and U21826 (N_21826,N_21445,N_21295);
xor U21827 (N_21827,N_21134,N_21326);
xnor U21828 (N_21828,N_21443,N_21031);
or U21829 (N_21829,N_21188,N_21209);
xnor U21830 (N_21830,N_21356,N_21166);
xnor U21831 (N_21831,N_21218,N_21326);
and U21832 (N_21832,N_21353,N_21078);
and U21833 (N_21833,N_21386,N_21040);
nor U21834 (N_21834,N_21240,N_21173);
nand U21835 (N_21835,N_21421,N_21453);
nand U21836 (N_21836,N_21043,N_21419);
nand U21837 (N_21837,N_21458,N_21136);
nor U21838 (N_21838,N_21459,N_21282);
and U21839 (N_21839,N_21378,N_21015);
nor U21840 (N_21840,N_21452,N_21351);
nand U21841 (N_21841,N_21191,N_21224);
nand U21842 (N_21842,N_21136,N_21365);
nand U21843 (N_21843,N_21135,N_21266);
and U21844 (N_21844,N_21210,N_21010);
nor U21845 (N_21845,N_21265,N_21213);
xor U21846 (N_21846,N_21291,N_21181);
xor U21847 (N_21847,N_21294,N_21059);
nor U21848 (N_21848,N_21044,N_21485);
nand U21849 (N_21849,N_21380,N_21452);
xnor U21850 (N_21850,N_21027,N_21209);
nor U21851 (N_21851,N_21448,N_21011);
or U21852 (N_21852,N_21390,N_21134);
or U21853 (N_21853,N_21325,N_21213);
or U21854 (N_21854,N_21342,N_21253);
nand U21855 (N_21855,N_21144,N_21135);
and U21856 (N_21856,N_21251,N_21010);
xnor U21857 (N_21857,N_21234,N_21180);
or U21858 (N_21858,N_21186,N_21108);
nand U21859 (N_21859,N_21403,N_21499);
or U21860 (N_21860,N_21456,N_21088);
or U21861 (N_21861,N_21322,N_21142);
xor U21862 (N_21862,N_21150,N_21200);
or U21863 (N_21863,N_21256,N_21371);
nand U21864 (N_21864,N_21332,N_21401);
nand U21865 (N_21865,N_21422,N_21174);
nand U21866 (N_21866,N_21493,N_21173);
nand U21867 (N_21867,N_21181,N_21467);
nor U21868 (N_21868,N_21326,N_21406);
nor U21869 (N_21869,N_21471,N_21316);
nor U21870 (N_21870,N_21493,N_21053);
or U21871 (N_21871,N_21035,N_21281);
xnor U21872 (N_21872,N_21140,N_21086);
xnor U21873 (N_21873,N_21361,N_21154);
and U21874 (N_21874,N_21130,N_21196);
xor U21875 (N_21875,N_21467,N_21092);
and U21876 (N_21876,N_21423,N_21310);
nor U21877 (N_21877,N_21251,N_21335);
nand U21878 (N_21878,N_21045,N_21062);
or U21879 (N_21879,N_21024,N_21077);
or U21880 (N_21880,N_21320,N_21092);
or U21881 (N_21881,N_21403,N_21399);
xnor U21882 (N_21882,N_21338,N_21299);
nor U21883 (N_21883,N_21222,N_21052);
or U21884 (N_21884,N_21075,N_21105);
xnor U21885 (N_21885,N_21057,N_21220);
or U21886 (N_21886,N_21378,N_21080);
nand U21887 (N_21887,N_21057,N_21370);
nand U21888 (N_21888,N_21074,N_21243);
nor U21889 (N_21889,N_21381,N_21416);
xor U21890 (N_21890,N_21340,N_21427);
or U21891 (N_21891,N_21386,N_21237);
or U21892 (N_21892,N_21087,N_21017);
xnor U21893 (N_21893,N_21439,N_21385);
and U21894 (N_21894,N_21275,N_21022);
and U21895 (N_21895,N_21208,N_21037);
xor U21896 (N_21896,N_21151,N_21029);
nor U21897 (N_21897,N_21204,N_21102);
nand U21898 (N_21898,N_21026,N_21459);
and U21899 (N_21899,N_21098,N_21019);
nor U21900 (N_21900,N_21239,N_21134);
or U21901 (N_21901,N_21214,N_21388);
nor U21902 (N_21902,N_21023,N_21065);
or U21903 (N_21903,N_21437,N_21153);
and U21904 (N_21904,N_21246,N_21301);
and U21905 (N_21905,N_21178,N_21372);
nor U21906 (N_21906,N_21188,N_21453);
and U21907 (N_21907,N_21317,N_21490);
xor U21908 (N_21908,N_21081,N_21098);
nor U21909 (N_21909,N_21349,N_21146);
xor U21910 (N_21910,N_21124,N_21251);
or U21911 (N_21911,N_21150,N_21167);
nor U21912 (N_21912,N_21420,N_21401);
xor U21913 (N_21913,N_21335,N_21205);
xor U21914 (N_21914,N_21448,N_21399);
and U21915 (N_21915,N_21437,N_21411);
nor U21916 (N_21916,N_21373,N_21148);
nor U21917 (N_21917,N_21396,N_21318);
nor U21918 (N_21918,N_21332,N_21366);
or U21919 (N_21919,N_21041,N_21458);
and U21920 (N_21920,N_21401,N_21151);
xor U21921 (N_21921,N_21387,N_21268);
xor U21922 (N_21922,N_21333,N_21390);
xnor U21923 (N_21923,N_21473,N_21269);
nand U21924 (N_21924,N_21305,N_21450);
nor U21925 (N_21925,N_21051,N_21249);
nor U21926 (N_21926,N_21297,N_21216);
or U21927 (N_21927,N_21156,N_21493);
xnor U21928 (N_21928,N_21437,N_21360);
or U21929 (N_21929,N_21064,N_21414);
xnor U21930 (N_21930,N_21150,N_21398);
or U21931 (N_21931,N_21205,N_21115);
nor U21932 (N_21932,N_21136,N_21303);
and U21933 (N_21933,N_21255,N_21458);
nand U21934 (N_21934,N_21292,N_21036);
xor U21935 (N_21935,N_21083,N_21068);
or U21936 (N_21936,N_21345,N_21320);
and U21937 (N_21937,N_21340,N_21148);
nor U21938 (N_21938,N_21165,N_21416);
nand U21939 (N_21939,N_21461,N_21148);
and U21940 (N_21940,N_21122,N_21183);
nand U21941 (N_21941,N_21406,N_21245);
or U21942 (N_21942,N_21094,N_21330);
and U21943 (N_21943,N_21178,N_21438);
and U21944 (N_21944,N_21146,N_21200);
nor U21945 (N_21945,N_21259,N_21255);
xnor U21946 (N_21946,N_21107,N_21426);
nand U21947 (N_21947,N_21479,N_21292);
xor U21948 (N_21948,N_21408,N_21377);
xnor U21949 (N_21949,N_21212,N_21096);
xor U21950 (N_21950,N_21384,N_21449);
nand U21951 (N_21951,N_21340,N_21070);
and U21952 (N_21952,N_21042,N_21018);
nand U21953 (N_21953,N_21432,N_21019);
xor U21954 (N_21954,N_21471,N_21168);
nor U21955 (N_21955,N_21420,N_21137);
xnor U21956 (N_21956,N_21285,N_21111);
and U21957 (N_21957,N_21465,N_21079);
xnor U21958 (N_21958,N_21029,N_21233);
or U21959 (N_21959,N_21131,N_21347);
and U21960 (N_21960,N_21060,N_21199);
or U21961 (N_21961,N_21373,N_21002);
nor U21962 (N_21962,N_21146,N_21257);
nor U21963 (N_21963,N_21122,N_21385);
nand U21964 (N_21964,N_21203,N_21085);
xnor U21965 (N_21965,N_21172,N_21192);
nor U21966 (N_21966,N_21367,N_21212);
or U21967 (N_21967,N_21319,N_21129);
xnor U21968 (N_21968,N_21207,N_21117);
nand U21969 (N_21969,N_21091,N_21415);
nor U21970 (N_21970,N_21176,N_21462);
nor U21971 (N_21971,N_21027,N_21357);
and U21972 (N_21972,N_21415,N_21031);
nor U21973 (N_21973,N_21333,N_21257);
or U21974 (N_21974,N_21473,N_21159);
nor U21975 (N_21975,N_21134,N_21175);
xor U21976 (N_21976,N_21491,N_21272);
xor U21977 (N_21977,N_21219,N_21436);
and U21978 (N_21978,N_21248,N_21243);
or U21979 (N_21979,N_21150,N_21136);
or U21980 (N_21980,N_21419,N_21402);
and U21981 (N_21981,N_21202,N_21311);
xnor U21982 (N_21982,N_21431,N_21140);
nor U21983 (N_21983,N_21426,N_21394);
nand U21984 (N_21984,N_21076,N_21472);
and U21985 (N_21985,N_21107,N_21097);
nor U21986 (N_21986,N_21169,N_21303);
nand U21987 (N_21987,N_21008,N_21098);
xnor U21988 (N_21988,N_21220,N_21424);
xor U21989 (N_21989,N_21116,N_21472);
nor U21990 (N_21990,N_21402,N_21006);
nand U21991 (N_21991,N_21135,N_21479);
or U21992 (N_21992,N_21178,N_21226);
nor U21993 (N_21993,N_21103,N_21218);
xor U21994 (N_21994,N_21141,N_21456);
xnor U21995 (N_21995,N_21079,N_21039);
and U21996 (N_21996,N_21197,N_21084);
xor U21997 (N_21997,N_21089,N_21021);
nor U21998 (N_21998,N_21353,N_21326);
nor U21999 (N_21999,N_21025,N_21371);
nand U22000 (N_22000,N_21807,N_21700);
and U22001 (N_22001,N_21933,N_21919);
and U22002 (N_22002,N_21934,N_21794);
or U22003 (N_22003,N_21860,N_21792);
nor U22004 (N_22004,N_21721,N_21825);
nor U22005 (N_22005,N_21908,N_21913);
xnor U22006 (N_22006,N_21902,N_21546);
or U22007 (N_22007,N_21517,N_21506);
and U22008 (N_22008,N_21885,N_21570);
nand U22009 (N_22009,N_21750,N_21822);
nand U22010 (N_22010,N_21630,N_21945);
nand U22011 (N_22011,N_21843,N_21552);
or U22012 (N_22012,N_21740,N_21952);
nor U22013 (N_22013,N_21884,N_21817);
and U22014 (N_22014,N_21679,N_21868);
or U22015 (N_22015,N_21767,N_21968);
and U22016 (N_22016,N_21705,N_21521);
nor U22017 (N_22017,N_21670,N_21806);
nor U22018 (N_22018,N_21802,N_21835);
or U22019 (N_22019,N_21882,N_21622);
or U22020 (N_22020,N_21975,N_21924);
xnor U22021 (N_22021,N_21909,N_21739);
and U22022 (N_22022,N_21626,N_21556);
and U22023 (N_22023,N_21980,N_21597);
and U22024 (N_22024,N_21501,N_21810);
xor U22025 (N_22025,N_21805,N_21686);
nor U22026 (N_22026,N_21972,N_21922);
or U22027 (N_22027,N_21808,N_21874);
xnor U22028 (N_22028,N_21624,N_21675);
nor U22029 (N_22029,N_21714,N_21731);
xor U22030 (N_22030,N_21708,N_21821);
and U22031 (N_22031,N_21725,N_21829);
or U22032 (N_22032,N_21666,N_21844);
or U22033 (N_22033,N_21702,N_21949);
nor U22034 (N_22034,N_21512,N_21753);
xor U22035 (N_22035,N_21732,N_21780);
xor U22036 (N_22036,N_21640,N_21538);
nor U22037 (N_22037,N_21967,N_21571);
and U22038 (N_22038,N_21607,N_21848);
or U22039 (N_22039,N_21717,N_21994);
nor U22040 (N_22040,N_21543,N_21923);
xnor U22041 (N_22041,N_21684,N_21921);
and U22042 (N_22042,N_21935,N_21855);
xnor U22043 (N_22043,N_21917,N_21639);
nor U22044 (N_22044,N_21950,N_21859);
nor U22045 (N_22045,N_21761,N_21531);
nor U22046 (N_22046,N_21911,N_21720);
nand U22047 (N_22047,N_21797,N_21615);
or U22048 (N_22048,N_21682,N_21891);
nor U22049 (N_22049,N_21567,N_21759);
or U22050 (N_22050,N_21789,N_21948);
xor U22051 (N_22051,N_21596,N_21937);
nand U22052 (N_22052,N_21943,N_21878);
or U22053 (N_22053,N_21809,N_21611);
xnor U22054 (N_22054,N_21656,N_21778);
xnor U22055 (N_22055,N_21730,N_21991);
and U22056 (N_22056,N_21635,N_21560);
and U22057 (N_22057,N_21602,N_21557);
nand U22058 (N_22058,N_21678,N_21838);
or U22059 (N_22059,N_21779,N_21986);
and U22060 (N_22060,N_21799,N_21654);
or U22061 (N_22061,N_21643,N_21852);
xnor U22062 (N_22062,N_21895,N_21625);
and U22063 (N_22063,N_21790,N_21582);
and U22064 (N_22064,N_21632,N_21513);
nor U22065 (N_22065,N_21925,N_21577);
nor U22066 (N_22066,N_21981,N_21566);
or U22067 (N_22067,N_21604,N_21685);
xor U22068 (N_22068,N_21853,N_21516);
nor U22069 (N_22069,N_21605,N_21926);
or U22070 (N_22070,N_21897,N_21992);
xnor U22071 (N_22071,N_21580,N_21875);
xor U22072 (N_22072,N_21849,N_21774);
and U22073 (N_22073,N_21545,N_21993);
and U22074 (N_22074,N_21770,N_21963);
nand U22075 (N_22075,N_21742,N_21827);
and U22076 (N_22076,N_21763,N_21573);
xnor U22077 (N_22077,N_21932,N_21749);
xor U22078 (N_22078,N_21649,N_21524);
nor U22079 (N_22079,N_21627,N_21757);
nand U22080 (N_22080,N_21520,N_21550);
or U22081 (N_22081,N_21508,N_21811);
nor U22082 (N_22082,N_21762,N_21578);
nand U22083 (N_22083,N_21969,N_21561);
nand U22084 (N_22084,N_21652,N_21540);
or U22085 (N_22085,N_21549,N_21537);
nor U22086 (N_22086,N_21965,N_21856);
xnor U22087 (N_22087,N_21687,N_21928);
xor U22088 (N_22088,N_21547,N_21947);
nor U22089 (N_22089,N_21648,N_21696);
or U22090 (N_22090,N_21754,N_21974);
nand U22091 (N_22091,N_21500,N_21766);
nand U22092 (N_22092,N_21608,N_21515);
and U22093 (N_22093,N_21988,N_21523);
or U22094 (N_22094,N_21833,N_21503);
nor U22095 (N_22095,N_21544,N_21658);
xnor U22096 (N_22096,N_21970,N_21647);
nor U22097 (N_22097,N_21709,N_21502);
and U22098 (N_22098,N_21959,N_21715);
nor U22099 (N_22099,N_21772,N_21636);
xnor U22100 (N_22100,N_21942,N_21575);
nor U22101 (N_22101,N_21755,N_21979);
and U22102 (N_22102,N_21542,N_21888);
xor U22103 (N_22103,N_21756,N_21866);
and U22104 (N_22104,N_21723,N_21744);
and U22105 (N_22105,N_21946,N_21941);
or U22106 (N_22106,N_21873,N_21938);
nand U22107 (N_22107,N_21769,N_21650);
nor U22108 (N_22108,N_21665,N_21514);
nand U22109 (N_22109,N_21701,N_21519);
xor U22110 (N_22110,N_21726,N_21834);
nand U22111 (N_22111,N_21631,N_21857);
nor U22112 (N_22112,N_21977,N_21601);
or U22113 (N_22113,N_21793,N_21846);
nand U22114 (N_22114,N_21893,N_21813);
nand U22115 (N_22115,N_21694,N_21579);
and U22116 (N_22116,N_21916,N_21870);
nand U22117 (N_22117,N_21837,N_21598);
and U22118 (N_22118,N_21592,N_21674);
nor U22119 (N_22119,N_21818,N_21534);
or U22120 (N_22120,N_21621,N_21655);
and U22121 (N_22121,N_21800,N_21747);
and U22122 (N_22122,N_21707,N_21619);
xnor U22123 (N_22123,N_21931,N_21782);
xor U22124 (N_22124,N_21990,N_21698);
xor U22125 (N_22125,N_21773,N_21783);
nand U22126 (N_22126,N_21828,N_21614);
and U22127 (N_22127,N_21664,N_21987);
xnor U22128 (N_22128,N_21613,N_21907);
and U22129 (N_22129,N_21691,N_21929);
nand U22130 (N_22130,N_21958,N_21847);
and U22131 (N_22131,N_21760,N_21668);
or U22132 (N_22132,N_21657,N_21905);
or U22133 (N_22133,N_21646,N_21940);
or U22134 (N_22134,N_21716,N_21999);
or U22135 (N_22135,N_21978,N_21927);
and U22136 (N_22136,N_21976,N_21826);
or U22137 (N_22137,N_21692,N_21661);
nor U22138 (N_22138,N_21889,N_21733);
nand U22139 (N_22139,N_21960,N_21953);
xnor U22140 (N_22140,N_21568,N_21997);
nand U22141 (N_22141,N_21877,N_21788);
nor U22142 (N_22142,N_21587,N_21962);
nor U22143 (N_22143,N_21588,N_21984);
or U22144 (N_22144,N_21681,N_21803);
nand U22145 (N_22145,N_21748,N_21971);
and U22146 (N_22146,N_21815,N_21659);
or U22147 (N_22147,N_21637,N_21886);
nor U22148 (N_22148,N_21900,N_21840);
nand U22149 (N_22149,N_21669,N_21936);
xnor U22150 (N_22150,N_21851,N_21594);
and U22151 (N_22151,N_21527,N_21558);
and U22152 (N_22152,N_21896,N_21536);
or U22153 (N_22153,N_21951,N_21583);
or U22154 (N_22154,N_21553,N_21585);
nor U22155 (N_22155,N_21738,N_21589);
nor U22156 (N_22156,N_21505,N_21559);
xnor U22157 (N_22157,N_21956,N_21955);
nor U22158 (N_22158,N_21528,N_21743);
or U22159 (N_22159,N_21871,N_21690);
nor U22160 (N_22160,N_21776,N_21982);
or U22161 (N_22161,N_21673,N_21939);
or U22162 (N_22162,N_21914,N_21819);
nor U22163 (N_22163,N_21576,N_21864);
nor U22164 (N_22164,N_21555,N_21676);
and U22165 (N_22165,N_21736,N_21966);
and U22166 (N_22166,N_21944,N_21904);
xor U22167 (N_22167,N_21541,N_21697);
and U22168 (N_22168,N_21795,N_21964);
xor U22169 (N_22169,N_21824,N_21710);
xnor U22170 (N_22170,N_21814,N_21603);
and U22171 (N_22171,N_21600,N_21644);
or U22172 (N_22172,N_21620,N_21973);
nand U22173 (N_22173,N_21645,N_21581);
or U22174 (N_22174,N_21504,N_21901);
and U22175 (N_22175,N_21812,N_21777);
nor U22176 (N_22176,N_21724,N_21737);
xor U22177 (N_22177,N_21862,N_21898);
xor U22178 (N_22178,N_21865,N_21641);
or U22179 (N_22179,N_21798,N_21839);
or U22180 (N_22180,N_21551,N_21689);
or U22181 (N_22181,N_21629,N_21998);
xnor U22182 (N_22182,N_21804,N_21518);
and U22183 (N_22183,N_21741,N_21768);
and U22184 (N_22184,N_21930,N_21775);
nor U22185 (N_22185,N_21718,N_21623);
and U22186 (N_22186,N_21683,N_21562);
nor U22187 (N_22187,N_21831,N_21554);
and U22188 (N_22188,N_21892,N_21910);
xnor U22189 (N_22189,N_21785,N_21734);
and U22190 (N_22190,N_21693,N_21918);
and U22191 (N_22191,N_21704,N_21662);
or U22192 (N_22192,N_21671,N_21784);
or U22193 (N_22193,N_21617,N_21699);
nor U22194 (N_22194,N_21703,N_21995);
xnor U22195 (N_22195,N_21660,N_21653);
and U22196 (N_22196,N_21539,N_21787);
and U22197 (N_22197,N_21510,N_21533);
or U22198 (N_22198,N_21565,N_21526);
xor U22199 (N_22199,N_21663,N_21595);
or U22200 (N_22200,N_21746,N_21876);
nor U22201 (N_22201,N_21564,N_21823);
and U22202 (N_22202,N_21507,N_21899);
nand U22203 (N_22203,N_21816,N_21548);
and U22204 (N_22204,N_21881,N_21961);
or U22205 (N_22205,N_21906,N_21529);
and U22206 (N_22206,N_21920,N_21719);
and U22207 (N_22207,N_21915,N_21688);
nand U22208 (N_22208,N_21532,N_21677);
nand U22209 (N_22209,N_21728,N_21863);
nor U22210 (N_22210,N_21854,N_21667);
or U22211 (N_22211,N_21879,N_21883);
nand U22212 (N_22212,N_21616,N_21609);
or U22213 (N_22213,N_21618,N_21985);
nand U22214 (N_22214,N_21634,N_21867);
or U22215 (N_22215,N_21712,N_21954);
and U22216 (N_22216,N_21996,N_21796);
and U22217 (N_22217,N_21752,N_21745);
xnor U22218 (N_22218,N_21572,N_21841);
xor U22219 (N_22219,N_21830,N_21989);
or U22220 (N_22220,N_21722,N_21832);
or U22221 (N_22221,N_21525,N_21599);
xnor U22222 (N_22222,N_21912,N_21845);
or U22223 (N_22223,N_21820,N_21591);
or U22224 (N_22224,N_21680,N_21706);
and U22225 (N_22225,N_21791,N_21861);
or U22226 (N_22226,N_21522,N_21638);
xor U22227 (N_22227,N_21530,N_21628);
xnor U22228 (N_22228,N_21610,N_21765);
xnor U22229 (N_22229,N_21887,N_21727);
or U22230 (N_22230,N_21590,N_21869);
nor U22231 (N_22231,N_21509,N_21786);
and U22232 (N_22232,N_21858,N_21584);
and U22233 (N_22233,N_21574,N_21729);
nand U22234 (N_22234,N_21957,N_21711);
nand U22235 (N_22235,N_21781,N_21801);
or U22236 (N_22236,N_21586,N_21764);
nand U22237 (N_22237,N_21903,N_21890);
nand U22238 (N_22238,N_21606,N_21569);
xor U22239 (N_22239,N_21651,N_21633);
and U22240 (N_22240,N_21894,N_21612);
nor U22241 (N_22241,N_21563,N_21672);
xor U22242 (N_22242,N_21511,N_21735);
nand U22243 (N_22243,N_21758,N_21872);
nor U22244 (N_22244,N_21850,N_21593);
and U22245 (N_22245,N_21751,N_21535);
and U22246 (N_22246,N_21695,N_21642);
nand U22247 (N_22247,N_21880,N_21842);
nor U22248 (N_22248,N_21771,N_21713);
or U22249 (N_22249,N_21836,N_21983);
nor U22250 (N_22250,N_21700,N_21652);
xor U22251 (N_22251,N_21732,N_21915);
or U22252 (N_22252,N_21878,N_21544);
or U22253 (N_22253,N_21588,N_21649);
or U22254 (N_22254,N_21962,N_21849);
or U22255 (N_22255,N_21968,N_21649);
and U22256 (N_22256,N_21651,N_21982);
xor U22257 (N_22257,N_21990,N_21895);
xor U22258 (N_22258,N_21567,N_21671);
nand U22259 (N_22259,N_21894,N_21754);
or U22260 (N_22260,N_21524,N_21812);
and U22261 (N_22261,N_21639,N_21625);
and U22262 (N_22262,N_21929,N_21962);
xnor U22263 (N_22263,N_21861,N_21911);
and U22264 (N_22264,N_21751,N_21861);
nand U22265 (N_22265,N_21867,N_21838);
nand U22266 (N_22266,N_21754,N_21913);
nor U22267 (N_22267,N_21515,N_21786);
xor U22268 (N_22268,N_21538,N_21659);
xnor U22269 (N_22269,N_21554,N_21532);
xnor U22270 (N_22270,N_21659,N_21655);
nor U22271 (N_22271,N_21973,N_21887);
nand U22272 (N_22272,N_21860,N_21874);
nand U22273 (N_22273,N_21525,N_21606);
xnor U22274 (N_22274,N_21950,N_21760);
and U22275 (N_22275,N_21841,N_21945);
and U22276 (N_22276,N_21896,N_21717);
xor U22277 (N_22277,N_21980,N_21820);
and U22278 (N_22278,N_21619,N_21750);
nand U22279 (N_22279,N_21564,N_21577);
xnor U22280 (N_22280,N_21831,N_21612);
xor U22281 (N_22281,N_21579,N_21875);
nand U22282 (N_22282,N_21899,N_21568);
and U22283 (N_22283,N_21525,N_21586);
and U22284 (N_22284,N_21850,N_21769);
xnor U22285 (N_22285,N_21905,N_21554);
and U22286 (N_22286,N_21915,N_21612);
xnor U22287 (N_22287,N_21828,N_21660);
and U22288 (N_22288,N_21785,N_21626);
nor U22289 (N_22289,N_21629,N_21597);
or U22290 (N_22290,N_21547,N_21641);
and U22291 (N_22291,N_21833,N_21605);
nand U22292 (N_22292,N_21592,N_21733);
nor U22293 (N_22293,N_21531,N_21836);
or U22294 (N_22294,N_21999,N_21514);
nand U22295 (N_22295,N_21807,N_21631);
xnor U22296 (N_22296,N_21736,N_21842);
xnor U22297 (N_22297,N_21598,N_21508);
xnor U22298 (N_22298,N_21579,N_21769);
or U22299 (N_22299,N_21965,N_21887);
nor U22300 (N_22300,N_21651,N_21854);
nor U22301 (N_22301,N_21580,N_21954);
nand U22302 (N_22302,N_21955,N_21913);
nand U22303 (N_22303,N_21913,N_21534);
nand U22304 (N_22304,N_21819,N_21810);
or U22305 (N_22305,N_21754,N_21706);
xnor U22306 (N_22306,N_21664,N_21866);
nor U22307 (N_22307,N_21917,N_21528);
nor U22308 (N_22308,N_21747,N_21848);
and U22309 (N_22309,N_21611,N_21928);
nand U22310 (N_22310,N_21637,N_21912);
nor U22311 (N_22311,N_21908,N_21956);
and U22312 (N_22312,N_21688,N_21604);
and U22313 (N_22313,N_21692,N_21763);
and U22314 (N_22314,N_21765,N_21565);
and U22315 (N_22315,N_21714,N_21517);
and U22316 (N_22316,N_21545,N_21539);
nand U22317 (N_22317,N_21705,N_21789);
and U22318 (N_22318,N_21745,N_21683);
and U22319 (N_22319,N_21975,N_21661);
and U22320 (N_22320,N_21769,N_21525);
or U22321 (N_22321,N_21571,N_21948);
nor U22322 (N_22322,N_21948,N_21695);
nor U22323 (N_22323,N_21693,N_21856);
or U22324 (N_22324,N_21855,N_21597);
xnor U22325 (N_22325,N_21849,N_21589);
and U22326 (N_22326,N_21981,N_21708);
or U22327 (N_22327,N_21608,N_21606);
and U22328 (N_22328,N_21966,N_21898);
xor U22329 (N_22329,N_21975,N_21920);
or U22330 (N_22330,N_21618,N_21862);
xor U22331 (N_22331,N_21525,N_21589);
nand U22332 (N_22332,N_21576,N_21540);
nor U22333 (N_22333,N_21952,N_21645);
nand U22334 (N_22334,N_21923,N_21760);
and U22335 (N_22335,N_21897,N_21531);
xnor U22336 (N_22336,N_21738,N_21651);
xnor U22337 (N_22337,N_21618,N_21851);
and U22338 (N_22338,N_21790,N_21672);
or U22339 (N_22339,N_21689,N_21816);
xor U22340 (N_22340,N_21749,N_21757);
or U22341 (N_22341,N_21787,N_21694);
or U22342 (N_22342,N_21962,N_21939);
xnor U22343 (N_22343,N_21505,N_21658);
and U22344 (N_22344,N_21820,N_21546);
xnor U22345 (N_22345,N_21849,N_21745);
nand U22346 (N_22346,N_21574,N_21639);
and U22347 (N_22347,N_21761,N_21852);
nand U22348 (N_22348,N_21738,N_21835);
nand U22349 (N_22349,N_21651,N_21899);
or U22350 (N_22350,N_21610,N_21532);
and U22351 (N_22351,N_21668,N_21767);
xor U22352 (N_22352,N_21671,N_21923);
or U22353 (N_22353,N_21571,N_21510);
and U22354 (N_22354,N_21642,N_21912);
nor U22355 (N_22355,N_21774,N_21936);
xnor U22356 (N_22356,N_21977,N_21867);
xnor U22357 (N_22357,N_21747,N_21530);
nor U22358 (N_22358,N_21608,N_21952);
nand U22359 (N_22359,N_21711,N_21730);
and U22360 (N_22360,N_21818,N_21665);
and U22361 (N_22361,N_21719,N_21702);
nor U22362 (N_22362,N_21976,N_21837);
and U22363 (N_22363,N_21705,N_21910);
nor U22364 (N_22364,N_21792,N_21893);
nand U22365 (N_22365,N_21552,N_21688);
nor U22366 (N_22366,N_21587,N_21971);
nor U22367 (N_22367,N_21687,N_21796);
nor U22368 (N_22368,N_21821,N_21599);
and U22369 (N_22369,N_21503,N_21882);
or U22370 (N_22370,N_21695,N_21889);
nand U22371 (N_22371,N_21827,N_21648);
or U22372 (N_22372,N_21909,N_21530);
nor U22373 (N_22373,N_21879,N_21786);
nand U22374 (N_22374,N_21537,N_21551);
nor U22375 (N_22375,N_21876,N_21921);
or U22376 (N_22376,N_21563,N_21633);
xnor U22377 (N_22377,N_21605,N_21915);
and U22378 (N_22378,N_21717,N_21639);
nor U22379 (N_22379,N_21639,N_21642);
xnor U22380 (N_22380,N_21979,N_21572);
nor U22381 (N_22381,N_21809,N_21529);
nand U22382 (N_22382,N_21516,N_21620);
or U22383 (N_22383,N_21959,N_21935);
nor U22384 (N_22384,N_21923,N_21827);
nor U22385 (N_22385,N_21612,N_21963);
nand U22386 (N_22386,N_21762,N_21521);
nor U22387 (N_22387,N_21845,N_21786);
and U22388 (N_22388,N_21607,N_21897);
nor U22389 (N_22389,N_21773,N_21610);
and U22390 (N_22390,N_21566,N_21886);
or U22391 (N_22391,N_21778,N_21945);
nor U22392 (N_22392,N_21897,N_21739);
xnor U22393 (N_22393,N_21569,N_21885);
nor U22394 (N_22394,N_21566,N_21859);
and U22395 (N_22395,N_21516,N_21962);
xor U22396 (N_22396,N_21678,N_21500);
nand U22397 (N_22397,N_21974,N_21728);
and U22398 (N_22398,N_21705,N_21842);
nand U22399 (N_22399,N_21664,N_21829);
nand U22400 (N_22400,N_21973,N_21811);
and U22401 (N_22401,N_21515,N_21851);
and U22402 (N_22402,N_21524,N_21976);
xnor U22403 (N_22403,N_21534,N_21622);
nor U22404 (N_22404,N_21776,N_21847);
and U22405 (N_22405,N_21532,N_21602);
or U22406 (N_22406,N_21726,N_21952);
nor U22407 (N_22407,N_21665,N_21836);
or U22408 (N_22408,N_21615,N_21779);
and U22409 (N_22409,N_21519,N_21887);
nor U22410 (N_22410,N_21624,N_21739);
and U22411 (N_22411,N_21800,N_21733);
nand U22412 (N_22412,N_21500,N_21726);
xor U22413 (N_22413,N_21780,N_21813);
nand U22414 (N_22414,N_21994,N_21661);
or U22415 (N_22415,N_21872,N_21606);
xor U22416 (N_22416,N_21549,N_21837);
nand U22417 (N_22417,N_21516,N_21915);
nor U22418 (N_22418,N_21962,N_21741);
xnor U22419 (N_22419,N_21912,N_21645);
and U22420 (N_22420,N_21758,N_21601);
nor U22421 (N_22421,N_21514,N_21619);
or U22422 (N_22422,N_21601,N_21660);
and U22423 (N_22423,N_21864,N_21869);
and U22424 (N_22424,N_21701,N_21928);
nand U22425 (N_22425,N_21530,N_21697);
nor U22426 (N_22426,N_21842,N_21903);
or U22427 (N_22427,N_21901,N_21906);
nor U22428 (N_22428,N_21802,N_21747);
or U22429 (N_22429,N_21754,N_21727);
nand U22430 (N_22430,N_21560,N_21667);
and U22431 (N_22431,N_21511,N_21683);
xnor U22432 (N_22432,N_21716,N_21777);
or U22433 (N_22433,N_21675,N_21877);
xnor U22434 (N_22434,N_21982,N_21543);
or U22435 (N_22435,N_21906,N_21995);
xnor U22436 (N_22436,N_21839,N_21935);
and U22437 (N_22437,N_21922,N_21919);
and U22438 (N_22438,N_21553,N_21872);
nand U22439 (N_22439,N_21736,N_21820);
and U22440 (N_22440,N_21611,N_21615);
and U22441 (N_22441,N_21723,N_21867);
nand U22442 (N_22442,N_21586,N_21938);
or U22443 (N_22443,N_21825,N_21835);
or U22444 (N_22444,N_21892,N_21674);
nor U22445 (N_22445,N_21659,N_21606);
or U22446 (N_22446,N_21771,N_21876);
nor U22447 (N_22447,N_21921,N_21841);
and U22448 (N_22448,N_21995,N_21986);
xnor U22449 (N_22449,N_21942,N_21591);
or U22450 (N_22450,N_21731,N_21904);
nor U22451 (N_22451,N_21539,N_21699);
nor U22452 (N_22452,N_21744,N_21890);
nand U22453 (N_22453,N_21506,N_21629);
and U22454 (N_22454,N_21806,N_21725);
and U22455 (N_22455,N_21855,N_21749);
xor U22456 (N_22456,N_21712,N_21806);
nor U22457 (N_22457,N_21689,N_21958);
or U22458 (N_22458,N_21675,N_21563);
and U22459 (N_22459,N_21954,N_21677);
xor U22460 (N_22460,N_21814,N_21959);
nand U22461 (N_22461,N_21959,N_21829);
nor U22462 (N_22462,N_21601,N_21894);
nand U22463 (N_22463,N_21670,N_21995);
xnor U22464 (N_22464,N_21709,N_21821);
nor U22465 (N_22465,N_21731,N_21718);
xor U22466 (N_22466,N_21641,N_21908);
nand U22467 (N_22467,N_21554,N_21668);
nand U22468 (N_22468,N_21696,N_21996);
nor U22469 (N_22469,N_21659,N_21552);
or U22470 (N_22470,N_21928,N_21857);
nand U22471 (N_22471,N_21704,N_21943);
nand U22472 (N_22472,N_21717,N_21893);
nand U22473 (N_22473,N_21525,N_21714);
or U22474 (N_22474,N_21523,N_21790);
and U22475 (N_22475,N_21764,N_21782);
nand U22476 (N_22476,N_21601,N_21859);
and U22477 (N_22477,N_21730,N_21789);
nor U22478 (N_22478,N_21790,N_21536);
xor U22479 (N_22479,N_21546,N_21815);
or U22480 (N_22480,N_21659,N_21526);
nand U22481 (N_22481,N_21601,N_21534);
nor U22482 (N_22482,N_21878,N_21879);
and U22483 (N_22483,N_21931,N_21790);
nand U22484 (N_22484,N_21686,N_21926);
or U22485 (N_22485,N_21860,N_21864);
and U22486 (N_22486,N_21942,N_21765);
and U22487 (N_22487,N_21995,N_21761);
or U22488 (N_22488,N_21680,N_21822);
and U22489 (N_22489,N_21760,N_21579);
or U22490 (N_22490,N_21682,N_21538);
and U22491 (N_22491,N_21834,N_21932);
and U22492 (N_22492,N_21918,N_21837);
xnor U22493 (N_22493,N_21695,N_21800);
xnor U22494 (N_22494,N_21825,N_21663);
nor U22495 (N_22495,N_21970,N_21547);
nor U22496 (N_22496,N_21538,N_21702);
nand U22497 (N_22497,N_21527,N_21979);
xor U22498 (N_22498,N_21538,N_21593);
and U22499 (N_22499,N_21972,N_21779);
nand U22500 (N_22500,N_22278,N_22121);
nand U22501 (N_22501,N_22248,N_22301);
xor U22502 (N_22502,N_22243,N_22101);
nand U22503 (N_22503,N_22283,N_22191);
xnor U22504 (N_22504,N_22181,N_22249);
nand U22505 (N_22505,N_22455,N_22001);
nor U22506 (N_22506,N_22317,N_22203);
xnor U22507 (N_22507,N_22465,N_22469);
or U22508 (N_22508,N_22263,N_22000);
and U22509 (N_22509,N_22076,N_22194);
nor U22510 (N_22510,N_22259,N_22485);
nor U22511 (N_22511,N_22160,N_22063);
xnor U22512 (N_22512,N_22175,N_22309);
nand U22513 (N_22513,N_22353,N_22190);
nand U22514 (N_22514,N_22406,N_22351);
or U22515 (N_22515,N_22024,N_22221);
nand U22516 (N_22516,N_22446,N_22449);
or U22517 (N_22517,N_22496,N_22339);
nor U22518 (N_22518,N_22111,N_22041);
or U22519 (N_22519,N_22039,N_22180);
or U22520 (N_22520,N_22021,N_22269);
nand U22521 (N_22521,N_22014,N_22102);
or U22522 (N_22522,N_22371,N_22226);
nand U22523 (N_22523,N_22489,N_22038);
and U22524 (N_22524,N_22238,N_22466);
and U22525 (N_22525,N_22133,N_22347);
xor U22526 (N_22526,N_22200,N_22186);
or U22527 (N_22527,N_22045,N_22064);
xnor U22528 (N_22528,N_22217,N_22373);
xnor U22529 (N_22529,N_22230,N_22428);
nor U22530 (N_22530,N_22116,N_22183);
nor U22531 (N_22531,N_22482,N_22320);
nor U22532 (N_22532,N_22222,N_22438);
or U22533 (N_22533,N_22372,N_22030);
xor U22534 (N_22534,N_22491,N_22058);
nand U22535 (N_22535,N_22486,N_22344);
nor U22536 (N_22536,N_22060,N_22197);
and U22537 (N_22537,N_22250,N_22313);
nor U22538 (N_22538,N_22098,N_22240);
or U22539 (N_22539,N_22042,N_22146);
nor U22540 (N_22540,N_22009,N_22336);
or U22541 (N_22541,N_22319,N_22450);
and U22542 (N_22542,N_22417,N_22052);
xnor U22543 (N_22543,N_22260,N_22077);
nor U22544 (N_22544,N_22171,N_22463);
or U22545 (N_22545,N_22280,N_22410);
or U22546 (N_22546,N_22059,N_22073);
nand U22547 (N_22547,N_22242,N_22147);
nor U22548 (N_22548,N_22342,N_22464);
nor U22549 (N_22549,N_22215,N_22376);
xor U22550 (N_22550,N_22108,N_22325);
nor U22551 (N_22551,N_22233,N_22007);
and U22552 (N_22552,N_22251,N_22369);
or U22553 (N_22553,N_22490,N_22026);
nand U22554 (N_22554,N_22433,N_22266);
nor U22555 (N_22555,N_22487,N_22214);
nor U22556 (N_22556,N_22182,N_22338);
xor U22557 (N_22557,N_22357,N_22131);
xnor U22558 (N_22558,N_22331,N_22389);
xnor U22559 (N_22559,N_22333,N_22168);
or U22560 (N_22560,N_22153,N_22154);
or U22561 (N_22561,N_22193,N_22177);
xnor U22562 (N_22562,N_22267,N_22361);
or U22563 (N_22563,N_22211,N_22151);
nor U22564 (N_22564,N_22341,N_22087);
or U22565 (N_22565,N_22397,N_22099);
nand U22566 (N_22566,N_22277,N_22481);
nor U22567 (N_22567,N_22055,N_22107);
nand U22568 (N_22568,N_22439,N_22396);
nor U22569 (N_22569,N_22235,N_22295);
nand U22570 (N_22570,N_22452,N_22126);
or U22571 (N_22571,N_22167,N_22460);
nand U22572 (N_22572,N_22299,N_22141);
and U22573 (N_22573,N_22327,N_22380);
nor U22574 (N_22574,N_22411,N_22425);
nand U22575 (N_22575,N_22286,N_22422);
and U22576 (N_22576,N_22326,N_22315);
or U22577 (N_22577,N_22148,N_22138);
nor U22578 (N_22578,N_22386,N_22470);
nor U22579 (N_22579,N_22314,N_22374);
or U22580 (N_22580,N_22002,N_22117);
xor U22581 (N_22581,N_22224,N_22401);
or U22582 (N_22582,N_22031,N_22231);
and U22583 (N_22583,N_22477,N_22252);
nand U22584 (N_22584,N_22135,N_22395);
nand U22585 (N_22585,N_22012,N_22441);
and U22586 (N_22586,N_22382,N_22174);
and U22587 (N_22587,N_22228,N_22213);
xor U22588 (N_22588,N_22409,N_22384);
xnor U22589 (N_22589,N_22364,N_22334);
nand U22590 (N_22590,N_22367,N_22311);
or U22591 (N_22591,N_22155,N_22069);
and U22592 (N_22592,N_22451,N_22285);
xnor U22593 (N_22593,N_22068,N_22127);
or U22594 (N_22594,N_22329,N_22156);
and U22595 (N_22595,N_22442,N_22343);
xor U22596 (N_22596,N_22322,N_22196);
nand U22597 (N_22597,N_22476,N_22236);
nor U22598 (N_22598,N_22400,N_22305);
or U22599 (N_22599,N_22208,N_22474);
or U22600 (N_22600,N_22037,N_22272);
xnor U22601 (N_22601,N_22142,N_22234);
nor U22602 (N_22602,N_22199,N_22070);
nor U22603 (N_22603,N_22348,N_22114);
and U22604 (N_22604,N_22275,N_22046);
xor U22605 (N_22605,N_22271,N_22444);
nor U22606 (N_22606,N_22276,N_22006);
nand U22607 (N_22607,N_22150,N_22247);
and U22608 (N_22608,N_22426,N_22015);
nand U22609 (N_22609,N_22293,N_22393);
and U22610 (N_22610,N_22381,N_22158);
xnor U22611 (N_22611,N_22404,N_22023);
or U22612 (N_22612,N_22443,N_22256);
and U22613 (N_22613,N_22051,N_22365);
xnor U22614 (N_22614,N_22048,N_22416);
nor U22615 (N_22615,N_22424,N_22090);
nand U22616 (N_22616,N_22094,N_22152);
or U22617 (N_22617,N_22494,N_22033);
nor U22618 (N_22618,N_22379,N_22005);
or U22619 (N_22619,N_22419,N_22284);
or U22620 (N_22620,N_22095,N_22316);
and U22621 (N_22621,N_22435,N_22436);
or U22622 (N_22622,N_22306,N_22209);
and U22623 (N_22623,N_22157,N_22165);
nor U22624 (N_22624,N_22169,N_22332);
or U22625 (N_22625,N_22270,N_22049);
and U22626 (N_22626,N_22420,N_22454);
or U22627 (N_22627,N_22223,N_22179);
nor U22628 (N_22628,N_22457,N_22349);
or U22629 (N_22629,N_22297,N_22407);
and U22630 (N_22630,N_22122,N_22300);
or U22631 (N_22631,N_22178,N_22136);
nor U22632 (N_22632,N_22020,N_22008);
or U22633 (N_22633,N_22066,N_22498);
nand U22634 (N_22634,N_22130,N_22262);
or U22635 (N_22635,N_22056,N_22140);
nor U22636 (N_22636,N_22461,N_22366);
nand U22637 (N_22637,N_22459,N_22447);
nand U22638 (N_22638,N_22370,N_22119);
nor U22639 (N_22639,N_22456,N_22291);
and U22640 (N_22640,N_22281,N_22050);
and U22641 (N_22641,N_22207,N_22134);
nor U22642 (N_22642,N_22375,N_22075);
xor U22643 (N_22643,N_22488,N_22472);
or U22644 (N_22644,N_22123,N_22053);
nor U22645 (N_22645,N_22081,N_22025);
or U22646 (N_22646,N_22378,N_22034);
and U22647 (N_22647,N_22054,N_22096);
nand U22648 (N_22648,N_22017,N_22377);
nor U22649 (N_22649,N_22368,N_22164);
xnor U22650 (N_22650,N_22354,N_22318);
or U22651 (N_22651,N_22398,N_22088);
and U22652 (N_22652,N_22307,N_22044);
or U22653 (N_22653,N_22478,N_22105);
xnor U22654 (N_22654,N_22337,N_22166);
nor U22655 (N_22655,N_22399,N_22359);
nor U22656 (N_22656,N_22387,N_22290);
xnor U22657 (N_22657,N_22360,N_22388);
or U22658 (N_22658,N_22479,N_22029);
nor U22659 (N_22659,N_22304,N_22018);
xnor U22660 (N_22660,N_22245,N_22061);
nor U22661 (N_22661,N_22161,N_22080);
or U22662 (N_22662,N_22071,N_22229);
and U22663 (N_22663,N_22057,N_22484);
and U22664 (N_22664,N_22279,N_22408);
nand U22665 (N_22665,N_22261,N_22427);
nor U22666 (N_22666,N_22218,N_22162);
or U22667 (N_22667,N_22145,N_22423);
or U22668 (N_22668,N_22074,N_22016);
or U22669 (N_22669,N_22072,N_22492);
and U22670 (N_22670,N_22363,N_22128);
nor U22671 (N_22671,N_22028,N_22144);
nor U22672 (N_22672,N_22324,N_22497);
nor U22673 (N_22673,N_22264,N_22198);
xor U22674 (N_22674,N_22091,N_22321);
nor U22675 (N_22675,N_22013,N_22458);
and U22676 (N_22676,N_22110,N_22113);
nor U22677 (N_22677,N_22184,N_22212);
nor U22678 (N_22678,N_22106,N_22083);
or U22679 (N_22679,N_22241,N_22085);
xor U22680 (N_22680,N_22067,N_22288);
nor U22681 (N_22681,N_22043,N_22204);
nor U22682 (N_22682,N_22129,N_22345);
xnor U22683 (N_22683,N_22210,N_22287);
xor U22684 (N_22684,N_22022,N_22092);
and U22685 (N_22685,N_22103,N_22468);
xnor U22686 (N_22686,N_22254,N_22019);
nor U22687 (N_22687,N_22172,N_22239);
or U22688 (N_22688,N_22244,N_22350);
xnor U22689 (N_22689,N_22232,N_22216);
or U22690 (N_22690,N_22298,N_22429);
or U22691 (N_22691,N_22453,N_22253);
nand U22692 (N_22692,N_22132,N_22473);
nor U22693 (N_22693,N_22035,N_22383);
or U22694 (N_22694,N_22202,N_22079);
and U22695 (N_22695,N_22414,N_22010);
nor U22696 (N_22696,N_22413,N_22405);
xnor U22697 (N_22697,N_22205,N_22330);
or U22698 (N_22698,N_22418,N_22206);
or U22699 (N_22699,N_22462,N_22137);
xnor U22700 (N_22700,N_22176,N_22445);
nor U22701 (N_22701,N_22340,N_22124);
nand U22702 (N_22702,N_22246,N_22475);
nand U22703 (N_22703,N_22187,N_22415);
nor U22704 (N_22704,N_22412,N_22036);
and U22705 (N_22705,N_22282,N_22084);
xor U22706 (N_22706,N_22163,N_22258);
and U22707 (N_22707,N_22294,N_22268);
nand U22708 (N_22708,N_22328,N_22255);
nor U22709 (N_22709,N_22225,N_22032);
nor U22710 (N_22710,N_22434,N_22403);
nand U22711 (N_22711,N_22352,N_22431);
and U22712 (N_22712,N_22220,N_22499);
and U22713 (N_22713,N_22335,N_22390);
or U22714 (N_22714,N_22089,N_22004);
nand U22715 (N_22715,N_22274,N_22118);
or U22716 (N_22716,N_22312,N_22011);
nor U22717 (N_22717,N_22362,N_22302);
and U22718 (N_22718,N_22385,N_22356);
and U22719 (N_22719,N_22391,N_22078);
or U22720 (N_22720,N_22237,N_22201);
nand U22721 (N_22721,N_22467,N_22109);
nor U22722 (N_22722,N_22392,N_22257);
nand U22723 (N_22723,N_22027,N_22308);
nand U22724 (N_22724,N_22047,N_22188);
or U22725 (N_22725,N_22432,N_22120);
and U22726 (N_22726,N_22003,N_22483);
or U22727 (N_22727,N_22358,N_22480);
nand U22728 (N_22728,N_22448,N_22104);
and U22729 (N_22729,N_22185,N_22402);
or U22730 (N_22730,N_22219,N_22394);
nand U22731 (N_22731,N_22040,N_22495);
or U22732 (N_22732,N_22440,N_22086);
nand U22733 (N_22733,N_22346,N_22355);
xnor U22734 (N_22734,N_22093,N_22143);
or U22735 (N_22735,N_22112,N_22192);
nand U22736 (N_22736,N_22323,N_22149);
nor U22737 (N_22737,N_22310,N_22065);
or U22738 (N_22738,N_22227,N_22159);
nand U22739 (N_22739,N_22437,N_22430);
nor U22740 (N_22740,N_22173,N_22097);
xnor U22741 (N_22741,N_22062,N_22100);
xor U22742 (N_22742,N_22195,N_22265);
or U22743 (N_22743,N_22139,N_22296);
nor U22744 (N_22744,N_22189,N_22115);
nand U22745 (N_22745,N_22273,N_22471);
xnor U22746 (N_22746,N_22082,N_22170);
nand U22747 (N_22747,N_22125,N_22421);
xor U22748 (N_22748,N_22289,N_22292);
or U22749 (N_22749,N_22303,N_22493);
nand U22750 (N_22750,N_22447,N_22395);
nand U22751 (N_22751,N_22367,N_22217);
nand U22752 (N_22752,N_22351,N_22320);
or U22753 (N_22753,N_22104,N_22313);
xnor U22754 (N_22754,N_22265,N_22053);
and U22755 (N_22755,N_22427,N_22132);
xor U22756 (N_22756,N_22300,N_22389);
nor U22757 (N_22757,N_22088,N_22413);
nor U22758 (N_22758,N_22253,N_22324);
nand U22759 (N_22759,N_22013,N_22245);
xnor U22760 (N_22760,N_22086,N_22407);
xor U22761 (N_22761,N_22016,N_22110);
nand U22762 (N_22762,N_22459,N_22354);
and U22763 (N_22763,N_22150,N_22200);
or U22764 (N_22764,N_22253,N_22459);
nand U22765 (N_22765,N_22459,N_22164);
or U22766 (N_22766,N_22197,N_22199);
and U22767 (N_22767,N_22266,N_22074);
and U22768 (N_22768,N_22173,N_22323);
or U22769 (N_22769,N_22274,N_22407);
nor U22770 (N_22770,N_22075,N_22297);
or U22771 (N_22771,N_22367,N_22498);
and U22772 (N_22772,N_22079,N_22176);
nand U22773 (N_22773,N_22236,N_22343);
xor U22774 (N_22774,N_22418,N_22437);
xnor U22775 (N_22775,N_22115,N_22264);
and U22776 (N_22776,N_22181,N_22070);
and U22777 (N_22777,N_22258,N_22254);
xor U22778 (N_22778,N_22242,N_22111);
and U22779 (N_22779,N_22152,N_22026);
nand U22780 (N_22780,N_22137,N_22151);
xnor U22781 (N_22781,N_22081,N_22165);
and U22782 (N_22782,N_22112,N_22108);
nand U22783 (N_22783,N_22426,N_22093);
nand U22784 (N_22784,N_22070,N_22379);
xor U22785 (N_22785,N_22492,N_22446);
and U22786 (N_22786,N_22254,N_22058);
nand U22787 (N_22787,N_22397,N_22257);
nor U22788 (N_22788,N_22356,N_22118);
xnor U22789 (N_22789,N_22051,N_22396);
and U22790 (N_22790,N_22297,N_22363);
xnor U22791 (N_22791,N_22176,N_22048);
xnor U22792 (N_22792,N_22127,N_22047);
nor U22793 (N_22793,N_22425,N_22307);
and U22794 (N_22794,N_22106,N_22393);
nor U22795 (N_22795,N_22328,N_22383);
and U22796 (N_22796,N_22241,N_22133);
or U22797 (N_22797,N_22012,N_22176);
xnor U22798 (N_22798,N_22194,N_22125);
nor U22799 (N_22799,N_22413,N_22205);
or U22800 (N_22800,N_22127,N_22420);
or U22801 (N_22801,N_22096,N_22107);
and U22802 (N_22802,N_22406,N_22004);
nand U22803 (N_22803,N_22329,N_22171);
and U22804 (N_22804,N_22171,N_22223);
nand U22805 (N_22805,N_22089,N_22232);
nor U22806 (N_22806,N_22287,N_22079);
nor U22807 (N_22807,N_22201,N_22485);
xnor U22808 (N_22808,N_22147,N_22257);
xnor U22809 (N_22809,N_22427,N_22214);
or U22810 (N_22810,N_22134,N_22368);
xnor U22811 (N_22811,N_22306,N_22288);
or U22812 (N_22812,N_22090,N_22169);
nor U22813 (N_22813,N_22229,N_22099);
nor U22814 (N_22814,N_22332,N_22012);
xor U22815 (N_22815,N_22251,N_22471);
or U22816 (N_22816,N_22312,N_22069);
or U22817 (N_22817,N_22364,N_22036);
nand U22818 (N_22818,N_22259,N_22281);
nand U22819 (N_22819,N_22427,N_22089);
and U22820 (N_22820,N_22120,N_22037);
nor U22821 (N_22821,N_22381,N_22309);
or U22822 (N_22822,N_22247,N_22136);
nand U22823 (N_22823,N_22458,N_22065);
nor U22824 (N_22824,N_22376,N_22254);
or U22825 (N_22825,N_22329,N_22443);
or U22826 (N_22826,N_22410,N_22348);
or U22827 (N_22827,N_22413,N_22179);
xor U22828 (N_22828,N_22279,N_22032);
xnor U22829 (N_22829,N_22374,N_22356);
xnor U22830 (N_22830,N_22062,N_22485);
nor U22831 (N_22831,N_22129,N_22251);
and U22832 (N_22832,N_22027,N_22358);
nor U22833 (N_22833,N_22380,N_22084);
nor U22834 (N_22834,N_22499,N_22256);
or U22835 (N_22835,N_22265,N_22138);
nor U22836 (N_22836,N_22440,N_22315);
nor U22837 (N_22837,N_22426,N_22455);
nand U22838 (N_22838,N_22454,N_22376);
nor U22839 (N_22839,N_22242,N_22117);
nor U22840 (N_22840,N_22432,N_22142);
nor U22841 (N_22841,N_22067,N_22086);
nand U22842 (N_22842,N_22384,N_22013);
and U22843 (N_22843,N_22138,N_22139);
or U22844 (N_22844,N_22178,N_22404);
and U22845 (N_22845,N_22175,N_22360);
and U22846 (N_22846,N_22155,N_22067);
nand U22847 (N_22847,N_22059,N_22497);
nand U22848 (N_22848,N_22090,N_22484);
and U22849 (N_22849,N_22169,N_22281);
xor U22850 (N_22850,N_22095,N_22370);
or U22851 (N_22851,N_22281,N_22380);
nand U22852 (N_22852,N_22492,N_22212);
nand U22853 (N_22853,N_22273,N_22468);
or U22854 (N_22854,N_22190,N_22125);
and U22855 (N_22855,N_22346,N_22284);
and U22856 (N_22856,N_22076,N_22308);
or U22857 (N_22857,N_22439,N_22156);
or U22858 (N_22858,N_22377,N_22389);
nand U22859 (N_22859,N_22397,N_22004);
and U22860 (N_22860,N_22395,N_22151);
and U22861 (N_22861,N_22392,N_22058);
and U22862 (N_22862,N_22035,N_22430);
xor U22863 (N_22863,N_22330,N_22073);
xor U22864 (N_22864,N_22301,N_22023);
nor U22865 (N_22865,N_22031,N_22143);
nor U22866 (N_22866,N_22291,N_22269);
or U22867 (N_22867,N_22395,N_22270);
nand U22868 (N_22868,N_22306,N_22026);
xnor U22869 (N_22869,N_22113,N_22045);
and U22870 (N_22870,N_22313,N_22145);
nand U22871 (N_22871,N_22494,N_22152);
xnor U22872 (N_22872,N_22353,N_22040);
xnor U22873 (N_22873,N_22160,N_22104);
nand U22874 (N_22874,N_22254,N_22492);
xnor U22875 (N_22875,N_22187,N_22276);
nand U22876 (N_22876,N_22002,N_22005);
nor U22877 (N_22877,N_22185,N_22142);
xnor U22878 (N_22878,N_22080,N_22498);
and U22879 (N_22879,N_22176,N_22267);
nor U22880 (N_22880,N_22245,N_22238);
and U22881 (N_22881,N_22099,N_22086);
or U22882 (N_22882,N_22246,N_22301);
or U22883 (N_22883,N_22016,N_22028);
nand U22884 (N_22884,N_22392,N_22015);
and U22885 (N_22885,N_22038,N_22448);
nand U22886 (N_22886,N_22168,N_22008);
nand U22887 (N_22887,N_22224,N_22084);
nand U22888 (N_22888,N_22489,N_22068);
nand U22889 (N_22889,N_22060,N_22455);
or U22890 (N_22890,N_22359,N_22317);
xor U22891 (N_22891,N_22293,N_22468);
or U22892 (N_22892,N_22214,N_22420);
and U22893 (N_22893,N_22442,N_22054);
xor U22894 (N_22894,N_22476,N_22177);
nor U22895 (N_22895,N_22141,N_22330);
xnor U22896 (N_22896,N_22010,N_22062);
nand U22897 (N_22897,N_22079,N_22475);
and U22898 (N_22898,N_22170,N_22363);
nand U22899 (N_22899,N_22037,N_22496);
and U22900 (N_22900,N_22192,N_22208);
and U22901 (N_22901,N_22310,N_22432);
nand U22902 (N_22902,N_22391,N_22070);
or U22903 (N_22903,N_22223,N_22021);
nand U22904 (N_22904,N_22077,N_22097);
nand U22905 (N_22905,N_22201,N_22055);
nor U22906 (N_22906,N_22063,N_22387);
and U22907 (N_22907,N_22323,N_22377);
nor U22908 (N_22908,N_22111,N_22318);
nor U22909 (N_22909,N_22075,N_22473);
xnor U22910 (N_22910,N_22438,N_22186);
xor U22911 (N_22911,N_22037,N_22490);
nand U22912 (N_22912,N_22445,N_22444);
and U22913 (N_22913,N_22364,N_22199);
nor U22914 (N_22914,N_22049,N_22483);
nor U22915 (N_22915,N_22098,N_22499);
nor U22916 (N_22916,N_22120,N_22184);
nand U22917 (N_22917,N_22400,N_22259);
nor U22918 (N_22918,N_22174,N_22106);
nor U22919 (N_22919,N_22026,N_22458);
and U22920 (N_22920,N_22313,N_22335);
xor U22921 (N_22921,N_22016,N_22050);
xnor U22922 (N_22922,N_22236,N_22021);
and U22923 (N_22923,N_22203,N_22136);
nor U22924 (N_22924,N_22396,N_22360);
nor U22925 (N_22925,N_22192,N_22491);
xor U22926 (N_22926,N_22478,N_22494);
or U22927 (N_22927,N_22462,N_22443);
and U22928 (N_22928,N_22252,N_22049);
xor U22929 (N_22929,N_22325,N_22478);
xnor U22930 (N_22930,N_22293,N_22048);
nand U22931 (N_22931,N_22259,N_22446);
nand U22932 (N_22932,N_22113,N_22379);
nor U22933 (N_22933,N_22457,N_22071);
nand U22934 (N_22934,N_22253,N_22416);
nor U22935 (N_22935,N_22459,N_22326);
or U22936 (N_22936,N_22367,N_22169);
or U22937 (N_22937,N_22015,N_22277);
and U22938 (N_22938,N_22287,N_22459);
xor U22939 (N_22939,N_22329,N_22068);
xor U22940 (N_22940,N_22235,N_22163);
nand U22941 (N_22941,N_22094,N_22171);
xnor U22942 (N_22942,N_22275,N_22335);
xor U22943 (N_22943,N_22101,N_22245);
nand U22944 (N_22944,N_22136,N_22242);
nor U22945 (N_22945,N_22133,N_22113);
xor U22946 (N_22946,N_22143,N_22121);
and U22947 (N_22947,N_22069,N_22173);
or U22948 (N_22948,N_22480,N_22499);
xor U22949 (N_22949,N_22037,N_22270);
xor U22950 (N_22950,N_22200,N_22280);
or U22951 (N_22951,N_22198,N_22063);
or U22952 (N_22952,N_22437,N_22060);
and U22953 (N_22953,N_22498,N_22007);
nand U22954 (N_22954,N_22274,N_22265);
or U22955 (N_22955,N_22127,N_22490);
nor U22956 (N_22956,N_22059,N_22417);
or U22957 (N_22957,N_22314,N_22088);
nand U22958 (N_22958,N_22278,N_22395);
and U22959 (N_22959,N_22146,N_22215);
or U22960 (N_22960,N_22063,N_22056);
xnor U22961 (N_22961,N_22427,N_22390);
or U22962 (N_22962,N_22309,N_22106);
and U22963 (N_22963,N_22351,N_22236);
nand U22964 (N_22964,N_22224,N_22126);
and U22965 (N_22965,N_22165,N_22115);
nand U22966 (N_22966,N_22401,N_22196);
nand U22967 (N_22967,N_22279,N_22291);
xor U22968 (N_22968,N_22315,N_22284);
xor U22969 (N_22969,N_22101,N_22434);
nor U22970 (N_22970,N_22436,N_22129);
nor U22971 (N_22971,N_22067,N_22201);
and U22972 (N_22972,N_22297,N_22252);
and U22973 (N_22973,N_22005,N_22433);
or U22974 (N_22974,N_22132,N_22411);
nor U22975 (N_22975,N_22477,N_22151);
nor U22976 (N_22976,N_22247,N_22447);
nand U22977 (N_22977,N_22428,N_22100);
nor U22978 (N_22978,N_22275,N_22012);
xor U22979 (N_22979,N_22299,N_22448);
or U22980 (N_22980,N_22462,N_22192);
and U22981 (N_22981,N_22223,N_22227);
and U22982 (N_22982,N_22323,N_22337);
xor U22983 (N_22983,N_22319,N_22300);
nand U22984 (N_22984,N_22062,N_22172);
or U22985 (N_22985,N_22185,N_22025);
or U22986 (N_22986,N_22462,N_22165);
nor U22987 (N_22987,N_22110,N_22346);
or U22988 (N_22988,N_22120,N_22035);
nor U22989 (N_22989,N_22000,N_22175);
nand U22990 (N_22990,N_22481,N_22214);
and U22991 (N_22991,N_22217,N_22145);
or U22992 (N_22992,N_22363,N_22109);
xor U22993 (N_22993,N_22022,N_22159);
nor U22994 (N_22994,N_22005,N_22415);
nand U22995 (N_22995,N_22034,N_22051);
or U22996 (N_22996,N_22240,N_22471);
nor U22997 (N_22997,N_22463,N_22471);
or U22998 (N_22998,N_22087,N_22017);
xor U22999 (N_22999,N_22388,N_22321);
nand U23000 (N_23000,N_22871,N_22525);
nor U23001 (N_23001,N_22734,N_22612);
nor U23002 (N_23002,N_22873,N_22717);
nor U23003 (N_23003,N_22941,N_22546);
or U23004 (N_23004,N_22945,N_22649);
nor U23005 (N_23005,N_22549,N_22831);
nand U23006 (N_23006,N_22564,N_22622);
or U23007 (N_23007,N_22597,N_22804);
nor U23008 (N_23008,N_22962,N_22805);
or U23009 (N_23009,N_22872,N_22868);
nand U23010 (N_23010,N_22814,N_22757);
nand U23011 (N_23011,N_22981,N_22802);
nor U23012 (N_23012,N_22664,N_22931);
xnor U23013 (N_23013,N_22613,N_22551);
nand U23014 (N_23014,N_22921,N_22808);
nand U23015 (N_23015,N_22889,N_22663);
and U23016 (N_23016,N_22771,N_22654);
and U23017 (N_23017,N_22997,N_22798);
or U23018 (N_23018,N_22888,N_22518);
or U23019 (N_23019,N_22595,N_22932);
xor U23020 (N_23020,N_22676,N_22530);
xor U23021 (N_23021,N_22956,N_22630);
nor U23022 (N_23022,N_22965,N_22503);
xnor U23023 (N_23023,N_22538,N_22713);
and U23024 (N_23024,N_22540,N_22864);
and U23025 (N_23025,N_22780,N_22898);
nand U23026 (N_23026,N_22502,N_22510);
and U23027 (N_23027,N_22924,N_22995);
nor U23028 (N_23028,N_22821,N_22991);
nor U23029 (N_23029,N_22883,N_22841);
xnor U23030 (N_23030,N_22903,N_22854);
nand U23031 (N_23031,N_22975,N_22812);
or U23032 (N_23032,N_22880,N_22671);
nand U23033 (N_23033,N_22770,N_22838);
xnor U23034 (N_23034,N_22970,N_22759);
nor U23035 (N_23035,N_22547,N_22543);
xnor U23036 (N_23036,N_22886,N_22857);
and U23037 (N_23037,N_22747,N_22588);
nor U23038 (N_23038,N_22946,N_22721);
and U23039 (N_23039,N_22665,N_22755);
nor U23040 (N_23040,N_22837,N_22668);
and U23041 (N_23041,N_22620,N_22811);
nor U23042 (N_23042,N_22901,N_22840);
or U23043 (N_23043,N_22876,N_22983);
or U23044 (N_23044,N_22650,N_22586);
xor U23045 (N_23045,N_22528,N_22603);
xor U23046 (N_23046,N_22777,N_22584);
xor U23047 (N_23047,N_22589,N_22992);
nand U23048 (N_23048,N_22590,N_22953);
nand U23049 (N_23049,N_22714,N_22509);
and U23050 (N_23050,N_22527,N_22977);
nand U23051 (N_23051,N_22646,N_22516);
xnor U23052 (N_23052,N_22940,N_22591);
nand U23053 (N_23053,N_22918,N_22716);
or U23054 (N_23054,N_22958,N_22756);
nor U23055 (N_23055,N_22675,N_22696);
nand U23056 (N_23056,N_22938,N_22627);
or U23057 (N_23057,N_22999,N_22881);
or U23058 (N_23058,N_22596,N_22608);
nor U23059 (N_23059,N_22673,N_22599);
or U23060 (N_23060,N_22715,N_22799);
xnor U23061 (N_23061,N_22643,N_22521);
nand U23062 (N_23062,N_22925,N_22775);
nand U23063 (N_23063,N_22683,N_22951);
nand U23064 (N_23064,N_22607,N_22763);
nor U23065 (N_23065,N_22842,N_22849);
xor U23066 (N_23066,N_22576,N_22916);
nor U23067 (N_23067,N_22519,N_22574);
and U23068 (N_23068,N_22582,N_22762);
nor U23069 (N_23069,N_22993,N_22619);
and U23070 (N_23070,N_22726,N_22966);
and U23071 (N_23071,N_22973,N_22667);
xnor U23072 (N_23072,N_22990,N_22691);
xor U23073 (N_23073,N_22797,N_22542);
and U23074 (N_23074,N_22895,N_22557);
nand U23075 (N_23075,N_22988,N_22580);
and U23076 (N_23076,N_22978,N_22768);
and U23077 (N_23077,N_22861,N_22955);
and U23078 (N_23078,N_22526,N_22602);
xor U23079 (N_23079,N_22501,N_22642);
nand U23080 (N_23080,N_22529,N_22891);
xnor U23081 (N_23081,N_22754,N_22570);
and U23082 (N_23082,N_22915,N_22740);
or U23083 (N_23083,N_22606,N_22855);
xor U23084 (N_23084,N_22885,N_22914);
nand U23085 (N_23085,N_22897,N_22534);
xor U23086 (N_23086,N_22954,N_22784);
nand U23087 (N_23087,N_22820,N_22893);
or U23088 (N_23088,N_22567,N_22609);
nor U23089 (N_23089,N_22523,N_22611);
and U23090 (N_23090,N_22677,N_22544);
or U23091 (N_23091,N_22794,N_22823);
nand U23092 (N_23092,N_22745,N_22628);
xor U23093 (N_23093,N_22598,N_22593);
nor U23094 (N_23094,N_22929,N_22658);
nor U23095 (N_23095,N_22578,N_22760);
nand U23096 (N_23096,N_22749,N_22788);
xnor U23097 (N_23097,N_22877,N_22692);
nand U23098 (N_23098,N_22682,N_22699);
nor U23099 (N_23099,N_22847,N_22653);
and U23100 (N_23100,N_22919,N_22987);
and U23101 (N_23101,N_22913,N_22552);
or U23102 (N_23102,N_22651,N_22824);
nand U23103 (N_23103,N_22670,N_22566);
or U23104 (N_23104,N_22739,N_22979);
and U23105 (N_23105,N_22513,N_22705);
or U23106 (N_23106,N_22936,N_22697);
nand U23107 (N_23107,N_22884,N_22875);
nand U23108 (N_23108,N_22656,N_22907);
xnor U23109 (N_23109,N_22772,N_22822);
or U23110 (N_23110,N_22944,N_22695);
or U23111 (N_23111,N_22927,N_22985);
and U23112 (N_23112,N_22815,N_22569);
and U23113 (N_23113,N_22894,N_22572);
or U23114 (N_23114,N_22746,N_22900);
and U23115 (N_23115,N_22718,N_22594);
or U23116 (N_23116,N_22581,N_22935);
nand U23117 (N_23117,N_22563,N_22730);
or U23118 (N_23118,N_22723,N_22733);
nand U23119 (N_23119,N_22912,N_22700);
nor U23120 (N_23120,N_22774,N_22605);
nand U23121 (N_23121,N_22858,N_22865);
or U23122 (N_23122,N_22910,N_22843);
nor U23123 (N_23123,N_22948,N_22867);
nand U23124 (N_23124,N_22905,N_22852);
or U23125 (N_23125,N_22947,N_22752);
nor U23126 (N_23126,N_22618,N_22790);
or U23127 (N_23127,N_22796,N_22587);
nand U23128 (N_23128,N_22922,N_22565);
nor U23129 (N_23129,N_22920,N_22636);
and U23130 (N_23130,N_22982,N_22748);
or U23131 (N_23131,N_22556,N_22735);
and U23132 (N_23132,N_22681,N_22825);
xnor U23133 (N_23133,N_22785,N_22960);
xnor U23134 (N_23134,N_22522,N_22737);
nand U23135 (N_23135,N_22728,N_22515);
xor U23136 (N_23136,N_22698,N_22614);
nand U23137 (N_23137,N_22952,N_22776);
nand U23138 (N_23138,N_22839,N_22917);
xor U23139 (N_23139,N_22629,N_22537);
xor U23140 (N_23140,N_22809,N_22957);
nand U23141 (N_23141,N_22610,N_22583);
or U23142 (N_23142,N_22719,N_22859);
nor U23143 (N_23143,N_22517,N_22701);
and U23144 (N_23144,N_22795,N_22791);
and U23145 (N_23145,N_22703,N_22866);
nor U23146 (N_23146,N_22758,N_22661);
and U23147 (N_23147,N_22638,N_22617);
nor U23148 (N_23148,N_22689,N_22783);
nand U23149 (N_23149,N_22626,N_22647);
or U23150 (N_23150,N_22835,N_22878);
nor U23151 (N_23151,N_22833,N_22969);
xnor U23152 (N_23152,N_22856,N_22562);
or U23153 (N_23153,N_22706,N_22555);
xnor U23154 (N_23154,N_22633,N_22694);
nand U23155 (N_23155,N_22744,N_22887);
nor U23156 (N_23156,N_22961,N_22813);
nor U23157 (N_23157,N_22819,N_22968);
xnor U23158 (N_23158,N_22624,N_22686);
or U23159 (N_23159,N_22707,N_22926);
nor U23160 (N_23160,N_22980,N_22666);
and U23161 (N_23161,N_22687,N_22906);
nand U23162 (N_23162,N_22964,N_22950);
xnor U23163 (N_23163,N_22930,N_22680);
and U23164 (N_23164,N_22769,N_22976);
nor U23165 (N_23165,N_22767,N_22817);
xor U23166 (N_23166,N_22635,N_22967);
and U23167 (N_23167,N_22939,N_22810);
and U23168 (N_23168,N_22800,N_22508);
and U23169 (N_23169,N_22781,N_22934);
and U23170 (N_23170,N_22690,N_22787);
or U23171 (N_23171,N_22807,N_22520);
or U23172 (N_23172,N_22826,N_22545);
or U23173 (N_23173,N_22860,N_22933);
or U23174 (N_23174,N_22848,N_22585);
or U23175 (N_23175,N_22688,N_22778);
xnor U23176 (N_23176,N_22550,N_22561);
nand U23177 (N_23177,N_22674,N_22908);
xor U23178 (N_23178,N_22616,N_22773);
xnor U23179 (N_23179,N_22869,N_22601);
nand U23180 (N_23180,N_22725,N_22644);
nor U23181 (N_23181,N_22986,N_22657);
and U23182 (N_23182,N_22829,N_22511);
and U23183 (N_23183,N_22577,N_22949);
nor U23184 (N_23184,N_22963,N_22732);
or U23185 (N_23185,N_22604,N_22500);
or U23186 (N_23186,N_22684,N_22766);
or U23187 (N_23187,N_22708,N_22792);
nor U23188 (N_23188,N_22803,N_22742);
nor U23189 (N_23189,N_22853,N_22937);
or U23190 (N_23190,N_22789,N_22539);
nand U23191 (N_23191,N_22541,N_22729);
and U23192 (N_23192,N_22532,N_22892);
or U23193 (N_23193,N_22943,N_22558);
and U23194 (N_23194,N_22669,N_22846);
or U23195 (N_23195,N_22724,N_22639);
or U23196 (N_23196,N_22720,N_22514);
nand U23197 (N_23197,N_22998,N_22709);
or U23198 (N_23198,N_22712,N_22896);
nand U23199 (N_23199,N_22631,N_22959);
and U23200 (N_23200,N_22652,N_22818);
nand U23201 (N_23201,N_22641,N_22524);
or U23202 (N_23202,N_22575,N_22710);
and U23203 (N_23203,N_22989,N_22984);
or U23204 (N_23204,N_22994,N_22904);
nor U23205 (N_23205,N_22844,N_22659);
xnor U23206 (N_23206,N_22909,N_22816);
nor U23207 (N_23207,N_22573,N_22741);
or U23208 (N_23208,N_22743,N_22648);
nor U23209 (N_23209,N_22506,N_22996);
nor U23210 (N_23210,N_22579,N_22536);
nand U23211 (N_23211,N_22704,N_22793);
and U23212 (N_23212,N_22640,N_22874);
and U23213 (N_23213,N_22764,N_22902);
or U23214 (N_23214,N_22890,N_22845);
xor U23215 (N_23215,N_22685,N_22702);
nor U23216 (N_23216,N_22751,N_22850);
xnor U23217 (N_23217,N_22834,N_22832);
nand U23218 (N_23218,N_22634,N_22899);
or U23219 (N_23219,N_22600,N_22806);
nor U23220 (N_23220,N_22801,N_22731);
nor U23221 (N_23221,N_22559,N_22779);
and U23222 (N_23222,N_22554,N_22765);
nand U23223 (N_23223,N_22882,N_22851);
nand U23224 (N_23224,N_22753,N_22655);
nand U23225 (N_23225,N_22660,N_22507);
nand U23226 (N_23226,N_22782,N_22828);
nand U23227 (N_23227,N_22531,N_22974);
and U23228 (N_23228,N_22879,N_22727);
nand U23229 (N_23229,N_22592,N_22560);
or U23230 (N_23230,N_22911,N_22662);
nand U23231 (N_23231,N_22533,N_22693);
xor U23232 (N_23232,N_22711,N_22645);
nor U23233 (N_23233,N_22615,N_22568);
nand U23234 (N_23234,N_22571,N_22722);
nor U23235 (N_23235,N_22621,N_22761);
nor U23236 (N_23236,N_22971,N_22827);
xor U23237 (N_23237,N_22870,N_22830);
or U23238 (N_23238,N_22862,N_22679);
nor U23239 (N_23239,N_22625,N_22863);
and U23240 (N_23240,N_22942,N_22672);
or U23241 (N_23241,N_22623,N_22535);
or U23242 (N_23242,N_22928,N_22738);
nand U23243 (N_23243,N_22750,N_22512);
or U23244 (N_23244,N_22637,N_22736);
and U23245 (N_23245,N_22836,N_22786);
and U23246 (N_23246,N_22678,N_22632);
and U23247 (N_23247,N_22504,N_22923);
and U23248 (N_23248,N_22553,N_22548);
xor U23249 (N_23249,N_22505,N_22972);
or U23250 (N_23250,N_22690,N_22765);
or U23251 (N_23251,N_22555,N_22750);
nor U23252 (N_23252,N_22857,N_22539);
xor U23253 (N_23253,N_22969,N_22979);
nand U23254 (N_23254,N_22720,N_22896);
or U23255 (N_23255,N_22896,N_22657);
xnor U23256 (N_23256,N_22695,N_22595);
xor U23257 (N_23257,N_22962,N_22637);
or U23258 (N_23258,N_22764,N_22659);
and U23259 (N_23259,N_22820,N_22689);
nor U23260 (N_23260,N_22857,N_22893);
nor U23261 (N_23261,N_22596,N_22593);
or U23262 (N_23262,N_22586,N_22564);
nand U23263 (N_23263,N_22721,N_22954);
and U23264 (N_23264,N_22954,N_22812);
xnor U23265 (N_23265,N_22969,N_22769);
or U23266 (N_23266,N_22640,N_22623);
xor U23267 (N_23267,N_22623,N_22674);
or U23268 (N_23268,N_22513,N_22525);
or U23269 (N_23269,N_22802,N_22999);
and U23270 (N_23270,N_22876,N_22523);
nor U23271 (N_23271,N_22816,N_22566);
xnor U23272 (N_23272,N_22863,N_22739);
nor U23273 (N_23273,N_22575,N_22719);
xor U23274 (N_23274,N_22632,N_22656);
xnor U23275 (N_23275,N_22544,N_22821);
and U23276 (N_23276,N_22966,N_22676);
xnor U23277 (N_23277,N_22724,N_22515);
and U23278 (N_23278,N_22665,N_22824);
and U23279 (N_23279,N_22592,N_22672);
and U23280 (N_23280,N_22552,N_22664);
and U23281 (N_23281,N_22585,N_22836);
and U23282 (N_23282,N_22937,N_22730);
or U23283 (N_23283,N_22910,N_22914);
nor U23284 (N_23284,N_22702,N_22929);
and U23285 (N_23285,N_22504,N_22875);
nand U23286 (N_23286,N_22958,N_22683);
nor U23287 (N_23287,N_22989,N_22877);
or U23288 (N_23288,N_22759,N_22840);
xnor U23289 (N_23289,N_22916,N_22636);
or U23290 (N_23290,N_22676,N_22577);
or U23291 (N_23291,N_22779,N_22858);
and U23292 (N_23292,N_22996,N_22744);
and U23293 (N_23293,N_22614,N_22521);
or U23294 (N_23294,N_22931,N_22750);
nor U23295 (N_23295,N_22640,N_22787);
or U23296 (N_23296,N_22710,N_22950);
nor U23297 (N_23297,N_22852,N_22615);
nand U23298 (N_23298,N_22588,N_22974);
xor U23299 (N_23299,N_22543,N_22581);
or U23300 (N_23300,N_22854,N_22500);
xnor U23301 (N_23301,N_22762,N_22540);
xnor U23302 (N_23302,N_22802,N_22709);
xnor U23303 (N_23303,N_22609,N_22977);
xnor U23304 (N_23304,N_22945,N_22519);
xor U23305 (N_23305,N_22622,N_22562);
xor U23306 (N_23306,N_22882,N_22667);
nor U23307 (N_23307,N_22994,N_22808);
and U23308 (N_23308,N_22975,N_22925);
nor U23309 (N_23309,N_22523,N_22930);
and U23310 (N_23310,N_22877,N_22603);
nand U23311 (N_23311,N_22800,N_22519);
nand U23312 (N_23312,N_22847,N_22596);
xnor U23313 (N_23313,N_22964,N_22927);
nand U23314 (N_23314,N_22821,N_22739);
nor U23315 (N_23315,N_22820,N_22880);
and U23316 (N_23316,N_22601,N_22773);
and U23317 (N_23317,N_22851,N_22810);
xor U23318 (N_23318,N_22549,N_22888);
and U23319 (N_23319,N_22706,N_22678);
or U23320 (N_23320,N_22936,N_22563);
nor U23321 (N_23321,N_22763,N_22603);
and U23322 (N_23322,N_22529,N_22904);
and U23323 (N_23323,N_22544,N_22772);
nor U23324 (N_23324,N_22587,N_22694);
nor U23325 (N_23325,N_22611,N_22609);
or U23326 (N_23326,N_22827,N_22818);
xnor U23327 (N_23327,N_22620,N_22614);
xnor U23328 (N_23328,N_22945,N_22687);
and U23329 (N_23329,N_22961,N_22823);
or U23330 (N_23330,N_22872,N_22867);
and U23331 (N_23331,N_22626,N_22838);
nor U23332 (N_23332,N_22729,N_22721);
nand U23333 (N_23333,N_22634,N_22927);
or U23334 (N_23334,N_22520,N_22577);
xnor U23335 (N_23335,N_22706,N_22631);
nand U23336 (N_23336,N_22842,N_22781);
xnor U23337 (N_23337,N_22619,N_22605);
or U23338 (N_23338,N_22548,N_22593);
nor U23339 (N_23339,N_22608,N_22652);
and U23340 (N_23340,N_22747,N_22580);
xor U23341 (N_23341,N_22723,N_22939);
nand U23342 (N_23342,N_22944,N_22612);
nand U23343 (N_23343,N_22993,N_22505);
nor U23344 (N_23344,N_22928,N_22982);
and U23345 (N_23345,N_22714,N_22844);
nand U23346 (N_23346,N_22501,N_22620);
and U23347 (N_23347,N_22609,N_22985);
xnor U23348 (N_23348,N_22641,N_22807);
nand U23349 (N_23349,N_22683,N_22751);
and U23350 (N_23350,N_22854,N_22912);
nand U23351 (N_23351,N_22511,N_22985);
and U23352 (N_23352,N_22859,N_22587);
xor U23353 (N_23353,N_22999,N_22565);
or U23354 (N_23354,N_22700,N_22751);
xnor U23355 (N_23355,N_22647,N_22697);
and U23356 (N_23356,N_22583,N_22910);
nand U23357 (N_23357,N_22742,N_22738);
or U23358 (N_23358,N_22785,N_22852);
and U23359 (N_23359,N_22630,N_22796);
nand U23360 (N_23360,N_22556,N_22716);
or U23361 (N_23361,N_22989,N_22708);
nand U23362 (N_23362,N_22522,N_22947);
nor U23363 (N_23363,N_22580,N_22937);
xor U23364 (N_23364,N_22770,N_22707);
nand U23365 (N_23365,N_22790,N_22839);
and U23366 (N_23366,N_22774,N_22942);
and U23367 (N_23367,N_22794,N_22645);
xnor U23368 (N_23368,N_22946,N_22829);
nor U23369 (N_23369,N_22826,N_22556);
nor U23370 (N_23370,N_22850,N_22642);
nand U23371 (N_23371,N_22522,N_22876);
xor U23372 (N_23372,N_22687,N_22555);
nor U23373 (N_23373,N_22725,N_22960);
nor U23374 (N_23374,N_22974,N_22983);
or U23375 (N_23375,N_22764,N_22816);
and U23376 (N_23376,N_22826,N_22536);
or U23377 (N_23377,N_22721,N_22936);
or U23378 (N_23378,N_22942,N_22814);
nand U23379 (N_23379,N_22530,N_22809);
or U23380 (N_23380,N_22972,N_22900);
and U23381 (N_23381,N_22710,N_22824);
or U23382 (N_23382,N_22897,N_22617);
nand U23383 (N_23383,N_22602,N_22684);
nand U23384 (N_23384,N_22690,N_22830);
nand U23385 (N_23385,N_22877,N_22627);
nand U23386 (N_23386,N_22661,N_22560);
xnor U23387 (N_23387,N_22550,N_22620);
and U23388 (N_23388,N_22560,N_22790);
nand U23389 (N_23389,N_22637,N_22558);
xor U23390 (N_23390,N_22584,N_22612);
nand U23391 (N_23391,N_22814,N_22789);
xnor U23392 (N_23392,N_22500,N_22658);
nor U23393 (N_23393,N_22777,N_22925);
and U23394 (N_23394,N_22637,N_22565);
nand U23395 (N_23395,N_22835,N_22652);
or U23396 (N_23396,N_22690,N_22653);
nand U23397 (N_23397,N_22872,N_22642);
or U23398 (N_23398,N_22835,N_22651);
or U23399 (N_23399,N_22552,N_22926);
or U23400 (N_23400,N_22797,N_22742);
or U23401 (N_23401,N_22583,N_22619);
or U23402 (N_23402,N_22528,N_22784);
nor U23403 (N_23403,N_22742,N_22599);
nor U23404 (N_23404,N_22863,N_22798);
nor U23405 (N_23405,N_22966,N_22865);
or U23406 (N_23406,N_22591,N_22826);
and U23407 (N_23407,N_22722,N_22945);
nand U23408 (N_23408,N_22962,N_22927);
or U23409 (N_23409,N_22753,N_22653);
xor U23410 (N_23410,N_22676,N_22513);
xnor U23411 (N_23411,N_22714,N_22864);
or U23412 (N_23412,N_22790,N_22519);
xnor U23413 (N_23413,N_22514,N_22984);
or U23414 (N_23414,N_22788,N_22592);
nor U23415 (N_23415,N_22985,N_22545);
xor U23416 (N_23416,N_22683,N_22586);
or U23417 (N_23417,N_22889,N_22530);
or U23418 (N_23418,N_22988,N_22668);
or U23419 (N_23419,N_22720,N_22775);
nor U23420 (N_23420,N_22751,N_22702);
nand U23421 (N_23421,N_22655,N_22820);
or U23422 (N_23422,N_22866,N_22628);
xnor U23423 (N_23423,N_22829,N_22539);
and U23424 (N_23424,N_22764,N_22585);
and U23425 (N_23425,N_22555,N_22534);
nand U23426 (N_23426,N_22614,N_22579);
nand U23427 (N_23427,N_22948,N_22816);
or U23428 (N_23428,N_22652,N_22568);
nand U23429 (N_23429,N_22564,N_22874);
and U23430 (N_23430,N_22595,N_22580);
or U23431 (N_23431,N_22787,N_22546);
or U23432 (N_23432,N_22805,N_22508);
nand U23433 (N_23433,N_22931,N_22955);
nand U23434 (N_23434,N_22996,N_22726);
nand U23435 (N_23435,N_22824,N_22628);
xor U23436 (N_23436,N_22527,N_22652);
nor U23437 (N_23437,N_22751,N_22640);
and U23438 (N_23438,N_22608,N_22973);
nand U23439 (N_23439,N_22923,N_22690);
nor U23440 (N_23440,N_22571,N_22636);
or U23441 (N_23441,N_22874,N_22989);
nand U23442 (N_23442,N_22967,N_22984);
nand U23443 (N_23443,N_22601,N_22833);
xnor U23444 (N_23444,N_22538,N_22652);
or U23445 (N_23445,N_22785,N_22887);
nand U23446 (N_23446,N_22627,N_22930);
nand U23447 (N_23447,N_22886,N_22778);
xor U23448 (N_23448,N_22861,N_22792);
nor U23449 (N_23449,N_22853,N_22753);
xor U23450 (N_23450,N_22869,N_22622);
nand U23451 (N_23451,N_22594,N_22520);
nand U23452 (N_23452,N_22540,N_22901);
and U23453 (N_23453,N_22861,N_22982);
and U23454 (N_23454,N_22717,N_22516);
and U23455 (N_23455,N_22811,N_22885);
and U23456 (N_23456,N_22987,N_22582);
nand U23457 (N_23457,N_22757,N_22564);
xor U23458 (N_23458,N_22890,N_22588);
nand U23459 (N_23459,N_22676,N_22954);
xor U23460 (N_23460,N_22657,N_22995);
and U23461 (N_23461,N_22710,N_22971);
nor U23462 (N_23462,N_22655,N_22971);
nand U23463 (N_23463,N_22856,N_22602);
and U23464 (N_23464,N_22775,N_22954);
xnor U23465 (N_23465,N_22741,N_22998);
xnor U23466 (N_23466,N_22539,N_22827);
and U23467 (N_23467,N_22600,N_22543);
and U23468 (N_23468,N_22699,N_22795);
and U23469 (N_23469,N_22625,N_22900);
nor U23470 (N_23470,N_22760,N_22721);
or U23471 (N_23471,N_22833,N_22719);
xnor U23472 (N_23472,N_22641,N_22635);
and U23473 (N_23473,N_22954,N_22853);
nor U23474 (N_23474,N_22510,N_22557);
nor U23475 (N_23475,N_22930,N_22737);
and U23476 (N_23476,N_22964,N_22577);
or U23477 (N_23477,N_22832,N_22625);
xnor U23478 (N_23478,N_22971,N_22599);
nor U23479 (N_23479,N_22723,N_22894);
or U23480 (N_23480,N_22775,N_22560);
or U23481 (N_23481,N_22541,N_22687);
nand U23482 (N_23482,N_22918,N_22523);
nor U23483 (N_23483,N_22620,N_22877);
nor U23484 (N_23484,N_22875,N_22724);
xor U23485 (N_23485,N_22748,N_22967);
xor U23486 (N_23486,N_22587,N_22880);
xnor U23487 (N_23487,N_22881,N_22687);
nor U23488 (N_23488,N_22889,N_22571);
nand U23489 (N_23489,N_22796,N_22570);
nand U23490 (N_23490,N_22567,N_22764);
and U23491 (N_23491,N_22694,N_22900);
xnor U23492 (N_23492,N_22834,N_22601);
nand U23493 (N_23493,N_22538,N_22643);
and U23494 (N_23494,N_22689,N_22620);
or U23495 (N_23495,N_22895,N_22901);
and U23496 (N_23496,N_22649,N_22583);
nor U23497 (N_23497,N_22640,N_22895);
nand U23498 (N_23498,N_22784,N_22516);
nor U23499 (N_23499,N_22588,N_22791);
xor U23500 (N_23500,N_23498,N_23153);
xor U23501 (N_23501,N_23390,N_23227);
nand U23502 (N_23502,N_23010,N_23269);
nand U23503 (N_23503,N_23161,N_23294);
and U23504 (N_23504,N_23168,N_23473);
and U23505 (N_23505,N_23011,N_23013);
nor U23506 (N_23506,N_23411,N_23214);
or U23507 (N_23507,N_23148,N_23375);
and U23508 (N_23508,N_23014,N_23402);
and U23509 (N_23509,N_23379,N_23271);
xnor U23510 (N_23510,N_23196,N_23239);
nor U23511 (N_23511,N_23453,N_23490);
nor U23512 (N_23512,N_23458,N_23325);
xnor U23513 (N_23513,N_23179,N_23219);
nor U23514 (N_23514,N_23349,N_23182);
xnor U23515 (N_23515,N_23064,N_23306);
and U23516 (N_23516,N_23039,N_23202);
nand U23517 (N_23517,N_23494,N_23304);
xor U23518 (N_23518,N_23472,N_23491);
xor U23519 (N_23519,N_23287,N_23428);
and U23520 (N_23520,N_23160,N_23144);
and U23521 (N_23521,N_23436,N_23055);
and U23522 (N_23522,N_23059,N_23340);
or U23523 (N_23523,N_23067,N_23429);
and U23524 (N_23524,N_23025,N_23001);
nand U23525 (N_23525,N_23215,N_23417);
nor U23526 (N_23526,N_23102,N_23074);
or U23527 (N_23527,N_23298,N_23286);
xor U23528 (N_23528,N_23437,N_23370);
nor U23529 (N_23529,N_23068,N_23103);
and U23530 (N_23530,N_23289,N_23145);
or U23531 (N_23531,N_23335,N_23203);
nand U23532 (N_23532,N_23445,N_23091);
and U23533 (N_23533,N_23254,N_23365);
nand U23534 (N_23534,N_23079,N_23044);
and U23535 (N_23535,N_23303,N_23112);
xnor U23536 (N_23536,N_23355,N_23328);
or U23537 (N_23537,N_23108,N_23166);
and U23538 (N_23538,N_23190,N_23308);
nor U23539 (N_23539,N_23027,N_23272);
nand U23540 (N_23540,N_23213,N_23047);
and U23541 (N_23541,N_23075,N_23195);
or U23542 (N_23542,N_23018,N_23362);
and U23543 (N_23543,N_23493,N_23406);
nand U23544 (N_23544,N_23371,N_23261);
xor U23545 (N_23545,N_23101,N_23149);
and U23546 (N_23546,N_23206,N_23124);
nor U23547 (N_23547,N_23095,N_23357);
xor U23548 (N_23548,N_23348,N_23209);
xnor U23549 (N_23549,N_23127,N_23433);
nor U23550 (N_23550,N_23143,N_23031);
xor U23551 (N_23551,N_23255,N_23300);
nor U23552 (N_23552,N_23360,N_23029);
nor U23553 (N_23553,N_23016,N_23041);
or U23554 (N_23554,N_23235,N_23457);
nor U23555 (N_23555,N_23356,N_23056);
xor U23556 (N_23556,N_23481,N_23234);
xor U23557 (N_23557,N_23434,N_23169);
nand U23558 (N_23558,N_23109,N_23054);
nor U23559 (N_23559,N_23183,N_23412);
nor U23560 (N_23560,N_23347,N_23447);
nor U23561 (N_23561,N_23024,N_23497);
or U23562 (N_23562,N_23307,N_23413);
or U23563 (N_23563,N_23464,N_23021);
nand U23564 (N_23564,N_23045,N_23023);
nand U23565 (N_23565,N_23084,N_23291);
or U23566 (N_23566,N_23345,N_23346);
xor U23567 (N_23567,N_23042,N_23100);
nand U23568 (N_23568,N_23443,N_23128);
and U23569 (N_23569,N_23057,N_23053);
nor U23570 (N_23570,N_23488,N_23405);
or U23571 (N_23571,N_23009,N_23086);
xor U23572 (N_23572,N_23185,N_23270);
nor U23573 (N_23573,N_23395,N_23380);
nand U23574 (N_23574,N_23164,N_23050);
xor U23575 (N_23575,N_23142,N_23424);
xor U23576 (N_23576,N_23275,N_23006);
or U23577 (N_23577,N_23394,N_23423);
or U23578 (N_23578,N_23430,N_23341);
or U23579 (N_23579,N_23118,N_23043);
nor U23580 (N_23580,N_23037,N_23425);
nor U23581 (N_23581,N_23312,N_23337);
xnor U23582 (N_23582,N_23281,N_23140);
xnor U23583 (N_23583,N_23333,N_23094);
nor U23584 (N_23584,N_23225,N_23210);
or U23585 (N_23585,N_23163,N_23280);
and U23586 (N_23586,N_23061,N_23125);
and U23587 (N_23587,N_23080,N_23354);
and U23588 (N_23588,N_23141,N_23276);
or U23589 (N_23589,N_23231,N_23301);
nor U23590 (N_23590,N_23454,N_23052);
xor U23591 (N_23591,N_23237,N_23197);
or U23592 (N_23592,N_23320,N_23489);
and U23593 (N_23593,N_23176,N_23478);
or U23594 (N_23594,N_23186,N_23066);
nor U23595 (N_23595,N_23322,N_23422);
and U23596 (N_23596,N_23170,N_23278);
and U23597 (N_23597,N_23022,N_23463);
nor U23598 (N_23598,N_23465,N_23191);
nand U23599 (N_23599,N_23116,N_23381);
and U23600 (N_23600,N_23477,N_23093);
nand U23601 (N_23601,N_23467,N_23321);
nor U23602 (N_23602,N_23104,N_23446);
nor U23603 (N_23603,N_23073,N_23189);
and U23604 (N_23604,N_23482,N_23266);
nand U23605 (N_23605,N_23311,N_23373);
nand U23606 (N_23606,N_23499,N_23288);
nor U23607 (N_23607,N_23028,N_23290);
nor U23608 (N_23608,N_23442,N_23076);
or U23609 (N_23609,N_23327,N_23259);
xnor U23610 (N_23610,N_23096,N_23441);
and U23611 (N_23611,N_23451,N_23343);
nor U23612 (N_23612,N_23211,N_23462);
nor U23613 (N_23613,N_23178,N_23471);
and U23614 (N_23614,N_23263,N_23257);
nand U23615 (N_23615,N_23426,N_23097);
and U23616 (N_23616,N_23363,N_23245);
nand U23617 (N_23617,N_23172,N_23344);
or U23618 (N_23618,N_23366,N_23331);
and U23619 (N_23619,N_23040,N_23114);
nand U23620 (N_23620,N_23194,N_23297);
nand U23621 (N_23621,N_23110,N_23299);
xnor U23622 (N_23622,N_23469,N_23475);
xnor U23623 (N_23623,N_23256,N_23049);
and U23624 (N_23624,N_23087,N_23158);
nor U23625 (N_23625,N_23285,N_23393);
nor U23626 (N_23626,N_23089,N_23435);
xnor U23627 (N_23627,N_23032,N_23007);
xnor U23628 (N_23628,N_23200,N_23199);
nor U23629 (N_23629,N_23000,N_23217);
or U23630 (N_23630,N_23247,N_23338);
and U23631 (N_23631,N_23487,N_23420);
xnor U23632 (N_23632,N_23293,N_23137);
nand U23633 (N_23633,N_23175,N_23314);
nand U23634 (N_23634,N_23171,N_23106);
nand U23635 (N_23635,N_23008,N_23419);
and U23636 (N_23636,N_23051,N_23132);
or U23637 (N_23637,N_23192,N_23407);
xor U23638 (N_23638,N_23408,N_23174);
and U23639 (N_23639,N_23358,N_23483);
nor U23640 (N_23640,N_23479,N_23250);
nor U23641 (N_23641,N_23019,N_23427);
xor U23642 (N_23642,N_23155,N_23099);
or U23643 (N_23643,N_23310,N_23083);
xnor U23644 (N_23644,N_23034,N_23085);
xnor U23645 (N_23645,N_23070,N_23332);
nand U23646 (N_23646,N_23005,N_23440);
nor U23647 (N_23647,N_23150,N_23004);
xor U23648 (N_23648,N_23156,N_23167);
nand U23649 (N_23649,N_23136,N_23377);
xor U23650 (N_23650,N_23410,N_23267);
nand U23651 (N_23651,N_23212,N_23165);
nor U23652 (N_23652,N_23246,N_23220);
nor U23653 (N_23653,N_23404,N_23260);
nor U23654 (N_23654,N_23113,N_23369);
xor U23655 (N_23655,N_23223,N_23351);
and U23656 (N_23656,N_23432,N_23459);
nand U23657 (N_23657,N_23207,N_23374);
and U23658 (N_23658,N_23204,N_23461);
and U23659 (N_23659,N_23466,N_23252);
nor U23660 (N_23660,N_23228,N_23180);
nor U23661 (N_23661,N_23030,N_23268);
nor U23662 (N_23662,N_23081,N_23273);
nand U23663 (N_23663,N_23386,N_23262);
nand U23664 (N_23664,N_23216,N_23396);
nor U23665 (N_23665,N_23229,N_23002);
and U23666 (N_23666,N_23316,N_23058);
and U23667 (N_23667,N_23431,N_23240);
and U23668 (N_23668,N_23414,N_23361);
and U23669 (N_23669,N_23378,N_23060);
or U23670 (N_23670,N_23352,N_23065);
and U23671 (N_23671,N_23495,N_23038);
xor U23672 (N_23672,N_23205,N_23444);
xor U23673 (N_23673,N_23305,N_23035);
xnor U23674 (N_23674,N_23221,N_23193);
nand U23675 (N_23675,N_23339,N_23418);
or U23676 (N_23676,N_23324,N_23242);
or U23677 (N_23677,N_23224,N_23090);
and U23678 (N_23678,N_23474,N_23492);
and U23679 (N_23679,N_23376,N_23387);
nand U23680 (N_23680,N_23382,N_23152);
xnor U23681 (N_23681,N_23201,N_23123);
nor U23682 (N_23682,N_23198,N_23456);
nand U23683 (N_23683,N_23455,N_23181);
and U23684 (N_23684,N_23470,N_23115);
and U23685 (N_23685,N_23026,N_23313);
xor U23686 (N_23686,N_23364,N_23284);
nor U23687 (N_23687,N_23063,N_23389);
nor U23688 (N_23688,N_23449,N_23184);
nand U23689 (N_23689,N_23319,N_23372);
xnor U23690 (N_23690,N_23485,N_23020);
xor U23691 (N_23691,N_23069,N_23135);
xor U23692 (N_23692,N_23230,N_23077);
and U23693 (N_23693,N_23134,N_23107);
nand U23694 (N_23694,N_23468,N_23253);
nand U23695 (N_23695,N_23036,N_23249);
nor U23696 (N_23696,N_23342,N_23309);
xor U23697 (N_23697,N_23438,N_23484);
or U23698 (N_23698,N_23138,N_23062);
nor U23699 (N_23699,N_23258,N_23460);
or U23700 (N_23700,N_23277,N_23385);
xor U23701 (N_23701,N_23399,N_23048);
xor U23702 (N_23702,N_23046,N_23119);
and U23703 (N_23703,N_23336,N_23302);
and U23704 (N_23704,N_23088,N_23098);
nand U23705 (N_23705,N_23105,N_23151);
nand U23706 (N_23706,N_23480,N_23439);
nor U23707 (N_23707,N_23177,N_23383);
xnor U23708 (N_23708,N_23241,N_23264);
xor U23709 (N_23709,N_23283,N_23222);
nand U23710 (N_23710,N_23232,N_23323);
nor U23711 (N_23711,N_23448,N_23295);
nor U23712 (N_23712,N_23353,N_23330);
and U23713 (N_23713,N_23359,N_23071);
and U23714 (N_23714,N_23236,N_23012);
nor U23715 (N_23715,N_23318,N_23147);
xor U23716 (N_23716,N_23401,N_23122);
or U23717 (N_23717,N_23078,N_23126);
nor U23718 (N_23718,N_23092,N_23133);
xor U23719 (N_23719,N_23120,N_23486);
nand U23720 (N_23720,N_23244,N_23173);
nor U23721 (N_23721,N_23121,N_23188);
nor U23722 (N_23722,N_23218,N_23452);
nor U23723 (N_23723,N_23326,N_23292);
and U23724 (N_23724,N_23279,N_23282);
xor U23725 (N_23725,N_23238,N_23400);
and U23726 (N_23726,N_23117,N_23274);
nand U23727 (N_23727,N_23317,N_23392);
nor U23728 (N_23728,N_23162,N_23157);
and U23729 (N_23729,N_23003,N_23421);
nand U23730 (N_23730,N_23017,N_23233);
and U23731 (N_23731,N_23139,N_23251);
nor U23732 (N_23732,N_23111,N_23082);
nor U23733 (N_23733,N_23131,N_23398);
nor U23734 (N_23734,N_23415,N_23208);
xnor U23735 (N_23735,N_23130,N_23450);
nor U23736 (N_23736,N_23367,N_23416);
nor U23737 (N_23737,N_23072,N_23409);
nor U23738 (N_23738,N_23296,N_23248);
and U23739 (N_23739,N_23129,N_23315);
and U23740 (N_23740,N_23496,N_23476);
xor U23741 (N_23741,N_23033,N_23368);
or U23742 (N_23742,N_23384,N_23159);
xor U23743 (N_23743,N_23403,N_23350);
nor U23744 (N_23744,N_23334,N_23388);
and U23745 (N_23745,N_23154,N_23243);
nand U23746 (N_23746,N_23226,N_23015);
or U23747 (N_23747,N_23391,N_23397);
and U23748 (N_23748,N_23265,N_23187);
xor U23749 (N_23749,N_23146,N_23329);
and U23750 (N_23750,N_23452,N_23232);
nor U23751 (N_23751,N_23471,N_23219);
nor U23752 (N_23752,N_23237,N_23352);
and U23753 (N_23753,N_23339,N_23199);
nor U23754 (N_23754,N_23070,N_23127);
xor U23755 (N_23755,N_23139,N_23026);
and U23756 (N_23756,N_23445,N_23227);
or U23757 (N_23757,N_23244,N_23249);
or U23758 (N_23758,N_23034,N_23360);
or U23759 (N_23759,N_23121,N_23466);
xnor U23760 (N_23760,N_23191,N_23296);
and U23761 (N_23761,N_23204,N_23201);
and U23762 (N_23762,N_23441,N_23190);
xnor U23763 (N_23763,N_23441,N_23475);
nand U23764 (N_23764,N_23438,N_23401);
xor U23765 (N_23765,N_23061,N_23138);
or U23766 (N_23766,N_23470,N_23318);
and U23767 (N_23767,N_23306,N_23266);
nand U23768 (N_23768,N_23195,N_23210);
nand U23769 (N_23769,N_23211,N_23126);
or U23770 (N_23770,N_23141,N_23249);
xor U23771 (N_23771,N_23160,N_23202);
nor U23772 (N_23772,N_23282,N_23422);
xor U23773 (N_23773,N_23427,N_23183);
nand U23774 (N_23774,N_23338,N_23116);
nand U23775 (N_23775,N_23395,N_23391);
nor U23776 (N_23776,N_23035,N_23256);
nor U23777 (N_23777,N_23054,N_23019);
or U23778 (N_23778,N_23402,N_23427);
nand U23779 (N_23779,N_23388,N_23473);
or U23780 (N_23780,N_23195,N_23378);
xnor U23781 (N_23781,N_23217,N_23243);
and U23782 (N_23782,N_23390,N_23245);
nand U23783 (N_23783,N_23203,N_23044);
nand U23784 (N_23784,N_23247,N_23052);
or U23785 (N_23785,N_23353,N_23386);
nor U23786 (N_23786,N_23158,N_23003);
nor U23787 (N_23787,N_23438,N_23282);
nor U23788 (N_23788,N_23466,N_23324);
and U23789 (N_23789,N_23404,N_23096);
xor U23790 (N_23790,N_23281,N_23293);
or U23791 (N_23791,N_23215,N_23498);
nand U23792 (N_23792,N_23376,N_23341);
and U23793 (N_23793,N_23168,N_23238);
and U23794 (N_23794,N_23289,N_23118);
xnor U23795 (N_23795,N_23024,N_23478);
or U23796 (N_23796,N_23360,N_23088);
and U23797 (N_23797,N_23165,N_23432);
or U23798 (N_23798,N_23261,N_23198);
xor U23799 (N_23799,N_23467,N_23085);
and U23800 (N_23800,N_23330,N_23478);
and U23801 (N_23801,N_23257,N_23163);
or U23802 (N_23802,N_23399,N_23129);
nor U23803 (N_23803,N_23325,N_23300);
xnor U23804 (N_23804,N_23084,N_23088);
nand U23805 (N_23805,N_23312,N_23033);
nand U23806 (N_23806,N_23349,N_23445);
nor U23807 (N_23807,N_23157,N_23089);
or U23808 (N_23808,N_23247,N_23447);
or U23809 (N_23809,N_23355,N_23061);
and U23810 (N_23810,N_23461,N_23165);
or U23811 (N_23811,N_23005,N_23381);
and U23812 (N_23812,N_23128,N_23429);
nand U23813 (N_23813,N_23108,N_23204);
nand U23814 (N_23814,N_23145,N_23081);
or U23815 (N_23815,N_23032,N_23370);
nand U23816 (N_23816,N_23207,N_23174);
and U23817 (N_23817,N_23181,N_23019);
nor U23818 (N_23818,N_23082,N_23205);
and U23819 (N_23819,N_23461,N_23236);
or U23820 (N_23820,N_23083,N_23498);
and U23821 (N_23821,N_23491,N_23368);
and U23822 (N_23822,N_23053,N_23179);
and U23823 (N_23823,N_23339,N_23217);
xnor U23824 (N_23824,N_23007,N_23360);
or U23825 (N_23825,N_23237,N_23481);
and U23826 (N_23826,N_23462,N_23046);
nand U23827 (N_23827,N_23116,N_23237);
xor U23828 (N_23828,N_23320,N_23031);
xor U23829 (N_23829,N_23253,N_23085);
or U23830 (N_23830,N_23039,N_23364);
nor U23831 (N_23831,N_23234,N_23155);
nand U23832 (N_23832,N_23137,N_23006);
nor U23833 (N_23833,N_23001,N_23383);
and U23834 (N_23834,N_23004,N_23106);
or U23835 (N_23835,N_23000,N_23202);
nand U23836 (N_23836,N_23177,N_23040);
nor U23837 (N_23837,N_23206,N_23399);
nor U23838 (N_23838,N_23396,N_23097);
nor U23839 (N_23839,N_23293,N_23031);
nor U23840 (N_23840,N_23490,N_23388);
nand U23841 (N_23841,N_23096,N_23289);
or U23842 (N_23842,N_23321,N_23439);
nand U23843 (N_23843,N_23122,N_23372);
nand U23844 (N_23844,N_23229,N_23413);
and U23845 (N_23845,N_23204,N_23371);
nand U23846 (N_23846,N_23217,N_23317);
and U23847 (N_23847,N_23478,N_23357);
and U23848 (N_23848,N_23078,N_23301);
nand U23849 (N_23849,N_23412,N_23170);
nor U23850 (N_23850,N_23245,N_23087);
xor U23851 (N_23851,N_23181,N_23313);
nor U23852 (N_23852,N_23480,N_23264);
nand U23853 (N_23853,N_23267,N_23299);
or U23854 (N_23854,N_23010,N_23460);
or U23855 (N_23855,N_23237,N_23060);
and U23856 (N_23856,N_23352,N_23476);
nor U23857 (N_23857,N_23365,N_23094);
nor U23858 (N_23858,N_23357,N_23155);
or U23859 (N_23859,N_23164,N_23038);
and U23860 (N_23860,N_23280,N_23057);
nand U23861 (N_23861,N_23118,N_23301);
nand U23862 (N_23862,N_23194,N_23363);
xor U23863 (N_23863,N_23294,N_23375);
nor U23864 (N_23864,N_23143,N_23257);
or U23865 (N_23865,N_23198,N_23045);
and U23866 (N_23866,N_23288,N_23068);
nor U23867 (N_23867,N_23209,N_23297);
or U23868 (N_23868,N_23222,N_23226);
xor U23869 (N_23869,N_23199,N_23496);
xor U23870 (N_23870,N_23173,N_23416);
and U23871 (N_23871,N_23337,N_23452);
xnor U23872 (N_23872,N_23472,N_23416);
xor U23873 (N_23873,N_23369,N_23380);
nor U23874 (N_23874,N_23142,N_23496);
nor U23875 (N_23875,N_23382,N_23307);
nor U23876 (N_23876,N_23494,N_23197);
nand U23877 (N_23877,N_23220,N_23170);
nor U23878 (N_23878,N_23241,N_23155);
and U23879 (N_23879,N_23219,N_23050);
and U23880 (N_23880,N_23277,N_23436);
nor U23881 (N_23881,N_23125,N_23002);
nor U23882 (N_23882,N_23271,N_23480);
or U23883 (N_23883,N_23372,N_23158);
and U23884 (N_23884,N_23362,N_23254);
nor U23885 (N_23885,N_23332,N_23052);
nor U23886 (N_23886,N_23216,N_23211);
xnor U23887 (N_23887,N_23273,N_23413);
and U23888 (N_23888,N_23252,N_23383);
nand U23889 (N_23889,N_23478,N_23040);
nor U23890 (N_23890,N_23222,N_23200);
nand U23891 (N_23891,N_23179,N_23005);
xor U23892 (N_23892,N_23073,N_23003);
nor U23893 (N_23893,N_23480,N_23079);
nor U23894 (N_23894,N_23258,N_23362);
nor U23895 (N_23895,N_23202,N_23401);
or U23896 (N_23896,N_23221,N_23265);
nand U23897 (N_23897,N_23333,N_23029);
or U23898 (N_23898,N_23306,N_23394);
nand U23899 (N_23899,N_23278,N_23462);
and U23900 (N_23900,N_23296,N_23194);
or U23901 (N_23901,N_23262,N_23295);
nor U23902 (N_23902,N_23348,N_23051);
nor U23903 (N_23903,N_23074,N_23292);
xor U23904 (N_23904,N_23349,N_23215);
or U23905 (N_23905,N_23022,N_23402);
nand U23906 (N_23906,N_23240,N_23399);
or U23907 (N_23907,N_23076,N_23220);
and U23908 (N_23908,N_23391,N_23242);
or U23909 (N_23909,N_23294,N_23263);
nor U23910 (N_23910,N_23080,N_23320);
xor U23911 (N_23911,N_23060,N_23035);
nor U23912 (N_23912,N_23027,N_23068);
nor U23913 (N_23913,N_23345,N_23340);
nand U23914 (N_23914,N_23221,N_23164);
nand U23915 (N_23915,N_23212,N_23377);
nor U23916 (N_23916,N_23350,N_23374);
and U23917 (N_23917,N_23005,N_23233);
and U23918 (N_23918,N_23217,N_23346);
or U23919 (N_23919,N_23117,N_23200);
xnor U23920 (N_23920,N_23237,N_23204);
nor U23921 (N_23921,N_23067,N_23496);
nor U23922 (N_23922,N_23217,N_23292);
nand U23923 (N_23923,N_23311,N_23067);
and U23924 (N_23924,N_23470,N_23058);
xor U23925 (N_23925,N_23304,N_23175);
nor U23926 (N_23926,N_23110,N_23010);
or U23927 (N_23927,N_23388,N_23088);
xor U23928 (N_23928,N_23159,N_23206);
nand U23929 (N_23929,N_23146,N_23388);
or U23930 (N_23930,N_23432,N_23162);
xnor U23931 (N_23931,N_23481,N_23462);
nand U23932 (N_23932,N_23171,N_23260);
xor U23933 (N_23933,N_23181,N_23273);
nor U23934 (N_23934,N_23347,N_23064);
nor U23935 (N_23935,N_23118,N_23115);
xnor U23936 (N_23936,N_23365,N_23464);
nor U23937 (N_23937,N_23467,N_23309);
or U23938 (N_23938,N_23292,N_23027);
and U23939 (N_23939,N_23028,N_23098);
xnor U23940 (N_23940,N_23237,N_23350);
xnor U23941 (N_23941,N_23284,N_23196);
xnor U23942 (N_23942,N_23364,N_23225);
nor U23943 (N_23943,N_23331,N_23278);
nand U23944 (N_23944,N_23080,N_23449);
and U23945 (N_23945,N_23129,N_23207);
nand U23946 (N_23946,N_23427,N_23184);
and U23947 (N_23947,N_23248,N_23229);
nand U23948 (N_23948,N_23267,N_23255);
nor U23949 (N_23949,N_23462,N_23366);
nor U23950 (N_23950,N_23271,N_23150);
and U23951 (N_23951,N_23050,N_23422);
or U23952 (N_23952,N_23366,N_23394);
nand U23953 (N_23953,N_23398,N_23361);
nand U23954 (N_23954,N_23073,N_23324);
nor U23955 (N_23955,N_23049,N_23060);
nand U23956 (N_23956,N_23340,N_23411);
and U23957 (N_23957,N_23272,N_23117);
and U23958 (N_23958,N_23156,N_23399);
or U23959 (N_23959,N_23480,N_23450);
and U23960 (N_23960,N_23336,N_23490);
nand U23961 (N_23961,N_23470,N_23204);
nand U23962 (N_23962,N_23097,N_23129);
and U23963 (N_23963,N_23258,N_23317);
and U23964 (N_23964,N_23028,N_23233);
nand U23965 (N_23965,N_23016,N_23408);
and U23966 (N_23966,N_23442,N_23408);
and U23967 (N_23967,N_23323,N_23483);
xor U23968 (N_23968,N_23179,N_23065);
xnor U23969 (N_23969,N_23490,N_23278);
nor U23970 (N_23970,N_23334,N_23143);
and U23971 (N_23971,N_23388,N_23135);
nor U23972 (N_23972,N_23144,N_23081);
or U23973 (N_23973,N_23121,N_23393);
xor U23974 (N_23974,N_23336,N_23359);
nor U23975 (N_23975,N_23480,N_23483);
xnor U23976 (N_23976,N_23276,N_23080);
and U23977 (N_23977,N_23237,N_23109);
xnor U23978 (N_23978,N_23224,N_23028);
nand U23979 (N_23979,N_23134,N_23429);
nand U23980 (N_23980,N_23161,N_23195);
nand U23981 (N_23981,N_23050,N_23252);
nor U23982 (N_23982,N_23006,N_23127);
nand U23983 (N_23983,N_23241,N_23186);
nand U23984 (N_23984,N_23458,N_23390);
or U23985 (N_23985,N_23410,N_23423);
nor U23986 (N_23986,N_23112,N_23008);
or U23987 (N_23987,N_23095,N_23070);
nor U23988 (N_23988,N_23406,N_23184);
or U23989 (N_23989,N_23287,N_23183);
nor U23990 (N_23990,N_23338,N_23324);
xor U23991 (N_23991,N_23494,N_23279);
and U23992 (N_23992,N_23421,N_23315);
and U23993 (N_23993,N_23458,N_23011);
or U23994 (N_23994,N_23271,N_23233);
or U23995 (N_23995,N_23027,N_23099);
xnor U23996 (N_23996,N_23222,N_23098);
and U23997 (N_23997,N_23297,N_23103);
xor U23998 (N_23998,N_23246,N_23330);
or U23999 (N_23999,N_23328,N_23379);
xnor U24000 (N_24000,N_23863,N_23591);
nand U24001 (N_24001,N_23546,N_23949);
nor U24002 (N_24002,N_23535,N_23727);
and U24003 (N_24003,N_23929,N_23987);
and U24004 (N_24004,N_23556,N_23585);
xnor U24005 (N_24005,N_23653,N_23892);
xnor U24006 (N_24006,N_23910,N_23924);
nand U24007 (N_24007,N_23715,N_23971);
or U24008 (N_24008,N_23852,N_23554);
or U24009 (N_24009,N_23531,N_23505);
nand U24010 (N_24010,N_23921,N_23918);
nor U24011 (N_24011,N_23595,N_23826);
xnor U24012 (N_24012,N_23940,N_23795);
or U24013 (N_24013,N_23741,N_23822);
and U24014 (N_24014,N_23763,N_23661);
or U24015 (N_24015,N_23509,N_23537);
and U24016 (N_24016,N_23835,N_23866);
xor U24017 (N_24017,N_23520,N_23856);
xor U24018 (N_24018,N_23854,N_23790);
and U24019 (N_24019,N_23736,N_23885);
xnor U24020 (N_24020,N_23791,N_23550);
nand U24021 (N_24021,N_23700,N_23858);
nand U24022 (N_24022,N_23686,N_23620);
nand U24023 (N_24023,N_23525,N_23806);
xnor U24024 (N_24024,N_23658,N_23528);
nor U24025 (N_24025,N_23983,N_23702);
nor U24026 (N_24026,N_23538,N_23769);
nand U24027 (N_24027,N_23568,N_23503);
nor U24028 (N_24028,N_23845,N_23884);
nand U24029 (N_24029,N_23708,N_23926);
and U24030 (N_24030,N_23840,N_23996);
xnor U24031 (N_24031,N_23621,N_23991);
nand U24032 (N_24032,N_23523,N_23733);
or U24033 (N_24033,N_23747,N_23757);
xnor U24034 (N_24034,N_23697,N_23812);
and U24035 (N_24035,N_23931,N_23985);
or U24036 (N_24036,N_23802,N_23792);
nor U24037 (N_24037,N_23848,N_23911);
nand U24038 (N_24038,N_23909,N_23824);
xor U24039 (N_24039,N_23842,N_23850);
and U24040 (N_24040,N_23682,N_23969);
xor U24041 (N_24041,N_23579,N_23994);
nor U24042 (N_24042,N_23603,N_23742);
nand U24043 (N_24043,N_23735,N_23617);
xnor U24044 (N_24044,N_23916,N_23714);
nand U24045 (N_24045,N_23978,N_23589);
and U24046 (N_24046,N_23560,N_23897);
and U24047 (N_24047,N_23734,N_23743);
or U24048 (N_24048,N_23646,N_23820);
and U24049 (N_24049,N_23879,N_23615);
or U24050 (N_24050,N_23865,N_23526);
nor U24051 (N_24051,N_23624,N_23542);
nand U24052 (N_24052,N_23610,N_23593);
nor U24053 (N_24053,N_23811,N_23974);
nand U24054 (N_24054,N_23712,N_23573);
xor U24055 (N_24055,N_23775,N_23794);
or U24056 (N_24056,N_23645,N_23684);
nor U24057 (N_24057,N_23776,N_23789);
nand U24058 (N_24058,N_23563,N_23547);
nand U24059 (N_24059,N_23860,N_23847);
xor U24060 (N_24060,N_23687,N_23740);
nand U24061 (N_24061,N_23631,N_23659);
nor U24062 (N_24062,N_23944,N_23670);
nor U24063 (N_24063,N_23504,N_23711);
and U24064 (N_24064,N_23606,N_23957);
xnor U24065 (N_24065,N_23951,N_23968);
xor U24066 (N_24066,N_23915,N_23512);
or U24067 (N_24067,N_23704,N_23594);
xor U24068 (N_24068,N_23752,N_23799);
nand U24069 (N_24069,N_23750,N_23638);
xnor U24070 (N_24070,N_23507,N_23696);
and U24071 (N_24071,N_23914,N_23644);
or U24072 (N_24072,N_23846,N_23693);
or U24073 (N_24073,N_23590,N_23730);
nor U24074 (N_24074,N_23995,N_23954);
and U24075 (N_24075,N_23518,N_23724);
or U24076 (N_24076,N_23936,N_23583);
or U24077 (N_24077,N_23864,N_23880);
or U24078 (N_24078,N_23908,N_23816);
xnor U24079 (N_24079,N_23514,N_23829);
nand U24080 (N_24080,N_23975,N_23899);
nand U24081 (N_24081,N_23521,N_23770);
or U24082 (N_24082,N_23642,N_23828);
nand U24083 (N_24083,N_23762,N_23689);
nand U24084 (N_24084,N_23731,N_23699);
xor U24085 (N_24085,N_23887,N_23785);
or U24086 (N_24086,N_23705,N_23643);
nand U24087 (N_24087,N_23541,N_23746);
nand U24088 (N_24088,N_23511,N_23559);
nand U24089 (N_24089,N_23849,N_23683);
and U24090 (N_24090,N_23764,N_23510);
xnor U24091 (N_24091,N_23600,N_23576);
and U24092 (N_24092,N_23758,N_23989);
and U24093 (N_24093,N_23797,N_23901);
xnor U24094 (N_24094,N_23906,N_23959);
and U24095 (N_24095,N_23649,N_23793);
nand U24096 (N_24096,N_23986,N_23925);
nor U24097 (N_24097,N_23932,N_23834);
xnor U24098 (N_24098,N_23647,N_23961);
or U24099 (N_24099,N_23891,N_23713);
xor U24100 (N_24100,N_23553,N_23722);
xor U24101 (N_24101,N_23946,N_23571);
xor U24102 (N_24102,N_23876,N_23656);
nor U24103 (N_24103,N_23941,N_23823);
and U24104 (N_24104,N_23552,N_23753);
nor U24105 (N_24105,N_23695,N_23934);
or U24106 (N_24106,N_23871,N_23611);
nor U24107 (N_24107,N_23868,N_23597);
or U24108 (N_24108,N_23601,N_23830);
or U24109 (N_24109,N_23979,N_23572);
and U24110 (N_24110,N_23582,N_23536);
xnor U24111 (N_24111,N_23774,N_23955);
nor U24112 (N_24112,N_23577,N_23663);
nor U24113 (N_24113,N_23922,N_23737);
and U24114 (N_24114,N_23965,N_23632);
nor U24115 (N_24115,N_23506,N_23804);
nand U24116 (N_24116,N_23913,N_23878);
nor U24117 (N_24117,N_23558,N_23657);
xnor U24118 (N_24118,N_23655,N_23673);
and U24119 (N_24119,N_23841,N_23927);
xor U24120 (N_24120,N_23751,N_23990);
and U24121 (N_24121,N_23588,N_23718);
nor U24122 (N_24122,N_23818,N_23780);
nand U24123 (N_24123,N_23896,N_23500);
nand U24124 (N_24124,N_23609,N_23534);
nor U24125 (N_24125,N_23709,N_23960);
nand U24126 (N_24126,N_23729,N_23933);
and U24127 (N_24127,N_23947,N_23973);
nand U24128 (N_24128,N_23636,N_23679);
nand U24129 (N_24129,N_23798,N_23516);
nand U24130 (N_24130,N_23873,N_23787);
or U24131 (N_24131,N_23905,N_23626);
nor U24132 (N_24132,N_23888,N_23964);
xor U24133 (N_24133,N_23800,N_23666);
and U24134 (N_24134,N_23667,N_23981);
or U24135 (N_24135,N_23972,N_23681);
nor U24136 (N_24136,N_23977,N_23529);
and U24137 (N_24137,N_23853,N_23710);
nand U24138 (N_24138,N_23814,N_23928);
xnor U24139 (N_24139,N_23773,N_23997);
and U24140 (N_24140,N_23599,N_23781);
nand U24141 (N_24141,N_23627,N_23721);
nand U24142 (N_24142,N_23907,N_23832);
or U24143 (N_24143,N_23540,N_23825);
nand U24144 (N_24144,N_23945,N_23570);
and U24145 (N_24145,N_23651,N_23935);
nor U24146 (N_24146,N_23508,N_23650);
and U24147 (N_24147,N_23574,N_23567);
or U24148 (N_24148,N_23754,N_23779);
xnor U24149 (N_24149,N_23665,N_23950);
nand U24150 (N_24150,N_23839,N_23889);
nor U24151 (N_24151,N_23634,N_23859);
nor U24152 (N_24152,N_23584,N_23630);
xnor U24153 (N_24153,N_23904,N_23988);
nand U24154 (N_24154,N_23843,N_23675);
and U24155 (N_24155,N_23970,N_23691);
and U24156 (N_24156,N_23629,N_23917);
and U24157 (N_24157,N_23628,N_23819);
xnor U24158 (N_24158,N_23707,N_23519);
or U24159 (N_24159,N_23719,N_23575);
and U24160 (N_24160,N_23855,N_23676);
and U24161 (N_24161,N_23838,N_23527);
xnor U24162 (N_24162,N_23903,N_23677);
nor U24163 (N_24163,N_23532,N_23761);
nor U24164 (N_24164,N_23652,N_23557);
or U24165 (N_24165,N_23694,N_23966);
nand U24166 (N_24166,N_23772,N_23613);
nor U24167 (N_24167,N_23998,N_23956);
or U24168 (N_24168,N_23618,N_23706);
and U24169 (N_24169,N_23883,N_23720);
xnor U24170 (N_24170,N_23783,N_23524);
nand U24171 (N_24171,N_23616,N_23544);
and U24172 (N_24172,N_23680,N_23768);
xor U24173 (N_24173,N_23662,N_23827);
xor U24174 (N_24174,N_23895,N_23723);
or U24175 (N_24175,N_23633,N_23614);
xnor U24176 (N_24176,N_23596,N_23958);
xor U24177 (N_24177,N_23566,N_23501);
nand U24178 (N_24178,N_23703,N_23569);
or U24179 (N_24179,N_23555,N_23851);
and U24180 (N_24180,N_23767,N_23837);
nand U24181 (N_24181,N_23796,N_23598);
nand U24182 (N_24182,N_23672,N_23886);
nor U24183 (N_24183,N_23821,N_23999);
and U24184 (N_24184,N_23875,N_23759);
and U24185 (N_24185,N_23522,N_23664);
xor U24186 (N_24186,N_23639,N_23831);
or U24187 (N_24187,N_23900,N_23561);
or U24188 (N_24188,N_23619,N_23898);
and U24189 (N_24189,N_23623,N_23912);
and U24190 (N_24190,N_23605,N_23882);
or U24191 (N_24191,N_23813,N_23877);
and U24192 (N_24192,N_23738,N_23760);
or U24193 (N_24193,N_23817,N_23660);
nor U24194 (N_24194,N_23515,N_23602);
nand U24195 (N_24195,N_23942,N_23668);
or U24196 (N_24196,N_23953,N_23671);
xnor U24197 (N_24197,N_23564,N_23867);
nor U24198 (N_24198,N_23801,N_23739);
or U24199 (N_24199,N_23543,N_23716);
xor U24200 (N_24200,N_23893,N_23782);
xnor U24201 (N_24201,N_23874,N_23530);
xor U24202 (N_24202,N_23777,N_23586);
or U24203 (N_24203,N_23692,N_23744);
or U24204 (N_24204,N_23635,N_23805);
nand U24205 (N_24205,N_23967,N_23786);
xnor U24206 (N_24206,N_23533,N_23612);
xnor U24207 (N_24207,N_23920,N_23578);
nand U24208 (N_24208,N_23562,N_23622);
xnor U24209 (N_24209,N_23565,N_23766);
and U24210 (N_24210,N_23963,N_23807);
nor U24211 (N_24211,N_23833,N_23604);
xor U24212 (N_24212,N_23517,N_23784);
nor U24213 (N_24213,N_23725,N_23688);
xor U24214 (N_24214,N_23788,N_23690);
xnor U24215 (N_24215,N_23992,N_23755);
or U24216 (N_24216,N_23698,N_23771);
and U24217 (N_24217,N_23939,N_23669);
and U24218 (N_24218,N_23592,N_23587);
nor U24219 (N_24219,N_23640,N_23948);
or U24220 (N_24220,N_23872,N_23756);
nor U24221 (N_24221,N_23902,N_23728);
or U24222 (N_24222,N_23982,N_23607);
and U24223 (N_24223,N_23861,N_23732);
nand U24224 (N_24224,N_23844,N_23938);
or U24225 (N_24225,N_23648,N_23952);
and U24226 (N_24226,N_23749,N_23923);
xor U24227 (N_24227,N_23513,N_23881);
nand U24228 (N_24228,N_23862,N_23937);
nand U24229 (N_24229,N_23980,N_23976);
and U24230 (N_24230,N_23869,N_23870);
nand U24231 (N_24231,N_23836,N_23748);
xnor U24232 (N_24232,N_23502,N_23548);
or U24233 (N_24233,N_23717,N_23803);
nand U24234 (N_24234,N_23810,N_23943);
and U24235 (N_24235,N_23654,N_23625);
or U24236 (N_24236,N_23608,N_23539);
and U24237 (N_24237,N_23745,N_23778);
or U24238 (N_24238,N_23857,N_23809);
nand U24239 (N_24239,N_23894,N_23815);
or U24240 (N_24240,N_23545,N_23962);
and U24241 (N_24241,N_23678,N_23637);
nor U24242 (N_24242,N_23726,N_23919);
xnor U24243 (N_24243,N_23701,N_23890);
and U24244 (N_24244,N_23808,N_23551);
xnor U24245 (N_24245,N_23765,N_23984);
xnor U24246 (N_24246,N_23581,N_23580);
nor U24247 (N_24247,N_23930,N_23549);
and U24248 (N_24248,N_23685,N_23641);
nor U24249 (N_24249,N_23993,N_23674);
nor U24250 (N_24250,N_23883,N_23904);
xor U24251 (N_24251,N_23785,N_23987);
and U24252 (N_24252,N_23702,N_23909);
nand U24253 (N_24253,N_23779,N_23947);
or U24254 (N_24254,N_23564,N_23560);
or U24255 (N_24255,N_23773,N_23977);
xor U24256 (N_24256,N_23647,N_23681);
nand U24257 (N_24257,N_23844,N_23572);
nand U24258 (N_24258,N_23508,N_23780);
xor U24259 (N_24259,N_23619,N_23750);
or U24260 (N_24260,N_23582,N_23564);
and U24261 (N_24261,N_23915,N_23961);
xor U24262 (N_24262,N_23722,N_23654);
or U24263 (N_24263,N_23697,N_23663);
nor U24264 (N_24264,N_23906,N_23772);
nand U24265 (N_24265,N_23554,N_23763);
and U24266 (N_24266,N_23703,N_23598);
nor U24267 (N_24267,N_23877,N_23706);
nand U24268 (N_24268,N_23957,N_23750);
nor U24269 (N_24269,N_23998,N_23673);
nor U24270 (N_24270,N_23583,N_23548);
nor U24271 (N_24271,N_23845,N_23589);
or U24272 (N_24272,N_23856,N_23723);
or U24273 (N_24273,N_23790,N_23880);
nor U24274 (N_24274,N_23717,N_23933);
or U24275 (N_24275,N_23552,N_23943);
and U24276 (N_24276,N_23902,N_23607);
xnor U24277 (N_24277,N_23732,N_23584);
nor U24278 (N_24278,N_23531,N_23562);
nor U24279 (N_24279,N_23664,N_23592);
nand U24280 (N_24280,N_23844,N_23661);
xnor U24281 (N_24281,N_23720,N_23625);
and U24282 (N_24282,N_23987,N_23517);
and U24283 (N_24283,N_23876,N_23710);
xor U24284 (N_24284,N_23919,N_23568);
or U24285 (N_24285,N_23777,N_23545);
nor U24286 (N_24286,N_23526,N_23516);
nand U24287 (N_24287,N_23503,N_23565);
and U24288 (N_24288,N_23688,N_23870);
or U24289 (N_24289,N_23827,N_23573);
xnor U24290 (N_24290,N_23682,N_23986);
nor U24291 (N_24291,N_23622,N_23909);
and U24292 (N_24292,N_23594,N_23845);
nand U24293 (N_24293,N_23882,N_23681);
xor U24294 (N_24294,N_23784,N_23773);
nor U24295 (N_24295,N_23582,N_23808);
and U24296 (N_24296,N_23884,N_23849);
nor U24297 (N_24297,N_23764,N_23689);
nor U24298 (N_24298,N_23964,N_23512);
nor U24299 (N_24299,N_23589,N_23585);
and U24300 (N_24300,N_23927,N_23504);
nand U24301 (N_24301,N_23679,N_23515);
or U24302 (N_24302,N_23984,N_23952);
nor U24303 (N_24303,N_23688,N_23654);
nand U24304 (N_24304,N_23581,N_23999);
nor U24305 (N_24305,N_23823,N_23930);
nor U24306 (N_24306,N_23749,N_23621);
xnor U24307 (N_24307,N_23800,N_23843);
or U24308 (N_24308,N_23747,N_23764);
and U24309 (N_24309,N_23894,N_23965);
nand U24310 (N_24310,N_23934,N_23618);
nor U24311 (N_24311,N_23608,N_23830);
and U24312 (N_24312,N_23779,N_23764);
nor U24313 (N_24313,N_23712,N_23901);
or U24314 (N_24314,N_23902,N_23801);
nand U24315 (N_24315,N_23611,N_23953);
nand U24316 (N_24316,N_23779,N_23641);
nor U24317 (N_24317,N_23757,N_23979);
nand U24318 (N_24318,N_23708,N_23516);
nand U24319 (N_24319,N_23913,N_23529);
nor U24320 (N_24320,N_23977,N_23926);
or U24321 (N_24321,N_23885,N_23831);
or U24322 (N_24322,N_23593,N_23889);
xnor U24323 (N_24323,N_23848,N_23516);
or U24324 (N_24324,N_23609,N_23559);
and U24325 (N_24325,N_23830,N_23681);
nor U24326 (N_24326,N_23956,N_23557);
nand U24327 (N_24327,N_23545,N_23935);
and U24328 (N_24328,N_23936,N_23705);
and U24329 (N_24329,N_23684,N_23603);
nor U24330 (N_24330,N_23519,N_23597);
nand U24331 (N_24331,N_23703,N_23798);
nor U24332 (N_24332,N_23822,N_23564);
xor U24333 (N_24333,N_23531,N_23884);
nand U24334 (N_24334,N_23962,N_23864);
nand U24335 (N_24335,N_23915,N_23802);
or U24336 (N_24336,N_23960,N_23631);
xnor U24337 (N_24337,N_23854,N_23550);
and U24338 (N_24338,N_23547,N_23798);
xnor U24339 (N_24339,N_23795,N_23870);
and U24340 (N_24340,N_23938,N_23974);
and U24341 (N_24341,N_23580,N_23784);
nand U24342 (N_24342,N_23930,N_23705);
nand U24343 (N_24343,N_23594,N_23962);
nand U24344 (N_24344,N_23961,N_23772);
or U24345 (N_24345,N_23846,N_23546);
nand U24346 (N_24346,N_23852,N_23753);
and U24347 (N_24347,N_23849,N_23936);
xor U24348 (N_24348,N_23780,N_23989);
nand U24349 (N_24349,N_23966,N_23700);
xnor U24350 (N_24350,N_23746,N_23762);
or U24351 (N_24351,N_23722,N_23983);
xor U24352 (N_24352,N_23557,N_23586);
or U24353 (N_24353,N_23751,N_23582);
nand U24354 (N_24354,N_23919,N_23669);
xnor U24355 (N_24355,N_23552,N_23947);
xnor U24356 (N_24356,N_23701,N_23682);
xor U24357 (N_24357,N_23596,N_23626);
nand U24358 (N_24358,N_23987,N_23789);
nand U24359 (N_24359,N_23781,N_23836);
or U24360 (N_24360,N_23597,N_23874);
nand U24361 (N_24361,N_23760,N_23984);
or U24362 (N_24362,N_23905,N_23502);
xor U24363 (N_24363,N_23813,N_23516);
nor U24364 (N_24364,N_23861,N_23646);
nand U24365 (N_24365,N_23768,N_23548);
and U24366 (N_24366,N_23624,N_23533);
nor U24367 (N_24367,N_23772,N_23893);
nor U24368 (N_24368,N_23654,N_23956);
and U24369 (N_24369,N_23780,N_23632);
nand U24370 (N_24370,N_23760,N_23776);
nor U24371 (N_24371,N_23951,N_23740);
nor U24372 (N_24372,N_23535,N_23782);
nor U24373 (N_24373,N_23843,N_23500);
nand U24374 (N_24374,N_23877,N_23965);
nor U24375 (N_24375,N_23780,N_23720);
or U24376 (N_24376,N_23667,N_23828);
nor U24377 (N_24377,N_23651,N_23822);
nor U24378 (N_24378,N_23963,N_23986);
or U24379 (N_24379,N_23656,N_23867);
nand U24380 (N_24380,N_23544,N_23689);
nor U24381 (N_24381,N_23975,N_23611);
or U24382 (N_24382,N_23897,N_23620);
nor U24383 (N_24383,N_23547,N_23748);
xor U24384 (N_24384,N_23633,N_23862);
xor U24385 (N_24385,N_23696,N_23937);
xnor U24386 (N_24386,N_23674,N_23570);
nor U24387 (N_24387,N_23612,N_23656);
and U24388 (N_24388,N_23515,N_23760);
and U24389 (N_24389,N_23963,N_23513);
nand U24390 (N_24390,N_23508,N_23844);
or U24391 (N_24391,N_23536,N_23709);
nor U24392 (N_24392,N_23603,N_23999);
or U24393 (N_24393,N_23940,N_23627);
nor U24394 (N_24394,N_23550,N_23761);
and U24395 (N_24395,N_23509,N_23560);
nand U24396 (N_24396,N_23957,N_23655);
xnor U24397 (N_24397,N_23627,N_23531);
nand U24398 (N_24398,N_23696,N_23770);
or U24399 (N_24399,N_23944,N_23613);
nor U24400 (N_24400,N_23932,N_23938);
nor U24401 (N_24401,N_23859,N_23697);
nand U24402 (N_24402,N_23666,N_23992);
and U24403 (N_24403,N_23865,N_23519);
or U24404 (N_24404,N_23801,N_23798);
nand U24405 (N_24405,N_23670,N_23793);
nor U24406 (N_24406,N_23644,N_23831);
xor U24407 (N_24407,N_23697,N_23748);
nand U24408 (N_24408,N_23655,N_23587);
nand U24409 (N_24409,N_23838,N_23557);
nor U24410 (N_24410,N_23659,N_23747);
nand U24411 (N_24411,N_23801,N_23768);
nor U24412 (N_24412,N_23632,N_23550);
or U24413 (N_24413,N_23631,N_23544);
xnor U24414 (N_24414,N_23960,N_23722);
xor U24415 (N_24415,N_23810,N_23584);
xnor U24416 (N_24416,N_23966,N_23946);
or U24417 (N_24417,N_23552,N_23668);
xor U24418 (N_24418,N_23547,N_23814);
xor U24419 (N_24419,N_23549,N_23862);
nand U24420 (N_24420,N_23651,N_23787);
xor U24421 (N_24421,N_23988,N_23681);
nand U24422 (N_24422,N_23951,N_23651);
nor U24423 (N_24423,N_23866,N_23771);
nand U24424 (N_24424,N_23575,N_23537);
or U24425 (N_24425,N_23663,N_23979);
or U24426 (N_24426,N_23625,N_23627);
and U24427 (N_24427,N_23612,N_23666);
or U24428 (N_24428,N_23960,N_23548);
nor U24429 (N_24429,N_23585,N_23576);
and U24430 (N_24430,N_23665,N_23879);
and U24431 (N_24431,N_23880,N_23952);
nand U24432 (N_24432,N_23649,N_23509);
nand U24433 (N_24433,N_23896,N_23957);
nor U24434 (N_24434,N_23841,N_23934);
xor U24435 (N_24435,N_23834,N_23682);
and U24436 (N_24436,N_23559,N_23929);
nor U24437 (N_24437,N_23853,N_23791);
nor U24438 (N_24438,N_23969,N_23956);
or U24439 (N_24439,N_23558,N_23777);
nand U24440 (N_24440,N_23701,N_23934);
or U24441 (N_24441,N_23974,N_23659);
xnor U24442 (N_24442,N_23706,N_23775);
or U24443 (N_24443,N_23869,N_23501);
and U24444 (N_24444,N_23932,N_23551);
or U24445 (N_24445,N_23536,N_23948);
or U24446 (N_24446,N_23922,N_23774);
nand U24447 (N_24447,N_23531,N_23814);
and U24448 (N_24448,N_23735,N_23813);
or U24449 (N_24449,N_23907,N_23572);
or U24450 (N_24450,N_23805,N_23605);
xor U24451 (N_24451,N_23720,N_23908);
or U24452 (N_24452,N_23920,N_23818);
xor U24453 (N_24453,N_23547,N_23651);
and U24454 (N_24454,N_23808,N_23771);
and U24455 (N_24455,N_23525,N_23907);
xor U24456 (N_24456,N_23700,N_23816);
nor U24457 (N_24457,N_23750,N_23520);
or U24458 (N_24458,N_23811,N_23771);
xor U24459 (N_24459,N_23918,N_23639);
or U24460 (N_24460,N_23516,N_23504);
nor U24461 (N_24461,N_23802,N_23670);
nand U24462 (N_24462,N_23602,N_23557);
xor U24463 (N_24463,N_23833,N_23867);
or U24464 (N_24464,N_23708,N_23568);
nand U24465 (N_24465,N_23901,N_23992);
nor U24466 (N_24466,N_23702,N_23612);
nand U24467 (N_24467,N_23645,N_23580);
xnor U24468 (N_24468,N_23830,N_23762);
or U24469 (N_24469,N_23999,N_23639);
nand U24470 (N_24470,N_23536,N_23600);
nand U24471 (N_24471,N_23874,N_23963);
and U24472 (N_24472,N_23532,N_23978);
xnor U24473 (N_24473,N_23779,N_23984);
nand U24474 (N_24474,N_23991,N_23603);
nand U24475 (N_24475,N_23554,N_23640);
and U24476 (N_24476,N_23834,N_23914);
xor U24477 (N_24477,N_23518,N_23954);
and U24478 (N_24478,N_23770,N_23628);
nor U24479 (N_24479,N_23721,N_23797);
and U24480 (N_24480,N_23679,N_23936);
nand U24481 (N_24481,N_23789,N_23920);
nand U24482 (N_24482,N_23953,N_23898);
and U24483 (N_24483,N_23617,N_23837);
nand U24484 (N_24484,N_23806,N_23605);
nand U24485 (N_24485,N_23810,N_23521);
xnor U24486 (N_24486,N_23740,N_23636);
or U24487 (N_24487,N_23602,N_23824);
or U24488 (N_24488,N_23534,N_23854);
nor U24489 (N_24489,N_23935,N_23619);
nor U24490 (N_24490,N_23725,N_23532);
or U24491 (N_24491,N_23641,N_23536);
or U24492 (N_24492,N_23953,N_23842);
nand U24493 (N_24493,N_23760,N_23822);
nor U24494 (N_24494,N_23975,N_23628);
nand U24495 (N_24495,N_23642,N_23928);
xnor U24496 (N_24496,N_23555,N_23953);
nand U24497 (N_24497,N_23745,N_23818);
or U24498 (N_24498,N_23982,N_23540);
nor U24499 (N_24499,N_23780,N_23663);
nand U24500 (N_24500,N_24061,N_24277);
and U24501 (N_24501,N_24269,N_24083);
nand U24502 (N_24502,N_24263,N_24383);
xnor U24503 (N_24503,N_24321,N_24444);
xnor U24504 (N_24504,N_24424,N_24062);
or U24505 (N_24505,N_24100,N_24177);
or U24506 (N_24506,N_24226,N_24485);
and U24507 (N_24507,N_24435,N_24139);
nand U24508 (N_24508,N_24481,N_24000);
or U24509 (N_24509,N_24106,N_24386);
and U24510 (N_24510,N_24251,N_24264);
and U24511 (N_24511,N_24146,N_24215);
nor U24512 (N_24512,N_24153,N_24340);
and U24513 (N_24513,N_24302,N_24471);
and U24514 (N_24514,N_24312,N_24316);
or U24515 (N_24515,N_24461,N_24410);
or U24516 (N_24516,N_24474,N_24466);
nor U24517 (N_24517,N_24325,N_24469);
nor U24518 (N_24518,N_24246,N_24040);
and U24519 (N_24519,N_24067,N_24261);
nand U24520 (N_24520,N_24016,N_24237);
or U24521 (N_24521,N_24494,N_24479);
nor U24522 (N_24522,N_24433,N_24206);
nand U24523 (N_24523,N_24252,N_24274);
nor U24524 (N_24524,N_24378,N_24279);
nand U24525 (N_24525,N_24331,N_24356);
nand U24526 (N_24526,N_24462,N_24431);
or U24527 (N_24527,N_24432,N_24046);
xnor U24528 (N_24528,N_24381,N_24349);
nor U24529 (N_24529,N_24006,N_24289);
nor U24530 (N_24530,N_24370,N_24256);
nor U24531 (N_24531,N_24114,N_24449);
nor U24532 (N_24532,N_24079,N_24074);
xor U24533 (N_24533,N_24218,N_24398);
and U24534 (N_24534,N_24232,N_24049);
and U24535 (N_24535,N_24484,N_24166);
xnor U24536 (N_24536,N_24475,N_24291);
nor U24537 (N_24537,N_24089,N_24160);
and U24538 (N_24538,N_24082,N_24286);
and U24539 (N_24539,N_24224,N_24360);
or U24540 (N_24540,N_24297,N_24280);
nand U24541 (N_24541,N_24488,N_24158);
and U24542 (N_24542,N_24311,N_24119);
xor U24543 (N_24543,N_24450,N_24318);
xnor U24544 (N_24544,N_24339,N_24303);
or U24545 (N_24545,N_24394,N_24404);
or U24546 (N_24546,N_24014,N_24362);
nand U24547 (N_24547,N_24292,N_24487);
xnor U24548 (N_24548,N_24497,N_24168);
and U24549 (N_24549,N_24384,N_24017);
and U24550 (N_24550,N_24405,N_24030);
xnor U24551 (N_24551,N_24343,N_24140);
or U24552 (N_24552,N_24313,N_24464);
xnor U24553 (N_24553,N_24396,N_24392);
xnor U24554 (N_24554,N_24233,N_24094);
nand U24555 (N_24555,N_24024,N_24068);
and U24556 (N_24556,N_24162,N_24171);
or U24557 (N_24557,N_24273,N_24283);
xnor U24558 (N_24558,N_24380,N_24376);
xnor U24559 (N_24559,N_24472,N_24365);
xnor U24560 (N_24560,N_24029,N_24188);
nor U24561 (N_24561,N_24086,N_24127);
and U24562 (N_24562,N_24217,N_24178);
nor U24563 (N_24563,N_24077,N_24480);
and U24564 (N_24564,N_24451,N_24369);
xor U24565 (N_24565,N_24042,N_24421);
xor U24566 (N_24566,N_24097,N_24195);
xnor U24567 (N_24567,N_24141,N_24330);
and U24568 (N_24568,N_24336,N_24457);
xnor U24569 (N_24569,N_24212,N_24281);
nand U24570 (N_24570,N_24323,N_24348);
nor U24571 (N_24571,N_24441,N_24193);
nor U24572 (N_24572,N_24422,N_24131);
xor U24573 (N_24573,N_24058,N_24107);
xnor U24574 (N_24574,N_24148,N_24197);
nand U24575 (N_24575,N_24492,N_24064);
xnor U24576 (N_24576,N_24257,N_24309);
or U24577 (N_24577,N_24105,N_24467);
xnor U24578 (N_24578,N_24282,N_24142);
and U24579 (N_24579,N_24004,N_24041);
nor U24580 (N_24580,N_24242,N_24144);
or U24581 (N_24581,N_24183,N_24020);
and U24582 (N_24582,N_24254,N_24425);
xnor U24583 (N_24583,N_24163,N_24184);
or U24584 (N_24584,N_24181,N_24138);
nand U24585 (N_24585,N_24011,N_24034);
or U24586 (N_24586,N_24448,N_24123);
nor U24587 (N_24587,N_24081,N_24440);
or U24588 (N_24588,N_24335,N_24473);
nand U24589 (N_24589,N_24387,N_24495);
nand U24590 (N_24590,N_24373,N_24222);
nor U24591 (N_24591,N_24436,N_24416);
and U24592 (N_24592,N_24229,N_24021);
and U24593 (N_24593,N_24262,N_24445);
and U24594 (N_24594,N_24293,N_24203);
nand U24595 (N_24595,N_24391,N_24388);
and U24596 (N_24596,N_24057,N_24124);
xnor U24597 (N_24597,N_24287,N_24327);
xor U24598 (N_24598,N_24120,N_24334);
or U24599 (N_24599,N_24275,N_24428);
or U24600 (N_24600,N_24230,N_24361);
nand U24601 (N_24601,N_24109,N_24301);
or U24602 (N_24602,N_24096,N_24447);
nand U24603 (N_24603,N_24156,N_24368);
xor U24604 (N_24604,N_24374,N_24414);
or U24605 (N_24605,N_24491,N_24413);
nor U24606 (N_24606,N_24255,N_24266);
xnor U24607 (N_24607,N_24152,N_24434);
and U24608 (N_24608,N_24250,N_24202);
or U24609 (N_24609,N_24442,N_24265);
and U24610 (N_24610,N_24132,N_24400);
nand U24611 (N_24611,N_24031,N_24213);
nor U24612 (N_24612,N_24051,N_24055);
or U24613 (N_24613,N_24128,N_24458);
nand U24614 (N_24614,N_24243,N_24438);
or U24615 (N_24615,N_24452,N_24320);
xnor U24616 (N_24616,N_24110,N_24375);
or U24617 (N_24617,N_24003,N_24054);
nor U24618 (N_24618,N_24276,N_24117);
nor U24619 (N_24619,N_24008,N_24239);
xor U24620 (N_24620,N_24308,N_24231);
nand U24621 (N_24621,N_24399,N_24052);
and U24622 (N_24622,N_24066,N_24085);
nor U24623 (N_24623,N_24092,N_24121);
or U24624 (N_24624,N_24102,N_24043);
and U24625 (N_24625,N_24322,N_24379);
and U24626 (N_24626,N_24403,N_24084);
nor U24627 (N_24627,N_24352,N_24151);
nor U24628 (N_24628,N_24048,N_24078);
xnor U24629 (N_24629,N_24337,N_24395);
nand U24630 (N_24630,N_24182,N_24039);
nand U24631 (N_24631,N_24167,N_24354);
nand U24632 (N_24632,N_24198,N_24045);
nor U24633 (N_24633,N_24406,N_24227);
nor U24634 (N_24634,N_24377,N_24498);
nand U24635 (N_24635,N_24366,N_24463);
or U24636 (N_24636,N_24133,N_24259);
and U24637 (N_24637,N_24022,N_24268);
nand U24638 (N_24638,N_24290,N_24341);
or U24639 (N_24639,N_24023,N_24499);
and U24640 (N_24640,N_24284,N_24482);
nor U24641 (N_24641,N_24036,N_24207);
and U24642 (N_24642,N_24346,N_24001);
nor U24643 (N_24643,N_24372,N_24430);
nand U24644 (N_24644,N_24345,N_24018);
nor U24645 (N_24645,N_24098,N_24111);
nor U24646 (N_24646,N_24407,N_24314);
and U24647 (N_24647,N_24032,N_24216);
nor U24648 (N_24648,N_24260,N_24172);
nor U24649 (N_24649,N_24477,N_24355);
xor U24650 (N_24650,N_24186,N_24214);
or U24651 (N_24651,N_24192,N_24417);
nand U24652 (N_24652,N_24317,N_24053);
or U24653 (N_24653,N_24103,N_24219);
xor U24654 (N_24654,N_24056,N_24208);
nand U24655 (N_24655,N_24429,N_24267);
or U24656 (N_24656,N_24190,N_24069);
xnor U24657 (N_24657,N_24357,N_24490);
and U24658 (N_24658,N_24415,N_24143);
nor U24659 (N_24659,N_24409,N_24200);
xor U24660 (N_24660,N_24154,N_24095);
xor U24661 (N_24661,N_24459,N_24118);
xor U24662 (N_24662,N_24187,N_24328);
and U24663 (N_24663,N_24306,N_24411);
or U24664 (N_24664,N_24446,N_24122);
or U24665 (N_24665,N_24221,N_24271);
nor U24666 (N_24666,N_24070,N_24175);
or U24667 (N_24667,N_24326,N_24179);
or U24668 (N_24668,N_24165,N_24324);
or U24669 (N_24669,N_24389,N_24059);
xnor U24670 (N_24670,N_24244,N_24135);
and U24671 (N_24671,N_24087,N_24363);
or U24672 (N_24672,N_24390,N_24228);
nand U24673 (N_24673,N_24236,N_24385);
or U24674 (N_24674,N_24199,N_24397);
or U24675 (N_24675,N_24382,N_24329);
xor U24676 (N_24676,N_24272,N_24465);
or U24677 (N_24677,N_24205,N_24235);
or U24678 (N_24678,N_24364,N_24358);
or U24679 (N_24679,N_24402,N_24115);
nand U24680 (N_24680,N_24468,N_24027);
nor U24681 (N_24681,N_24307,N_24393);
nand U24682 (N_24682,N_24113,N_24025);
and U24683 (N_24683,N_24159,N_24130);
nand U24684 (N_24684,N_24496,N_24420);
and U24685 (N_24685,N_24426,N_24170);
xor U24686 (N_24686,N_24136,N_24012);
xnor U24687 (N_24687,N_24174,N_24101);
nand U24688 (N_24688,N_24253,N_24093);
nand U24689 (N_24689,N_24155,N_24478);
nor U24690 (N_24690,N_24249,N_24408);
or U24691 (N_24691,N_24035,N_24300);
or U24692 (N_24692,N_24238,N_24104);
xnor U24693 (N_24693,N_24285,N_24112);
xnor U24694 (N_24694,N_24033,N_24088);
xor U24695 (N_24695,N_24240,N_24419);
nor U24696 (N_24696,N_24412,N_24245);
nand U24697 (N_24697,N_24191,N_24248);
or U24698 (N_24698,N_24220,N_24125);
nor U24699 (N_24699,N_24173,N_24028);
nand U24700 (N_24700,N_24296,N_24013);
nor U24701 (N_24701,N_24169,N_24427);
xnor U24702 (N_24702,N_24367,N_24189);
or U24703 (N_24703,N_24060,N_24304);
or U24704 (N_24704,N_24489,N_24476);
nor U24705 (N_24705,N_24423,N_24439);
xnor U24706 (N_24706,N_24299,N_24147);
nand U24707 (N_24707,N_24196,N_24209);
or U24708 (N_24708,N_24176,N_24332);
nor U24709 (N_24709,N_24371,N_24164);
or U24710 (N_24710,N_24129,N_24108);
nand U24711 (N_24711,N_24470,N_24149);
or U24712 (N_24712,N_24443,N_24005);
nand U24713 (N_24713,N_24270,N_24063);
xor U24714 (N_24714,N_24211,N_24072);
or U24715 (N_24715,N_24038,N_24298);
xnor U24716 (N_24716,N_24047,N_24455);
or U24717 (N_24717,N_24453,N_24315);
xor U24718 (N_24718,N_24009,N_24456);
nor U24719 (N_24719,N_24241,N_24294);
xor U24720 (N_24720,N_24247,N_24099);
xor U24721 (N_24721,N_24210,N_24026);
and U24722 (N_24722,N_24145,N_24007);
nor U24723 (N_24723,N_24493,N_24185);
or U24724 (N_24724,N_24418,N_24201);
nand U24725 (N_24725,N_24037,N_24310);
nand U24726 (N_24726,N_24234,N_24180);
and U24727 (N_24727,N_24454,N_24161);
nand U24728 (N_24728,N_24075,N_24080);
and U24729 (N_24729,N_24090,N_24204);
nor U24730 (N_24730,N_24116,N_24134);
nand U24731 (N_24731,N_24333,N_24137);
xnor U24732 (N_24732,N_24225,N_24338);
nor U24733 (N_24733,N_24359,N_24050);
nor U24734 (N_24734,N_24350,N_24091);
and U24735 (N_24735,N_24319,N_24076);
and U24736 (N_24736,N_24305,N_24486);
nor U24737 (N_24737,N_24065,N_24295);
or U24738 (N_24738,N_24019,N_24460);
nor U24739 (N_24739,N_24010,N_24288);
nor U24740 (N_24740,N_24437,N_24223);
xnor U24741 (N_24741,N_24258,N_24347);
and U24742 (N_24742,N_24073,N_24157);
and U24743 (N_24743,N_24126,N_24278);
nor U24744 (N_24744,N_24015,N_24401);
and U24745 (N_24745,N_24353,N_24044);
and U24746 (N_24746,N_24002,N_24351);
and U24747 (N_24747,N_24483,N_24342);
nor U24748 (N_24748,N_24150,N_24071);
or U24749 (N_24749,N_24194,N_24344);
nor U24750 (N_24750,N_24245,N_24334);
or U24751 (N_24751,N_24127,N_24121);
or U24752 (N_24752,N_24427,N_24117);
and U24753 (N_24753,N_24318,N_24256);
or U24754 (N_24754,N_24104,N_24243);
and U24755 (N_24755,N_24353,N_24222);
and U24756 (N_24756,N_24230,N_24383);
xnor U24757 (N_24757,N_24248,N_24103);
nor U24758 (N_24758,N_24122,N_24167);
nor U24759 (N_24759,N_24114,N_24208);
nand U24760 (N_24760,N_24093,N_24110);
nor U24761 (N_24761,N_24092,N_24153);
or U24762 (N_24762,N_24059,N_24077);
and U24763 (N_24763,N_24102,N_24136);
nand U24764 (N_24764,N_24164,N_24455);
or U24765 (N_24765,N_24125,N_24442);
nor U24766 (N_24766,N_24044,N_24370);
nand U24767 (N_24767,N_24249,N_24236);
and U24768 (N_24768,N_24334,N_24084);
and U24769 (N_24769,N_24242,N_24046);
and U24770 (N_24770,N_24239,N_24406);
or U24771 (N_24771,N_24355,N_24465);
and U24772 (N_24772,N_24073,N_24394);
nand U24773 (N_24773,N_24216,N_24223);
nand U24774 (N_24774,N_24195,N_24475);
nor U24775 (N_24775,N_24282,N_24188);
nand U24776 (N_24776,N_24415,N_24170);
xor U24777 (N_24777,N_24120,N_24445);
nor U24778 (N_24778,N_24297,N_24483);
nand U24779 (N_24779,N_24323,N_24334);
nor U24780 (N_24780,N_24141,N_24438);
nand U24781 (N_24781,N_24476,N_24218);
xor U24782 (N_24782,N_24111,N_24277);
xor U24783 (N_24783,N_24481,N_24213);
nand U24784 (N_24784,N_24407,N_24091);
nor U24785 (N_24785,N_24430,N_24075);
xnor U24786 (N_24786,N_24203,N_24488);
nand U24787 (N_24787,N_24461,N_24298);
or U24788 (N_24788,N_24092,N_24125);
and U24789 (N_24789,N_24181,N_24360);
xnor U24790 (N_24790,N_24403,N_24195);
nor U24791 (N_24791,N_24004,N_24470);
xor U24792 (N_24792,N_24423,N_24333);
or U24793 (N_24793,N_24185,N_24134);
nand U24794 (N_24794,N_24028,N_24427);
xor U24795 (N_24795,N_24418,N_24371);
or U24796 (N_24796,N_24298,N_24287);
nand U24797 (N_24797,N_24073,N_24453);
or U24798 (N_24798,N_24276,N_24224);
and U24799 (N_24799,N_24276,N_24048);
xor U24800 (N_24800,N_24297,N_24047);
nor U24801 (N_24801,N_24235,N_24064);
and U24802 (N_24802,N_24147,N_24195);
xnor U24803 (N_24803,N_24407,N_24271);
nor U24804 (N_24804,N_24161,N_24397);
nor U24805 (N_24805,N_24313,N_24234);
and U24806 (N_24806,N_24072,N_24022);
or U24807 (N_24807,N_24385,N_24498);
or U24808 (N_24808,N_24470,N_24394);
nand U24809 (N_24809,N_24387,N_24317);
or U24810 (N_24810,N_24083,N_24410);
nand U24811 (N_24811,N_24290,N_24374);
nor U24812 (N_24812,N_24189,N_24018);
xnor U24813 (N_24813,N_24141,N_24255);
nor U24814 (N_24814,N_24181,N_24314);
or U24815 (N_24815,N_24223,N_24117);
and U24816 (N_24816,N_24310,N_24274);
or U24817 (N_24817,N_24135,N_24316);
or U24818 (N_24818,N_24413,N_24425);
xor U24819 (N_24819,N_24421,N_24221);
nor U24820 (N_24820,N_24322,N_24198);
nor U24821 (N_24821,N_24021,N_24216);
or U24822 (N_24822,N_24033,N_24490);
and U24823 (N_24823,N_24029,N_24014);
nor U24824 (N_24824,N_24398,N_24227);
xor U24825 (N_24825,N_24330,N_24227);
and U24826 (N_24826,N_24432,N_24356);
nor U24827 (N_24827,N_24317,N_24460);
nand U24828 (N_24828,N_24282,N_24440);
nand U24829 (N_24829,N_24321,N_24391);
and U24830 (N_24830,N_24386,N_24440);
and U24831 (N_24831,N_24294,N_24475);
nand U24832 (N_24832,N_24339,N_24356);
and U24833 (N_24833,N_24449,N_24020);
nand U24834 (N_24834,N_24304,N_24241);
nor U24835 (N_24835,N_24059,N_24299);
xor U24836 (N_24836,N_24411,N_24378);
nor U24837 (N_24837,N_24249,N_24272);
or U24838 (N_24838,N_24223,N_24014);
nor U24839 (N_24839,N_24139,N_24312);
or U24840 (N_24840,N_24231,N_24155);
and U24841 (N_24841,N_24330,N_24354);
nor U24842 (N_24842,N_24130,N_24298);
or U24843 (N_24843,N_24051,N_24384);
and U24844 (N_24844,N_24491,N_24245);
xor U24845 (N_24845,N_24242,N_24141);
xnor U24846 (N_24846,N_24476,N_24214);
nor U24847 (N_24847,N_24324,N_24457);
and U24848 (N_24848,N_24244,N_24004);
and U24849 (N_24849,N_24276,N_24329);
and U24850 (N_24850,N_24094,N_24131);
nand U24851 (N_24851,N_24408,N_24063);
xnor U24852 (N_24852,N_24458,N_24145);
or U24853 (N_24853,N_24192,N_24435);
and U24854 (N_24854,N_24119,N_24163);
xnor U24855 (N_24855,N_24222,N_24098);
or U24856 (N_24856,N_24101,N_24095);
xor U24857 (N_24857,N_24428,N_24127);
or U24858 (N_24858,N_24321,N_24387);
nor U24859 (N_24859,N_24183,N_24346);
and U24860 (N_24860,N_24194,N_24492);
and U24861 (N_24861,N_24167,N_24423);
nor U24862 (N_24862,N_24232,N_24473);
nand U24863 (N_24863,N_24336,N_24470);
nand U24864 (N_24864,N_24001,N_24297);
or U24865 (N_24865,N_24262,N_24194);
and U24866 (N_24866,N_24461,N_24127);
and U24867 (N_24867,N_24435,N_24197);
nor U24868 (N_24868,N_24259,N_24093);
or U24869 (N_24869,N_24409,N_24395);
nand U24870 (N_24870,N_24252,N_24424);
nor U24871 (N_24871,N_24153,N_24254);
xnor U24872 (N_24872,N_24374,N_24150);
or U24873 (N_24873,N_24117,N_24001);
nor U24874 (N_24874,N_24103,N_24067);
nor U24875 (N_24875,N_24485,N_24106);
xnor U24876 (N_24876,N_24334,N_24121);
nor U24877 (N_24877,N_24028,N_24389);
and U24878 (N_24878,N_24098,N_24189);
nor U24879 (N_24879,N_24196,N_24483);
xor U24880 (N_24880,N_24096,N_24076);
nand U24881 (N_24881,N_24222,N_24397);
nor U24882 (N_24882,N_24142,N_24415);
nor U24883 (N_24883,N_24118,N_24372);
nor U24884 (N_24884,N_24392,N_24446);
nor U24885 (N_24885,N_24382,N_24121);
or U24886 (N_24886,N_24083,N_24009);
and U24887 (N_24887,N_24249,N_24092);
and U24888 (N_24888,N_24016,N_24408);
nand U24889 (N_24889,N_24442,N_24278);
xor U24890 (N_24890,N_24438,N_24403);
and U24891 (N_24891,N_24339,N_24322);
xor U24892 (N_24892,N_24270,N_24227);
or U24893 (N_24893,N_24319,N_24453);
xor U24894 (N_24894,N_24178,N_24448);
nand U24895 (N_24895,N_24262,N_24238);
nand U24896 (N_24896,N_24231,N_24457);
and U24897 (N_24897,N_24480,N_24358);
nor U24898 (N_24898,N_24039,N_24196);
xnor U24899 (N_24899,N_24386,N_24338);
and U24900 (N_24900,N_24281,N_24381);
xnor U24901 (N_24901,N_24347,N_24483);
nor U24902 (N_24902,N_24360,N_24272);
xnor U24903 (N_24903,N_24117,N_24101);
nor U24904 (N_24904,N_24247,N_24123);
xnor U24905 (N_24905,N_24090,N_24410);
nand U24906 (N_24906,N_24034,N_24167);
xor U24907 (N_24907,N_24111,N_24411);
and U24908 (N_24908,N_24282,N_24411);
and U24909 (N_24909,N_24134,N_24462);
or U24910 (N_24910,N_24276,N_24479);
xnor U24911 (N_24911,N_24038,N_24485);
nor U24912 (N_24912,N_24304,N_24192);
or U24913 (N_24913,N_24293,N_24431);
nand U24914 (N_24914,N_24043,N_24126);
nor U24915 (N_24915,N_24379,N_24462);
nor U24916 (N_24916,N_24414,N_24283);
nand U24917 (N_24917,N_24183,N_24094);
nand U24918 (N_24918,N_24259,N_24136);
xnor U24919 (N_24919,N_24117,N_24030);
or U24920 (N_24920,N_24405,N_24323);
nand U24921 (N_24921,N_24485,N_24138);
or U24922 (N_24922,N_24253,N_24078);
xor U24923 (N_24923,N_24320,N_24103);
xnor U24924 (N_24924,N_24356,N_24463);
xor U24925 (N_24925,N_24181,N_24482);
and U24926 (N_24926,N_24203,N_24474);
and U24927 (N_24927,N_24142,N_24396);
nor U24928 (N_24928,N_24270,N_24401);
and U24929 (N_24929,N_24037,N_24129);
and U24930 (N_24930,N_24056,N_24499);
xor U24931 (N_24931,N_24249,N_24489);
or U24932 (N_24932,N_24307,N_24240);
nor U24933 (N_24933,N_24326,N_24294);
nand U24934 (N_24934,N_24093,N_24414);
or U24935 (N_24935,N_24314,N_24043);
nand U24936 (N_24936,N_24042,N_24206);
xor U24937 (N_24937,N_24308,N_24044);
nor U24938 (N_24938,N_24240,N_24286);
xor U24939 (N_24939,N_24326,N_24255);
or U24940 (N_24940,N_24382,N_24210);
nand U24941 (N_24941,N_24228,N_24090);
nor U24942 (N_24942,N_24285,N_24281);
or U24943 (N_24943,N_24163,N_24180);
and U24944 (N_24944,N_24361,N_24089);
xnor U24945 (N_24945,N_24194,N_24010);
nand U24946 (N_24946,N_24158,N_24028);
or U24947 (N_24947,N_24301,N_24034);
nand U24948 (N_24948,N_24237,N_24331);
xnor U24949 (N_24949,N_24192,N_24266);
xnor U24950 (N_24950,N_24002,N_24142);
nand U24951 (N_24951,N_24201,N_24127);
nand U24952 (N_24952,N_24073,N_24046);
and U24953 (N_24953,N_24213,N_24103);
and U24954 (N_24954,N_24060,N_24083);
xor U24955 (N_24955,N_24452,N_24209);
nor U24956 (N_24956,N_24403,N_24042);
xnor U24957 (N_24957,N_24228,N_24191);
nand U24958 (N_24958,N_24038,N_24483);
nor U24959 (N_24959,N_24463,N_24178);
nor U24960 (N_24960,N_24458,N_24432);
xnor U24961 (N_24961,N_24307,N_24292);
nor U24962 (N_24962,N_24212,N_24438);
nand U24963 (N_24963,N_24478,N_24267);
nand U24964 (N_24964,N_24008,N_24009);
xor U24965 (N_24965,N_24443,N_24074);
nor U24966 (N_24966,N_24478,N_24376);
nand U24967 (N_24967,N_24252,N_24245);
nor U24968 (N_24968,N_24183,N_24164);
and U24969 (N_24969,N_24181,N_24347);
or U24970 (N_24970,N_24223,N_24086);
nor U24971 (N_24971,N_24075,N_24336);
nand U24972 (N_24972,N_24483,N_24399);
nand U24973 (N_24973,N_24220,N_24100);
nor U24974 (N_24974,N_24075,N_24495);
xnor U24975 (N_24975,N_24400,N_24200);
and U24976 (N_24976,N_24157,N_24144);
xnor U24977 (N_24977,N_24170,N_24186);
xnor U24978 (N_24978,N_24138,N_24047);
and U24979 (N_24979,N_24131,N_24040);
xnor U24980 (N_24980,N_24398,N_24147);
nand U24981 (N_24981,N_24096,N_24115);
or U24982 (N_24982,N_24127,N_24256);
and U24983 (N_24983,N_24199,N_24378);
nor U24984 (N_24984,N_24187,N_24045);
nor U24985 (N_24985,N_24179,N_24057);
nor U24986 (N_24986,N_24021,N_24494);
and U24987 (N_24987,N_24433,N_24299);
and U24988 (N_24988,N_24383,N_24155);
and U24989 (N_24989,N_24412,N_24210);
and U24990 (N_24990,N_24270,N_24135);
or U24991 (N_24991,N_24490,N_24086);
nor U24992 (N_24992,N_24470,N_24362);
and U24993 (N_24993,N_24054,N_24094);
or U24994 (N_24994,N_24298,N_24472);
nor U24995 (N_24995,N_24455,N_24495);
and U24996 (N_24996,N_24312,N_24052);
nor U24997 (N_24997,N_24234,N_24297);
or U24998 (N_24998,N_24103,N_24004);
or U24999 (N_24999,N_24300,N_24091);
or UO_0 (O_0,N_24673,N_24772);
or UO_1 (O_1,N_24680,N_24573);
xor UO_2 (O_2,N_24524,N_24933);
or UO_3 (O_3,N_24890,N_24813);
and UO_4 (O_4,N_24523,N_24920);
or UO_5 (O_5,N_24674,N_24941);
nor UO_6 (O_6,N_24939,N_24762);
xnor UO_7 (O_7,N_24575,N_24820);
xnor UO_8 (O_8,N_24553,N_24634);
and UO_9 (O_9,N_24924,N_24932);
nand UO_10 (O_10,N_24990,N_24823);
or UO_11 (O_11,N_24861,N_24842);
nor UO_12 (O_12,N_24669,N_24899);
xor UO_13 (O_13,N_24878,N_24819);
nand UO_14 (O_14,N_24963,N_24697);
nor UO_15 (O_15,N_24522,N_24914);
nor UO_16 (O_16,N_24504,N_24738);
nand UO_17 (O_17,N_24798,N_24649);
nand UO_18 (O_18,N_24507,N_24721);
and UO_19 (O_19,N_24921,N_24646);
or UO_20 (O_20,N_24824,N_24994);
and UO_21 (O_21,N_24836,N_24537);
and UO_22 (O_22,N_24527,N_24544);
nor UO_23 (O_23,N_24767,N_24759);
and UO_24 (O_24,N_24949,N_24539);
or UO_25 (O_25,N_24644,N_24833);
or UO_26 (O_26,N_24911,N_24708);
or UO_27 (O_27,N_24663,N_24962);
and UO_28 (O_28,N_24538,N_24734);
and UO_29 (O_29,N_24615,N_24934);
and UO_30 (O_30,N_24901,N_24714);
and UO_31 (O_31,N_24750,N_24791);
or UO_32 (O_32,N_24966,N_24935);
and UO_33 (O_33,N_24642,N_24672);
xor UO_34 (O_34,N_24923,N_24886);
nor UO_35 (O_35,N_24943,N_24979);
nor UO_36 (O_36,N_24690,N_24591);
xnor UO_37 (O_37,N_24752,N_24853);
nand UO_38 (O_38,N_24597,N_24509);
xor UO_39 (O_39,N_24554,N_24908);
and UO_40 (O_40,N_24992,N_24518);
xnor UO_41 (O_41,N_24582,N_24927);
nor UO_42 (O_42,N_24800,N_24787);
or UO_43 (O_43,N_24816,N_24916);
and UO_44 (O_44,N_24756,N_24684);
xor UO_45 (O_45,N_24747,N_24955);
xor UO_46 (O_46,N_24892,N_24797);
xnor UO_47 (O_47,N_24803,N_24789);
xor UO_48 (O_48,N_24661,N_24694);
xor UO_49 (O_49,N_24725,N_24884);
and UO_50 (O_50,N_24530,N_24698);
nor UO_51 (O_51,N_24712,N_24980);
xnor UO_52 (O_52,N_24792,N_24560);
or UO_53 (O_53,N_24691,N_24814);
or UO_54 (O_54,N_24766,N_24810);
and UO_55 (O_55,N_24862,N_24993);
xnor UO_56 (O_56,N_24894,N_24961);
or UO_57 (O_57,N_24952,N_24975);
nand UO_58 (O_58,N_24811,N_24818);
xnor UO_59 (O_59,N_24701,N_24964);
or UO_60 (O_60,N_24865,N_24840);
nand UO_61 (O_61,N_24540,N_24568);
nand UO_62 (O_62,N_24586,N_24867);
nand UO_63 (O_63,N_24802,N_24874);
xor UO_64 (O_64,N_24793,N_24545);
nand UO_65 (O_65,N_24854,N_24928);
nand UO_66 (O_66,N_24631,N_24531);
nor UO_67 (O_67,N_24667,N_24877);
xor UO_68 (O_68,N_24559,N_24757);
or UO_69 (O_69,N_24898,N_24706);
or UO_70 (O_70,N_24957,N_24751);
or UO_71 (O_71,N_24781,N_24724);
nor UO_72 (O_72,N_24536,N_24740);
nand UO_73 (O_73,N_24623,N_24737);
nand UO_74 (O_74,N_24906,N_24900);
nor UO_75 (O_75,N_24543,N_24780);
nand UO_76 (O_76,N_24645,N_24577);
nor UO_77 (O_77,N_24557,N_24600);
nand UO_78 (O_78,N_24825,N_24610);
nor UO_79 (O_79,N_24655,N_24918);
nor UO_80 (O_80,N_24958,N_24891);
and UO_81 (O_81,N_24729,N_24775);
xnor UO_82 (O_82,N_24930,N_24718);
and UO_83 (O_83,N_24686,N_24777);
nand UO_84 (O_84,N_24913,N_24670);
nor UO_85 (O_85,N_24850,N_24859);
xor UO_86 (O_86,N_24965,N_24685);
nor UO_87 (O_87,N_24972,N_24513);
or UO_88 (O_88,N_24728,N_24774);
xnor UO_89 (O_89,N_24950,N_24960);
and UO_90 (O_90,N_24720,N_24662);
or UO_91 (O_91,N_24815,N_24681);
nand UO_92 (O_92,N_24755,N_24984);
xnor UO_93 (O_93,N_24657,N_24956);
nand UO_94 (O_94,N_24974,N_24709);
and UO_95 (O_95,N_24599,N_24566);
xnor UO_96 (O_96,N_24576,N_24648);
xnor UO_97 (O_97,N_24748,N_24977);
or UO_98 (O_98,N_24754,N_24804);
nand UO_99 (O_99,N_24883,N_24969);
nor UO_100 (O_100,N_24640,N_24936);
or UO_101 (O_101,N_24940,N_24598);
and UO_102 (O_102,N_24567,N_24562);
or UO_103 (O_103,N_24506,N_24564);
nor UO_104 (O_104,N_24746,N_24660);
nand UO_105 (O_105,N_24594,N_24851);
or UO_106 (O_106,N_24502,N_24919);
nor UO_107 (O_107,N_24753,N_24547);
nand UO_108 (O_108,N_24786,N_24593);
or UO_109 (O_109,N_24666,N_24585);
and UO_110 (O_110,N_24639,N_24702);
xnor UO_111 (O_111,N_24745,N_24589);
nand UO_112 (O_112,N_24839,N_24832);
nand UO_113 (O_113,N_24583,N_24882);
nand UO_114 (O_114,N_24696,N_24596);
nand UO_115 (O_115,N_24528,N_24864);
or UO_116 (O_116,N_24959,N_24711);
xor UO_117 (O_117,N_24852,N_24855);
nand UO_118 (O_118,N_24574,N_24616);
and UO_119 (O_119,N_24693,N_24622);
xor UO_120 (O_120,N_24595,N_24733);
and UO_121 (O_121,N_24907,N_24809);
and UO_122 (O_122,N_24510,N_24749);
xnor UO_123 (O_123,N_24739,N_24659);
and UO_124 (O_124,N_24532,N_24905);
nand UO_125 (O_125,N_24703,N_24873);
nor UO_126 (O_126,N_24870,N_24763);
nor UO_127 (O_127,N_24863,N_24876);
nor UO_128 (O_128,N_24525,N_24550);
nor UO_129 (O_129,N_24570,N_24727);
xor UO_130 (O_130,N_24500,N_24846);
nor UO_131 (O_131,N_24571,N_24501);
nor UO_132 (O_132,N_24604,N_24779);
nand UO_133 (O_133,N_24587,N_24700);
nand UO_134 (O_134,N_24904,N_24627);
nand UO_135 (O_135,N_24967,N_24869);
nor UO_136 (O_136,N_24770,N_24997);
and UO_137 (O_137,N_24618,N_24954);
nor UO_138 (O_138,N_24687,N_24893);
nand UO_139 (O_139,N_24879,N_24794);
and UO_140 (O_140,N_24871,N_24989);
xnor UO_141 (O_141,N_24704,N_24834);
and UO_142 (O_142,N_24603,N_24505);
nor UO_143 (O_143,N_24665,N_24785);
and UO_144 (O_144,N_24735,N_24563);
nand UO_145 (O_145,N_24581,N_24926);
or UO_146 (O_146,N_24608,N_24971);
or UO_147 (O_147,N_24512,N_24897);
or UO_148 (O_148,N_24719,N_24641);
nor UO_149 (O_149,N_24533,N_24849);
or UO_150 (O_150,N_24601,N_24716);
and UO_151 (O_151,N_24866,N_24812);
or UO_152 (O_152,N_24881,N_24722);
xnor UO_153 (O_153,N_24679,N_24529);
xor UO_154 (O_154,N_24590,N_24534);
xnor UO_155 (O_155,N_24678,N_24847);
or UO_156 (O_156,N_24912,N_24808);
xor UO_157 (O_157,N_24982,N_24713);
and UO_158 (O_158,N_24860,N_24784);
nand UO_159 (O_159,N_24676,N_24925);
xor UO_160 (O_160,N_24683,N_24555);
nor UO_161 (O_161,N_24710,N_24773);
nor UO_162 (O_162,N_24742,N_24895);
xnor UO_163 (O_163,N_24858,N_24541);
or UO_164 (O_164,N_24625,N_24788);
nor UO_165 (O_165,N_24743,N_24584);
nand UO_166 (O_166,N_24986,N_24896);
nor UO_167 (O_167,N_24831,N_24732);
nand UO_168 (O_168,N_24931,N_24771);
nand UO_169 (O_169,N_24668,N_24613);
nor UO_170 (O_170,N_24572,N_24658);
or UO_171 (O_171,N_24736,N_24845);
xor UO_172 (O_172,N_24768,N_24611);
xnor UO_173 (O_173,N_24580,N_24947);
and UO_174 (O_174,N_24826,N_24519);
and UO_175 (O_175,N_24985,N_24602);
and UO_176 (O_176,N_24948,N_24558);
nand UO_177 (O_177,N_24548,N_24880);
or UO_178 (O_178,N_24546,N_24841);
or UO_179 (O_179,N_24782,N_24689);
nor UO_180 (O_180,N_24579,N_24652);
or UO_181 (O_181,N_24744,N_24795);
nand UO_182 (O_182,N_24664,N_24692);
nand UO_183 (O_183,N_24910,N_24717);
or UO_184 (O_184,N_24817,N_24838);
xor UO_185 (O_185,N_24723,N_24621);
nand UO_186 (O_186,N_24628,N_24612);
xor UO_187 (O_187,N_24677,N_24760);
or UO_188 (O_188,N_24856,N_24758);
nand UO_189 (O_189,N_24614,N_24636);
nand UO_190 (O_190,N_24903,N_24868);
xnor UO_191 (O_191,N_24629,N_24801);
or UO_192 (O_192,N_24695,N_24857);
nand UO_193 (O_193,N_24549,N_24592);
xnor UO_194 (O_194,N_24624,N_24671);
and UO_195 (O_195,N_24726,N_24938);
nand UO_196 (O_196,N_24578,N_24635);
or UO_197 (O_197,N_24520,N_24828);
nor UO_198 (O_198,N_24973,N_24796);
or UO_199 (O_199,N_24968,N_24633);
nand UO_200 (O_200,N_24656,N_24556);
and UO_201 (O_201,N_24805,N_24630);
or UO_202 (O_202,N_24511,N_24945);
xnor UO_203 (O_203,N_24607,N_24799);
xor UO_204 (O_204,N_24915,N_24761);
xnor UO_205 (O_205,N_24978,N_24552);
or UO_206 (O_206,N_24561,N_24970);
xnor UO_207 (O_207,N_24829,N_24843);
nand UO_208 (O_208,N_24705,N_24688);
xnor UO_209 (O_209,N_24889,N_24606);
nand UO_210 (O_210,N_24515,N_24551);
and UO_211 (O_211,N_24917,N_24517);
xor UO_212 (O_212,N_24643,N_24998);
or UO_213 (O_213,N_24741,N_24944);
nand UO_214 (O_214,N_24776,N_24875);
or UO_215 (O_215,N_24764,N_24647);
and UO_216 (O_216,N_24508,N_24707);
nor UO_217 (O_217,N_24922,N_24765);
nor UO_218 (O_218,N_24996,N_24991);
xor UO_219 (O_219,N_24617,N_24731);
and UO_220 (O_220,N_24999,N_24885);
or UO_221 (O_221,N_24844,N_24682);
or UO_222 (O_222,N_24783,N_24542);
or UO_223 (O_223,N_24637,N_24827);
nand UO_224 (O_224,N_24951,N_24942);
or UO_225 (O_225,N_24806,N_24987);
and UO_226 (O_226,N_24675,N_24699);
and UO_227 (O_227,N_24653,N_24983);
nand UO_228 (O_228,N_24848,N_24929);
or UO_229 (O_229,N_24807,N_24516);
or UO_230 (O_230,N_24514,N_24769);
xnor UO_231 (O_231,N_24837,N_24946);
nor UO_232 (O_232,N_24620,N_24888);
and UO_233 (O_233,N_24588,N_24651);
xnor UO_234 (O_234,N_24976,N_24650);
or UO_235 (O_235,N_24821,N_24503);
xor UO_236 (O_236,N_24730,N_24605);
xnor UO_237 (O_237,N_24790,N_24981);
xnor UO_238 (O_238,N_24822,N_24638);
or UO_239 (O_239,N_24715,N_24569);
nor UO_240 (O_240,N_24626,N_24835);
or UO_241 (O_241,N_24654,N_24619);
or UO_242 (O_242,N_24937,N_24521);
nand UO_243 (O_243,N_24632,N_24535);
and UO_244 (O_244,N_24609,N_24872);
and UO_245 (O_245,N_24830,N_24526);
or UO_246 (O_246,N_24887,N_24995);
nand UO_247 (O_247,N_24988,N_24778);
and UO_248 (O_248,N_24565,N_24909);
and UO_249 (O_249,N_24953,N_24902);
and UO_250 (O_250,N_24770,N_24901);
nand UO_251 (O_251,N_24792,N_24877);
or UO_252 (O_252,N_24742,N_24885);
nor UO_253 (O_253,N_24530,N_24549);
or UO_254 (O_254,N_24886,N_24974);
nand UO_255 (O_255,N_24867,N_24825);
and UO_256 (O_256,N_24801,N_24609);
nand UO_257 (O_257,N_24796,N_24979);
nand UO_258 (O_258,N_24894,N_24727);
nand UO_259 (O_259,N_24508,N_24600);
and UO_260 (O_260,N_24966,N_24997);
nand UO_261 (O_261,N_24956,N_24986);
and UO_262 (O_262,N_24723,N_24887);
and UO_263 (O_263,N_24888,N_24965);
and UO_264 (O_264,N_24933,N_24871);
xnor UO_265 (O_265,N_24959,N_24534);
xor UO_266 (O_266,N_24539,N_24777);
nand UO_267 (O_267,N_24881,N_24809);
and UO_268 (O_268,N_24613,N_24511);
nor UO_269 (O_269,N_24763,N_24810);
xor UO_270 (O_270,N_24956,N_24678);
nor UO_271 (O_271,N_24944,N_24738);
or UO_272 (O_272,N_24649,N_24537);
nor UO_273 (O_273,N_24769,N_24534);
or UO_274 (O_274,N_24634,N_24641);
or UO_275 (O_275,N_24735,N_24822);
or UO_276 (O_276,N_24503,N_24740);
nor UO_277 (O_277,N_24857,N_24916);
and UO_278 (O_278,N_24809,N_24644);
nor UO_279 (O_279,N_24860,N_24507);
or UO_280 (O_280,N_24515,N_24964);
nand UO_281 (O_281,N_24935,N_24854);
and UO_282 (O_282,N_24940,N_24777);
nor UO_283 (O_283,N_24767,N_24766);
nor UO_284 (O_284,N_24538,N_24725);
and UO_285 (O_285,N_24785,N_24585);
nor UO_286 (O_286,N_24723,N_24637);
and UO_287 (O_287,N_24689,N_24976);
xnor UO_288 (O_288,N_24772,N_24832);
and UO_289 (O_289,N_24691,N_24652);
or UO_290 (O_290,N_24585,N_24523);
or UO_291 (O_291,N_24920,N_24700);
nand UO_292 (O_292,N_24582,N_24538);
xnor UO_293 (O_293,N_24761,N_24800);
nand UO_294 (O_294,N_24550,N_24947);
or UO_295 (O_295,N_24662,N_24625);
nand UO_296 (O_296,N_24835,N_24569);
or UO_297 (O_297,N_24526,N_24543);
or UO_298 (O_298,N_24536,N_24585);
xnor UO_299 (O_299,N_24729,N_24844);
nor UO_300 (O_300,N_24887,N_24926);
nor UO_301 (O_301,N_24837,N_24632);
nor UO_302 (O_302,N_24823,N_24704);
and UO_303 (O_303,N_24534,N_24898);
nor UO_304 (O_304,N_24705,N_24728);
and UO_305 (O_305,N_24756,N_24722);
xnor UO_306 (O_306,N_24546,N_24677);
nand UO_307 (O_307,N_24702,N_24752);
nor UO_308 (O_308,N_24999,N_24500);
nor UO_309 (O_309,N_24922,N_24974);
nor UO_310 (O_310,N_24636,N_24950);
xnor UO_311 (O_311,N_24508,N_24847);
nand UO_312 (O_312,N_24858,N_24884);
and UO_313 (O_313,N_24549,N_24938);
xor UO_314 (O_314,N_24673,N_24904);
nor UO_315 (O_315,N_24974,N_24724);
nand UO_316 (O_316,N_24665,N_24599);
nand UO_317 (O_317,N_24597,N_24644);
and UO_318 (O_318,N_24743,N_24824);
and UO_319 (O_319,N_24853,N_24584);
nand UO_320 (O_320,N_24610,N_24633);
xnor UO_321 (O_321,N_24644,N_24571);
and UO_322 (O_322,N_24618,N_24503);
xnor UO_323 (O_323,N_24506,N_24898);
nor UO_324 (O_324,N_24950,N_24558);
and UO_325 (O_325,N_24603,N_24662);
nor UO_326 (O_326,N_24803,N_24623);
xnor UO_327 (O_327,N_24951,N_24577);
nor UO_328 (O_328,N_24690,N_24511);
nand UO_329 (O_329,N_24936,N_24641);
nand UO_330 (O_330,N_24515,N_24686);
xor UO_331 (O_331,N_24919,N_24554);
nand UO_332 (O_332,N_24663,N_24553);
nor UO_333 (O_333,N_24544,N_24824);
and UO_334 (O_334,N_24657,N_24929);
or UO_335 (O_335,N_24964,N_24948);
xnor UO_336 (O_336,N_24980,N_24880);
nor UO_337 (O_337,N_24600,N_24591);
xnor UO_338 (O_338,N_24507,N_24787);
nor UO_339 (O_339,N_24896,N_24526);
and UO_340 (O_340,N_24965,N_24597);
nor UO_341 (O_341,N_24506,N_24531);
nand UO_342 (O_342,N_24615,N_24630);
xnor UO_343 (O_343,N_24703,N_24599);
and UO_344 (O_344,N_24538,N_24833);
and UO_345 (O_345,N_24695,N_24829);
or UO_346 (O_346,N_24800,N_24974);
nor UO_347 (O_347,N_24893,N_24606);
or UO_348 (O_348,N_24842,N_24940);
or UO_349 (O_349,N_24777,N_24745);
or UO_350 (O_350,N_24528,N_24504);
or UO_351 (O_351,N_24911,N_24843);
nand UO_352 (O_352,N_24951,N_24627);
or UO_353 (O_353,N_24861,N_24887);
or UO_354 (O_354,N_24956,N_24602);
or UO_355 (O_355,N_24658,N_24770);
and UO_356 (O_356,N_24646,N_24946);
nand UO_357 (O_357,N_24605,N_24900);
or UO_358 (O_358,N_24987,N_24962);
or UO_359 (O_359,N_24620,N_24644);
or UO_360 (O_360,N_24768,N_24575);
xor UO_361 (O_361,N_24517,N_24943);
xor UO_362 (O_362,N_24612,N_24743);
or UO_363 (O_363,N_24878,N_24717);
xor UO_364 (O_364,N_24974,N_24642);
and UO_365 (O_365,N_24563,N_24811);
and UO_366 (O_366,N_24750,N_24988);
nor UO_367 (O_367,N_24624,N_24646);
xor UO_368 (O_368,N_24707,N_24787);
or UO_369 (O_369,N_24713,N_24784);
nand UO_370 (O_370,N_24929,N_24631);
and UO_371 (O_371,N_24728,N_24698);
or UO_372 (O_372,N_24830,N_24855);
or UO_373 (O_373,N_24797,N_24513);
nand UO_374 (O_374,N_24890,N_24825);
nor UO_375 (O_375,N_24699,N_24859);
xor UO_376 (O_376,N_24536,N_24595);
nand UO_377 (O_377,N_24894,N_24614);
and UO_378 (O_378,N_24704,N_24878);
xor UO_379 (O_379,N_24937,N_24958);
nor UO_380 (O_380,N_24899,N_24800);
nand UO_381 (O_381,N_24708,N_24808);
nand UO_382 (O_382,N_24961,N_24917);
and UO_383 (O_383,N_24839,N_24982);
nor UO_384 (O_384,N_24623,N_24587);
nand UO_385 (O_385,N_24629,N_24674);
nor UO_386 (O_386,N_24757,N_24526);
nor UO_387 (O_387,N_24774,N_24906);
xor UO_388 (O_388,N_24696,N_24921);
nor UO_389 (O_389,N_24910,N_24880);
nor UO_390 (O_390,N_24552,N_24727);
nand UO_391 (O_391,N_24543,N_24858);
and UO_392 (O_392,N_24646,N_24564);
or UO_393 (O_393,N_24518,N_24566);
or UO_394 (O_394,N_24882,N_24786);
xnor UO_395 (O_395,N_24745,N_24616);
nand UO_396 (O_396,N_24665,N_24683);
nor UO_397 (O_397,N_24754,N_24747);
or UO_398 (O_398,N_24759,N_24565);
nand UO_399 (O_399,N_24839,N_24970);
nand UO_400 (O_400,N_24622,N_24955);
nor UO_401 (O_401,N_24553,N_24848);
nand UO_402 (O_402,N_24667,N_24514);
nor UO_403 (O_403,N_24990,N_24791);
or UO_404 (O_404,N_24843,N_24515);
nor UO_405 (O_405,N_24743,N_24789);
xor UO_406 (O_406,N_24699,N_24617);
nor UO_407 (O_407,N_24926,N_24596);
nor UO_408 (O_408,N_24648,N_24849);
or UO_409 (O_409,N_24611,N_24642);
or UO_410 (O_410,N_24588,N_24643);
xnor UO_411 (O_411,N_24976,N_24541);
nor UO_412 (O_412,N_24565,N_24796);
nand UO_413 (O_413,N_24526,N_24800);
and UO_414 (O_414,N_24749,N_24877);
and UO_415 (O_415,N_24550,N_24935);
xnor UO_416 (O_416,N_24733,N_24753);
or UO_417 (O_417,N_24822,N_24720);
nand UO_418 (O_418,N_24640,N_24863);
nand UO_419 (O_419,N_24857,N_24933);
nor UO_420 (O_420,N_24863,N_24572);
or UO_421 (O_421,N_24518,N_24811);
and UO_422 (O_422,N_24625,N_24846);
nand UO_423 (O_423,N_24900,N_24781);
nand UO_424 (O_424,N_24869,N_24740);
and UO_425 (O_425,N_24959,N_24589);
and UO_426 (O_426,N_24511,N_24857);
and UO_427 (O_427,N_24708,N_24693);
nand UO_428 (O_428,N_24921,N_24743);
nand UO_429 (O_429,N_24766,N_24990);
xnor UO_430 (O_430,N_24661,N_24863);
and UO_431 (O_431,N_24526,N_24797);
nand UO_432 (O_432,N_24633,N_24916);
or UO_433 (O_433,N_24887,N_24692);
and UO_434 (O_434,N_24733,N_24867);
nand UO_435 (O_435,N_24951,N_24985);
or UO_436 (O_436,N_24580,N_24648);
nor UO_437 (O_437,N_24573,N_24619);
nor UO_438 (O_438,N_24661,N_24686);
nor UO_439 (O_439,N_24923,N_24931);
and UO_440 (O_440,N_24684,N_24809);
and UO_441 (O_441,N_24740,N_24647);
and UO_442 (O_442,N_24618,N_24922);
xnor UO_443 (O_443,N_24651,N_24521);
nor UO_444 (O_444,N_24954,N_24573);
xnor UO_445 (O_445,N_24619,N_24966);
or UO_446 (O_446,N_24897,N_24715);
xor UO_447 (O_447,N_24592,N_24772);
nand UO_448 (O_448,N_24864,N_24608);
nor UO_449 (O_449,N_24890,N_24538);
xnor UO_450 (O_450,N_24600,N_24916);
nand UO_451 (O_451,N_24615,N_24952);
and UO_452 (O_452,N_24622,N_24516);
nand UO_453 (O_453,N_24596,N_24955);
nand UO_454 (O_454,N_24915,N_24521);
nor UO_455 (O_455,N_24584,N_24939);
or UO_456 (O_456,N_24573,N_24920);
or UO_457 (O_457,N_24514,N_24948);
xnor UO_458 (O_458,N_24535,N_24777);
and UO_459 (O_459,N_24746,N_24510);
xor UO_460 (O_460,N_24912,N_24592);
nand UO_461 (O_461,N_24847,N_24988);
xor UO_462 (O_462,N_24809,N_24734);
or UO_463 (O_463,N_24719,N_24911);
or UO_464 (O_464,N_24571,N_24822);
or UO_465 (O_465,N_24586,N_24621);
nand UO_466 (O_466,N_24504,N_24701);
nand UO_467 (O_467,N_24779,N_24551);
nand UO_468 (O_468,N_24525,N_24855);
nand UO_469 (O_469,N_24518,N_24845);
and UO_470 (O_470,N_24956,N_24850);
or UO_471 (O_471,N_24703,N_24692);
nand UO_472 (O_472,N_24806,N_24871);
nor UO_473 (O_473,N_24866,N_24873);
nand UO_474 (O_474,N_24794,N_24637);
nor UO_475 (O_475,N_24584,N_24813);
nand UO_476 (O_476,N_24878,N_24628);
nor UO_477 (O_477,N_24662,N_24709);
nand UO_478 (O_478,N_24810,N_24537);
nor UO_479 (O_479,N_24801,N_24831);
nand UO_480 (O_480,N_24504,N_24554);
or UO_481 (O_481,N_24509,N_24853);
nor UO_482 (O_482,N_24637,N_24709);
and UO_483 (O_483,N_24755,N_24670);
nand UO_484 (O_484,N_24586,N_24629);
or UO_485 (O_485,N_24649,N_24894);
nand UO_486 (O_486,N_24885,N_24906);
xor UO_487 (O_487,N_24724,N_24666);
or UO_488 (O_488,N_24873,N_24617);
nand UO_489 (O_489,N_24524,N_24886);
nand UO_490 (O_490,N_24546,N_24693);
xnor UO_491 (O_491,N_24739,N_24854);
nor UO_492 (O_492,N_24786,N_24944);
and UO_493 (O_493,N_24588,N_24545);
nand UO_494 (O_494,N_24896,N_24578);
nor UO_495 (O_495,N_24804,N_24794);
or UO_496 (O_496,N_24557,N_24884);
nor UO_497 (O_497,N_24865,N_24633);
and UO_498 (O_498,N_24997,N_24700);
nand UO_499 (O_499,N_24626,N_24585);
nor UO_500 (O_500,N_24715,N_24584);
nand UO_501 (O_501,N_24722,N_24911);
and UO_502 (O_502,N_24851,N_24781);
or UO_503 (O_503,N_24589,N_24684);
and UO_504 (O_504,N_24949,N_24926);
nand UO_505 (O_505,N_24541,N_24677);
xnor UO_506 (O_506,N_24565,N_24813);
or UO_507 (O_507,N_24824,N_24874);
and UO_508 (O_508,N_24762,N_24803);
nand UO_509 (O_509,N_24828,N_24560);
or UO_510 (O_510,N_24672,N_24685);
and UO_511 (O_511,N_24925,N_24645);
xor UO_512 (O_512,N_24918,N_24865);
xnor UO_513 (O_513,N_24858,N_24910);
or UO_514 (O_514,N_24800,N_24573);
xnor UO_515 (O_515,N_24700,N_24709);
or UO_516 (O_516,N_24603,N_24624);
nor UO_517 (O_517,N_24614,N_24862);
nor UO_518 (O_518,N_24960,N_24876);
nor UO_519 (O_519,N_24691,N_24816);
xor UO_520 (O_520,N_24696,N_24743);
nor UO_521 (O_521,N_24524,N_24552);
or UO_522 (O_522,N_24940,N_24641);
nand UO_523 (O_523,N_24703,N_24854);
nor UO_524 (O_524,N_24859,N_24508);
nand UO_525 (O_525,N_24670,N_24732);
or UO_526 (O_526,N_24854,N_24895);
xnor UO_527 (O_527,N_24799,N_24825);
and UO_528 (O_528,N_24507,N_24793);
or UO_529 (O_529,N_24787,N_24599);
or UO_530 (O_530,N_24559,N_24568);
xnor UO_531 (O_531,N_24637,N_24940);
xnor UO_532 (O_532,N_24571,N_24711);
or UO_533 (O_533,N_24894,N_24757);
and UO_534 (O_534,N_24886,N_24804);
and UO_535 (O_535,N_24778,N_24969);
xor UO_536 (O_536,N_24612,N_24719);
nor UO_537 (O_537,N_24716,N_24614);
and UO_538 (O_538,N_24704,N_24530);
nor UO_539 (O_539,N_24659,N_24902);
xnor UO_540 (O_540,N_24825,N_24677);
nor UO_541 (O_541,N_24747,N_24597);
nor UO_542 (O_542,N_24699,N_24759);
xnor UO_543 (O_543,N_24818,N_24535);
nor UO_544 (O_544,N_24654,N_24657);
nor UO_545 (O_545,N_24880,N_24649);
nand UO_546 (O_546,N_24834,N_24996);
and UO_547 (O_547,N_24566,N_24822);
nand UO_548 (O_548,N_24766,N_24846);
nor UO_549 (O_549,N_24612,N_24853);
nand UO_550 (O_550,N_24770,N_24921);
or UO_551 (O_551,N_24903,N_24941);
xnor UO_552 (O_552,N_24892,N_24880);
nor UO_553 (O_553,N_24525,N_24980);
and UO_554 (O_554,N_24899,N_24641);
nor UO_555 (O_555,N_24679,N_24782);
or UO_556 (O_556,N_24911,N_24569);
or UO_557 (O_557,N_24655,N_24699);
nand UO_558 (O_558,N_24581,N_24858);
nand UO_559 (O_559,N_24901,N_24560);
xnor UO_560 (O_560,N_24627,N_24945);
nand UO_561 (O_561,N_24930,N_24641);
and UO_562 (O_562,N_24537,N_24647);
nor UO_563 (O_563,N_24603,N_24805);
xor UO_564 (O_564,N_24518,N_24657);
xnor UO_565 (O_565,N_24712,N_24707);
or UO_566 (O_566,N_24938,N_24511);
nor UO_567 (O_567,N_24872,N_24884);
and UO_568 (O_568,N_24679,N_24553);
or UO_569 (O_569,N_24882,N_24986);
and UO_570 (O_570,N_24518,N_24938);
nand UO_571 (O_571,N_24857,N_24614);
and UO_572 (O_572,N_24590,N_24683);
nand UO_573 (O_573,N_24500,N_24844);
nand UO_574 (O_574,N_24943,N_24952);
or UO_575 (O_575,N_24970,N_24516);
nand UO_576 (O_576,N_24772,N_24746);
nor UO_577 (O_577,N_24550,N_24598);
and UO_578 (O_578,N_24988,N_24928);
and UO_579 (O_579,N_24828,N_24834);
nand UO_580 (O_580,N_24788,N_24924);
nor UO_581 (O_581,N_24914,N_24540);
nand UO_582 (O_582,N_24542,N_24501);
or UO_583 (O_583,N_24919,N_24878);
nor UO_584 (O_584,N_24909,N_24568);
nand UO_585 (O_585,N_24634,N_24653);
nor UO_586 (O_586,N_24798,N_24981);
or UO_587 (O_587,N_24500,N_24623);
nor UO_588 (O_588,N_24870,N_24596);
or UO_589 (O_589,N_24766,N_24909);
or UO_590 (O_590,N_24815,N_24907);
and UO_591 (O_591,N_24888,N_24757);
and UO_592 (O_592,N_24611,N_24508);
nor UO_593 (O_593,N_24750,N_24868);
and UO_594 (O_594,N_24748,N_24605);
nor UO_595 (O_595,N_24900,N_24768);
nand UO_596 (O_596,N_24945,N_24574);
nor UO_597 (O_597,N_24954,N_24692);
and UO_598 (O_598,N_24659,N_24519);
xor UO_599 (O_599,N_24888,N_24600);
or UO_600 (O_600,N_24624,N_24568);
nand UO_601 (O_601,N_24722,N_24648);
nand UO_602 (O_602,N_24894,N_24898);
nor UO_603 (O_603,N_24630,N_24832);
nor UO_604 (O_604,N_24829,N_24906);
and UO_605 (O_605,N_24546,N_24981);
nor UO_606 (O_606,N_24568,N_24768);
nand UO_607 (O_607,N_24712,N_24776);
and UO_608 (O_608,N_24837,N_24649);
nor UO_609 (O_609,N_24661,N_24774);
nand UO_610 (O_610,N_24758,N_24688);
nor UO_611 (O_611,N_24548,N_24850);
nor UO_612 (O_612,N_24735,N_24983);
nor UO_613 (O_613,N_24635,N_24696);
xnor UO_614 (O_614,N_24731,N_24898);
and UO_615 (O_615,N_24901,N_24960);
nor UO_616 (O_616,N_24521,N_24893);
nand UO_617 (O_617,N_24743,N_24588);
xor UO_618 (O_618,N_24849,N_24926);
or UO_619 (O_619,N_24848,N_24871);
and UO_620 (O_620,N_24673,N_24547);
xor UO_621 (O_621,N_24528,N_24706);
nor UO_622 (O_622,N_24941,N_24628);
or UO_623 (O_623,N_24788,N_24536);
or UO_624 (O_624,N_24741,N_24644);
or UO_625 (O_625,N_24790,N_24713);
nor UO_626 (O_626,N_24604,N_24826);
or UO_627 (O_627,N_24648,N_24989);
nor UO_628 (O_628,N_24838,N_24714);
and UO_629 (O_629,N_24822,N_24876);
nor UO_630 (O_630,N_24971,N_24773);
and UO_631 (O_631,N_24982,N_24781);
nand UO_632 (O_632,N_24535,N_24995);
nand UO_633 (O_633,N_24954,N_24911);
or UO_634 (O_634,N_24752,N_24997);
or UO_635 (O_635,N_24542,N_24869);
and UO_636 (O_636,N_24758,N_24956);
nor UO_637 (O_637,N_24907,N_24919);
xor UO_638 (O_638,N_24663,N_24851);
or UO_639 (O_639,N_24669,N_24940);
and UO_640 (O_640,N_24611,N_24551);
xnor UO_641 (O_641,N_24727,N_24560);
nor UO_642 (O_642,N_24508,N_24767);
or UO_643 (O_643,N_24704,N_24750);
and UO_644 (O_644,N_24571,N_24540);
or UO_645 (O_645,N_24923,N_24544);
or UO_646 (O_646,N_24715,N_24779);
nor UO_647 (O_647,N_24628,N_24552);
xor UO_648 (O_648,N_24890,N_24563);
nand UO_649 (O_649,N_24745,N_24697);
nor UO_650 (O_650,N_24873,N_24648);
and UO_651 (O_651,N_24622,N_24931);
nand UO_652 (O_652,N_24867,N_24739);
and UO_653 (O_653,N_24598,N_24745);
nand UO_654 (O_654,N_24552,N_24988);
xnor UO_655 (O_655,N_24633,N_24842);
xnor UO_656 (O_656,N_24569,N_24638);
and UO_657 (O_657,N_24848,N_24820);
nand UO_658 (O_658,N_24810,N_24592);
or UO_659 (O_659,N_24934,N_24782);
nand UO_660 (O_660,N_24765,N_24833);
or UO_661 (O_661,N_24812,N_24618);
nand UO_662 (O_662,N_24573,N_24643);
nand UO_663 (O_663,N_24681,N_24993);
or UO_664 (O_664,N_24675,N_24545);
nor UO_665 (O_665,N_24677,N_24702);
nor UO_666 (O_666,N_24911,N_24585);
or UO_667 (O_667,N_24610,N_24733);
and UO_668 (O_668,N_24629,N_24994);
xor UO_669 (O_669,N_24676,N_24638);
xnor UO_670 (O_670,N_24766,N_24985);
and UO_671 (O_671,N_24963,N_24502);
nor UO_672 (O_672,N_24997,N_24563);
nand UO_673 (O_673,N_24848,N_24523);
and UO_674 (O_674,N_24584,N_24640);
nor UO_675 (O_675,N_24502,N_24684);
nor UO_676 (O_676,N_24910,N_24891);
xor UO_677 (O_677,N_24859,N_24781);
nand UO_678 (O_678,N_24866,N_24861);
or UO_679 (O_679,N_24963,N_24854);
and UO_680 (O_680,N_24523,N_24630);
xnor UO_681 (O_681,N_24748,N_24691);
or UO_682 (O_682,N_24645,N_24998);
and UO_683 (O_683,N_24523,N_24853);
or UO_684 (O_684,N_24674,N_24807);
nand UO_685 (O_685,N_24713,N_24570);
nor UO_686 (O_686,N_24939,N_24951);
and UO_687 (O_687,N_24721,N_24855);
nand UO_688 (O_688,N_24573,N_24712);
nand UO_689 (O_689,N_24786,N_24555);
or UO_690 (O_690,N_24666,N_24811);
or UO_691 (O_691,N_24774,N_24616);
xor UO_692 (O_692,N_24787,N_24556);
nand UO_693 (O_693,N_24851,N_24595);
nor UO_694 (O_694,N_24886,N_24634);
nand UO_695 (O_695,N_24615,N_24980);
nor UO_696 (O_696,N_24688,N_24829);
and UO_697 (O_697,N_24967,N_24604);
xnor UO_698 (O_698,N_24508,N_24963);
and UO_699 (O_699,N_24919,N_24977);
nor UO_700 (O_700,N_24580,N_24641);
nand UO_701 (O_701,N_24658,N_24974);
xnor UO_702 (O_702,N_24878,N_24727);
or UO_703 (O_703,N_24542,N_24938);
and UO_704 (O_704,N_24757,N_24723);
xnor UO_705 (O_705,N_24693,N_24946);
or UO_706 (O_706,N_24598,N_24733);
nand UO_707 (O_707,N_24734,N_24726);
nor UO_708 (O_708,N_24706,N_24742);
nor UO_709 (O_709,N_24772,N_24508);
nand UO_710 (O_710,N_24732,N_24506);
xnor UO_711 (O_711,N_24656,N_24790);
or UO_712 (O_712,N_24768,N_24672);
and UO_713 (O_713,N_24544,N_24899);
and UO_714 (O_714,N_24773,N_24610);
nand UO_715 (O_715,N_24903,N_24740);
nor UO_716 (O_716,N_24929,N_24790);
xnor UO_717 (O_717,N_24888,N_24569);
nand UO_718 (O_718,N_24930,N_24666);
xor UO_719 (O_719,N_24933,N_24692);
nor UO_720 (O_720,N_24589,N_24647);
xnor UO_721 (O_721,N_24582,N_24532);
nand UO_722 (O_722,N_24981,N_24926);
nor UO_723 (O_723,N_24646,N_24580);
xnor UO_724 (O_724,N_24600,N_24810);
or UO_725 (O_725,N_24530,N_24994);
or UO_726 (O_726,N_24976,N_24982);
nand UO_727 (O_727,N_24654,N_24524);
xnor UO_728 (O_728,N_24540,N_24637);
xnor UO_729 (O_729,N_24732,N_24905);
or UO_730 (O_730,N_24799,N_24966);
nand UO_731 (O_731,N_24794,N_24712);
or UO_732 (O_732,N_24649,N_24675);
xor UO_733 (O_733,N_24739,N_24907);
or UO_734 (O_734,N_24679,N_24519);
nand UO_735 (O_735,N_24560,N_24503);
or UO_736 (O_736,N_24753,N_24986);
nand UO_737 (O_737,N_24849,N_24701);
nor UO_738 (O_738,N_24503,N_24878);
nor UO_739 (O_739,N_24577,N_24775);
or UO_740 (O_740,N_24628,N_24682);
xor UO_741 (O_741,N_24618,N_24585);
or UO_742 (O_742,N_24920,N_24871);
nor UO_743 (O_743,N_24912,N_24626);
or UO_744 (O_744,N_24602,N_24975);
nor UO_745 (O_745,N_24691,N_24932);
nand UO_746 (O_746,N_24607,N_24519);
nand UO_747 (O_747,N_24886,N_24881);
xnor UO_748 (O_748,N_24917,N_24795);
or UO_749 (O_749,N_24977,N_24776);
nand UO_750 (O_750,N_24766,N_24986);
and UO_751 (O_751,N_24953,N_24991);
nor UO_752 (O_752,N_24578,N_24933);
xor UO_753 (O_753,N_24513,N_24712);
nand UO_754 (O_754,N_24824,N_24972);
or UO_755 (O_755,N_24827,N_24661);
xor UO_756 (O_756,N_24944,N_24540);
or UO_757 (O_757,N_24856,N_24579);
and UO_758 (O_758,N_24954,N_24598);
nor UO_759 (O_759,N_24779,N_24844);
or UO_760 (O_760,N_24796,N_24718);
nand UO_761 (O_761,N_24767,N_24972);
or UO_762 (O_762,N_24799,N_24609);
nand UO_763 (O_763,N_24967,N_24805);
or UO_764 (O_764,N_24650,N_24619);
and UO_765 (O_765,N_24856,N_24994);
nor UO_766 (O_766,N_24752,N_24897);
and UO_767 (O_767,N_24668,N_24816);
or UO_768 (O_768,N_24630,N_24651);
nor UO_769 (O_769,N_24768,N_24899);
nor UO_770 (O_770,N_24742,N_24528);
xor UO_771 (O_771,N_24579,N_24679);
and UO_772 (O_772,N_24564,N_24928);
nand UO_773 (O_773,N_24661,N_24943);
and UO_774 (O_774,N_24735,N_24624);
xnor UO_775 (O_775,N_24725,N_24881);
nand UO_776 (O_776,N_24510,N_24743);
or UO_777 (O_777,N_24836,N_24805);
nand UO_778 (O_778,N_24612,N_24629);
or UO_779 (O_779,N_24908,N_24512);
nand UO_780 (O_780,N_24863,N_24524);
nor UO_781 (O_781,N_24736,N_24702);
nand UO_782 (O_782,N_24794,N_24808);
nand UO_783 (O_783,N_24825,N_24817);
or UO_784 (O_784,N_24983,N_24656);
or UO_785 (O_785,N_24652,N_24695);
xnor UO_786 (O_786,N_24923,N_24707);
and UO_787 (O_787,N_24980,N_24698);
nand UO_788 (O_788,N_24829,N_24631);
or UO_789 (O_789,N_24912,N_24552);
or UO_790 (O_790,N_24817,N_24967);
and UO_791 (O_791,N_24716,N_24776);
nor UO_792 (O_792,N_24602,N_24571);
nor UO_793 (O_793,N_24633,N_24991);
xnor UO_794 (O_794,N_24624,N_24732);
xnor UO_795 (O_795,N_24727,N_24606);
nor UO_796 (O_796,N_24750,N_24989);
nand UO_797 (O_797,N_24563,N_24976);
xnor UO_798 (O_798,N_24571,N_24528);
xor UO_799 (O_799,N_24706,N_24950);
nand UO_800 (O_800,N_24650,N_24582);
nand UO_801 (O_801,N_24932,N_24603);
xor UO_802 (O_802,N_24845,N_24667);
nor UO_803 (O_803,N_24579,N_24854);
nor UO_804 (O_804,N_24735,N_24579);
nand UO_805 (O_805,N_24601,N_24953);
nor UO_806 (O_806,N_24759,N_24912);
and UO_807 (O_807,N_24539,N_24758);
nor UO_808 (O_808,N_24741,N_24822);
xnor UO_809 (O_809,N_24961,N_24933);
xor UO_810 (O_810,N_24910,N_24838);
nand UO_811 (O_811,N_24629,N_24790);
and UO_812 (O_812,N_24767,N_24861);
and UO_813 (O_813,N_24952,N_24801);
and UO_814 (O_814,N_24926,N_24959);
nor UO_815 (O_815,N_24685,N_24682);
nand UO_816 (O_816,N_24833,N_24776);
xnor UO_817 (O_817,N_24613,N_24948);
or UO_818 (O_818,N_24640,N_24868);
nor UO_819 (O_819,N_24855,N_24518);
nor UO_820 (O_820,N_24835,N_24513);
xnor UO_821 (O_821,N_24637,N_24775);
nand UO_822 (O_822,N_24802,N_24940);
or UO_823 (O_823,N_24661,N_24826);
nand UO_824 (O_824,N_24763,N_24684);
or UO_825 (O_825,N_24570,N_24862);
nor UO_826 (O_826,N_24812,N_24630);
nand UO_827 (O_827,N_24990,N_24931);
nand UO_828 (O_828,N_24597,N_24673);
xnor UO_829 (O_829,N_24868,N_24533);
and UO_830 (O_830,N_24888,N_24843);
nand UO_831 (O_831,N_24938,N_24585);
xnor UO_832 (O_832,N_24583,N_24547);
nor UO_833 (O_833,N_24710,N_24831);
or UO_834 (O_834,N_24960,N_24898);
nor UO_835 (O_835,N_24667,N_24788);
nand UO_836 (O_836,N_24762,N_24649);
and UO_837 (O_837,N_24623,N_24745);
nor UO_838 (O_838,N_24900,N_24713);
or UO_839 (O_839,N_24658,N_24883);
xor UO_840 (O_840,N_24543,N_24627);
nor UO_841 (O_841,N_24884,N_24576);
nand UO_842 (O_842,N_24741,N_24993);
nand UO_843 (O_843,N_24699,N_24837);
xor UO_844 (O_844,N_24988,N_24904);
xor UO_845 (O_845,N_24641,N_24815);
nand UO_846 (O_846,N_24801,N_24752);
and UO_847 (O_847,N_24579,N_24547);
and UO_848 (O_848,N_24769,N_24913);
nor UO_849 (O_849,N_24586,N_24832);
xor UO_850 (O_850,N_24672,N_24844);
or UO_851 (O_851,N_24737,N_24533);
nor UO_852 (O_852,N_24993,N_24912);
nor UO_853 (O_853,N_24792,N_24830);
or UO_854 (O_854,N_24987,N_24849);
nor UO_855 (O_855,N_24894,N_24600);
or UO_856 (O_856,N_24634,N_24968);
nand UO_857 (O_857,N_24694,N_24958);
or UO_858 (O_858,N_24830,N_24864);
nand UO_859 (O_859,N_24972,N_24557);
nand UO_860 (O_860,N_24975,N_24726);
nand UO_861 (O_861,N_24864,N_24781);
nand UO_862 (O_862,N_24732,N_24536);
and UO_863 (O_863,N_24908,N_24605);
and UO_864 (O_864,N_24532,N_24849);
and UO_865 (O_865,N_24934,N_24952);
and UO_866 (O_866,N_24620,N_24756);
nand UO_867 (O_867,N_24913,N_24895);
xor UO_868 (O_868,N_24527,N_24726);
nand UO_869 (O_869,N_24800,N_24514);
nand UO_870 (O_870,N_24565,N_24853);
or UO_871 (O_871,N_24960,N_24988);
nand UO_872 (O_872,N_24887,N_24844);
xor UO_873 (O_873,N_24716,N_24777);
nand UO_874 (O_874,N_24562,N_24939);
nor UO_875 (O_875,N_24939,N_24701);
and UO_876 (O_876,N_24898,N_24635);
or UO_877 (O_877,N_24888,N_24848);
or UO_878 (O_878,N_24552,N_24619);
and UO_879 (O_879,N_24612,N_24757);
or UO_880 (O_880,N_24644,N_24500);
and UO_881 (O_881,N_24900,N_24686);
nand UO_882 (O_882,N_24924,N_24506);
xnor UO_883 (O_883,N_24524,N_24927);
or UO_884 (O_884,N_24641,N_24790);
and UO_885 (O_885,N_24733,N_24819);
nor UO_886 (O_886,N_24941,N_24945);
xor UO_887 (O_887,N_24607,N_24835);
or UO_888 (O_888,N_24932,N_24888);
or UO_889 (O_889,N_24780,N_24529);
nand UO_890 (O_890,N_24651,N_24726);
nand UO_891 (O_891,N_24936,N_24859);
and UO_892 (O_892,N_24692,N_24592);
and UO_893 (O_893,N_24549,N_24948);
and UO_894 (O_894,N_24793,N_24944);
xor UO_895 (O_895,N_24539,N_24598);
nand UO_896 (O_896,N_24969,N_24748);
xnor UO_897 (O_897,N_24921,N_24501);
nor UO_898 (O_898,N_24791,N_24687);
nand UO_899 (O_899,N_24815,N_24728);
xor UO_900 (O_900,N_24680,N_24800);
or UO_901 (O_901,N_24645,N_24573);
nand UO_902 (O_902,N_24686,N_24517);
nor UO_903 (O_903,N_24868,N_24659);
and UO_904 (O_904,N_24921,N_24876);
or UO_905 (O_905,N_24854,N_24617);
and UO_906 (O_906,N_24654,N_24847);
xor UO_907 (O_907,N_24512,N_24779);
and UO_908 (O_908,N_24680,N_24526);
nor UO_909 (O_909,N_24521,N_24702);
nor UO_910 (O_910,N_24793,N_24681);
and UO_911 (O_911,N_24894,N_24721);
or UO_912 (O_912,N_24823,N_24546);
nand UO_913 (O_913,N_24648,N_24766);
xor UO_914 (O_914,N_24986,N_24911);
xor UO_915 (O_915,N_24631,N_24564);
nand UO_916 (O_916,N_24938,N_24729);
nor UO_917 (O_917,N_24955,N_24661);
nand UO_918 (O_918,N_24737,N_24618);
nand UO_919 (O_919,N_24845,N_24622);
or UO_920 (O_920,N_24686,N_24595);
xor UO_921 (O_921,N_24762,N_24520);
nor UO_922 (O_922,N_24905,N_24603);
or UO_923 (O_923,N_24804,N_24752);
nand UO_924 (O_924,N_24650,N_24728);
and UO_925 (O_925,N_24911,N_24851);
or UO_926 (O_926,N_24672,N_24906);
xnor UO_927 (O_927,N_24914,N_24963);
or UO_928 (O_928,N_24540,N_24975);
nand UO_929 (O_929,N_24770,N_24816);
xnor UO_930 (O_930,N_24746,N_24662);
nor UO_931 (O_931,N_24776,N_24798);
nand UO_932 (O_932,N_24920,N_24588);
nand UO_933 (O_933,N_24526,N_24787);
xnor UO_934 (O_934,N_24795,N_24637);
nor UO_935 (O_935,N_24761,N_24842);
nor UO_936 (O_936,N_24948,N_24520);
nor UO_937 (O_937,N_24628,N_24549);
or UO_938 (O_938,N_24680,N_24555);
nor UO_939 (O_939,N_24646,N_24504);
xor UO_940 (O_940,N_24652,N_24615);
nor UO_941 (O_941,N_24998,N_24768);
xnor UO_942 (O_942,N_24676,N_24662);
nor UO_943 (O_943,N_24800,N_24777);
nor UO_944 (O_944,N_24565,N_24871);
nand UO_945 (O_945,N_24697,N_24557);
or UO_946 (O_946,N_24704,N_24954);
xnor UO_947 (O_947,N_24652,N_24869);
or UO_948 (O_948,N_24902,N_24840);
and UO_949 (O_949,N_24946,N_24913);
nand UO_950 (O_950,N_24678,N_24687);
xnor UO_951 (O_951,N_24636,N_24671);
and UO_952 (O_952,N_24827,N_24511);
xor UO_953 (O_953,N_24601,N_24567);
nand UO_954 (O_954,N_24771,N_24951);
or UO_955 (O_955,N_24589,N_24978);
and UO_956 (O_956,N_24507,N_24695);
xnor UO_957 (O_957,N_24787,N_24920);
nand UO_958 (O_958,N_24528,N_24668);
or UO_959 (O_959,N_24547,N_24729);
and UO_960 (O_960,N_24510,N_24582);
xor UO_961 (O_961,N_24809,N_24802);
or UO_962 (O_962,N_24864,N_24943);
or UO_963 (O_963,N_24922,N_24533);
xnor UO_964 (O_964,N_24946,N_24649);
or UO_965 (O_965,N_24621,N_24502);
nand UO_966 (O_966,N_24728,N_24991);
or UO_967 (O_967,N_24869,N_24983);
nor UO_968 (O_968,N_24716,N_24663);
nor UO_969 (O_969,N_24742,N_24556);
nand UO_970 (O_970,N_24772,N_24793);
xor UO_971 (O_971,N_24989,N_24591);
xnor UO_972 (O_972,N_24669,N_24762);
nand UO_973 (O_973,N_24960,N_24725);
nand UO_974 (O_974,N_24542,N_24563);
xor UO_975 (O_975,N_24840,N_24788);
or UO_976 (O_976,N_24533,N_24763);
and UO_977 (O_977,N_24870,N_24959);
and UO_978 (O_978,N_24958,N_24583);
xnor UO_979 (O_979,N_24510,N_24647);
nand UO_980 (O_980,N_24759,N_24638);
xnor UO_981 (O_981,N_24580,N_24933);
xor UO_982 (O_982,N_24893,N_24905);
xnor UO_983 (O_983,N_24810,N_24832);
nand UO_984 (O_984,N_24957,N_24811);
xnor UO_985 (O_985,N_24676,N_24852);
xor UO_986 (O_986,N_24551,N_24855);
nor UO_987 (O_987,N_24795,N_24683);
or UO_988 (O_988,N_24879,N_24620);
xor UO_989 (O_989,N_24745,N_24902);
and UO_990 (O_990,N_24961,N_24952);
or UO_991 (O_991,N_24788,N_24971);
and UO_992 (O_992,N_24948,N_24949);
xnor UO_993 (O_993,N_24767,N_24708);
and UO_994 (O_994,N_24644,N_24780);
xnor UO_995 (O_995,N_24818,N_24921);
or UO_996 (O_996,N_24874,N_24576);
and UO_997 (O_997,N_24972,N_24525);
and UO_998 (O_998,N_24516,N_24987);
and UO_999 (O_999,N_24688,N_24653);
xnor UO_1000 (O_1000,N_24813,N_24590);
xnor UO_1001 (O_1001,N_24704,N_24661);
or UO_1002 (O_1002,N_24910,N_24882);
or UO_1003 (O_1003,N_24608,N_24957);
nor UO_1004 (O_1004,N_24524,N_24761);
xor UO_1005 (O_1005,N_24884,N_24531);
and UO_1006 (O_1006,N_24849,N_24905);
or UO_1007 (O_1007,N_24738,N_24567);
xor UO_1008 (O_1008,N_24651,N_24550);
or UO_1009 (O_1009,N_24503,N_24759);
or UO_1010 (O_1010,N_24796,N_24582);
and UO_1011 (O_1011,N_24875,N_24907);
xor UO_1012 (O_1012,N_24766,N_24707);
nor UO_1013 (O_1013,N_24679,N_24885);
or UO_1014 (O_1014,N_24592,N_24585);
nor UO_1015 (O_1015,N_24963,N_24624);
and UO_1016 (O_1016,N_24817,N_24546);
nand UO_1017 (O_1017,N_24663,N_24567);
or UO_1018 (O_1018,N_24893,N_24596);
nor UO_1019 (O_1019,N_24555,N_24516);
xnor UO_1020 (O_1020,N_24829,N_24895);
or UO_1021 (O_1021,N_24792,N_24743);
or UO_1022 (O_1022,N_24527,N_24755);
xor UO_1023 (O_1023,N_24814,N_24563);
nand UO_1024 (O_1024,N_24617,N_24747);
nor UO_1025 (O_1025,N_24638,N_24623);
and UO_1026 (O_1026,N_24998,N_24600);
or UO_1027 (O_1027,N_24600,N_24983);
nand UO_1028 (O_1028,N_24627,N_24833);
nor UO_1029 (O_1029,N_24942,N_24917);
nor UO_1030 (O_1030,N_24847,N_24822);
xor UO_1031 (O_1031,N_24828,N_24635);
nand UO_1032 (O_1032,N_24633,N_24528);
nand UO_1033 (O_1033,N_24566,N_24747);
nor UO_1034 (O_1034,N_24906,N_24743);
xor UO_1035 (O_1035,N_24857,N_24737);
or UO_1036 (O_1036,N_24515,N_24597);
xnor UO_1037 (O_1037,N_24822,N_24840);
nand UO_1038 (O_1038,N_24775,N_24752);
or UO_1039 (O_1039,N_24560,N_24927);
nor UO_1040 (O_1040,N_24665,N_24862);
or UO_1041 (O_1041,N_24894,N_24810);
xor UO_1042 (O_1042,N_24553,N_24502);
nand UO_1043 (O_1043,N_24686,N_24918);
and UO_1044 (O_1044,N_24696,N_24931);
and UO_1045 (O_1045,N_24663,N_24747);
and UO_1046 (O_1046,N_24997,N_24538);
nand UO_1047 (O_1047,N_24531,N_24507);
xnor UO_1048 (O_1048,N_24519,N_24765);
or UO_1049 (O_1049,N_24591,N_24833);
xor UO_1050 (O_1050,N_24738,N_24726);
and UO_1051 (O_1051,N_24966,N_24825);
or UO_1052 (O_1052,N_24944,N_24906);
and UO_1053 (O_1053,N_24501,N_24746);
and UO_1054 (O_1054,N_24534,N_24893);
and UO_1055 (O_1055,N_24598,N_24655);
nand UO_1056 (O_1056,N_24650,N_24523);
nand UO_1057 (O_1057,N_24798,N_24951);
nand UO_1058 (O_1058,N_24538,N_24517);
or UO_1059 (O_1059,N_24875,N_24970);
nand UO_1060 (O_1060,N_24893,N_24765);
nand UO_1061 (O_1061,N_24872,N_24844);
xor UO_1062 (O_1062,N_24816,N_24789);
xor UO_1063 (O_1063,N_24620,N_24551);
nand UO_1064 (O_1064,N_24548,N_24865);
or UO_1065 (O_1065,N_24618,N_24947);
nand UO_1066 (O_1066,N_24655,N_24937);
nand UO_1067 (O_1067,N_24899,N_24975);
and UO_1068 (O_1068,N_24989,N_24926);
xor UO_1069 (O_1069,N_24721,N_24991);
xnor UO_1070 (O_1070,N_24871,N_24832);
xnor UO_1071 (O_1071,N_24975,N_24534);
and UO_1072 (O_1072,N_24905,N_24815);
nor UO_1073 (O_1073,N_24762,N_24756);
nor UO_1074 (O_1074,N_24967,N_24576);
and UO_1075 (O_1075,N_24757,N_24832);
nand UO_1076 (O_1076,N_24898,N_24664);
nor UO_1077 (O_1077,N_24572,N_24639);
or UO_1078 (O_1078,N_24657,N_24650);
or UO_1079 (O_1079,N_24664,N_24708);
nand UO_1080 (O_1080,N_24888,N_24962);
or UO_1081 (O_1081,N_24608,N_24564);
xnor UO_1082 (O_1082,N_24649,N_24858);
and UO_1083 (O_1083,N_24928,N_24888);
or UO_1084 (O_1084,N_24548,N_24672);
and UO_1085 (O_1085,N_24639,N_24560);
nand UO_1086 (O_1086,N_24607,N_24548);
and UO_1087 (O_1087,N_24770,N_24920);
or UO_1088 (O_1088,N_24817,N_24664);
xor UO_1089 (O_1089,N_24504,N_24638);
xnor UO_1090 (O_1090,N_24643,N_24595);
xor UO_1091 (O_1091,N_24769,N_24541);
and UO_1092 (O_1092,N_24640,N_24676);
or UO_1093 (O_1093,N_24746,N_24799);
nand UO_1094 (O_1094,N_24797,N_24783);
nand UO_1095 (O_1095,N_24592,N_24758);
or UO_1096 (O_1096,N_24960,N_24900);
xnor UO_1097 (O_1097,N_24553,N_24804);
and UO_1098 (O_1098,N_24833,N_24884);
and UO_1099 (O_1099,N_24733,N_24602);
nor UO_1100 (O_1100,N_24740,N_24885);
nor UO_1101 (O_1101,N_24730,N_24656);
xnor UO_1102 (O_1102,N_24680,N_24779);
or UO_1103 (O_1103,N_24511,N_24736);
nor UO_1104 (O_1104,N_24718,N_24987);
or UO_1105 (O_1105,N_24643,N_24959);
xor UO_1106 (O_1106,N_24539,N_24697);
or UO_1107 (O_1107,N_24888,N_24975);
and UO_1108 (O_1108,N_24984,N_24742);
nor UO_1109 (O_1109,N_24799,N_24965);
xor UO_1110 (O_1110,N_24783,N_24917);
and UO_1111 (O_1111,N_24753,N_24724);
nor UO_1112 (O_1112,N_24777,N_24672);
or UO_1113 (O_1113,N_24967,N_24534);
xnor UO_1114 (O_1114,N_24688,N_24672);
and UO_1115 (O_1115,N_24924,N_24529);
nor UO_1116 (O_1116,N_24641,N_24564);
and UO_1117 (O_1117,N_24942,N_24859);
and UO_1118 (O_1118,N_24708,N_24882);
xor UO_1119 (O_1119,N_24734,N_24738);
nand UO_1120 (O_1120,N_24558,N_24623);
and UO_1121 (O_1121,N_24795,N_24578);
or UO_1122 (O_1122,N_24852,N_24712);
or UO_1123 (O_1123,N_24709,N_24514);
nand UO_1124 (O_1124,N_24954,N_24754);
nor UO_1125 (O_1125,N_24532,N_24658);
nor UO_1126 (O_1126,N_24946,N_24629);
xnor UO_1127 (O_1127,N_24587,N_24641);
nor UO_1128 (O_1128,N_24738,N_24654);
xor UO_1129 (O_1129,N_24822,N_24600);
xor UO_1130 (O_1130,N_24794,N_24757);
nor UO_1131 (O_1131,N_24862,N_24576);
or UO_1132 (O_1132,N_24872,N_24652);
nor UO_1133 (O_1133,N_24930,N_24625);
or UO_1134 (O_1134,N_24583,N_24602);
xor UO_1135 (O_1135,N_24669,N_24960);
nand UO_1136 (O_1136,N_24790,N_24624);
xor UO_1137 (O_1137,N_24639,N_24723);
nand UO_1138 (O_1138,N_24550,N_24503);
xor UO_1139 (O_1139,N_24938,N_24652);
or UO_1140 (O_1140,N_24720,N_24579);
nor UO_1141 (O_1141,N_24757,N_24616);
nand UO_1142 (O_1142,N_24761,N_24897);
or UO_1143 (O_1143,N_24907,N_24790);
and UO_1144 (O_1144,N_24572,N_24921);
and UO_1145 (O_1145,N_24522,N_24911);
nor UO_1146 (O_1146,N_24664,N_24744);
or UO_1147 (O_1147,N_24692,N_24979);
nor UO_1148 (O_1148,N_24784,N_24885);
or UO_1149 (O_1149,N_24969,N_24946);
or UO_1150 (O_1150,N_24910,N_24547);
nor UO_1151 (O_1151,N_24983,N_24512);
nor UO_1152 (O_1152,N_24676,N_24623);
and UO_1153 (O_1153,N_24623,N_24951);
nor UO_1154 (O_1154,N_24655,N_24877);
xnor UO_1155 (O_1155,N_24836,N_24683);
nor UO_1156 (O_1156,N_24831,N_24643);
or UO_1157 (O_1157,N_24761,N_24781);
xor UO_1158 (O_1158,N_24704,N_24695);
and UO_1159 (O_1159,N_24824,N_24693);
nor UO_1160 (O_1160,N_24558,N_24815);
nor UO_1161 (O_1161,N_24955,N_24535);
nand UO_1162 (O_1162,N_24909,N_24968);
or UO_1163 (O_1163,N_24703,N_24718);
and UO_1164 (O_1164,N_24683,N_24753);
nand UO_1165 (O_1165,N_24632,N_24707);
and UO_1166 (O_1166,N_24948,N_24570);
or UO_1167 (O_1167,N_24533,N_24764);
or UO_1168 (O_1168,N_24673,N_24745);
nor UO_1169 (O_1169,N_24922,N_24695);
nor UO_1170 (O_1170,N_24516,N_24852);
nand UO_1171 (O_1171,N_24912,N_24630);
or UO_1172 (O_1172,N_24511,N_24870);
nor UO_1173 (O_1173,N_24733,N_24885);
nor UO_1174 (O_1174,N_24847,N_24526);
nor UO_1175 (O_1175,N_24846,N_24524);
nor UO_1176 (O_1176,N_24933,N_24633);
xor UO_1177 (O_1177,N_24953,N_24777);
nand UO_1178 (O_1178,N_24553,N_24904);
nor UO_1179 (O_1179,N_24581,N_24840);
or UO_1180 (O_1180,N_24661,N_24761);
nand UO_1181 (O_1181,N_24591,N_24557);
nand UO_1182 (O_1182,N_24949,N_24688);
xnor UO_1183 (O_1183,N_24513,N_24647);
and UO_1184 (O_1184,N_24781,N_24610);
and UO_1185 (O_1185,N_24753,N_24857);
nand UO_1186 (O_1186,N_24977,N_24575);
or UO_1187 (O_1187,N_24672,N_24547);
and UO_1188 (O_1188,N_24579,N_24659);
nand UO_1189 (O_1189,N_24895,N_24567);
or UO_1190 (O_1190,N_24597,N_24904);
nand UO_1191 (O_1191,N_24928,N_24859);
nand UO_1192 (O_1192,N_24513,N_24509);
and UO_1193 (O_1193,N_24505,N_24679);
nor UO_1194 (O_1194,N_24790,N_24992);
and UO_1195 (O_1195,N_24580,N_24829);
xor UO_1196 (O_1196,N_24585,N_24576);
or UO_1197 (O_1197,N_24860,N_24961);
or UO_1198 (O_1198,N_24974,N_24891);
and UO_1199 (O_1199,N_24545,N_24821);
or UO_1200 (O_1200,N_24569,N_24806);
or UO_1201 (O_1201,N_24693,N_24748);
nor UO_1202 (O_1202,N_24987,N_24554);
and UO_1203 (O_1203,N_24629,N_24546);
and UO_1204 (O_1204,N_24721,N_24665);
nand UO_1205 (O_1205,N_24788,N_24849);
xor UO_1206 (O_1206,N_24754,N_24677);
or UO_1207 (O_1207,N_24769,N_24701);
and UO_1208 (O_1208,N_24720,N_24980);
nor UO_1209 (O_1209,N_24660,N_24629);
xnor UO_1210 (O_1210,N_24622,N_24512);
and UO_1211 (O_1211,N_24849,N_24892);
or UO_1212 (O_1212,N_24915,N_24782);
nand UO_1213 (O_1213,N_24781,N_24798);
or UO_1214 (O_1214,N_24864,N_24530);
nand UO_1215 (O_1215,N_24959,N_24566);
xor UO_1216 (O_1216,N_24846,N_24905);
and UO_1217 (O_1217,N_24801,N_24504);
xnor UO_1218 (O_1218,N_24579,N_24969);
nand UO_1219 (O_1219,N_24589,N_24587);
or UO_1220 (O_1220,N_24885,N_24896);
nor UO_1221 (O_1221,N_24903,N_24861);
nand UO_1222 (O_1222,N_24560,N_24800);
nand UO_1223 (O_1223,N_24762,N_24751);
nand UO_1224 (O_1224,N_24797,N_24821);
or UO_1225 (O_1225,N_24849,N_24779);
nor UO_1226 (O_1226,N_24994,N_24835);
or UO_1227 (O_1227,N_24600,N_24768);
xnor UO_1228 (O_1228,N_24678,N_24581);
xnor UO_1229 (O_1229,N_24886,N_24759);
or UO_1230 (O_1230,N_24723,N_24835);
nor UO_1231 (O_1231,N_24910,N_24716);
nor UO_1232 (O_1232,N_24825,N_24594);
nand UO_1233 (O_1233,N_24690,N_24619);
nor UO_1234 (O_1234,N_24592,N_24681);
xor UO_1235 (O_1235,N_24590,N_24859);
xnor UO_1236 (O_1236,N_24916,N_24640);
and UO_1237 (O_1237,N_24599,N_24508);
xnor UO_1238 (O_1238,N_24895,N_24630);
nor UO_1239 (O_1239,N_24685,N_24803);
and UO_1240 (O_1240,N_24572,N_24782);
and UO_1241 (O_1241,N_24521,N_24953);
nand UO_1242 (O_1242,N_24617,N_24683);
xor UO_1243 (O_1243,N_24850,N_24594);
nand UO_1244 (O_1244,N_24805,N_24916);
xnor UO_1245 (O_1245,N_24599,N_24576);
xor UO_1246 (O_1246,N_24667,N_24713);
and UO_1247 (O_1247,N_24563,N_24712);
or UO_1248 (O_1248,N_24571,N_24850);
xor UO_1249 (O_1249,N_24756,N_24833);
nand UO_1250 (O_1250,N_24725,N_24750);
nand UO_1251 (O_1251,N_24733,N_24925);
nand UO_1252 (O_1252,N_24777,N_24915);
xor UO_1253 (O_1253,N_24937,N_24853);
nor UO_1254 (O_1254,N_24564,N_24921);
and UO_1255 (O_1255,N_24739,N_24628);
nor UO_1256 (O_1256,N_24513,N_24827);
or UO_1257 (O_1257,N_24619,N_24647);
and UO_1258 (O_1258,N_24845,N_24919);
nor UO_1259 (O_1259,N_24730,N_24549);
or UO_1260 (O_1260,N_24661,N_24941);
nand UO_1261 (O_1261,N_24929,N_24880);
or UO_1262 (O_1262,N_24963,N_24626);
and UO_1263 (O_1263,N_24881,N_24939);
nor UO_1264 (O_1264,N_24949,N_24805);
or UO_1265 (O_1265,N_24914,N_24644);
and UO_1266 (O_1266,N_24556,N_24785);
and UO_1267 (O_1267,N_24671,N_24779);
nor UO_1268 (O_1268,N_24914,N_24854);
and UO_1269 (O_1269,N_24566,N_24889);
or UO_1270 (O_1270,N_24717,N_24598);
or UO_1271 (O_1271,N_24636,N_24662);
or UO_1272 (O_1272,N_24631,N_24954);
nor UO_1273 (O_1273,N_24694,N_24773);
or UO_1274 (O_1274,N_24960,N_24617);
or UO_1275 (O_1275,N_24606,N_24720);
xnor UO_1276 (O_1276,N_24510,N_24515);
and UO_1277 (O_1277,N_24537,N_24527);
or UO_1278 (O_1278,N_24655,N_24661);
xor UO_1279 (O_1279,N_24657,N_24503);
and UO_1280 (O_1280,N_24550,N_24938);
nand UO_1281 (O_1281,N_24703,N_24881);
and UO_1282 (O_1282,N_24524,N_24607);
xor UO_1283 (O_1283,N_24631,N_24845);
nand UO_1284 (O_1284,N_24744,N_24887);
xnor UO_1285 (O_1285,N_24618,N_24675);
or UO_1286 (O_1286,N_24800,N_24694);
and UO_1287 (O_1287,N_24726,N_24519);
and UO_1288 (O_1288,N_24630,N_24948);
nand UO_1289 (O_1289,N_24891,N_24836);
nor UO_1290 (O_1290,N_24807,N_24942);
xnor UO_1291 (O_1291,N_24967,N_24975);
or UO_1292 (O_1292,N_24941,N_24776);
xor UO_1293 (O_1293,N_24958,N_24837);
nor UO_1294 (O_1294,N_24893,N_24814);
and UO_1295 (O_1295,N_24718,N_24985);
and UO_1296 (O_1296,N_24536,N_24856);
nand UO_1297 (O_1297,N_24846,N_24769);
xor UO_1298 (O_1298,N_24547,N_24572);
nor UO_1299 (O_1299,N_24808,N_24684);
xnor UO_1300 (O_1300,N_24512,N_24828);
nor UO_1301 (O_1301,N_24576,N_24719);
nand UO_1302 (O_1302,N_24591,N_24797);
or UO_1303 (O_1303,N_24899,N_24712);
nor UO_1304 (O_1304,N_24813,N_24652);
and UO_1305 (O_1305,N_24769,N_24955);
xnor UO_1306 (O_1306,N_24546,N_24967);
nor UO_1307 (O_1307,N_24553,N_24893);
xor UO_1308 (O_1308,N_24765,N_24503);
nor UO_1309 (O_1309,N_24581,N_24969);
nand UO_1310 (O_1310,N_24979,N_24899);
xor UO_1311 (O_1311,N_24589,N_24772);
and UO_1312 (O_1312,N_24606,N_24745);
and UO_1313 (O_1313,N_24981,N_24500);
nor UO_1314 (O_1314,N_24842,N_24776);
xor UO_1315 (O_1315,N_24555,N_24545);
xnor UO_1316 (O_1316,N_24753,N_24672);
and UO_1317 (O_1317,N_24855,N_24943);
and UO_1318 (O_1318,N_24509,N_24706);
or UO_1319 (O_1319,N_24739,N_24904);
nor UO_1320 (O_1320,N_24838,N_24934);
nand UO_1321 (O_1321,N_24587,N_24762);
and UO_1322 (O_1322,N_24862,N_24651);
xor UO_1323 (O_1323,N_24513,N_24743);
or UO_1324 (O_1324,N_24708,N_24530);
nand UO_1325 (O_1325,N_24924,N_24534);
and UO_1326 (O_1326,N_24817,N_24683);
or UO_1327 (O_1327,N_24711,N_24801);
or UO_1328 (O_1328,N_24994,N_24559);
nor UO_1329 (O_1329,N_24934,N_24695);
and UO_1330 (O_1330,N_24608,N_24650);
nor UO_1331 (O_1331,N_24771,N_24738);
and UO_1332 (O_1332,N_24838,N_24673);
or UO_1333 (O_1333,N_24535,N_24951);
and UO_1334 (O_1334,N_24566,N_24664);
or UO_1335 (O_1335,N_24844,N_24737);
or UO_1336 (O_1336,N_24708,N_24949);
nor UO_1337 (O_1337,N_24602,N_24991);
and UO_1338 (O_1338,N_24760,N_24903);
xor UO_1339 (O_1339,N_24936,N_24528);
and UO_1340 (O_1340,N_24684,N_24590);
xnor UO_1341 (O_1341,N_24544,N_24564);
xor UO_1342 (O_1342,N_24804,N_24890);
nor UO_1343 (O_1343,N_24530,N_24766);
nand UO_1344 (O_1344,N_24650,N_24970);
nand UO_1345 (O_1345,N_24721,N_24965);
xnor UO_1346 (O_1346,N_24753,N_24784);
and UO_1347 (O_1347,N_24625,N_24677);
xor UO_1348 (O_1348,N_24597,N_24635);
xnor UO_1349 (O_1349,N_24505,N_24502);
nand UO_1350 (O_1350,N_24941,N_24614);
nand UO_1351 (O_1351,N_24993,N_24544);
nor UO_1352 (O_1352,N_24538,N_24790);
nand UO_1353 (O_1353,N_24626,N_24988);
nand UO_1354 (O_1354,N_24583,N_24650);
and UO_1355 (O_1355,N_24540,N_24763);
nand UO_1356 (O_1356,N_24543,N_24701);
nand UO_1357 (O_1357,N_24992,N_24564);
xor UO_1358 (O_1358,N_24706,N_24818);
and UO_1359 (O_1359,N_24895,N_24638);
nand UO_1360 (O_1360,N_24659,N_24505);
or UO_1361 (O_1361,N_24576,N_24727);
and UO_1362 (O_1362,N_24644,N_24944);
and UO_1363 (O_1363,N_24711,N_24527);
and UO_1364 (O_1364,N_24533,N_24843);
nor UO_1365 (O_1365,N_24689,N_24613);
nor UO_1366 (O_1366,N_24946,N_24593);
nor UO_1367 (O_1367,N_24585,N_24852);
nand UO_1368 (O_1368,N_24629,N_24694);
nand UO_1369 (O_1369,N_24500,N_24732);
nand UO_1370 (O_1370,N_24751,N_24536);
or UO_1371 (O_1371,N_24876,N_24873);
nor UO_1372 (O_1372,N_24762,N_24545);
nor UO_1373 (O_1373,N_24796,N_24505);
nor UO_1374 (O_1374,N_24891,N_24952);
nor UO_1375 (O_1375,N_24961,N_24791);
nand UO_1376 (O_1376,N_24799,N_24649);
nor UO_1377 (O_1377,N_24872,N_24886);
and UO_1378 (O_1378,N_24987,N_24519);
or UO_1379 (O_1379,N_24869,N_24758);
nor UO_1380 (O_1380,N_24558,N_24691);
nor UO_1381 (O_1381,N_24556,N_24681);
or UO_1382 (O_1382,N_24712,N_24788);
and UO_1383 (O_1383,N_24622,N_24728);
or UO_1384 (O_1384,N_24915,N_24945);
xnor UO_1385 (O_1385,N_24868,N_24788);
nand UO_1386 (O_1386,N_24946,N_24534);
xor UO_1387 (O_1387,N_24852,N_24865);
and UO_1388 (O_1388,N_24562,N_24580);
or UO_1389 (O_1389,N_24933,N_24852);
and UO_1390 (O_1390,N_24807,N_24928);
or UO_1391 (O_1391,N_24969,N_24641);
xnor UO_1392 (O_1392,N_24887,N_24563);
or UO_1393 (O_1393,N_24648,N_24615);
nand UO_1394 (O_1394,N_24574,N_24895);
nor UO_1395 (O_1395,N_24670,N_24924);
and UO_1396 (O_1396,N_24559,N_24553);
or UO_1397 (O_1397,N_24880,N_24702);
and UO_1398 (O_1398,N_24901,N_24793);
nand UO_1399 (O_1399,N_24752,N_24792);
and UO_1400 (O_1400,N_24811,N_24601);
xnor UO_1401 (O_1401,N_24836,N_24564);
nor UO_1402 (O_1402,N_24852,N_24558);
and UO_1403 (O_1403,N_24565,N_24569);
nand UO_1404 (O_1404,N_24804,N_24563);
xor UO_1405 (O_1405,N_24692,N_24959);
and UO_1406 (O_1406,N_24770,N_24628);
nand UO_1407 (O_1407,N_24754,N_24988);
nand UO_1408 (O_1408,N_24861,N_24598);
or UO_1409 (O_1409,N_24683,N_24646);
nand UO_1410 (O_1410,N_24820,N_24512);
xnor UO_1411 (O_1411,N_24877,N_24819);
or UO_1412 (O_1412,N_24873,N_24639);
and UO_1413 (O_1413,N_24799,N_24554);
or UO_1414 (O_1414,N_24982,N_24855);
nor UO_1415 (O_1415,N_24933,N_24792);
nor UO_1416 (O_1416,N_24982,N_24767);
nand UO_1417 (O_1417,N_24795,N_24770);
nand UO_1418 (O_1418,N_24920,N_24660);
nand UO_1419 (O_1419,N_24862,N_24925);
nand UO_1420 (O_1420,N_24752,N_24732);
xnor UO_1421 (O_1421,N_24512,N_24515);
and UO_1422 (O_1422,N_24726,N_24615);
nand UO_1423 (O_1423,N_24827,N_24992);
nor UO_1424 (O_1424,N_24558,N_24567);
nand UO_1425 (O_1425,N_24827,N_24836);
nor UO_1426 (O_1426,N_24962,N_24720);
nand UO_1427 (O_1427,N_24680,N_24605);
and UO_1428 (O_1428,N_24618,N_24918);
nor UO_1429 (O_1429,N_24993,N_24788);
and UO_1430 (O_1430,N_24818,N_24520);
nor UO_1431 (O_1431,N_24515,N_24672);
xnor UO_1432 (O_1432,N_24907,N_24824);
nor UO_1433 (O_1433,N_24861,N_24570);
xnor UO_1434 (O_1434,N_24873,N_24782);
and UO_1435 (O_1435,N_24892,N_24506);
xor UO_1436 (O_1436,N_24634,N_24737);
and UO_1437 (O_1437,N_24698,N_24661);
or UO_1438 (O_1438,N_24614,N_24539);
nand UO_1439 (O_1439,N_24892,N_24925);
nand UO_1440 (O_1440,N_24739,N_24750);
nor UO_1441 (O_1441,N_24670,N_24795);
or UO_1442 (O_1442,N_24913,N_24623);
or UO_1443 (O_1443,N_24864,N_24599);
nor UO_1444 (O_1444,N_24783,N_24516);
and UO_1445 (O_1445,N_24605,N_24800);
xor UO_1446 (O_1446,N_24572,N_24674);
nor UO_1447 (O_1447,N_24701,N_24745);
and UO_1448 (O_1448,N_24565,N_24945);
xor UO_1449 (O_1449,N_24925,N_24908);
or UO_1450 (O_1450,N_24994,N_24590);
xnor UO_1451 (O_1451,N_24805,N_24986);
or UO_1452 (O_1452,N_24847,N_24666);
and UO_1453 (O_1453,N_24646,N_24714);
nor UO_1454 (O_1454,N_24600,N_24514);
xnor UO_1455 (O_1455,N_24609,N_24906);
nor UO_1456 (O_1456,N_24758,N_24580);
nand UO_1457 (O_1457,N_24610,N_24757);
nand UO_1458 (O_1458,N_24724,N_24686);
nand UO_1459 (O_1459,N_24792,N_24501);
and UO_1460 (O_1460,N_24949,N_24653);
or UO_1461 (O_1461,N_24826,N_24771);
and UO_1462 (O_1462,N_24904,N_24671);
or UO_1463 (O_1463,N_24513,N_24771);
and UO_1464 (O_1464,N_24957,N_24804);
nor UO_1465 (O_1465,N_24649,N_24591);
xnor UO_1466 (O_1466,N_24649,N_24835);
or UO_1467 (O_1467,N_24572,N_24621);
or UO_1468 (O_1468,N_24860,N_24681);
nand UO_1469 (O_1469,N_24858,N_24701);
nor UO_1470 (O_1470,N_24714,N_24835);
xor UO_1471 (O_1471,N_24893,N_24757);
nand UO_1472 (O_1472,N_24685,N_24678);
xnor UO_1473 (O_1473,N_24581,N_24532);
nand UO_1474 (O_1474,N_24681,N_24501);
or UO_1475 (O_1475,N_24968,N_24775);
nor UO_1476 (O_1476,N_24506,N_24876);
xnor UO_1477 (O_1477,N_24939,N_24658);
xnor UO_1478 (O_1478,N_24693,N_24661);
and UO_1479 (O_1479,N_24500,N_24715);
xnor UO_1480 (O_1480,N_24884,N_24616);
nor UO_1481 (O_1481,N_24918,N_24656);
and UO_1482 (O_1482,N_24826,N_24769);
or UO_1483 (O_1483,N_24579,N_24820);
nor UO_1484 (O_1484,N_24888,N_24607);
or UO_1485 (O_1485,N_24658,N_24545);
xor UO_1486 (O_1486,N_24813,N_24669);
xor UO_1487 (O_1487,N_24839,N_24581);
nor UO_1488 (O_1488,N_24513,N_24918);
xor UO_1489 (O_1489,N_24976,N_24507);
and UO_1490 (O_1490,N_24550,N_24728);
nand UO_1491 (O_1491,N_24747,N_24581);
and UO_1492 (O_1492,N_24993,N_24936);
nor UO_1493 (O_1493,N_24832,N_24628);
or UO_1494 (O_1494,N_24980,N_24638);
nor UO_1495 (O_1495,N_24908,N_24760);
xor UO_1496 (O_1496,N_24744,N_24999);
nor UO_1497 (O_1497,N_24864,N_24619);
nor UO_1498 (O_1498,N_24621,N_24885);
or UO_1499 (O_1499,N_24870,N_24530);
or UO_1500 (O_1500,N_24612,N_24765);
or UO_1501 (O_1501,N_24515,N_24842);
or UO_1502 (O_1502,N_24607,N_24798);
and UO_1503 (O_1503,N_24630,N_24564);
nor UO_1504 (O_1504,N_24962,N_24516);
or UO_1505 (O_1505,N_24749,N_24583);
nand UO_1506 (O_1506,N_24596,N_24917);
and UO_1507 (O_1507,N_24788,N_24960);
nand UO_1508 (O_1508,N_24964,N_24736);
xor UO_1509 (O_1509,N_24665,N_24834);
xnor UO_1510 (O_1510,N_24685,N_24998);
nand UO_1511 (O_1511,N_24719,N_24615);
xnor UO_1512 (O_1512,N_24602,N_24639);
nand UO_1513 (O_1513,N_24961,N_24506);
and UO_1514 (O_1514,N_24727,N_24567);
xnor UO_1515 (O_1515,N_24542,N_24592);
nand UO_1516 (O_1516,N_24594,N_24773);
nor UO_1517 (O_1517,N_24929,N_24732);
and UO_1518 (O_1518,N_24666,N_24853);
or UO_1519 (O_1519,N_24792,N_24871);
or UO_1520 (O_1520,N_24875,N_24716);
xor UO_1521 (O_1521,N_24685,N_24647);
nor UO_1522 (O_1522,N_24690,N_24509);
nor UO_1523 (O_1523,N_24564,N_24904);
or UO_1524 (O_1524,N_24587,N_24704);
and UO_1525 (O_1525,N_24567,N_24930);
or UO_1526 (O_1526,N_24681,N_24576);
xnor UO_1527 (O_1527,N_24523,N_24804);
xnor UO_1528 (O_1528,N_24573,N_24931);
and UO_1529 (O_1529,N_24740,N_24823);
nor UO_1530 (O_1530,N_24564,N_24975);
or UO_1531 (O_1531,N_24574,N_24750);
xnor UO_1532 (O_1532,N_24676,N_24989);
xor UO_1533 (O_1533,N_24926,N_24541);
xor UO_1534 (O_1534,N_24980,N_24557);
nor UO_1535 (O_1535,N_24650,N_24868);
or UO_1536 (O_1536,N_24630,N_24781);
nand UO_1537 (O_1537,N_24758,N_24926);
or UO_1538 (O_1538,N_24695,N_24778);
nand UO_1539 (O_1539,N_24531,N_24575);
nor UO_1540 (O_1540,N_24924,N_24548);
and UO_1541 (O_1541,N_24897,N_24950);
or UO_1542 (O_1542,N_24668,N_24858);
or UO_1543 (O_1543,N_24887,N_24791);
xor UO_1544 (O_1544,N_24916,N_24821);
nand UO_1545 (O_1545,N_24923,N_24979);
nor UO_1546 (O_1546,N_24736,N_24846);
xnor UO_1547 (O_1547,N_24815,N_24664);
nor UO_1548 (O_1548,N_24867,N_24816);
nor UO_1549 (O_1549,N_24568,N_24736);
nand UO_1550 (O_1550,N_24873,N_24878);
xnor UO_1551 (O_1551,N_24748,N_24612);
nand UO_1552 (O_1552,N_24952,N_24574);
nor UO_1553 (O_1553,N_24691,N_24651);
or UO_1554 (O_1554,N_24661,N_24783);
nand UO_1555 (O_1555,N_24613,N_24522);
nand UO_1556 (O_1556,N_24890,N_24556);
nor UO_1557 (O_1557,N_24913,N_24580);
nor UO_1558 (O_1558,N_24716,N_24771);
xor UO_1559 (O_1559,N_24518,N_24567);
and UO_1560 (O_1560,N_24794,N_24687);
nand UO_1561 (O_1561,N_24973,N_24767);
nand UO_1562 (O_1562,N_24876,N_24982);
nor UO_1563 (O_1563,N_24981,N_24792);
nor UO_1564 (O_1564,N_24926,N_24525);
and UO_1565 (O_1565,N_24521,N_24894);
and UO_1566 (O_1566,N_24593,N_24912);
nand UO_1567 (O_1567,N_24580,N_24864);
nor UO_1568 (O_1568,N_24989,N_24628);
xor UO_1569 (O_1569,N_24755,N_24612);
nand UO_1570 (O_1570,N_24759,N_24875);
and UO_1571 (O_1571,N_24665,N_24767);
xnor UO_1572 (O_1572,N_24982,N_24596);
nor UO_1573 (O_1573,N_24734,N_24978);
nor UO_1574 (O_1574,N_24936,N_24879);
and UO_1575 (O_1575,N_24970,N_24873);
nor UO_1576 (O_1576,N_24950,N_24871);
or UO_1577 (O_1577,N_24814,N_24886);
nand UO_1578 (O_1578,N_24998,N_24785);
or UO_1579 (O_1579,N_24746,N_24607);
or UO_1580 (O_1580,N_24975,N_24966);
xor UO_1581 (O_1581,N_24532,N_24627);
xor UO_1582 (O_1582,N_24647,N_24867);
nand UO_1583 (O_1583,N_24528,N_24717);
nand UO_1584 (O_1584,N_24934,N_24668);
nor UO_1585 (O_1585,N_24870,N_24599);
and UO_1586 (O_1586,N_24579,N_24630);
nand UO_1587 (O_1587,N_24997,N_24692);
or UO_1588 (O_1588,N_24900,N_24659);
nand UO_1589 (O_1589,N_24792,N_24632);
nand UO_1590 (O_1590,N_24747,N_24702);
nand UO_1591 (O_1591,N_24958,N_24839);
xnor UO_1592 (O_1592,N_24564,N_24765);
nor UO_1593 (O_1593,N_24719,N_24980);
xnor UO_1594 (O_1594,N_24523,N_24623);
nor UO_1595 (O_1595,N_24759,N_24993);
or UO_1596 (O_1596,N_24654,N_24547);
or UO_1597 (O_1597,N_24506,N_24538);
nand UO_1598 (O_1598,N_24554,N_24773);
nor UO_1599 (O_1599,N_24715,N_24708);
and UO_1600 (O_1600,N_24503,N_24999);
xnor UO_1601 (O_1601,N_24564,N_24539);
nor UO_1602 (O_1602,N_24721,N_24806);
or UO_1603 (O_1603,N_24587,N_24545);
nor UO_1604 (O_1604,N_24895,N_24614);
xnor UO_1605 (O_1605,N_24937,N_24776);
nand UO_1606 (O_1606,N_24984,N_24798);
nor UO_1607 (O_1607,N_24942,N_24730);
or UO_1608 (O_1608,N_24782,N_24837);
nand UO_1609 (O_1609,N_24995,N_24965);
xnor UO_1610 (O_1610,N_24569,N_24560);
or UO_1611 (O_1611,N_24808,N_24945);
or UO_1612 (O_1612,N_24738,N_24636);
xnor UO_1613 (O_1613,N_24647,N_24886);
and UO_1614 (O_1614,N_24924,N_24682);
xor UO_1615 (O_1615,N_24792,N_24885);
nor UO_1616 (O_1616,N_24589,N_24707);
or UO_1617 (O_1617,N_24754,N_24678);
and UO_1618 (O_1618,N_24778,N_24976);
xor UO_1619 (O_1619,N_24993,N_24665);
nand UO_1620 (O_1620,N_24953,N_24918);
and UO_1621 (O_1621,N_24940,N_24661);
xor UO_1622 (O_1622,N_24635,N_24718);
nor UO_1623 (O_1623,N_24943,N_24918);
nand UO_1624 (O_1624,N_24906,N_24602);
nand UO_1625 (O_1625,N_24538,N_24971);
xor UO_1626 (O_1626,N_24791,N_24717);
or UO_1627 (O_1627,N_24739,N_24619);
and UO_1628 (O_1628,N_24713,N_24903);
and UO_1629 (O_1629,N_24931,N_24635);
nand UO_1630 (O_1630,N_24787,N_24824);
nor UO_1631 (O_1631,N_24621,N_24591);
nor UO_1632 (O_1632,N_24754,N_24653);
nor UO_1633 (O_1633,N_24786,N_24738);
nor UO_1634 (O_1634,N_24591,N_24685);
nand UO_1635 (O_1635,N_24556,N_24662);
and UO_1636 (O_1636,N_24635,N_24701);
xor UO_1637 (O_1637,N_24595,N_24778);
nand UO_1638 (O_1638,N_24589,N_24708);
nor UO_1639 (O_1639,N_24883,N_24891);
xor UO_1640 (O_1640,N_24961,N_24990);
nand UO_1641 (O_1641,N_24949,N_24576);
or UO_1642 (O_1642,N_24845,N_24675);
nor UO_1643 (O_1643,N_24699,N_24851);
or UO_1644 (O_1644,N_24843,N_24976);
nor UO_1645 (O_1645,N_24648,N_24966);
nor UO_1646 (O_1646,N_24946,N_24835);
and UO_1647 (O_1647,N_24606,N_24624);
and UO_1648 (O_1648,N_24764,N_24962);
nand UO_1649 (O_1649,N_24950,N_24863);
or UO_1650 (O_1650,N_24567,N_24755);
and UO_1651 (O_1651,N_24789,N_24829);
nor UO_1652 (O_1652,N_24687,N_24507);
and UO_1653 (O_1653,N_24765,N_24956);
nand UO_1654 (O_1654,N_24728,N_24723);
nor UO_1655 (O_1655,N_24632,N_24559);
nand UO_1656 (O_1656,N_24571,N_24888);
nand UO_1657 (O_1657,N_24675,N_24697);
and UO_1658 (O_1658,N_24681,N_24854);
xnor UO_1659 (O_1659,N_24694,N_24670);
or UO_1660 (O_1660,N_24782,N_24590);
or UO_1661 (O_1661,N_24927,N_24585);
nor UO_1662 (O_1662,N_24671,N_24880);
nand UO_1663 (O_1663,N_24812,N_24676);
xor UO_1664 (O_1664,N_24616,N_24668);
nand UO_1665 (O_1665,N_24503,N_24512);
and UO_1666 (O_1666,N_24806,N_24581);
nor UO_1667 (O_1667,N_24792,N_24565);
nand UO_1668 (O_1668,N_24913,N_24800);
and UO_1669 (O_1669,N_24963,N_24820);
xnor UO_1670 (O_1670,N_24613,N_24923);
nor UO_1671 (O_1671,N_24608,N_24975);
nand UO_1672 (O_1672,N_24873,N_24932);
or UO_1673 (O_1673,N_24852,N_24894);
and UO_1674 (O_1674,N_24549,N_24695);
or UO_1675 (O_1675,N_24621,N_24556);
or UO_1676 (O_1676,N_24960,N_24582);
and UO_1677 (O_1677,N_24814,N_24601);
xor UO_1678 (O_1678,N_24614,N_24813);
and UO_1679 (O_1679,N_24520,N_24876);
and UO_1680 (O_1680,N_24946,N_24941);
and UO_1681 (O_1681,N_24633,N_24613);
nand UO_1682 (O_1682,N_24694,N_24833);
and UO_1683 (O_1683,N_24769,N_24524);
and UO_1684 (O_1684,N_24672,N_24650);
and UO_1685 (O_1685,N_24737,N_24572);
xor UO_1686 (O_1686,N_24812,N_24649);
nand UO_1687 (O_1687,N_24590,N_24748);
xor UO_1688 (O_1688,N_24526,N_24714);
nand UO_1689 (O_1689,N_24932,N_24975);
nor UO_1690 (O_1690,N_24918,N_24675);
and UO_1691 (O_1691,N_24674,N_24747);
nor UO_1692 (O_1692,N_24805,N_24969);
and UO_1693 (O_1693,N_24887,N_24762);
or UO_1694 (O_1694,N_24759,N_24867);
or UO_1695 (O_1695,N_24869,N_24538);
xnor UO_1696 (O_1696,N_24677,N_24610);
xnor UO_1697 (O_1697,N_24938,N_24619);
or UO_1698 (O_1698,N_24590,N_24733);
nor UO_1699 (O_1699,N_24826,N_24978);
and UO_1700 (O_1700,N_24813,N_24615);
xor UO_1701 (O_1701,N_24604,N_24762);
xnor UO_1702 (O_1702,N_24800,N_24813);
xor UO_1703 (O_1703,N_24504,N_24989);
nand UO_1704 (O_1704,N_24793,N_24817);
xnor UO_1705 (O_1705,N_24916,N_24839);
xor UO_1706 (O_1706,N_24596,N_24788);
nor UO_1707 (O_1707,N_24557,N_24630);
or UO_1708 (O_1708,N_24914,N_24772);
xor UO_1709 (O_1709,N_24668,N_24716);
nor UO_1710 (O_1710,N_24829,N_24910);
xnor UO_1711 (O_1711,N_24665,N_24775);
and UO_1712 (O_1712,N_24912,N_24744);
and UO_1713 (O_1713,N_24575,N_24948);
or UO_1714 (O_1714,N_24707,N_24560);
nor UO_1715 (O_1715,N_24767,N_24573);
or UO_1716 (O_1716,N_24573,N_24577);
nand UO_1717 (O_1717,N_24613,N_24752);
nand UO_1718 (O_1718,N_24599,N_24951);
nand UO_1719 (O_1719,N_24904,N_24670);
or UO_1720 (O_1720,N_24673,N_24549);
nand UO_1721 (O_1721,N_24579,N_24777);
and UO_1722 (O_1722,N_24640,N_24813);
and UO_1723 (O_1723,N_24599,N_24862);
nor UO_1724 (O_1724,N_24596,N_24797);
nor UO_1725 (O_1725,N_24593,N_24704);
or UO_1726 (O_1726,N_24749,N_24797);
nand UO_1727 (O_1727,N_24902,N_24599);
and UO_1728 (O_1728,N_24959,N_24949);
xnor UO_1729 (O_1729,N_24545,N_24519);
and UO_1730 (O_1730,N_24564,N_24617);
xor UO_1731 (O_1731,N_24962,N_24722);
and UO_1732 (O_1732,N_24550,N_24901);
xnor UO_1733 (O_1733,N_24813,N_24983);
and UO_1734 (O_1734,N_24825,N_24732);
and UO_1735 (O_1735,N_24613,N_24548);
xnor UO_1736 (O_1736,N_24529,N_24710);
nand UO_1737 (O_1737,N_24559,N_24500);
and UO_1738 (O_1738,N_24676,N_24959);
or UO_1739 (O_1739,N_24556,N_24901);
and UO_1740 (O_1740,N_24510,N_24590);
nor UO_1741 (O_1741,N_24748,N_24980);
or UO_1742 (O_1742,N_24696,N_24576);
and UO_1743 (O_1743,N_24652,N_24633);
nand UO_1744 (O_1744,N_24957,N_24634);
xnor UO_1745 (O_1745,N_24803,N_24907);
xor UO_1746 (O_1746,N_24914,N_24719);
nand UO_1747 (O_1747,N_24726,N_24545);
nand UO_1748 (O_1748,N_24851,N_24756);
and UO_1749 (O_1749,N_24601,N_24535);
and UO_1750 (O_1750,N_24855,N_24865);
and UO_1751 (O_1751,N_24899,N_24743);
and UO_1752 (O_1752,N_24907,N_24584);
nor UO_1753 (O_1753,N_24532,N_24730);
and UO_1754 (O_1754,N_24520,N_24649);
or UO_1755 (O_1755,N_24935,N_24613);
nand UO_1756 (O_1756,N_24724,N_24872);
nor UO_1757 (O_1757,N_24753,N_24865);
xnor UO_1758 (O_1758,N_24846,N_24537);
or UO_1759 (O_1759,N_24577,N_24627);
nor UO_1760 (O_1760,N_24789,N_24767);
and UO_1761 (O_1761,N_24849,N_24873);
nor UO_1762 (O_1762,N_24534,N_24807);
xor UO_1763 (O_1763,N_24661,N_24580);
nor UO_1764 (O_1764,N_24703,N_24607);
xnor UO_1765 (O_1765,N_24779,N_24598);
nor UO_1766 (O_1766,N_24585,N_24554);
or UO_1767 (O_1767,N_24544,N_24696);
nand UO_1768 (O_1768,N_24765,N_24822);
and UO_1769 (O_1769,N_24880,N_24689);
xor UO_1770 (O_1770,N_24504,N_24532);
xnor UO_1771 (O_1771,N_24653,N_24950);
nor UO_1772 (O_1772,N_24860,N_24799);
and UO_1773 (O_1773,N_24698,N_24747);
nand UO_1774 (O_1774,N_24884,N_24755);
nand UO_1775 (O_1775,N_24967,N_24673);
nor UO_1776 (O_1776,N_24591,N_24897);
or UO_1777 (O_1777,N_24843,N_24935);
and UO_1778 (O_1778,N_24865,N_24680);
nor UO_1779 (O_1779,N_24993,N_24801);
nand UO_1780 (O_1780,N_24734,N_24919);
nand UO_1781 (O_1781,N_24931,N_24742);
and UO_1782 (O_1782,N_24524,N_24930);
or UO_1783 (O_1783,N_24904,N_24632);
nand UO_1784 (O_1784,N_24719,N_24676);
nand UO_1785 (O_1785,N_24721,N_24994);
xnor UO_1786 (O_1786,N_24827,N_24902);
or UO_1787 (O_1787,N_24958,N_24707);
and UO_1788 (O_1788,N_24979,N_24763);
and UO_1789 (O_1789,N_24547,N_24798);
xor UO_1790 (O_1790,N_24960,N_24501);
nand UO_1791 (O_1791,N_24735,N_24725);
nand UO_1792 (O_1792,N_24787,N_24904);
xor UO_1793 (O_1793,N_24834,N_24654);
or UO_1794 (O_1794,N_24859,N_24644);
nand UO_1795 (O_1795,N_24962,N_24818);
nor UO_1796 (O_1796,N_24544,N_24608);
nand UO_1797 (O_1797,N_24872,N_24973);
xnor UO_1798 (O_1798,N_24506,N_24964);
and UO_1799 (O_1799,N_24934,N_24667);
nor UO_1800 (O_1800,N_24846,N_24598);
xor UO_1801 (O_1801,N_24971,N_24556);
nor UO_1802 (O_1802,N_24591,N_24749);
and UO_1803 (O_1803,N_24600,N_24662);
or UO_1804 (O_1804,N_24671,N_24888);
and UO_1805 (O_1805,N_24647,N_24840);
nor UO_1806 (O_1806,N_24827,N_24996);
nand UO_1807 (O_1807,N_24583,N_24873);
and UO_1808 (O_1808,N_24850,N_24741);
and UO_1809 (O_1809,N_24611,N_24664);
or UO_1810 (O_1810,N_24672,N_24975);
nor UO_1811 (O_1811,N_24852,N_24916);
or UO_1812 (O_1812,N_24883,N_24672);
xnor UO_1813 (O_1813,N_24809,N_24738);
xnor UO_1814 (O_1814,N_24805,N_24605);
or UO_1815 (O_1815,N_24755,N_24846);
nor UO_1816 (O_1816,N_24647,N_24623);
nor UO_1817 (O_1817,N_24542,N_24887);
xnor UO_1818 (O_1818,N_24619,N_24688);
nand UO_1819 (O_1819,N_24920,N_24610);
and UO_1820 (O_1820,N_24677,N_24758);
xor UO_1821 (O_1821,N_24617,N_24975);
or UO_1822 (O_1822,N_24868,N_24816);
nor UO_1823 (O_1823,N_24728,N_24578);
and UO_1824 (O_1824,N_24977,N_24944);
or UO_1825 (O_1825,N_24855,N_24586);
nor UO_1826 (O_1826,N_24949,N_24538);
nand UO_1827 (O_1827,N_24787,N_24649);
xnor UO_1828 (O_1828,N_24996,N_24714);
and UO_1829 (O_1829,N_24621,N_24875);
nor UO_1830 (O_1830,N_24922,N_24953);
nor UO_1831 (O_1831,N_24968,N_24613);
xor UO_1832 (O_1832,N_24593,N_24922);
nor UO_1833 (O_1833,N_24782,N_24697);
nand UO_1834 (O_1834,N_24544,N_24868);
and UO_1835 (O_1835,N_24691,N_24628);
or UO_1836 (O_1836,N_24523,N_24948);
nand UO_1837 (O_1837,N_24994,N_24867);
nand UO_1838 (O_1838,N_24940,N_24789);
or UO_1839 (O_1839,N_24567,N_24671);
and UO_1840 (O_1840,N_24915,N_24983);
nor UO_1841 (O_1841,N_24527,N_24836);
and UO_1842 (O_1842,N_24795,N_24897);
or UO_1843 (O_1843,N_24552,N_24721);
and UO_1844 (O_1844,N_24697,N_24955);
and UO_1845 (O_1845,N_24976,N_24988);
nand UO_1846 (O_1846,N_24823,N_24597);
nor UO_1847 (O_1847,N_24903,N_24787);
nand UO_1848 (O_1848,N_24746,N_24588);
or UO_1849 (O_1849,N_24752,N_24779);
or UO_1850 (O_1850,N_24523,N_24760);
nand UO_1851 (O_1851,N_24501,N_24836);
nand UO_1852 (O_1852,N_24904,N_24825);
and UO_1853 (O_1853,N_24733,N_24796);
or UO_1854 (O_1854,N_24518,N_24591);
and UO_1855 (O_1855,N_24754,N_24860);
xnor UO_1856 (O_1856,N_24882,N_24617);
xor UO_1857 (O_1857,N_24931,N_24831);
xnor UO_1858 (O_1858,N_24963,N_24893);
nor UO_1859 (O_1859,N_24702,N_24795);
or UO_1860 (O_1860,N_24674,N_24958);
nand UO_1861 (O_1861,N_24906,N_24881);
and UO_1862 (O_1862,N_24707,N_24995);
nor UO_1863 (O_1863,N_24644,N_24934);
nor UO_1864 (O_1864,N_24868,N_24542);
and UO_1865 (O_1865,N_24963,N_24758);
xnor UO_1866 (O_1866,N_24841,N_24752);
nor UO_1867 (O_1867,N_24697,N_24503);
and UO_1868 (O_1868,N_24875,N_24973);
or UO_1869 (O_1869,N_24819,N_24719);
xnor UO_1870 (O_1870,N_24563,N_24701);
nand UO_1871 (O_1871,N_24835,N_24878);
or UO_1872 (O_1872,N_24583,N_24999);
nor UO_1873 (O_1873,N_24707,N_24956);
xnor UO_1874 (O_1874,N_24641,N_24671);
or UO_1875 (O_1875,N_24593,N_24595);
nor UO_1876 (O_1876,N_24853,N_24929);
and UO_1877 (O_1877,N_24882,N_24719);
nand UO_1878 (O_1878,N_24776,N_24674);
and UO_1879 (O_1879,N_24938,N_24933);
or UO_1880 (O_1880,N_24720,N_24828);
nor UO_1881 (O_1881,N_24756,N_24934);
nand UO_1882 (O_1882,N_24847,N_24892);
nand UO_1883 (O_1883,N_24931,N_24798);
nand UO_1884 (O_1884,N_24558,N_24947);
or UO_1885 (O_1885,N_24891,N_24877);
and UO_1886 (O_1886,N_24525,N_24876);
and UO_1887 (O_1887,N_24902,N_24783);
or UO_1888 (O_1888,N_24951,N_24680);
and UO_1889 (O_1889,N_24840,N_24504);
nor UO_1890 (O_1890,N_24824,N_24932);
and UO_1891 (O_1891,N_24854,N_24853);
xor UO_1892 (O_1892,N_24872,N_24938);
and UO_1893 (O_1893,N_24612,N_24849);
nor UO_1894 (O_1894,N_24905,N_24695);
or UO_1895 (O_1895,N_24796,N_24826);
nand UO_1896 (O_1896,N_24791,N_24540);
and UO_1897 (O_1897,N_24722,N_24693);
nor UO_1898 (O_1898,N_24511,N_24810);
nor UO_1899 (O_1899,N_24846,N_24641);
nand UO_1900 (O_1900,N_24762,N_24884);
or UO_1901 (O_1901,N_24805,N_24591);
nand UO_1902 (O_1902,N_24898,N_24687);
nor UO_1903 (O_1903,N_24921,N_24609);
nand UO_1904 (O_1904,N_24831,N_24573);
nor UO_1905 (O_1905,N_24511,N_24882);
nand UO_1906 (O_1906,N_24902,N_24882);
and UO_1907 (O_1907,N_24618,N_24604);
and UO_1908 (O_1908,N_24555,N_24724);
and UO_1909 (O_1909,N_24744,N_24804);
nand UO_1910 (O_1910,N_24785,N_24643);
or UO_1911 (O_1911,N_24664,N_24812);
xnor UO_1912 (O_1912,N_24719,N_24608);
nand UO_1913 (O_1913,N_24511,N_24530);
nor UO_1914 (O_1914,N_24543,N_24808);
nand UO_1915 (O_1915,N_24955,N_24920);
or UO_1916 (O_1916,N_24907,N_24812);
and UO_1917 (O_1917,N_24998,N_24959);
nand UO_1918 (O_1918,N_24720,N_24703);
nand UO_1919 (O_1919,N_24742,N_24701);
or UO_1920 (O_1920,N_24921,N_24942);
and UO_1921 (O_1921,N_24813,N_24956);
xnor UO_1922 (O_1922,N_24900,N_24561);
and UO_1923 (O_1923,N_24858,N_24869);
nand UO_1924 (O_1924,N_24504,N_24871);
nor UO_1925 (O_1925,N_24645,N_24884);
nor UO_1926 (O_1926,N_24702,N_24817);
nand UO_1927 (O_1927,N_24557,N_24601);
xnor UO_1928 (O_1928,N_24526,N_24668);
xor UO_1929 (O_1929,N_24904,N_24681);
or UO_1930 (O_1930,N_24939,N_24515);
nand UO_1931 (O_1931,N_24986,N_24714);
nor UO_1932 (O_1932,N_24539,N_24596);
nand UO_1933 (O_1933,N_24849,N_24694);
and UO_1934 (O_1934,N_24590,N_24973);
nand UO_1935 (O_1935,N_24684,N_24851);
nand UO_1936 (O_1936,N_24669,N_24534);
and UO_1937 (O_1937,N_24637,N_24629);
xnor UO_1938 (O_1938,N_24865,N_24987);
nand UO_1939 (O_1939,N_24771,N_24769);
or UO_1940 (O_1940,N_24975,N_24575);
nor UO_1941 (O_1941,N_24623,N_24817);
and UO_1942 (O_1942,N_24687,N_24836);
and UO_1943 (O_1943,N_24952,N_24544);
nor UO_1944 (O_1944,N_24635,N_24651);
xnor UO_1945 (O_1945,N_24774,N_24731);
xor UO_1946 (O_1946,N_24561,N_24595);
and UO_1947 (O_1947,N_24926,N_24977);
xor UO_1948 (O_1948,N_24505,N_24753);
xor UO_1949 (O_1949,N_24714,N_24554);
nand UO_1950 (O_1950,N_24766,N_24785);
nor UO_1951 (O_1951,N_24650,N_24779);
xnor UO_1952 (O_1952,N_24534,N_24983);
and UO_1953 (O_1953,N_24684,N_24943);
or UO_1954 (O_1954,N_24880,N_24810);
xor UO_1955 (O_1955,N_24848,N_24877);
xor UO_1956 (O_1956,N_24697,N_24645);
and UO_1957 (O_1957,N_24640,N_24767);
or UO_1958 (O_1958,N_24970,N_24505);
and UO_1959 (O_1959,N_24752,N_24784);
and UO_1960 (O_1960,N_24616,N_24525);
and UO_1961 (O_1961,N_24809,N_24992);
xor UO_1962 (O_1962,N_24820,N_24710);
nor UO_1963 (O_1963,N_24891,N_24871);
and UO_1964 (O_1964,N_24643,N_24576);
or UO_1965 (O_1965,N_24902,N_24586);
and UO_1966 (O_1966,N_24694,N_24501);
nor UO_1967 (O_1967,N_24686,N_24538);
or UO_1968 (O_1968,N_24953,N_24730);
nand UO_1969 (O_1969,N_24809,N_24882);
or UO_1970 (O_1970,N_24878,N_24932);
or UO_1971 (O_1971,N_24642,N_24887);
xor UO_1972 (O_1972,N_24741,N_24590);
and UO_1973 (O_1973,N_24781,N_24745);
nor UO_1974 (O_1974,N_24827,N_24911);
and UO_1975 (O_1975,N_24792,N_24709);
nor UO_1976 (O_1976,N_24801,N_24657);
and UO_1977 (O_1977,N_24540,N_24717);
nor UO_1978 (O_1978,N_24976,N_24525);
xor UO_1979 (O_1979,N_24818,N_24644);
xor UO_1980 (O_1980,N_24997,N_24840);
xor UO_1981 (O_1981,N_24736,N_24700);
nand UO_1982 (O_1982,N_24589,N_24926);
nor UO_1983 (O_1983,N_24819,N_24996);
nor UO_1984 (O_1984,N_24848,N_24902);
or UO_1985 (O_1985,N_24854,N_24698);
xnor UO_1986 (O_1986,N_24750,N_24999);
nand UO_1987 (O_1987,N_24783,N_24515);
xor UO_1988 (O_1988,N_24626,N_24699);
nor UO_1989 (O_1989,N_24990,N_24750);
nand UO_1990 (O_1990,N_24726,N_24623);
xor UO_1991 (O_1991,N_24751,N_24794);
and UO_1992 (O_1992,N_24997,N_24917);
nor UO_1993 (O_1993,N_24578,N_24548);
and UO_1994 (O_1994,N_24885,N_24579);
xnor UO_1995 (O_1995,N_24562,N_24830);
or UO_1996 (O_1996,N_24963,N_24625);
or UO_1997 (O_1997,N_24615,N_24655);
nand UO_1998 (O_1998,N_24738,N_24796);
nand UO_1999 (O_1999,N_24865,N_24883);
or UO_2000 (O_2000,N_24714,N_24778);
or UO_2001 (O_2001,N_24538,N_24663);
and UO_2002 (O_2002,N_24823,N_24902);
and UO_2003 (O_2003,N_24832,N_24713);
and UO_2004 (O_2004,N_24848,N_24572);
xnor UO_2005 (O_2005,N_24929,N_24930);
nor UO_2006 (O_2006,N_24573,N_24729);
or UO_2007 (O_2007,N_24827,N_24575);
xnor UO_2008 (O_2008,N_24928,N_24881);
xor UO_2009 (O_2009,N_24565,N_24506);
xor UO_2010 (O_2010,N_24726,N_24504);
or UO_2011 (O_2011,N_24702,N_24606);
or UO_2012 (O_2012,N_24759,N_24964);
and UO_2013 (O_2013,N_24627,N_24718);
nand UO_2014 (O_2014,N_24675,N_24753);
xnor UO_2015 (O_2015,N_24516,N_24628);
nand UO_2016 (O_2016,N_24609,N_24562);
nor UO_2017 (O_2017,N_24791,N_24970);
nor UO_2018 (O_2018,N_24627,N_24962);
nor UO_2019 (O_2019,N_24657,N_24747);
xnor UO_2020 (O_2020,N_24667,N_24699);
nand UO_2021 (O_2021,N_24935,N_24512);
xor UO_2022 (O_2022,N_24547,N_24548);
xnor UO_2023 (O_2023,N_24842,N_24866);
nor UO_2024 (O_2024,N_24899,N_24615);
nand UO_2025 (O_2025,N_24591,N_24702);
or UO_2026 (O_2026,N_24992,N_24608);
and UO_2027 (O_2027,N_24611,N_24565);
xor UO_2028 (O_2028,N_24765,N_24573);
and UO_2029 (O_2029,N_24745,N_24882);
and UO_2030 (O_2030,N_24914,N_24663);
nor UO_2031 (O_2031,N_24608,N_24709);
nand UO_2032 (O_2032,N_24800,N_24849);
xor UO_2033 (O_2033,N_24508,N_24829);
nor UO_2034 (O_2034,N_24835,N_24688);
xor UO_2035 (O_2035,N_24616,N_24743);
nand UO_2036 (O_2036,N_24624,N_24889);
nor UO_2037 (O_2037,N_24699,N_24981);
nand UO_2038 (O_2038,N_24504,N_24715);
xnor UO_2039 (O_2039,N_24608,N_24787);
xor UO_2040 (O_2040,N_24769,N_24618);
nor UO_2041 (O_2041,N_24753,N_24874);
or UO_2042 (O_2042,N_24562,N_24793);
nand UO_2043 (O_2043,N_24990,N_24540);
and UO_2044 (O_2044,N_24516,N_24750);
and UO_2045 (O_2045,N_24521,N_24946);
xor UO_2046 (O_2046,N_24595,N_24554);
nand UO_2047 (O_2047,N_24988,N_24862);
and UO_2048 (O_2048,N_24704,N_24628);
nand UO_2049 (O_2049,N_24651,N_24939);
xnor UO_2050 (O_2050,N_24698,N_24535);
and UO_2051 (O_2051,N_24864,N_24700);
and UO_2052 (O_2052,N_24776,N_24781);
xnor UO_2053 (O_2053,N_24567,N_24737);
nor UO_2054 (O_2054,N_24739,N_24793);
and UO_2055 (O_2055,N_24768,N_24777);
or UO_2056 (O_2056,N_24924,N_24812);
or UO_2057 (O_2057,N_24789,N_24560);
and UO_2058 (O_2058,N_24959,N_24712);
nand UO_2059 (O_2059,N_24992,N_24654);
nand UO_2060 (O_2060,N_24505,N_24942);
nor UO_2061 (O_2061,N_24633,N_24751);
or UO_2062 (O_2062,N_24844,N_24896);
nand UO_2063 (O_2063,N_24790,N_24690);
or UO_2064 (O_2064,N_24503,N_24853);
or UO_2065 (O_2065,N_24715,N_24866);
or UO_2066 (O_2066,N_24510,N_24886);
nand UO_2067 (O_2067,N_24594,N_24823);
or UO_2068 (O_2068,N_24941,N_24914);
xnor UO_2069 (O_2069,N_24502,N_24666);
nand UO_2070 (O_2070,N_24667,N_24530);
and UO_2071 (O_2071,N_24559,N_24615);
nand UO_2072 (O_2072,N_24899,N_24812);
xor UO_2073 (O_2073,N_24532,N_24945);
nor UO_2074 (O_2074,N_24503,N_24872);
nand UO_2075 (O_2075,N_24837,N_24880);
and UO_2076 (O_2076,N_24597,N_24655);
xor UO_2077 (O_2077,N_24891,N_24610);
xor UO_2078 (O_2078,N_24570,N_24609);
and UO_2079 (O_2079,N_24837,N_24700);
xnor UO_2080 (O_2080,N_24842,N_24534);
and UO_2081 (O_2081,N_24825,N_24599);
xnor UO_2082 (O_2082,N_24818,N_24534);
or UO_2083 (O_2083,N_24977,N_24917);
and UO_2084 (O_2084,N_24719,N_24637);
or UO_2085 (O_2085,N_24652,N_24715);
xor UO_2086 (O_2086,N_24967,N_24608);
nand UO_2087 (O_2087,N_24754,N_24591);
nor UO_2088 (O_2088,N_24633,N_24686);
and UO_2089 (O_2089,N_24926,N_24609);
nor UO_2090 (O_2090,N_24796,N_24765);
nor UO_2091 (O_2091,N_24559,N_24881);
nor UO_2092 (O_2092,N_24948,N_24934);
xor UO_2093 (O_2093,N_24577,N_24611);
xnor UO_2094 (O_2094,N_24883,N_24508);
nand UO_2095 (O_2095,N_24523,N_24888);
xnor UO_2096 (O_2096,N_24669,N_24805);
and UO_2097 (O_2097,N_24968,N_24562);
and UO_2098 (O_2098,N_24909,N_24928);
nand UO_2099 (O_2099,N_24935,N_24769);
nand UO_2100 (O_2100,N_24794,N_24960);
or UO_2101 (O_2101,N_24792,N_24854);
xnor UO_2102 (O_2102,N_24875,N_24712);
or UO_2103 (O_2103,N_24826,N_24613);
and UO_2104 (O_2104,N_24532,N_24891);
xnor UO_2105 (O_2105,N_24504,N_24879);
xnor UO_2106 (O_2106,N_24593,N_24540);
nor UO_2107 (O_2107,N_24775,N_24513);
xnor UO_2108 (O_2108,N_24572,N_24635);
nor UO_2109 (O_2109,N_24847,N_24946);
or UO_2110 (O_2110,N_24913,N_24854);
nor UO_2111 (O_2111,N_24752,N_24515);
nand UO_2112 (O_2112,N_24934,N_24915);
and UO_2113 (O_2113,N_24724,N_24645);
xor UO_2114 (O_2114,N_24648,N_24574);
xnor UO_2115 (O_2115,N_24870,N_24649);
or UO_2116 (O_2116,N_24915,N_24866);
xnor UO_2117 (O_2117,N_24601,N_24692);
xor UO_2118 (O_2118,N_24722,N_24631);
nand UO_2119 (O_2119,N_24992,N_24886);
nor UO_2120 (O_2120,N_24537,N_24830);
or UO_2121 (O_2121,N_24639,N_24942);
nand UO_2122 (O_2122,N_24693,N_24685);
xor UO_2123 (O_2123,N_24583,N_24805);
xnor UO_2124 (O_2124,N_24600,N_24578);
nor UO_2125 (O_2125,N_24999,N_24824);
nor UO_2126 (O_2126,N_24545,N_24848);
nand UO_2127 (O_2127,N_24844,N_24822);
or UO_2128 (O_2128,N_24899,N_24658);
or UO_2129 (O_2129,N_24765,N_24818);
and UO_2130 (O_2130,N_24586,N_24811);
nand UO_2131 (O_2131,N_24849,N_24555);
xor UO_2132 (O_2132,N_24570,N_24625);
nor UO_2133 (O_2133,N_24688,N_24524);
nand UO_2134 (O_2134,N_24542,N_24508);
nor UO_2135 (O_2135,N_24884,N_24814);
and UO_2136 (O_2136,N_24648,N_24935);
nand UO_2137 (O_2137,N_24673,N_24878);
nand UO_2138 (O_2138,N_24989,N_24819);
xor UO_2139 (O_2139,N_24676,N_24804);
nand UO_2140 (O_2140,N_24555,N_24831);
nor UO_2141 (O_2141,N_24648,N_24713);
xor UO_2142 (O_2142,N_24827,N_24832);
and UO_2143 (O_2143,N_24576,N_24788);
nor UO_2144 (O_2144,N_24716,N_24582);
xor UO_2145 (O_2145,N_24541,N_24680);
and UO_2146 (O_2146,N_24689,N_24705);
or UO_2147 (O_2147,N_24505,N_24833);
or UO_2148 (O_2148,N_24742,N_24582);
or UO_2149 (O_2149,N_24777,N_24606);
or UO_2150 (O_2150,N_24637,N_24660);
or UO_2151 (O_2151,N_24927,N_24900);
nand UO_2152 (O_2152,N_24586,N_24583);
nand UO_2153 (O_2153,N_24610,N_24720);
xor UO_2154 (O_2154,N_24704,N_24674);
xor UO_2155 (O_2155,N_24872,N_24977);
xnor UO_2156 (O_2156,N_24674,N_24838);
nand UO_2157 (O_2157,N_24824,N_24556);
or UO_2158 (O_2158,N_24951,N_24792);
xnor UO_2159 (O_2159,N_24962,N_24956);
nor UO_2160 (O_2160,N_24541,N_24788);
or UO_2161 (O_2161,N_24706,N_24712);
or UO_2162 (O_2162,N_24738,N_24912);
and UO_2163 (O_2163,N_24792,N_24844);
xnor UO_2164 (O_2164,N_24619,N_24695);
nor UO_2165 (O_2165,N_24677,N_24939);
nand UO_2166 (O_2166,N_24536,N_24532);
nor UO_2167 (O_2167,N_24849,N_24994);
nor UO_2168 (O_2168,N_24936,N_24542);
nor UO_2169 (O_2169,N_24654,N_24927);
nor UO_2170 (O_2170,N_24670,N_24765);
nand UO_2171 (O_2171,N_24874,N_24934);
and UO_2172 (O_2172,N_24725,N_24563);
xnor UO_2173 (O_2173,N_24700,N_24744);
or UO_2174 (O_2174,N_24788,N_24557);
xnor UO_2175 (O_2175,N_24760,N_24818);
and UO_2176 (O_2176,N_24847,N_24853);
xnor UO_2177 (O_2177,N_24523,N_24734);
nand UO_2178 (O_2178,N_24936,N_24739);
xnor UO_2179 (O_2179,N_24556,N_24977);
or UO_2180 (O_2180,N_24755,N_24643);
and UO_2181 (O_2181,N_24654,N_24764);
or UO_2182 (O_2182,N_24961,N_24932);
xor UO_2183 (O_2183,N_24574,N_24879);
nor UO_2184 (O_2184,N_24654,N_24753);
xor UO_2185 (O_2185,N_24507,N_24982);
and UO_2186 (O_2186,N_24764,N_24802);
and UO_2187 (O_2187,N_24992,N_24833);
xor UO_2188 (O_2188,N_24911,N_24580);
nor UO_2189 (O_2189,N_24525,N_24881);
nor UO_2190 (O_2190,N_24564,N_24628);
and UO_2191 (O_2191,N_24977,N_24576);
xor UO_2192 (O_2192,N_24687,N_24527);
nand UO_2193 (O_2193,N_24927,N_24556);
or UO_2194 (O_2194,N_24622,N_24856);
xnor UO_2195 (O_2195,N_24749,N_24993);
nor UO_2196 (O_2196,N_24600,N_24612);
xnor UO_2197 (O_2197,N_24671,N_24538);
xnor UO_2198 (O_2198,N_24752,N_24807);
nand UO_2199 (O_2199,N_24670,N_24711);
and UO_2200 (O_2200,N_24912,N_24775);
nand UO_2201 (O_2201,N_24781,N_24882);
or UO_2202 (O_2202,N_24788,N_24853);
nor UO_2203 (O_2203,N_24532,N_24855);
nand UO_2204 (O_2204,N_24735,N_24634);
xnor UO_2205 (O_2205,N_24605,N_24524);
xor UO_2206 (O_2206,N_24782,N_24832);
xnor UO_2207 (O_2207,N_24685,N_24761);
nand UO_2208 (O_2208,N_24976,N_24519);
or UO_2209 (O_2209,N_24656,N_24888);
nor UO_2210 (O_2210,N_24837,N_24743);
and UO_2211 (O_2211,N_24677,N_24930);
and UO_2212 (O_2212,N_24794,N_24796);
and UO_2213 (O_2213,N_24533,N_24705);
nand UO_2214 (O_2214,N_24961,N_24511);
nor UO_2215 (O_2215,N_24966,N_24902);
nor UO_2216 (O_2216,N_24736,N_24551);
nand UO_2217 (O_2217,N_24525,N_24795);
nand UO_2218 (O_2218,N_24535,N_24530);
xnor UO_2219 (O_2219,N_24552,N_24604);
nand UO_2220 (O_2220,N_24860,N_24629);
or UO_2221 (O_2221,N_24982,N_24908);
nor UO_2222 (O_2222,N_24942,N_24786);
nor UO_2223 (O_2223,N_24542,N_24561);
or UO_2224 (O_2224,N_24790,N_24803);
or UO_2225 (O_2225,N_24780,N_24530);
nor UO_2226 (O_2226,N_24947,N_24564);
nand UO_2227 (O_2227,N_24704,N_24710);
or UO_2228 (O_2228,N_24625,N_24903);
or UO_2229 (O_2229,N_24513,N_24689);
or UO_2230 (O_2230,N_24823,N_24728);
xnor UO_2231 (O_2231,N_24819,N_24586);
nand UO_2232 (O_2232,N_24811,N_24712);
xnor UO_2233 (O_2233,N_24515,N_24661);
xor UO_2234 (O_2234,N_24749,N_24805);
nand UO_2235 (O_2235,N_24628,N_24728);
or UO_2236 (O_2236,N_24904,N_24672);
xnor UO_2237 (O_2237,N_24792,N_24971);
and UO_2238 (O_2238,N_24943,N_24605);
or UO_2239 (O_2239,N_24849,N_24943);
nand UO_2240 (O_2240,N_24937,N_24794);
or UO_2241 (O_2241,N_24727,N_24705);
or UO_2242 (O_2242,N_24923,N_24918);
and UO_2243 (O_2243,N_24864,N_24811);
xnor UO_2244 (O_2244,N_24657,N_24660);
nand UO_2245 (O_2245,N_24723,N_24797);
xor UO_2246 (O_2246,N_24906,N_24713);
xor UO_2247 (O_2247,N_24806,N_24747);
nand UO_2248 (O_2248,N_24810,N_24764);
nor UO_2249 (O_2249,N_24517,N_24899);
or UO_2250 (O_2250,N_24801,N_24905);
and UO_2251 (O_2251,N_24895,N_24631);
xor UO_2252 (O_2252,N_24985,N_24643);
xnor UO_2253 (O_2253,N_24613,N_24640);
or UO_2254 (O_2254,N_24646,N_24975);
and UO_2255 (O_2255,N_24875,N_24990);
nand UO_2256 (O_2256,N_24985,N_24537);
or UO_2257 (O_2257,N_24788,N_24790);
xnor UO_2258 (O_2258,N_24896,N_24573);
nand UO_2259 (O_2259,N_24944,N_24694);
or UO_2260 (O_2260,N_24845,N_24586);
nor UO_2261 (O_2261,N_24799,N_24606);
or UO_2262 (O_2262,N_24903,N_24987);
xor UO_2263 (O_2263,N_24586,N_24831);
xnor UO_2264 (O_2264,N_24918,N_24748);
or UO_2265 (O_2265,N_24576,N_24759);
or UO_2266 (O_2266,N_24517,N_24968);
nand UO_2267 (O_2267,N_24544,N_24752);
or UO_2268 (O_2268,N_24600,N_24819);
nor UO_2269 (O_2269,N_24585,N_24777);
xnor UO_2270 (O_2270,N_24970,N_24915);
xor UO_2271 (O_2271,N_24853,N_24897);
nand UO_2272 (O_2272,N_24778,N_24674);
nand UO_2273 (O_2273,N_24998,N_24717);
and UO_2274 (O_2274,N_24688,N_24617);
xnor UO_2275 (O_2275,N_24725,N_24785);
xnor UO_2276 (O_2276,N_24952,N_24981);
or UO_2277 (O_2277,N_24717,N_24661);
xnor UO_2278 (O_2278,N_24522,N_24602);
and UO_2279 (O_2279,N_24761,N_24583);
xor UO_2280 (O_2280,N_24991,N_24880);
xnor UO_2281 (O_2281,N_24645,N_24788);
xor UO_2282 (O_2282,N_24649,N_24731);
nand UO_2283 (O_2283,N_24668,N_24992);
or UO_2284 (O_2284,N_24640,N_24603);
nand UO_2285 (O_2285,N_24854,N_24982);
or UO_2286 (O_2286,N_24612,N_24877);
or UO_2287 (O_2287,N_24991,N_24796);
or UO_2288 (O_2288,N_24918,N_24619);
nand UO_2289 (O_2289,N_24788,N_24703);
xnor UO_2290 (O_2290,N_24885,N_24747);
or UO_2291 (O_2291,N_24722,N_24516);
nor UO_2292 (O_2292,N_24976,N_24889);
nor UO_2293 (O_2293,N_24776,N_24960);
nand UO_2294 (O_2294,N_24522,N_24709);
nor UO_2295 (O_2295,N_24782,N_24742);
xnor UO_2296 (O_2296,N_24922,N_24716);
nor UO_2297 (O_2297,N_24906,N_24606);
nand UO_2298 (O_2298,N_24831,N_24852);
nor UO_2299 (O_2299,N_24803,N_24555);
and UO_2300 (O_2300,N_24601,N_24753);
and UO_2301 (O_2301,N_24727,N_24967);
xnor UO_2302 (O_2302,N_24690,N_24716);
xnor UO_2303 (O_2303,N_24804,N_24548);
or UO_2304 (O_2304,N_24538,N_24948);
or UO_2305 (O_2305,N_24639,N_24866);
xor UO_2306 (O_2306,N_24545,N_24611);
xor UO_2307 (O_2307,N_24789,N_24853);
nand UO_2308 (O_2308,N_24934,N_24504);
and UO_2309 (O_2309,N_24511,N_24843);
nand UO_2310 (O_2310,N_24815,N_24567);
nand UO_2311 (O_2311,N_24740,N_24846);
xnor UO_2312 (O_2312,N_24521,N_24696);
and UO_2313 (O_2313,N_24808,N_24790);
nand UO_2314 (O_2314,N_24900,N_24934);
nor UO_2315 (O_2315,N_24511,N_24865);
or UO_2316 (O_2316,N_24756,N_24966);
and UO_2317 (O_2317,N_24566,N_24521);
nor UO_2318 (O_2318,N_24634,N_24903);
and UO_2319 (O_2319,N_24779,N_24945);
nor UO_2320 (O_2320,N_24518,N_24881);
nand UO_2321 (O_2321,N_24786,N_24601);
nor UO_2322 (O_2322,N_24837,N_24608);
nand UO_2323 (O_2323,N_24849,N_24503);
xnor UO_2324 (O_2324,N_24835,N_24524);
nor UO_2325 (O_2325,N_24986,N_24689);
and UO_2326 (O_2326,N_24700,N_24817);
or UO_2327 (O_2327,N_24502,N_24722);
or UO_2328 (O_2328,N_24741,N_24578);
or UO_2329 (O_2329,N_24960,N_24658);
or UO_2330 (O_2330,N_24702,N_24664);
or UO_2331 (O_2331,N_24958,N_24718);
and UO_2332 (O_2332,N_24939,N_24578);
nor UO_2333 (O_2333,N_24977,N_24653);
xnor UO_2334 (O_2334,N_24653,N_24827);
nor UO_2335 (O_2335,N_24593,N_24898);
xnor UO_2336 (O_2336,N_24991,N_24656);
and UO_2337 (O_2337,N_24584,N_24745);
nand UO_2338 (O_2338,N_24594,N_24675);
nand UO_2339 (O_2339,N_24829,N_24849);
nor UO_2340 (O_2340,N_24638,N_24524);
nand UO_2341 (O_2341,N_24891,N_24882);
xnor UO_2342 (O_2342,N_24745,N_24675);
xnor UO_2343 (O_2343,N_24518,N_24715);
and UO_2344 (O_2344,N_24753,N_24536);
nand UO_2345 (O_2345,N_24796,N_24639);
or UO_2346 (O_2346,N_24544,N_24883);
and UO_2347 (O_2347,N_24969,N_24724);
and UO_2348 (O_2348,N_24503,N_24908);
nor UO_2349 (O_2349,N_24701,N_24653);
xor UO_2350 (O_2350,N_24521,N_24545);
and UO_2351 (O_2351,N_24529,N_24908);
nor UO_2352 (O_2352,N_24855,N_24931);
nor UO_2353 (O_2353,N_24889,N_24728);
xor UO_2354 (O_2354,N_24825,N_24988);
or UO_2355 (O_2355,N_24826,N_24773);
and UO_2356 (O_2356,N_24929,N_24546);
xnor UO_2357 (O_2357,N_24822,N_24687);
or UO_2358 (O_2358,N_24913,N_24891);
nand UO_2359 (O_2359,N_24790,N_24994);
xor UO_2360 (O_2360,N_24838,N_24542);
or UO_2361 (O_2361,N_24662,N_24863);
xor UO_2362 (O_2362,N_24640,N_24634);
and UO_2363 (O_2363,N_24970,N_24645);
and UO_2364 (O_2364,N_24748,N_24742);
nor UO_2365 (O_2365,N_24906,N_24968);
nand UO_2366 (O_2366,N_24692,N_24747);
or UO_2367 (O_2367,N_24923,N_24712);
nand UO_2368 (O_2368,N_24548,N_24656);
nor UO_2369 (O_2369,N_24801,N_24799);
nand UO_2370 (O_2370,N_24641,N_24625);
xnor UO_2371 (O_2371,N_24713,N_24745);
nor UO_2372 (O_2372,N_24665,N_24686);
or UO_2373 (O_2373,N_24844,N_24989);
and UO_2374 (O_2374,N_24662,N_24835);
nor UO_2375 (O_2375,N_24945,N_24553);
nand UO_2376 (O_2376,N_24794,N_24609);
nor UO_2377 (O_2377,N_24669,N_24903);
and UO_2378 (O_2378,N_24761,N_24679);
or UO_2379 (O_2379,N_24943,N_24653);
xnor UO_2380 (O_2380,N_24949,N_24618);
nor UO_2381 (O_2381,N_24946,N_24980);
nor UO_2382 (O_2382,N_24881,N_24993);
nand UO_2383 (O_2383,N_24644,N_24727);
xor UO_2384 (O_2384,N_24991,N_24521);
or UO_2385 (O_2385,N_24964,N_24983);
xor UO_2386 (O_2386,N_24608,N_24519);
nand UO_2387 (O_2387,N_24921,N_24829);
xor UO_2388 (O_2388,N_24814,N_24505);
and UO_2389 (O_2389,N_24606,N_24952);
nand UO_2390 (O_2390,N_24953,N_24523);
nand UO_2391 (O_2391,N_24668,N_24507);
xor UO_2392 (O_2392,N_24619,N_24517);
and UO_2393 (O_2393,N_24732,N_24999);
nand UO_2394 (O_2394,N_24765,N_24850);
nand UO_2395 (O_2395,N_24825,N_24730);
or UO_2396 (O_2396,N_24791,N_24811);
nand UO_2397 (O_2397,N_24657,N_24756);
or UO_2398 (O_2398,N_24898,N_24625);
nor UO_2399 (O_2399,N_24562,N_24855);
nand UO_2400 (O_2400,N_24742,N_24607);
or UO_2401 (O_2401,N_24690,N_24901);
or UO_2402 (O_2402,N_24501,N_24564);
nand UO_2403 (O_2403,N_24530,N_24911);
nor UO_2404 (O_2404,N_24640,N_24572);
nand UO_2405 (O_2405,N_24668,N_24654);
nand UO_2406 (O_2406,N_24699,N_24754);
nor UO_2407 (O_2407,N_24939,N_24796);
nor UO_2408 (O_2408,N_24971,N_24567);
nand UO_2409 (O_2409,N_24504,N_24945);
nor UO_2410 (O_2410,N_24944,N_24870);
xnor UO_2411 (O_2411,N_24945,N_24946);
nand UO_2412 (O_2412,N_24799,N_24774);
nand UO_2413 (O_2413,N_24729,N_24705);
and UO_2414 (O_2414,N_24940,N_24521);
or UO_2415 (O_2415,N_24529,N_24507);
or UO_2416 (O_2416,N_24943,N_24985);
nand UO_2417 (O_2417,N_24661,N_24576);
nor UO_2418 (O_2418,N_24782,N_24909);
and UO_2419 (O_2419,N_24826,N_24840);
nor UO_2420 (O_2420,N_24873,N_24727);
or UO_2421 (O_2421,N_24554,N_24566);
xor UO_2422 (O_2422,N_24723,N_24656);
xor UO_2423 (O_2423,N_24787,N_24902);
nand UO_2424 (O_2424,N_24739,N_24860);
xnor UO_2425 (O_2425,N_24975,N_24980);
xnor UO_2426 (O_2426,N_24994,N_24614);
nor UO_2427 (O_2427,N_24509,N_24760);
and UO_2428 (O_2428,N_24716,N_24527);
nor UO_2429 (O_2429,N_24727,N_24502);
or UO_2430 (O_2430,N_24639,N_24910);
nand UO_2431 (O_2431,N_24586,N_24808);
nand UO_2432 (O_2432,N_24950,N_24547);
xor UO_2433 (O_2433,N_24777,N_24661);
or UO_2434 (O_2434,N_24742,N_24904);
xnor UO_2435 (O_2435,N_24874,N_24571);
xnor UO_2436 (O_2436,N_24883,N_24746);
or UO_2437 (O_2437,N_24607,N_24646);
nor UO_2438 (O_2438,N_24665,N_24633);
xnor UO_2439 (O_2439,N_24577,N_24699);
nor UO_2440 (O_2440,N_24895,N_24743);
nand UO_2441 (O_2441,N_24815,N_24790);
xnor UO_2442 (O_2442,N_24710,N_24536);
and UO_2443 (O_2443,N_24662,N_24767);
or UO_2444 (O_2444,N_24778,N_24797);
nand UO_2445 (O_2445,N_24914,N_24796);
nand UO_2446 (O_2446,N_24503,N_24753);
or UO_2447 (O_2447,N_24972,N_24556);
and UO_2448 (O_2448,N_24783,N_24781);
nand UO_2449 (O_2449,N_24802,N_24839);
and UO_2450 (O_2450,N_24509,N_24926);
or UO_2451 (O_2451,N_24626,N_24703);
nor UO_2452 (O_2452,N_24630,N_24526);
and UO_2453 (O_2453,N_24753,N_24572);
and UO_2454 (O_2454,N_24786,N_24621);
or UO_2455 (O_2455,N_24588,N_24708);
nor UO_2456 (O_2456,N_24890,N_24582);
and UO_2457 (O_2457,N_24982,N_24600);
nand UO_2458 (O_2458,N_24647,N_24809);
and UO_2459 (O_2459,N_24831,N_24777);
nand UO_2460 (O_2460,N_24814,N_24947);
xor UO_2461 (O_2461,N_24560,N_24770);
and UO_2462 (O_2462,N_24807,N_24985);
nand UO_2463 (O_2463,N_24644,N_24584);
or UO_2464 (O_2464,N_24683,N_24750);
and UO_2465 (O_2465,N_24588,N_24658);
xnor UO_2466 (O_2466,N_24922,N_24638);
nand UO_2467 (O_2467,N_24957,N_24763);
nand UO_2468 (O_2468,N_24533,N_24903);
or UO_2469 (O_2469,N_24924,N_24765);
nor UO_2470 (O_2470,N_24865,N_24641);
nor UO_2471 (O_2471,N_24591,N_24615);
xor UO_2472 (O_2472,N_24574,N_24690);
xnor UO_2473 (O_2473,N_24534,N_24969);
or UO_2474 (O_2474,N_24876,N_24896);
or UO_2475 (O_2475,N_24915,N_24955);
or UO_2476 (O_2476,N_24919,N_24870);
nor UO_2477 (O_2477,N_24930,N_24848);
and UO_2478 (O_2478,N_24611,N_24882);
nor UO_2479 (O_2479,N_24825,N_24739);
xnor UO_2480 (O_2480,N_24975,N_24795);
nor UO_2481 (O_2481,N_24877,N_24908);
nand UO_2482 (O_2482,N_24760,N_24984);
nand UO_2483 (O_2483,N_24709,N_24938);
nand UO_2484 (O_2484,N_24504,N_24685);
nand UO_2485 (O_2485,N_24531,N_24552);
or UO_2486 (O_2486,N_24786,N_24787);
nand UO_2487 (O_2487,N_24697,N_24629);
xnor UO_2488 (O_2488,N_24794,N_24911);
or UO_2489 (O_2489,N_24502,N_24907);
nor UO_2490 (O_2490,N_24773,N_24785);
nand UO_2491 (O_2491,N_24819,N_24806);
nand UO_2492 (O_2492,N_24547,N_24890);
nand UO_2493 (O_2493,N_24588,N_24748);
xnor UO_2494 (O_2494,N_24594,N_24854);
nand UO_2495 (O_2495,N_24714,N_24780);
nor UO_2496 (O_2496,N_24817,N_24570);
nor UO_2497 (O_2497,N_24899,N_24677);
and UO_2498 (O_2498,N_24742,N_24958);
xor UO_2499 (O_2499,N_24607,N_24705);
and UO_2500 (O_2500,N_24639,N_24693);
nor UO_2501 (O_2501,N_24700,N_24561);
nor UO_2502 (O_2502,N_24641,N_24511);
xor UO_2503 (O_2503,N_24608,N_24936);
nand UO_2504 (O_2504,N_24709,N_24979);
or UO_2505 (O_2505,N_24647,N_24566);
nand UO_2506 (O_2506,N_24594,N_24752);
nor UO_2507 (O_2507,N_24844,N_24709);
nor UO_2508 (O_2508,N_24735,N_24663);
nor UO_2509 (O_2509,N_24649,N_24701);
nor UO_2510 (O_2510,N_24752,N_24839);
and UO_2511 (O_2511,N_24641,N_24629);
xnor UO_2512 (O_2512,N_24905,N_24879);
or UO_2513 (O_2513,N_24866,N_24534);
xor UO_2514 (O_2514,N_24565,N_24958);
and UO_2515 (O_2515,N_24825,N_24953);
or UO_2516 (O_2516,N_24673,N_24714);
or UO_2517 (O_2517,N_24979,N_24705);
or UO_2518 (O_2518,N_24743,N_24712);
nor UO_2519 (O_2519,N_24891,N_24604);
and UO_2520 (O_2520,N_24764,N_24901);
or UO_2521 (O_2521,N_24727,N_24816);
or UO_2522 (O_2522,N_24699,N_24615);
nand UO_2523 (O_2523,N_24868,N_24829);
nand UO_2524 (O_2524,N_24826,N_24836);
nand UO_2525 (O_2525,N_24592,N_24908);
or UO_2526 (O_2526,N_24939,N_24646);
nor UO_2527 (O_2527,N_24517,N_24628);
and UO_2528 (O_2528,N_24961,N_24502);
nor UO_2529 (O_2529,N_24862,N_24633);
nor UO_2530 (O_2530,N_24658,N_24937);
nor UO_2531 (O_2531,N_24619,N_24855);
nor UO_2532 (O_2532,N_24745,N_24805);
xnor UO_2533 (O_2533,N_24719,N_24788);
nand UO_2534 (O_2534,N_24885,N_24691);
xnor UO_2535 (O_2535,N_24975,N_24651);
or UO_2536 (O_2536,N_24627,N_24645);
nor UO_2537 (O_2537,N_24768,N_24889);
nor UO_2538 (O_2538,N_24803,N_24590);
nor UO_2539 (O_2539,N_24888,N_24771);
nand UO_2540 (O_2540,N_24973,N_24826);
xor UO_2541 (O_2541,N_24818,N_24931);
nand UO_2542 (O_2542,N_24838,N_24992);
nor UO_2543 (O_2543,N_24718,N_24971);
xnor UO_2544 (O_2544,N_24950,N_24937);
and UO_2545 (O_2545,N_24928,N_24502);
xor UO_2546 (O_2546,N_24990,N_24696);
and UO_2547 (O_2547,N_24638,N_24647);
and UO_2548 (O_2548,N_24775,N_24694);
or UO_2549 (O_2549,N_24938,N_24664);
nand UO_2550 (O_2550,N_24823,N_24864);
nand UO_2551 (O_2551,N_24854,N_24847);
xnor UO_2552 (O_2552,N_24613,N_24615);
and UO_2553 (O_2553,N_24558,N_24786);
and UO_2554 (O_2554,N_24831,N_24510);
nor UO_2555 (O_2555,N_24742,N_24688);
nor UO_2556 (O_2556,N_24951,N_24923);
nor UO_2557 (O_2557,N_24971,N_24969);
nor UO_2558 (O_2558,N_24703,N_24856);
and UO_2559 (O_2559,N_24672,N_24561);
or UO_2560 (O_2560,N_24556,N_24953);
or UO_2561 (O_2561,N_24793,N_24665);
and UO_2562 (O_2562,N_24933,N_24600);
or UO_2563 (O_2563,N_24980,N_24805);
nand UO_2564 (O_2564,N_24742,N_24655);
nor UO_2565 (O_2565,N_24810,N_24773);
xnor UO_2566 (O_2566,N_24576,N_24974);
xor UO_2567 (O_2567,N_24685,N_24535);
or UO_2568 (O_2568,N_24726,N_24667);
xnor UO_2569 (O_2569,N_24693,N_24827);
nor UO_2570 (O_2570,N_24899,N_24825);
nor UO_2571 (O_2571,N_24757,N_24645);
and UO_2572 (O_2572,N_24718,N_24972);
and UO_2573 (O_2573,N_24549,N_24856);
or UO_2574 (O_2574,N_24773,N_24725);
or UO_2575 (O_2575,N_24969,N_24808);
and UO_2576 (O_2576,N_24533,N_24506);
nand UO_2577 (O_2577,N_24501,N_24712);
nor UO_2578 (O_2578,N_24921,N_24511);
nor UO_2579 (O_2579,N_24827,N_24801);
xor UO_2580 (O_2580,N_24573,N_24690);
nand UO_2581 (O_2581,N_24899,N_24699);
nor UO_2582 (O_2582,N_24700,N_24521);
nand UO_2583 (O_2583,N_24997,N_24868);
nor UO_2584 (O_2584,N_24695,N_24518);
or UO_2585 (O_2585,N_24645,N_24789);
xnor UO_2586 (O_2586,N_24702,N_24855);
xor UO_2587 (O_2587,N_24820,N_24557);
and UO_2588 (O_2588,N_24618,N_24754);
or UO_2589 (O_2589,N_24615,N_24623);
or UO_2590 (O_2590,N_24651,N_24730);
xnor UO_2591 (O_2591,N_24880,N_24504);
nor UO_2592 (O_2592,N_24603,N_24512);
xnor UO_2593 (O_2593,N_24810,N_24723);
nor UO_2594 (O_2594,N_24652,N_24694);
and UO_2595 (O_2595,N_24716,N_24567);
or UO_2596 (O_2596,N_24891,N_24966);
nand UO_2597 (O_2597,N_24926,N_24565);
xnor UO_2598 (O_2598,N_24821,N_24755);
and UO_2599 (O_2599,N_24799,N_24758);
and UO_2600 (O_2600,N_24634,N_24512);
and UO_2601 (O_2601,N_24829,N_24928);
or UO_2602 (O_2602,N_24613,N_24669);
or UO_2603 (O_2603,N_24832,N_24867);
or UO_2604 (O_2604,N_24857,N_24568);
nand UO_2605 (O_2605,N_24538,N_24561);
xor UO_2606 (O_2606,N_24739,N_24605);
and UO_2607 (O_2607,N_24858,N_24848);
xnor UO_2608 (O_2608,N_24801,N_24661);
xor UO_2609 (O_2609,N_24875,N_24507);
and UO_2610 (O_2610,N_24599,N_24800);
nor UO_2611 (O_2611,N_24597,N_24709);
and UO_2612 (O_2612,N_24538,N_24800);
nor UO_2613 (O_2613,N_24857,N_24655);
xor UO_2614 (O_2614,N_24567,N_24651);
or UO_2615 (O_2615,N_24959,N_24532);
and UO_2616 (O_2616,N_24676,N_24625);
nor UO_2617 (O_2617,N_24501,N_24949);
nor UO_2618 (O_2618,N_24845,N_24528);
nor UO_2619 (O_2619,N_24693,N_24786);
nand UO_2620 (O_2620,N_24790,N_24912);
and UO_2621 (O_2621,N_24831,N_24590);
nor UO_2622 (O_2622,N_24794,N_24848);
nor UO_2623 (O_2623,N_24633,N_24997);
nand UO_2624 (O_2624,N_24753,N_24583);
and UO_2625 (O_2625,N_24765,N_24543);
or UO_2626 (O_2626,N_24555,N_24870);
and UO_2627 (O_2627,N_24587,N_24834);
xor UO_2628 (O_2628,N_24776,N_24534);
and UO_2629 (O_2629,N_24793,N_24872);
and UO_2630 (O_2630,N_24948,N_24851);
and UO_2631 (O_2631,N_24894,N_24629);
or UO_2632 (O_2632,N_24950,N_24956);
nor UO_2633 (O_2633,N_24547,N_24843);
nand UO_2634 (O_2634,N_24565,N_24582);
or UO_2635 (O_2635,N_24801,N_24995);
xor UO_2636 (O_2636,N_24507,N_24670);
nor UO_2637 (O_2637,N_24905,N_24627);
or UO_2638 (O_2638,N_24940,N_24624);
or UO_2639 (O_2639,N_24995,N_24551);
xnor UO_2640 (O_2640,N_24614,N_24774);
nor UO_2641 (O_2641,N_24709,N_24580);
nand UO_2642 (O_2642,N_24939,N_24916);
xor UO_2643 (O_2643,N_24546,N_24740);
nor UO_2644 (O_2644,N_24511,N_24777);
nand UO_2645 (O_2645,N_24541,N_24580);
xor UO_2646 (O_2646,N_24807,N_24853);
nand UO_2647 (O_2647,N_24891,N_24689);
and UO_2648 (O_2648,N_24766,N_24697);
and UO_2649 (O_2649,N_24619,N_24502);
xnor UO_2650 (O_2650,N_24921,N_24736);
nor UO_2651 (O_2651,N_24570,N_24882);
nor UO_2652 (O_2652,N_24823,N_24607);
and UO_2653 (O_2653,N_24843,N_24638);
nand UO_2654 (O_2654,N_24951,N_24518);
and UO_2655 (O_2655,N_24882,N_24641);
nand UO_2656 (O_2656,N_24958,N_24903);
or UO_2657 (O_2657,N_24523,N_24860);
nand UO_2658 (O_2658,N_24691,N_24716);
xnor UO_2659 (O_2659,N_24941,N_24545);
nand UO_2660 (O_2660,N_24803,N_24722);
xnor UO_2661 (O_2661,N_24775,N_24862);
and UO_2662 (O_2662,N_24800,N_24731);
or UO_2663 (O_2663,N_24915,N_24894);
or UO_2664 (O_2664,N_24561,N_24792);
or UO_2665 (O_2665,N_24701,N_24854);
nor UO_2666 (O_2666,N_24525,N_24877);
xor UO_2667 (O_2667,N_24804,N_24534);
nor UO_2668 (O_2668,N_24742,N_24671);
nand UO_2669 (O_2669,N_24840,N_24708);
nor UO_2670 (O_2670,N_24674,N_24991);
or UO_2671 (O_2671,N_24695,N_24993);
xor UO_2672 (O_2672,N_24532,N_24584);
or UO_2673 (O_2673,N_24718,N_24529);
nor UO_2674 (O_2674,N_24577,N_24630);
xnor UO_2675 (O_2675,N_24729,N_24665);
nand UO_2676 (O_2676,N_24941,N_24981);
or UO_2677 (O_2677,N_24751,N_24801);
xnor UO_2678 (O_2678,N_24868,N_24914);
nor UO_2679 (O_2679,N_24732,N_24822);
xnor UO_2680 (O_2680,N_24589,N_24508);
nor UO_2681 (O_2681,N_24771,N_24952);
or UO_2682 (O_2682,N_24539,N_24969);
xor UO_2683 (O_2683,N_24846,N_24917);
or UO_2684 (O_2684,N_24697,N_24749);
nor UO_2685 (O_2685,N_24776,N_24704);
or UO_2686 (O_2686,N_24664,N_24794);
and UO_2687 (O_2687,N_24882,N_24612);
and UO_2688 (O_2688,N_24576,N_24517);
nand UO_2689 (O_2689,N_24975,N_24838);
and UO_2690 (O_2690,N_24619,N_24655);
xor UO_2691 (O_2691,N_24780,N_24560);
nand UO_2692 (O_2692,N_24756,N_24973);
nor UO_2693 (O_2693,N_24507,N_24940);
and UO_2694 (O_2694,N_24831,N_24832);
xnor UO_2695 (O_2695,N_24978,N_24737);
or UO_2696 (O_2696,N_24767,N_24968);
nand UO_2697 (O_2697,N_24972,N_24599);
nand UO_2698 (O_2698,N_24789,N_24775);
or UO_2699 (O_2699,N_24881,N_24794);
xor UO_2700 (O_2700,N_24666,N_24700);
xnor UO_2701 (O_2701,N_24747,N_24618);
or UO_2702 (O_2702,N_24870,N_24635);
nor UO_2703 (O_2703,N_24528,N_24835);
and UO_2704 (O_2704,N_24786,N_24723);
and UO_2705 (O_2705,N_24793,N_24914);
nor UO_2706 (O_2706,N_24523,N_24667);
and UO_2707 (O_2707,N_24739,N_24704);
nand UO_2708 (O_2708,N_24783,N_24539);
nor UO_2709 (O_2709,N_24739,N_24757);
nand UO_2710 (O_2710,N_24506,N_24935);
nand UO_2711 (O_2711,N_24894,N_24662);
and UO_2712 (O_2712,N_24550,N_24696);
or UO_2713 (O_2713,N_24739,N_24698);
or UO_2714 (O_2714,N_24960,N_24529);
xnor UO_2715 (O_2715,N_24620,N_24946);
and UO_2716 (O_2716,N_24621,N_24784);
nand UO_2717 (O_2717,N_24584,N_24975);
and UO_2718 (O_2718,N_24747,N_24627);
nand UO_2719 (O_2719,N_24923,N_24715);
nor UO_2720 (O_2720,N_24896,N_24701);
xnor UO_2721 (O_2721,N_24562,N_24826);
and UO_2722 (O_2722,N_24700,N_24944);
nand UO_2723 (O_2723,N_24509,N_24697);
or UO_2724 (O_2724,N_24854,N_24546);
nor UO_2725 (O_2725,N_24599,N_24878);
or UO_2726 (O_2726,N_24856,N_24630);
and UO_2727 (O_2727,N_24850,N_24623);
or UO_2728 (O_2728,N_24712,N_24793);
nand UO_2729 (O_2729,N_24519,N_24956);
xnor UO_2730 (O_2730,N_24864,N_24570);
nand UO_2731 (O_2731,N_24951,N_24959);
or UO_2732 (O_2732,N_24662,N_24535);
nand UO_2733 (O_2733,N_24876,N_24957);
xor UO_2734 (O_2734,N_24735,N_24803);
nand UO_2735 (O_2735,N_24533,N_24772);
and UO_2736 (O_2736,N_24518,N_24884);
nand UO_2737 (O_2737,N_24791,N_24801);
nor UO_2738 (O_2738,N_24687,N_24663);
and UO_2739 (O_2739,N_24581,N_24931);
and UO_2740 (O_2740,N_24826,N_24785);
nor UO_2741 (O_2741,N_24964,N_24531);
and UO_2742 (O_2742,N_24549,N_24796);
nor UO_2743 (O_2743,N_24869,N_24729);
or UO_2744 (O_2744,N_24670,N_24867);
nor UO_2745 (O_2745,N_24699,N_24882);
xor UO_2746 (O_2746,N_24793,N_24582);
nor UO_2747 (O_2747,N_24558,N_24985);
nand UO_2748 (O_2748,N_24702,N_24561);
and UO_2749 (O_2749,N_24817,N_24985);
nand UO_2750 (O_2750,N_24514,N_24665);
nor UO_2751 (O_2751,N_24678,N_24600);
xor UO_2752 (O_2752,N_24577,N_24972);
or UO_2753 (O_2753,N_24581,N_24651);
and UO_2754 (O_2754,N_24575,N_24503);
xor UO_2755 (O_2755,N_24556,N_24584);
nand UO_2756 (O_2756,N_24738,N_24721);
or UO_2757 (O_2757,N_24790,N_24872);
and UO_2758 (O_2758,N_24573,N_24838);
nand UO_2759 (O_2759,N_24933,N_24513);
and UO_2760 (O_2760,N_24504,N_24962);
nand UO_2761 (O_2761,N_24729,N_24634);
nand UO_2762 (O_2762,N_24636,N_24846);
nand UO_2763 (O_2763,N_24659,N_24743);
and UO_2764 (O_2764,N_24941,N_24592);
xnor UO_2765 (O_2765,N_24973,N_24980);
xor UO_2766 (O_2766,N_24531,N_24834);
and UO_2767 (O_2767,N_24974,N_24640);
xnor UO_2768 (O_2768,N_24738,N_24952);
and UO_2769 (O_2769,N_24930,N_24682);
xnor UO_2770 (O_2770,N_24500,N_24876);
or UO_2771 (O_2771,N_24757,N_24809);
and UO_2772 (O_2772,N_24731,N_24912);
or UO_2773 (O_2773,N_24880,N_24510);
and UO_2774 (O_2774,N_24748,N_24774);
nor UO_2775 (O_2775,N_24877,N_24743);
and UO_2776 (O_2776,N_24830,N_24719);
nor UO_2777 (O_2777,N_24658,N_24982);
nand UO_2778 (O_2778,N_24925,N_24617);
nand UO_2779 (O_2779,N_24512,N_24526);
xor UO_2780 (O_2780,N_24810,N_24912);
or UO_2781 (O_2781,N_24908,N_24573);
xor UO_2782 (O_2782,N_24980,N_24910);
xnor UO_2783 (O_2783,N_24853,N_24568);
nand UO_2784 (O_2784,N_24907,N_24894);
nor UO_2785 (O_2785,N_24927,N_24736);
nand UO_2786 (O_2786,N_24624,N_24767);
xor UO_2787 (O_2787,N_24551,N_24723);
nor UO_2788 (O_2788,N_24946,N_24702);
xnor UO_2789 (O_2789,N_24855,N_24770);
and UO_2790 (O_2790,N_24776,N_24872);
xor UO_2791 (O_2791,N_24877,N_24695);
nor UO_2792 (O_2792,N_24680,N_24670);
xor UO_2793 (O_2793,N_24937,N_24721);
nand UO_2794 (O_2794,N_24712,N_24970);
and UO_2795 (O_2795,N_24596,N_24684);
nor UO_2796 (O_2796,N_24582,N_24533);
or UO_2797 (O_2797,N_24986,N_24796);
and UO_2798 (O_2798,N_24810,N_24654);
nand UO_2799 (O_2799,N_24923,N_24565);
and UO_2800 (O_2800,N_24882,N_24598);
and UO_2801 (O_2801,N_24983,N_24525);
nand UO_2802 (O_2802,N_24562,N_24839);
nand UO_2803 (O_2803,N_24653,N_24981);
nor UO_2804 (O_2804,N_24719,N_24814);
or UO_2805 (O_2805,N_24693,N_24711);
nor UO_2806 (O_2806,N_24548,N_24957);
or UO_2807 (O_2807,N_24656,N_24619);
and UO_2808 (O_2808,N_24692,N_24775);
and UO_2809 (O_2809,N_24628,N_24537);
nand UO_2810 (O_2810,N_24623,N_24800);
or UO_2811 (O_2811,N_24962,N_24822);
or UO_2812 (O_2812,N_24890,N_24516);
nor UO_2813 (O_2813,N_24897,N_24797);
or UO_2814 (O_2814,N_24670,N_24781);
or UO_2815 (O_2815,N_24952,N_24653);
xor UO_2816 (O_2816,N_24530,N_24654);
nor UO_2817 (O_2817,N_24748,N_24510);
nor UO_2818 (O_2818,N_24550,N_24695);
nand UO_2819 (O_2819,N_24635,N_24876);
nand UO_2820 (O_2820,N_24877,N_24677);
nand UO_2821 (O_2821,N_24658,N_24630);
nor UO_2822 (O_2822,N_24970,N_24586);
xor UO_2823 (O_2823,N_24685,N_24954);
nor UO_2824 (O_2824,N_24543,N_24573);
nand UO_2825 (O_2825,N_24615,N_24966);
nand UO_2826 (O_2826,N_24555,N_24758);
or UO_2827 (O_2827,N_24867,N_24600);
xor UO_2828 (O_2828,N_24727,N_24708);
or UO_2829 (O_2829,N_24785,N_24793);
nor UO_2830 (O_2830,N_24888,N_24719);
nor UO_2831 (O_2831,N_24579,N_24835);
and UO_2832 (O_2832,N_24652,N_24762);
and UO_2833 (O_2833,N_24671,N_24642);
xnor UO_2834 (O_2834,N_24862,N_24638);
xor UO_2835 (O_2835,N_24955,N_24916);
and UO_2836 (O_2836,N_24829,N_24754);
or UO_2837 (O_2837,N_24770,N_24726);
xnor UO_2838 (O_2838,N_24589,N_24652);
xor UO_2839 (O_2839,N_24733,N_24799);
or UO_2840 (O_2840,N_24634,N_24757);
and UO_2841 (O_2841,N_24869,N_24724);
nand UO_2842 (O_2842,N_24536,N_24750);
or UO_2843 (O_2843,N_24592,N_24738);
nand UO_2844 (O_2844,N_24593,N_24837);
nand UO_2845 (O_2845,N_24681,N_24898);
and UO_2846 (O_2846,N_24589,N_24731);
or UO_2847 (O_2847,N_24735,N_24717);
xnor UO_2848 (O_2848,N_24527,N_24853);
or UO_2849 (O_2849,N_24517,N_24608);
or UO_2850 (O_2850,N_24802,N_24626);
nor UO_2851 (O_2851,N_24591,N_24892);
xnor UO_2852 (O_2852,N_24643,N_24952);
nor UO_2853 (O_2853,N_24937,N_24897);
nor UO_2854 (O_2854,N_24812,N_24545);
nand UO_2855 (O_2855,N_24972,N_24609);
xnor UO_2856 (O_2856,N_24705,N_24930);
xor UO_2857 (O_2857,N_24607,N_24694);
or UO_2858 (O_2858,N_24968,N_24888);
nand UO_2859 (O_2859,N_24746,N_24590);
and UO_2860 (O_2860,N_24870,N_24710);
nor UO_2861 (O_2861,N_24797,N_24746);
nor UO_2862 (O_2862,N_24951,N_24679);
xor UO_2863 (O_2863,N_24857,N_24802);
xor UO_2864 (O_2864,N_24502,N_24515);
or UO_2865 (O_2865,N_24807,N_24882);
and UO_2866 (O_2866,N_24925,N_24828);
nand UO_2867 (O_2867,N_24850,N_24562);
nor UO_2868 (O_2868,N_24629,N_24553);
nand UO_2869 (O_2869,N_24963,N_24999);
nand UO_2870 (O_2870,N_24900,N_24534);
or UO_2871 (O_2871,N_24783,N_24568);
xor UO_2872 (O_2872,N_24517,N_24600);
xnor UO_2873 (O_2873,N_24679,N_24700);
nor UO_2874 (O_2874,N_24707,N_24940);
nand UO_2875 (O_2875,N_24531,N_24859);
nor UO_2876 (O_2876,N_24670,N_24537);
nor UO_2877 (O_2877,N_24961,N_24631);
and UO_2878 (O_2878,N_24585,N_24902);
xor UO_2879 (O_2879,N_24838,N_24748);
and UO_2880 (O_2880,N_24924,N_24773);
xor UO_2881 (O_2881,N_24522,N_24821);
xnor UO_2882 (O_2882,N_24969,N_24997);
or UO_2883 (O_2883,N_24809,N_24693);
nand UO_2884 (O_2884,N_24596,N_24724);
and UO_2885 (O_2885,N_24646,N_24566);
or UO_2886 (O_2886,N_24875,N_24585);
nand UO_2887 (O_2887,N_24609,N_24587);
nor UO_2888 (O_2888,N_24581,N_24689);
or UO_2889 (O_2889,N_24721,N_24643);
or UO_2890 (O_2890,N_24783,N_24778);
nand UO_2891 (O_2891,N_24926,N_24776);
nor UO_2892 (O_2892,N_24893,N_24510);
or UO_2893 (O_2893,N_24592,N_24617);
and UO_2894 (O_2894,N_24820,N_24707);
or UO_2895 (O_2895,N_24857,N_24626);
and UO_2896 (O_2896,N_24568,N_24605);
xnor UO_2897 (O_2897,N_24878,N_24663);
nor UO_2898 (O_2898,N_24915,N_24618);
xnor UO_2899 (O_2899,N_24863,N_24989);
xnor UO_2900 (O_2900,N_24506,N_24976);
and UO_2901 (O_2901,N_24649,N_24690);
xor UO_2902 (O_2902,N_24996,N_24610);
xnor UO_2903 (O_2903,N_24893,N_24745);
nand UO_2904 (O_2904,N_24716,N_24882);
nand UO_2905 (O_2905,N_24850,N_24613);
or UO_2906 (O_2906,N_24896,N_24613);
or UO_2907 (O_2907,N_24712,N_24730);
nand UO_2908 (O_2908,N_24814,N_24974);
nand UO_2909 (O_2909,N_24761,N_24977);
xor UO_2910 (O_2910,N_24886,N_24708);
or UO_2911 (O_2911,N_24544,N_24516);
and UO_2912 (O_2912,N_24938,N_24685);
and UO_2913 (O_2913,N_24948,N_24858);
nor UO_2914 (O_2914,N_24884,N_24928);
nand UO_2915 (O_2915,N_24675,N_24867);
or UO_2916 (O_2916,N_24503,N_24972);
xnor UO_2917 (O_2917,N_24732,N_24726);
nand UO_2918 (O_2918,N_24789,N_24733);
nor UO_2919 (O_2919,N_24542,N_24569);
xnor UO_2920 (O_2920,N_24962,N_24890);
nand UO_2921 (O_2921,N_24964,N_24914);
nand UO_2922 (O_2922,N_24657,N_24762);
or UO_2923 (O_2923,N_24897,N_24675);
and UO_2924 (O_2924,N_24955,N_24867);
and UO_2925 (O_2925,N_24619,N_24628);
or UO_2926 (O_2926,N_24739,N_24512);
xnor UO_2927 (O_2927,N_24557,N_24855);
and UO_2928 (O_2928,N_24822,N_24570);
nor UO_2929 (O_2929,N_24566,N_24823);
or UO_2930 (O_2930,N_24965,N_24697);
or UO_2931 (O_2931,N_24632,N_24543);
or UO_2932 (O_2932,N_24672,N_24735);
and UO_2933 (O_2933,N_24739,N_24800);
nand UO_2934 (O_2934,N_24796,N_24932);
and UO_2935 (O_2935,N_24910,N_24945);
and UO_2936 (O_2936,N_24799,N_24973);
nand UO_2937 (O_2937,N_24648,N_24737);
and UO_2938 (O_2938,N_24979,N_24636);
or UO_2939 (O_2939,N_24737,N_24956);
nor UO_2940 (O_2940,N_24668,N_24903);
or UO_2941 (O_2941,N_24633,N_24879);
nor UO_2942 (O_2942,N_24975,N_24957);
or UO_2943 (O_2943,N_24871,N_24873);
nor UO_2944 (O_2944,N_24719,N_24802);
or UO_2945 (O_2945,N_24729,N_24813);
xnor UO_2946 (O_2946,N_24565,N_24793);
xor UO_2947 (O_2947,N_24511,N_24805);
nor UO_2948 (O_2948,N_24626,N_24664);
and UO_2949 (O_2949,N_24766,N_24642);
xor UO_2950 (O_2950,N_24839,N_24695);
and UO_2951 (O_2951,N_24774,N_24969);
nor UO_2952 (O_2952,N_24990,N_24867);
or UO_2953 (O_2953,N_24985,N_24518);
and UO_2954 (O_2954,N_24879,N_24740);
xnor UO_2955 (O_2955,N_24881,N_24951);
xor UO_2956 (O_2956,N_24851,N_24703);
nor UO_2957 (O_2957,N_24535,N_24657);
and UO_2958 (O_2958,N_24713,N_24502);
and UO_2959 (O_2959,N_24923,N_24916);
or UO_2960 (O_2960,N_24585,N_24680);
nand UO_2961 (O_2961,N_24732,N_24846);
and UO_2962 (O_2962,N_24564,N_24557);
and UO_2963 (O_2963,N_24593,N_24680);
or UO_2964 (O_2964,N_24509,N_24650);
and UO_2965 (O_2965,N_24874,N_24716);
or UO_2966 (O_2966,N_24725,N_24994);
and UO_2967 (O_2967,N_24969,N_24933);
xnor UO_2968 (O_2968,N_24924,N_24951);
nand UO_2969 (O_2969,N_24995,N_24868);
and UO_2970 (O_2970,N_24538,N_24705);
and UO_2971 (O_2971,N_24956,N_24927);
nor UO_2972 (O_2972,N_24512,N_24735);
or UO_2973 (O_2973,N_24749,N_24818);
xor UO_2974 (O_2974,N_24963,N_24552);
and UO_2975 (O_2975,N_24784,N_24939);
nor UO_2976 (O_2976,N_24826,N_24793);
or UO_2977 (O_2977,N_24936,N_24930);
nand UO_2978 (O_2978,N_24674,N_24821);
or UO_2979 (O_2979,N_24694,N_24664);
or UO_2980 (O_2980,N_24659,N_24626);
or UO_2981 (O_2981,N_24832,N_24500);
xnor UO_2982 (O_2982,N_24646,N_24813);
and UO_2983 (O_2983,N_24816,N_24917);
nand UO_2984 (O_2984,N_24539,N_24737);
xor UO_2985 (O_2985,N_24920,N_24597);
or UO_2986 (O_2986,N_24732,N_24570);
and UO_2987 (O_2987,N_24635,N_24713);
nor UO_2988 (O_2988,N_24743,N_24739);
nor UO_2989 (O_2989,N_24597,N_24889);
xor UO_2990 (O_2990,N_24745,N_24792);
nor UO_2991 (O_2991,N_24772,N_24902);
nor UO_2992 (O_2992,N_24967,N_24544);
and UO_2993 (O_2993,N_24679,N_24759);
nand UO_2994 (O_2994,N_24714,N_24824);
nor UO_2995 (O_2995,N_24860,N_24624);
and UO_2996 (O_2996,N_24636,N_24835);
and UO_2997 (O_2997,N_24707,N_24728);
xnor UO_2998 (O_2998,N_24911,N_24605);
nor UO_2999 (O_2999,N_24999,N_24644);
endmodule