module basic_2500_25000_3000_40_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_554,In_2159);
or U1 (N_1,In_701,In_1931);
and U2 (N_2,In_911,In_2100);
and U3 (N_3,In_1677,In_797);
or U4 (N_4,In_1903,In_920);
nor U5 (N_5,In_591,In_251);
xnor U6 (N_6,In_21,In_418);
xnor U7 (N_7,In_966,In_129);
or U8 (N_8,In_1083,In_412);
and U9 (N_9,In_1587,In_2157);
nor U10 (N_10,In_1375,In_1978);
or U11 (N_11,In_1209,In_531);
nor U12 (N_12,In_1507,In_879);
or U13 (N_13,In_1013,In_803);
xnor U14 (N_14,In_700,In_115);
xnor U15 (N_15,In_2282,In_760);
nor U16 (N_16,In_465,In_1848);
nand U17 (N_17,In_961,In_1455);
and U18 (N_18,In_1658,In_271);
nand U19 (N_19,In_533,In_2148);
nand U20 (N_20,In_1258,In_854);
nand U21 (N_21,In_1488,In_574);
nor U22 (N_22,In_315,In_1502);
nand U23 (N_23,In_583,In_1065);
and U24 (N_24,In_990,In_1392);
or U25 (N_25,In_824,In_1665);
nand U26 (N_26,In_2306,In_1726);
and U27 (N_27,In_576,In_94);
xor U28 (N_28,In_11,In_1996);
nor U29 (N_29,In_681,In_230);
or U30 (N_30,In_1590,In_1128);
nor U31 (N_31,In_2010,In_643);
nor U32 (N_32,In_114,In_112);
or U33 (N_33,In_352,In_651);
nand U34 (N_34,In_1181,In_1780);
xor U35 (N_35,In_2228,In_620);
nand U36 (N_36,In_1490,In_1845);
nor U37 (N_37,In_1205,In_625);
nor U38 (N_38,In_2024,In_479);
xnor U39 (N_39,In_1698,In_1149);
and U40 (N_40,In_28,In_214);
nand U41 (N_41,In_227,In_2383);
nor U42 (N_42,In_798,In_1116);
or U43 (N_43,In_1480,In_424);
nand U44 (N_44,In_229,In_914);
or U45 (N_45,In_567,In_1654);
and U46 (N_46,In_2465,In_1496);
nand U47 (N_47,In_2393,In_2366);
or U48 (N_48,In_111,In_497);
and U49 (N_49,In_1533,In_1132);
nor U50 (N_50,In_1262,In_551);
and U51 (N_51,In_181,In_847);
nand U52 (N_52,In_2341,In_1023);
and U53 (N_53,In_516,In_718);
nor U54 (N_54,In_1693,In_663);
or U55 (N_55,In_239,In_2074);
nor U56 (N_56,In_1971,In_2006);
or U57 (N_57,In_1439,In_864);
nor U58 (N_58,In_2063,In_278);
nor U59 (N_59,In_2078,In_204);
nor U60 (N_60,In_811,In_2057);
or U61 (N_61,In_834,In_1521);
nand U62 (N_62,In_439,In_1112);
nor U63 (N_63,In_1129,In_1619);
nor U64 (N_64,In_2446,In_1454);
xor U65 (N_65,In_120,In_364);
nor U66 (N_66,In_1236,In_117);
nand U67 (N_67,In_1611,In_2033);
xor U68 (N_68,In_1015,In_1057);
xor U69 (N_69,In_637,In_664);
nor U70 (N_70,In_691,In_2182);
xor U71 (N_71,In_1373,In_746);
and U72 (N_72,In_1605,In_1636);
and U73 (N_73,In_1846,In_2233);
and U74 (N_74,In_1610,In_1667);
and U75 (N_75,In_279,In_130);
xnor U76 (N_76,In_897,In_585);
or U77 (N_77,In_2072,In_403);
nand U78 (N_78,In_2092,In_603);
xor U79 (N_79,In_1124,In_1643);
and U80 (N_80,In_2187,In_1855);
or U81 (N_81,In_2002,In_501);
nand U82 (N_82,In_1223,In_778);
xnor U83 (N_83,In_878,In_1084);
nor U84 (N_84,In_1680,In_1456);
xor U85 (N_85,In_2039,In_1625);
and U86 (N_86,In_1609,In_1301);
or U87 (N_87,In_2189,In_2464);
or U88 (N_88,In_2125,In_1305);
or U89 (N_89,In_2018,In_1442);
or U90 (N_90,In_432,In_674);
or U91 (N_91,In_816,In_50);
xor U92 (N_92,In_155,In_1217);
nand U93 (N_93,In_264,In_2376);
nand U94 (N_94,In_2483,In_578);
and U95 (N_95,In_869,In_1261);
or U96 (N_96,In_1429,In_517);
or U97 (N_97,In_1140,In_1346);
or U98 (N_98,In_571,In_17);
or U99 (N_99,In_2403,In_55);
nor U100 (N_100,In_1230,In_1661);
and U101 (N_101,In_893,In_132);
and U102 (N_102,In_2338,In_2008);
xnor U103 (N_103,In_1436,In_1806);
xnor U104 (N_104,In_2045,In_846);
or U105 (N_105,In_2271,In_431);
or U106 (N_106,In_174,In_1813);
nand U107 (N_107,In_1354,In_493);
nor U108 (N_108,In_2242,In_187);
nand U109 (N_109,In_40,In_2067);
or U110 (N_110,In_1544,In_225);
xnor U111 (N_111,In_324,In_286);
xnor U112 (N_112,In_1670,In_1341);
or U113 (N_113,In_2384,In_1127);
nand U114 (N_114,In_85,In_825);
nor U115 (N_115,In_548,In_1268);
and U116 (N_116,In_650,In_604);
and U117 (N_117,In_13,In_1842);
nor U118 (N_118,In_782,In_1561);
xor U119 (N_119,In_1388,In_2236);
or U120 (N_120,In_1571,In_1830);
nand U121 (N_121,In_447,In_581);
and U122 (N_122,In_858,In_1159);
and U123 (N_123,In_241,In_1434);
and U124 (N_124,In_175,In_290);
nand U125 (N_125,In_1486,In_1540);
xor U126 (N_126,In_526,In_1107);
xor U127 (N_127,In_1196,In_1990);
or U128 (N_128,In_2119,In_713);
and U129 (N_129,In_2268,In_1448);
xnor U130 (N_130,In_1071,In_2489);
nor U131 (N_131,In_1326,In_568);
xnor U132 (N_132,In_359,In_1573);
nand U133 (N_133,In_2053,In_1534);
nand U134 (N_134,In_1051,In_265);
or U135 (N_135,In_894,In_1225);
or U136 (N_136,In_2354,In_1130);
nand U137 (N_137,In_455,In_2260);
or U138 (N_138,In_2052,In_2280);
or U139 (N_139,In_92,In_1902);
xor U140 (N_140,In_304,In_889);
xor U141 (N_141,In_274,In_1515);
nand U142 (N_142,In_250,In_1936);
and U143 (N_143,In_1098,In_2192);
nand U144 (N_144,In_940,In_1954);
and U145 (N_145,In_610,In_228);
xor U146 (N_146,In_221,In_1001);
or U147 (N_147,In_2443,In_1361);
xnor U148 (N_148,In_950,In_1745);
xor U149 (N_149,In_2196,In_99);
nor U150 (N_150,In_440,In_1905);
and U151 (N_151,In_745,In_2162);
xor U152 (N_152,In_2474,In_1946);
or U153 (N_153,In_1061,In_2479);
or U154 (N_154,In_2205,In_464);
and U155 (N_155,In_2040,In_758);
nor U156 (N_156,In_1141,In_1876);
nand U157 (N_157,In_957,In_636);
nor U158 (N_158,In_2396,In_1912);
and U159 (N_159,In_633,In_618);
and U160 (N_160,In_495,In_425);
nand U161 (N_161,In_337,In_1761);
nand U162 (N_162,In_456,In_457);
and U163 (N_163,In_1329,In_1694);
nor U164 (N_164,In_329,In_1079);
nand U165 (N_165,In_2218,In_1401);
nor U166 (N_166,In_1073,In_1788);
xnor U167 (N_167,In_1920,In_1245);
and U168 (N_168,In_2153,In_477);
nor U169 (N_169,In_104,In_923);
or U170 (N_170,In_1606,In_1979);
nand U171 (N_171,In_1198,In_2166);
or U172 (N_172,In_135,In_1569);
nand U173 (N_173,In_2250,In_2031);
xor U174 (N_174,In_1190,In_1741);
or U175 (N_175,In_451,In_371);
nor U176 (N_176,In_1151,In_1046);
and U177 (N_177,In_792,In_1031);
nor U178 (N_178,In_2099,In_396);
nor U179 (N_179,In_1279,In_2324);
nand U180 (N_180,In_116,In_1052);
nor U181 (N_181,In_830,In_689);
xor U182 (N_182,In_1215,In_406);
and U183 (N_183,In_615,In_1019);
xnor U184 (N_184,In_461,In_2232);
nand U185 (N_185,In_960,In_419);
nor U186 (N_186,In_460,In_1782);
and U187 (N_187,In_247,In_109);
nor U188 (N_188,In_1591,In_392);
nand U189 (N_189,In_150,In_1169);
or U190 (N_190,In_1983,In_1438);
and U191 (N_191,In_381,In_781);
and U192 (N_192,In_1468,In_299);
xnor U193 (N_193,In_205,In_2430);
nor U194 (N_194,In_711,In_360);
nand U195 (N_195,In_1459,In_113);
nor U196 (N_196,In_1735,In_2310);
or U197 (N_197,In_269,In_390);
nor U198 (N_198,In_141,In_1150);
and U199 (N_199,In_1075,In_2113);
and U200 (N_200,In_146,In_1288);
and U201 (N_201,In_759,In_2132);
and U202 (N_202,In_833,In_2346);
nand U203 (N_203,In_199,In_1798);
nor U204 (N_204,In_764,In_257);
nor U205 (N_205,In_1030,In_679);
nand U206 (N_206,In_1307,In_1344);
and U207 (N_207,In_1357,In_2358);
nor U208 (N_208,In_2331,In_16);
xor U209 (N_209,In_1481,In_1479);
nand U210 (N_210,In_1405,In_1187);
nand U211 (N_211,In_1148,In_414);
or U212 (N_212,In_2178,In_949);
nor U213 (N_213,In_2284,In_1701);
xor U214 (N_214,In_1688,In_1856);
and U215 (N_215,In_318,In_1418);
xnor U216 (N_216,In_2406,In_1765);
or U217 (N_217,In_2440,In_273);
xnor U218 (N_218,In_918,In_236);
and U219 (N_219,In_1040,In_182);
xnor U220 (N_220,In_1647,In_1387);
nand U221 (N_221,In_2200,In_595);
nand U222 (N_222,In_1663,In_1220);
and U223 (N_223,In_442,In_47);
and U224 (N_224,In_2071,In_1781);
nor U225 (N_225,In_1282,In_165);
nor U226 (N_226,In_906,In_1907);
nor U227 (N_227,In_1547,In_875);
or U228 (N_228,In_1742,In_1968);
and U229 (N_229,In_634,In_993);
nor U230 (N_230,In_1558,In_1672);
xor U231 (N_231,In_1267,In_80);
nor U232 (N_232,In_346,In_487);
and U233 (N_233,In_1944,In_2226);
and U234 (N_234,In_1728,In_2313);
nor U235 (N_235,In_1241,In_2043);
xor U236 (N_236,In_890,In_1212);
and U237 (N_237,In_839,In_1251);
or U238 (N_238,In_1551,In_968);
nand U239 (N_239,In_1458,In_26);
or U240 (N_240,In_89,In_786);
nor U241 (N_241,In_380,In_586);
and U242 (N_242,In_142,In_532);
and U243 (N_243,In_1582,In_1634);
and U244 (N_244,In_123,In_33);
xor U245 (N_245,In_587,In_1003);
and U246 (N_246,In_1592,In_1089);
xor U247 (N_247,In_927,In_802);
xor U248 (N_248,In_2265,In_509);
nand U249 (N_249,In_563,In_812);
nor U250 (N_250,In_1249,In_919);
nand U251 (N_251,In_2266,In_1312);
xor U252 (N_252,In_1419,In_668);
and U253 (N_253,In_1376,In_874);
nor U254 (N_254,In_1064,In_156);
or U255 (N_255,In_964,In_1202);
nor U256 (N_256,In_1601,In_1185);
xnor U257 (N_257,In_606,In_2357);
nand U258 (N_258,In_1675,In_865);
nor U259 (N_259,In_1988,In_1894);
or U260 (N_260,In_1424,In_2272);
nor U261 (N_261,In_2229,In_810);
nand U262 (N_262,In_900,In_794);
nor U263 (N_263,In_952,In_1348);
or U264 (N_264,In_1340,In_1886);
and U265 (N_265,In_564,In_1171);
nor U266 (N_266,In_755,In_1254);
and U267 (N_267,In_1033,In_1519);
nor U268 (N_268,In_322,In_2134);
or U269 (N_269,In_1325,In_2296);
or U270 (N_270,In_1981,In_2077);
xnor U271 (N_271,In_1280,In_1412);
nor U272 (N_272,In_275,In_1914);
xor U273 (N_273,In_1339,In_2257);
or U274 (N_274,In_730,In_1449);
and U275 (N_275,In_2164,In_1685);
and U276 (N_276,In_2442,In_1565);
or U277 (N_277,In_2378,In_1749);
xor U278 (N_278,In_2314,In_492);
or U279 (N_279,In_1952,In_1021);
nor U280 (N_280,In_1633,In_1049);
nor U281 (N_281,In_2254,In_1447);
xor U282 (N_282,In_59,In_632);
nor U283 (N_283,In_2022,In_503);
and U284 (N_284,In_2356,In_1409);
nor U285 (N_285,In_1244,In_2460);
and U286 (N_286,In_1821,In_95);
or U287 (N_287,In_2299,In_1000);
xnor U288 (N_288,In_1531,In_747);
xor U289 (N_289,In_362,In_2351);
nand U290 (N_290,In_32,In_2319);
or U291 (N_291,In_791,In_2434);
or U292 (N_292,In_1650,In_1397);
and U293 (N_293,In_267,In_1602);
xor U294 (N_294,In_2048,In_1702);
xnor U295 (N_295,In_1441,In_262);
nand U296 (N_296,In_627,In_1967);
or U297 (N_297,In_169,In_242);
or U298 (N_298,In_2081,In_1377);
and U299 (N_299,In_774,In_453);
xor U300 (N_300,In_1414,In_1614);
or U301 (N_301,In_1690,In_52);
xnor U302 (N_302,In_703,In_1872);
and U303 (N_303,In_344,In_368);
nor U304 (N_304,In_1485,In_184);
nor U305 (N_305,In_1240,In_356);
and U306 (N_306,In_144,In_1527);
nand U307 (N_307,In_2094,In_829);
or U308 (N_308,In_48,In_1359);
nand U309 (N_309,In_584,In_1482);
xnor U310 (N_310,In_617,In_496);
nand U311 (N_311,In_147,In_1445);
xor U312 (N_312,In_2211,In_2207);
nor U313 (N_313,In_1997,In_1757);
nor U314 (N_314,In_1259,In_1417);
and U315 (N_315,In_1529,In_289);
and U316 (N_316,In_1933,In_2386);
nand U317 (N_317,In_2286,In_2424);
xor U318 (N_318,In_478,In_541);
nor U319 (N_319,In_1469,In_1002);
nand U320 (N_320,In_293,In_1594);
or U321 (N_321,In_1736,In_226);
nor U322 (N_322,In_1186,In_2097);
nor U323 (N_323,In_2120,In_1867);
and U324 (N_324,In_817,In_611);
or U325 (N_325,In_2288,In_385);
nand U326 (N_326,In_1777,In_410);
nor U327 (N_327,In_291,In_1972);
or U328 (N_328,In_671,In_1957);
xnor U329 (N_329,In_69,In_1564);
xor U330 (N_330,In_119,In_2297);
nand U331 (N_331,In_1134,In_849);
or U332 (N_332,In_300,In_306);
xnor U333 (N_333,In_305,In_167);
nand U334 (N_334,In_2420,In_612);
nor U335 (N_335,In_1165,In_378);
or U336 (N_336,In_2064,In_2124);
xor U337 (N_337,In_766,In_2234);
nand U338 (N_338,In_558,In_107);
or U339 (N_339,In_312,In_1353);
nand U340 (N_340,In_539,In_805);
or U341 (N_341,In_2075,In_892);
xor U342 (N_342,In_105,In_2397);
xor U343 (N_343,In_1380,In_1809);
nor U344 (N_344,In_692,In_943);
and U345 (N_345,In_1560,In_498);
xor U346 (N_346,In_1315,In_1404);
nand U347 (N_347,In_1110,In_789);
and U348 (N_348,In_1992,In_515);
xnor U349 (N_349,In_1466,In_1101);
nand U350 (N_350,In_2047,In_2417);
nand U351 (N_351,In_547,In_1960);
nor U352 (N_352,In_139,In_2385);
nor U353 (N_353,In_25,In_2432);
and U354 (N_354,In_1877,In_835);
and U355 (N_355,In_308,In_1970);
xnor U356 (N_356,In_1617,In_1657);
xnor U357 (N_357,In_2199,In_1965);
nand U358 (N_358,In_2410,In_969);
and U359 (N_359,In_423,In_1508);
or U360 (N_360,In_1514,In_1007);
and U361 (N_361,In_2051,In_720);
and U362 (N_362,In_1584,In_34);
nor U363 (N_363,In_46,In_2300);
nor U364 (N_364,In_2412,In_2058);
and U365 (N_365,In_1264,In_1208);
and U366 (N_366,In_1950,In_288);
xor U367 (N_367,In_1776,In_1382);
nor U368 (N_368,In_1498,In_2359);
or U369 (N_369,In_1369,In_2315);
or U370 (N_370,In_1801,In_1398);
and U371 (N_371,In_1752,In_1273);
xor U372 (N_372,In_1473,In_232);
nand U373 (N_373,In_446,In_2241);
and U374 (N_374,In_311,In_1520);
xnor U375 (N_375,In_697,In_215);
nor U376 (N_376,In_1281,In_832);
and U377 (N_377,In_2170,In_128);
nand U378 (N_378,In_2088,In_276);
nand U379 (N_379,In_1308,In_1106);
xnor U380 (N_380,In_1836,In_1495);
xor U381 (N_381,In_2144,In_2418);
or U382 (N_382,In_1389,In_2289);
xnor U383 (N_383,In_1006,In_2348);
xor U384 (N_384,In_913,In_1743);
and U385 (N_385,In_1464,In_1216);
and U386 (N_386,In_601,In_2447);
or U387 (N_387,In_282,In_2405);
and U388 (N_388,In_2480,In_1088);
nand U389 (N_389,In_1526,In_787);
and U390 (N_390,In_1095,In_813);
nor U391 (N_391,In_684,In_389);
and U392 (N_392,In_14,In_1969);
nor U393 (N_393,In_605,In_669);
nor U394 (N_394,In_1704,In_1713);
and U395 (N_395,In_1618,In_1093);
and U396 (N_396,In_482,In_192);
nor U397 (N_397,In_2353,In_928);
nor U398 (N_398,In_871,In_1717);
nor U399 (N_399,In_363,In_77);
nand U400 (N_400,In_1005,In_2290);
nor U401 (N_401,In_1627,In_770);
xnor U402 (N_402,In_1916,In_1746);
and U403 (N_403,In_243,In_1452);
or U404 (N_404,In_2334,In_1837);
xnor U405 (N_405,In_856,In_1462);
xnor U406 (N_406,In_153,In_1904);
and U407 (N_407,In_1974,In_1027);
xor U408 (N_408,In_102,In_2013);
or U409 (N_409,In_218,In_2349);
or U410 (N_410,In_145,In_2373);
nand U411 (N_411,In_2374,In_1503);
nand U412 (N_412,In_1237,In_866);
or U413 (N_413,In_1906,In_1541);
and U414 (N_414,In_799,In_1535);
xor U415 (N_415,In_725,In_1036);
xor U416 (N_416,In_1552,In_1194);
or U417 (N_417,In_249,In_922);
or U418 (N_418,In_1108,In_1949);
or U419 (N_419,In_197,In_1191);
or U420 (N_420,In_1797,In_399);
nor U421 (N_421,In_1980,In_1852);
nand U422 (N_422,In_398,In_1756);
or U423 (N_423,In_596,In_481);
xor U424 (N_424,In_1327,In_722);
xnor U425 (N_425,In_1117,In_74);
nand U426 (N_426,In_2118,In_2150);
and U427 (N_427,In_953,In_1668);
nor U428 (N_428,In_901,In_2050);
and U429 (N_429,In_2302,In_1180);
and U430 (N_430,In_1499,In_1120);
nor U431 (N_431,In_1425,In_1860);
nor U432 (N_432,In_1109,In_2259);
xnor U433 (N_433,In_435,In_1651);
xnor U434 (N_434,In_2247,In_1318);
nand U435 (N_435,In_1440,In_1334);
nand U436 (N_436,In_2176,In_2225);
xnor U437 (N_437,In_1175,In_925);
xnor U438 (N_438,In_2186,In_2491);
nor U439 (N_439,In_2169,In_1343);
or U440 (N_440,In_2437,In_676);
nand U441 (N_441,In_1286,In_1335);
and U442 (N_442,In_640,In_186);
or U443 (N_443,In_1632,In_1391);
xnor U444 (N_444,In_1630,In_1799);
nand U445 (N_445,In_1513,In_653);
or U446 (N_446,In_347,In_1599);
nor U447 (N_447,In_2165,In_1406);
or U448 (N_448,In_1067,In_1697);
xnor U449 (N_449,In_1768,In_194);
nand U450 (N_450,In_1841,In_2311);
and U451 (N_451,In_1638,In_106);
and U452 (N_452,In_2030,In_83);
or U453 (N_453,In_1292,In_31);
or U454 (N_454,In_1719,In_154);
nor U455 (N_455,In_2389,In_220);
nand U456 (N_456,In_1020,In_1200);
nand U457 (N_457,In_741,In_1682);
nand U458 (N_458,In_35,In_1784);
nand U459 (N_459,In_148,In_2401);
nand U460 (N_460,In_608,In_2111);
nand U461 (N_461,In_2012,In_2155);
xnor U462 (N_462,In_1909,In_1825);
and U463 (N_463,In_965,In_499);
nor U464 (N_464,In_724,In_2082);
and U465 (N_465,In_1378,In_1977);
or U466 (N_466,In_62,In_1770);
nand U467 (N_467,In_2476,In_2387);
nand U468 (N_468,In_349,In_2419);
and U469 (N_469,In_1839,In_1060);
xor U470 (N_470,In_639,In_628);
and U471 (N_471,In_24,In_426);
and U472 (N_472,In_1930,In_2275);
and U473 (N_473,In_60,In_1349);
xnor U474 (N_474,In_2453,In_848);
xnor U475 (N_475,In_280,In_2466);
and U476 (N_476,In_2127,In_1966);
xor U477 (N_477,In_2425,In_852);
xnor U478 (N_478,In_1231,In_1161);
xor U479 (N_479,In_2026,In_951);
or U480 (N_480,In_546,In_1707);
nand U481 (N_481,In_2493,In_2168);
nor U482 (N_482,In_1446,In_158);
and U483 (N_483,In_2,In_818);
xnor U484 (N_484,In_1371,In_1358);
and U485 (N_485,In_2347,In_1901);
xnor U486 (N_486,In_710,In_903);
or U487 (N_487,In_1125,In_1577);
nand U488 (N_488,In_2255,In_762);
nand U489 (N_489,In_804,In_2066);
xnor U490 (N_490,In_2038,In_1063);
and U491 (N_491,In_1812,In_127);
xnor U492 (N_492,In_2128,In_1008);
nand U493 (N_493,In_1999,In_1709);
xor U494 (N_494,In_510,In_2216);
or U495 (N_495,In_2364,In_2171);
xor U496 (N_496,In_2339,In_413);
and U497 (N_497,In_1900,In_4);
and U498 (N_498,In_1773,In_2003);
nor U499 (N_499,In_248,In_1879);
or U500 (N_500,In_1314,In_776);
or U501 (N_501,In_1238,In_947);
xnor U502 (N_502,In_1762,In_2046);
nor U503 (N_503,In_1476,In_1131);
xor U504 (N_504,In_659,In_1310);
or U505 (N_505,In_2343,In_2473);
or U506 (N_506,In_342,In_1524);
nor U507 (N_507,In_433,In_82);
nand U508 (N_508,In_1010,In_986);
or U509 (N_509,In_1925,In_2370);
and U510 (N_510,In_962,In_1077);
xnor U511 (N_511,In_1528,In_823);
nand U512 (N_512,In_740,In_428);
and U513 (N_513,In_1309,In_1976);
nor U514 (N_514,In_880,In_2469);
and U515 (N_515,In_989,In_1938);
or U516 (N_516,In_2321,In_544);
xnor U517 (N_517,In_198,In_727);
nand U518 (N_518,In_1228,In_485);
and U519 (N_519,In_2138,In_1684);
nand U520 (N_520,In_726,In_2471);
xor U521 (N_521,In_2151,In_2214);
and U522 (N_522,In_2152,In_559);
xor U523 (N_523,In_838,In_1229);
nand U524 (N_524,In_307,In_1234);
nor U525 (N_525,In_967,In_1162);
nand U526 (N_526,In_562,In_1199);
and U527 (N_527,In_2231,In_2243);
xnor U528 (N_528,In_600,In_1170);
xor U529 (N_529,In_1011,In_2298);
nand U530 (N_530,In_1311,In_945);
nand U531 (N_531,In_383,In_538);
nand U532 (N_532,In_37,In_592);
xnor U533 (N_533,In_886,In_1090);
or U534 (N_534,In_1332,In_1432);
and U535 (N_535,In_707,In_1635);
or U536 (N_536,In_1055,In_118);
nor U537 (N_537,In_2303,In_738);
xor U538 (N_538,In_882,In_2140);
nor U539 (N_539,In_301,In_873);
nor U540 (N_540,In_1700,In_1861);
xor U541 (N_541,In_38,In_891);
or U542 (N_542,In_1274,In_1642);
and U543 (N_543,In_837,In_2021);
nand U544 (N_544,In_2004,In_2457);
and U545 (N_545,In_626,In_2470);
and U546 (N_546,In_1484,In_1622);
nand U547 (N_547,In_330,In_2049);
or U548 (N_548,In_2459,In_160);
nor U549 (N_549,In_1753,In_1082);
xor U550 (N_550,In_1204,In_270);
or U551 (N_551,In_2246,In_334);
or U552 (N_552,In_462,In_377);
or U553 (N_553,In_1953,In_444);
nor U554 (N_554,In_2475,In_808);
or U555 (N_555,In_1631,In_235);
xor U556 (N_556,In_1875,In_1755);
nand U557 (N_557,In_2198,In_699);
and U558 (N_558,In_1430,In_206);
or U559 (N_559,In_1832,In_2485);
nor U560 (N_560,In_1100,In_2014);
nor U561 (N_561,In_619,In_1032);
or U562 (N_562,In_1850,In_589);
nand U563 (N_563,In_790,In_599);
and U564 (N_564,In_1143,In_328);
or U565 (N_565,In_715,In_1475);
nor U566 (N_566,In_490,In_1751);
and U567 (N_567,In_1509,In_472);
nor U568 (N_568,In_2342,In_1022);
and U569 (N_569,In_1539,In_2458);
nand U570 (N_570,In_1786,In_1955);
and U571 (N_571,In_954,In_1750);
nand U572 (N_572,In_1910,In_1119);
or U573 (N_573,In_81,In_895);
or U574 (N_574,In_1648,In_1580);
or U575 (N_575,In_1085,In_2145);
nor U576 (N_576,In_978,In_2495);
or U577 (N_577,In_1295,In_138);
xnor U578 (N_578,In_2454,In_298);
or U579 (N_579,In_2382,In_594);
nand U580 (N_580,In_1686,In_1807);
xnor U581 (N_581,In_845,In_63);
and U582 (N_582,In_1557,In_317);
xor U583 (N_583,In_941,In_1086);
nand U584 (N_584,In_1351,In_36);
nand U585 (N_585,In_463,In_827);
nor U586 (N_586,In_1350,In_1939);
or U587 (N_587,In_1422,In_670);
or U588 (N_588,In_1207,In_2456);
and U589 (N_589,In_974,In_183);
or U590 (N_590,In_1045,In_1862);
and U591 (N_591,In_2037,In_2173);
and U592 (N_592,In_1183,In_2279);
nor U593 (N_593,In_2167,In_1247);
xor U594 (N_594,In_365,In_644);
nand U595 (N_595,In_417,In_2112);
and U596 (N_596,In_2042,In_1028);
nand U597 (N_597,In_2154,In_1290);
or U598 (N_598,In_326,In_2224);
nand U599 (N_599,In_1621,In_121);
and U600 (N_600,In_51,In_168);
or U601 (N_601,In_1926,In_675);
and U602 (N_602,In_1298,In_1714);
nor U603 (N_603,In_1203,In_2015);
nor U604 (N_604,In_1945,In_1608);
nor U605 (N_605,In_887,In_1779);
nand U606 (N_606,In_1050,In_1122);
nor U607 (N_607,In_542,In_706);
and U608 (N_608,In_773,In_87);
or U609 (N_609,In_915,In_658);
and U610 (N_610,In_1004,In_1911);
nand U611 (N_611,In_434,In_545);
xnor U612 (N_612,In_2320,In_1104);
nand U613 (N_613,In_2494,In_2252);
nand U614 (N_614,In_244,In_2490);
nor U615 (N_615,In_217,In_2388);
xnor U616 (N_616,In_1616,In_688);
and U617 (N_617,In_2221,In_1164);
nand U618 (N_618,In_1087,In_1291);
or U619 (N_619,In_302,In_896);
or U620 (N_620,In_2307,In_2395);
or U621 (N_621,In_1177,In_2350);
or U622 (N_622,In_598,In_1623);
nor U623 (N_623,In_1477,In_2371);
nor U624 (N_624,In_2202,In_1710);
and U625 (N_625,In_2484,In_1637);
or U626 (N_626,In_573,N_487);
nor U627 (N_627,N_74,In_2486);
nand U628 (N_628,N_281,N_400);
or U629 (N_629,N_195,In_97);
and U630 (N_630,In_1184,N_84);
or U631 (N_631,N_36,N_273);
and U632 (N_632,In_1785,In_1853);
nor U633 (N_633,In_955,In_1897);
or U634 (N_634,In_1828,In_1330);
nand U635 (N_635,N_535,In_1081);
nand U636 (N_636,N_399,N_119);
xor U637 (N_637,In_795,N_450);
xnor U638 (N_638,In_2444,In_1523);
nand U639 (N_639,In_514,In_382);
nor U640 (N_640,In_1589,In_1029);
and U641 (N_641,In_126,N_243);
and U642 (N_642,N_40,N_567);
and U643 (N_643,In_742,In_751);
nand U644 (N_644,In_1364,N_253);
nand U645 (N_645,N_228,In_1263);
xnor U646 (N_646,N_527,In_500);
and U647 (N_647,N_28,N_390);
or U648 (N_648,In_1385,In_1210);
nand U649 (N_649,N_541,N_537);
nor U650 (N_650,In_246,In_736);
and U651 (N_651,In_931,N_144);
nor U652 (N_652,N_475,In_820);
xnor U653 (N_653,In_1789,In_1817);
nor U654 (N_654,In_7,N_22);
nor U655 (N_655,In_602,In_1306);
xnor U656 (N_656,In_2073,In_938);
nor U657 (N_657,In_100,N_32);
xnor U658 (N_658,In_237,In_45);
xor U659 (N_659,In_857,N_445);
nor U660 (N_660,In_863,In_647);
or U661 (N_661,N_240,In_1705);
nand U662 (N_662,In_1760,In_2184);
and U663 (N_663,In_959,In_694);
nor U664 (N_664,N_266,In_1126);
and U665 (N_665,In_1824,In_2235);
and U666 (N_666,N_470,In_124);
and U667 (N_667,In_2044,In_841);
or U668 (N_668,In_1718,In_2110);
xor U669 (N_669,In_872,In_1054);
nand U670 (N_670,In_1604,N_75);
nor U671 (N_671,In_391,N_424);
nand U672 (N_672,N_47,N_65);
nand U673 (N_673,In_672,In_916);
nand U674 (N_674,In_975,In_1666);
or U675 (N_675,In_409,In_1941);
or U676 (N_676,In_1586,In_1435);
nand U677 (N_677,In_173,N_208);
xnor U678 (N_678,In_140,N_582);
xnor U679 (N_679,N_446,N_161);
nor U680 (N_680,N_421,N_428);
xnor U681 (N_681,In_1596,In_2191);
nand U682 (N_682,In_513,In_2025);
and U683 (N_683,In_2499,In_876);
and U684 (N_684,In_822,N_596);
and U685 (N_685,In_1820,N_554);
nor U686 (N_686,In_1959,N_624);
nor U687 (N_687,In_1989,N_612);
nor U688 (N_688,N_297,In_1416);
or U689 (N_689,In_1266,In_777);
nor U690 (N_690,In_1393,N_66);
xnor U691 (N_691,In_2463,N_13);
xnor U692 (N_692,In_1899,In_19);
nor U693 (N_693,N_175,In_2201);
xor U694 (N_694,In_2143,In_687);
or U695 (N_695,In_88,In_96);
and U696 (N_696,N_210,In_630);
and U697 (N_697,N_447,N_29);
or U698 (N_698,N_418,In_924);
nand U699 (N_699,In_468,In_2245);
or U700 (N_700,N_62,In_454);
and U701 (N_701,N_443,In_1814);
nand U702 (N_702,N_511,In_702);
and U703 (N_703,N_518,In_2076);
or U704 (N_704,In_991,In_320);
nand U705 (N_705,In_1218,N_255);
and U706 (N_706,In_946,In_401);
nor U707 (N_707,N_335,In_1948);
or U708 (N_708,In_575,In_775);
nor U709 (N_709,N_101,N_285);
nand U710 (N_710,N_560,In_645);
and U711 (N_711,In_2123,In_1864);
nand U712 (N_712,N_482,N_153);
nor U713 (N_713,In_261,In_1068);
nor U714 (N_714,N_211,N_152);
or U715 (N_715,In_384,In_367);
and U716 (N_716,N_360,In_2482);
xnor U717 (N_717,In_2109,In_1868);
nand U718 (N_718,In_2365,N_381);
xor U719 (N_719,In_1849,N_486);
xnor U720 (N_720,N_455,In_860);
nand U721 (N_721,In_1166,In_609);
and U722 (N_722,N_603,In_2415);
xnor U723 (N_723,N_5,In_1581);
xor U724 (N_724,In_616,In_1320);
nand U725 (N_725,In_753,In_549);
or U726 (N_726,In_1835,In_2093);
xnor U727 (N_727,In_843,In_1878);
or U728 (N_728,In_2427,In_1744);
nand U729 (N_729,N_107,In_2360);
nor U730 (N_730,In_1211,In_157);
or U731 (N_731,In_1940,N_140);
or U732 (N_732,In_1411,In_193);
nand U733 (N_733,N_71,In_2114);
xnor U734 (N_734,In_1094,In_622);
and U735 (N_735,In_1347,In_2305);
or U736 (N_736,N_557,N_561);
nand U737 (N_737,N_224,In_86);
or U738 (N_738,N_367,In_486);
and U739 (N_739,In_1407,In_1870);
nor U740 (N_740,N_186,N_11);
and U741 (N_741,N_507,In_2102);
nor U742 (N_742,In_552,In_1711);
and U743 (N_743,N_597,N_383);
and U744 (N_744,N_415,In_397);
nor U745 (N_745,In_550,In_1958);
or U746 (N_746,In_277,N_307);
nor U747 (N_747,In_2253,In_883);
or U748 (N_748,N_436,N_478);
and U749 (N_749,In_2065,In_313);
and U750 (N_750,In_2029,In_765);
or U751 (N_751,In_79,N_198);
xnor U752 (N_752,In_540,In_1731);
and U753 (N_753,In_569,N_357);
or U754 (N_754,N_324,N_179);
xor U755 (N_755,In_801,N_112);
nor U756 (N_756,N_310,In_535);
and U757 (N_757,In_2263,In_2183);
xnor U758 (N_758,N_389,In_1739);
nand U759 (N_759,In_370,N_509);
and U760 (N_760,N_607,In_164);
or U761 (N_761,In_2269,In_1778);
or U762 (N_762,In_2344,In_1646);
or U763 (N_763,N_236,In_1792);
and U764 (N_764,In_1155,In_1555);
and U765 (N_765,In_1943,In_788);
xnor U766 (N_766,In_357,In_1138);
and U767 (N_767,In_885,N_239);
and U768 (N_768,In_2210,In_998);
nor U769 (N_769,N_578,In_18);
and U770 (N_770,In_739,In_2011);
and U771 (N_771,N_160,In_963);
nand U772 (N_772,In_1922,In_2107);
nor U773 (N_773,In_1908,N_336);
nand U774 (N_774,In_2292,N_246);
xnor U775 (N_775,In_1384,In_561);
nor U776 (N_776,N_353,N_466);
and U777 (N_777,N_81,In_905);
and U778 (N_778,N_279,In_1024);
or U779 (N_779,N_427,N_591);
xor U780 (N_780,In_984,In_331);
nor U781 (N_781,In_2195,In_1356);
nor U782 (N_782,N_86,In_2133);
or U783 (N_783,In_1365,In_1342);
and U784 (N_784,N_448,In_2276);
and U785 (N_785,In_1802,In_101);
xnor U786 (N_786,In_2041,N_177);
or U787 (N_787,N_277,In_2333);
xor U788 (N_788,In_908,In_415);
xnor U789 (N_789,In_2061,In_2105);
and U790 (N_790,In_1866,In_209);
nand U791 (N_791,In_1568,In_2027);
or U792 (N_792,N_373,In_734);
and U793 (N_793,N_370,In_593);
nor U794 (N_794,In_1471,In_2441);
and U795 (N_795,In_1819,In_1201);
or U796 (N_796,In_480,In_566);
nand U797 (N_797,In_8,In_1740);
or U798 (N_798,In_1712,In_210);
xnor U799 (N_799,In_1578,In_1328);
or U800 (N_800,In_404,In_1929);
and U801 (N_801,In_2188,In_2023);
nor U802 (N_802,N_109,In_2098);
nand U803 (N_803,In_2461,In_287);
and U804 (N_804,In_1896,In_1363);
nor U805 (N_805,In_2108,In_429);
and U806 (N_806,In_1296,In_253);
nor U807 (N_807,In_1396,In_1559);
nand U808 (N_808,N_69,In_369);
xor U809 (N_809,N_476,In_1562);
nor U810 (N_810,In_350,N_467);
nor U811 (N_811,N_407,N_282);
or U812 (N_812,In_988,In_1146);
or U813 (N_813,N_227,In_1829);
or U814 (N_814,In_1722,N_141);
nand U815 (N_815,N_380,N_245);
nor U816 (N_816,In_1383,In_2323);
nand U817 (N_817,N_20,In_2498);
nand U818 (N_818,N_150,N_120);
nor U819 (N_819,In_828,N_35);
and U820 (N_820,N_213,In_649);
or U821 (N_821,In_907,In_1679);
nand U822 (N_822,In_1891,N_406);
nor U823 (N_823,In_2361,In_2091);
nor U824 (N_824,In_2237,In_917);
nand U825 (N_825,In_170,N_519);
nor U826 (N_826,In_1355,In_2089);
or U827 (N_827,In_2209,In_162);
and U828 (N_828,N_572,In_68);
xor U829 (N_829,In_1078,N_404);
nor U830 (N_830,N_376,In_826);
xnor U831 (N_831,In_819,N_465);
xor U832 (N_832,In_807,In_1593);
nor U833 (N_833,In_2194,In_570);
and U834 (N_834,In_1874,N_102);
or U835 (N_835,In_53,N_372);
or U836 (N_836,In_1720,N_449);
and U837 (N_837,In_2267,In_200);
xnor U838 (N_838,In_1808,In_296);
or U839 (N_839,In_1612,In_1009);
xor U840 (N_840,In_1847,N_143);
or U841 (N_841,In_1695,In_333);
nand U842 (N_842,In_1293,N_7);
and U843 (N_843,In_2337,In_769);
xnor U844 (N_844,N_393,N_503);
and U845 (N_845,In_1600,In_2270);
xnor U846 (N_846,In_1641,In_2203);
nor U847 (N_847,In_2326,N_314);
xor U848 (N_848,N_419,In_712);
and U849 (N_849,In_255,In_1656);
nor U850 (N_850,In_520,In_2059);
nand U851 (N_851,In_376,N_480);
xor U852 (N_852,N_133,N_77);
or U853 (N_853,N_21,In_1);
nor U854 (N_854,In_1579,In_1158);
nor U855 (N_855,N_576,In_2492);
nand U856 (N_856,In_266,In_1048);
or U857 (N_857,In_2345,In_1195);
nand U858 (N_858,In_646,In_2019);
nor U859 (N_859,N_510,In_1451);
nor U860 (N_860,N_223,N_375);
or U861 (N_861,In_638,N_562);
xnor U862 (N_862,In_420,N_90);
and U863 (N_863,In_1113,N_87);
and U864 (N_864,In_2034,In_1224);
xnor U865 (N_865,In_263,In_1816);
nor U866 (N_866,N_88,In_1769);
xnor U867 (N_867,In_994,In_2467);
or U868 (N_868,In_2087,N_108);
xor U869 (N_869,In_1649,N_550);
and U870 (N_870,In_1795,In_853);
and U871 (N_871,In_1727,In_870);
and U872 (N_872,In_2135,In_325);
nand U873 (N_873,In_2391,In_1734);
nand U874 (N_874,N_283,In_1834);
and U875 (N_875,In_1213,In_1463);
xnor U876 (N_876,In_1550,N_197);
nand U877 (N_877,N_42,In_2126);
nor U878 (N_878,In_1928,In_2007);
nor U879 (N_879,In_110,N_587);
nor U880 (N_880,In_656,In_1444);
and U881 (N_881,N_350,N_39);
nand U882 (N_882,In_2472,In_2362);
and U883 (N_883,In_2070,In_1074);
and U884 (N_884,In_1260,In_1893);
and U885 (N_885,In_1607,N_565);
or U886 (N_886,In_1595,In_316);
and U887 (N_887,In_654,In_588);
nor U888 (N_888,In_2009,In_466);
xor U889 (N_889,In_151,In_2136);
nor U890 (N_890,In_1729,In_728);
or U891 (N_891,In_761,In_1640);
xor U892 (N_892,N_386,In_1892);
or U893 (N_893,In_1737,N_588);
and U894 (N_894,N_204,In_1689);
nor U895 (N_895,N_452,In_1287);
or U896 (N_896,In_2256,N_278);
nand U897 (N_897,In_652,In_629);
or U898 (N_898,N_432,In_353);
or U899 (N_899,In_5,In_1898);
nand U900 (N_900,In_2431,In_2301);
nand U901 (N_901,N_294,In_2174);
xor U902 (N_902,In_784,N_242);
nand U903 (N_903,In_698,In_1182);
nand U904 (N_904,In_1272,In_624);
or U905 (N_905,N_201,N_70);
xor U906 (N_906,N_458,In_2398);
and U907 (N_907,N_248,N_37);
and U908 (N_908,N_514,In_1935);
or U909 (N_909,In_2239,N_394);
and U910 (N_910,N_49,In_1927);
and U911 (N_911,In_1160,N_440);
nor U912 (N_912,N_520,In_416);
nor U913 (N_913,In_840,N_617);
xnor U914 (N_914,N_99,N_229);
or U915 (N_915,In_1747,N_181);
xor U916 (N_916,N_325,N_231);
or U917 (N_917,In_2197,N_60);
and U918 (N_918,N_493,In_693);
xor U919 (N_919,In_245,N_609);
xnor U920 (N_920,N_185,In_2101);
nor U921 (N_921,In_361,N_599);
nand U922 (N_922,N_199,In_1039);
nor U923 (N_923,In_884,In_2330);
xnor U924 (N_924,In_98,N_540);
nor U925 (N_925,In_997,In_1934);
nor U926 (N_926,N_358,N_9);
and U927 (N_927,In_1173,In_2028);
xnor U928 (N_928,N_530,In_1058);
and U929 (N_929,N_555,In_2309);
and U930 (N_930,N_276,N_291);
nor U931 (N_931,In_1624,In_2212);
xor U932 (N_932,In_1137,In_2095);
or U933 (N_933,N_516,In_1012);
or U934 (N_934,N_408,In_1394);
xnor U935 (N_935,In_1235,In_2287);
xor U936 (N_936,N_422,N_485);
xnor U937 (N_937,In_494,In_690);
nand U938 (N_938,In_1399,In_1652);
nand U939 (N_939,In_1536,In_216);
xnor U940 (N_940,N_524,In_577);
and U941 (N_941,N_365,In_1147);
xor U942 (N_942,In_1826,In_1366);
and U943 (N_943,In_1474,In_785);
nand U944 (N_944,In_285,In_374);
or U945 (N_945,In_556,In_131);
or U946 (N_946,In_2249,In_2449);
or U947 (N_947,N_462,N_352);
xor U948 (N_948,In_202,In_1337);
nor U949 (N_949,In_1133,In_303);
or U950 (N_950,In_2381,In_2177);
and U951 (N_951,N_176,N_63);
nand U952 (N_952,N_346,N_303);
or U953 (N_953,N_337,In_2294);
and U954 (N_954,N_543,In_735);
and U955 (N_955,In_929,In_2141);
xnor U956 (N_956,N_321,N_127);
xnor U957 (N_957,In_529,In_6);
nand U958 (N_958,N_581,In_2327);
nand U959 (N_959,In_1437,In_1153);
nand U960 (N_960,In_771,In_2404);
nand U961 (N_961,In_1034,In_2377);
xnor U962 (N_962,In_518,N_611);
xnor U963 (N_963,In_1549,In_1895);
xnor U964 (N_964,In_2426,In_1111);
xor U965 (N_965,In_1135,N_589);
or U966 (N_966,N_110,In_219);
nand U967 (N_967,In_661,In_159);
xor U968 (N_968,N_417,N_58);
nand U969 (N_969,In_2423,In_527);
nor U970 (N_970,In_1963,In_1510);
nor U971 (N_971,In_768,In_1472);
nand U972 (N_972,In_2413,In_972);
nor U973 (N_973,In_842,In_2264);
xor U974 (N_974,In_408,In_733);
or U975 (N_975,N_474,In_2285);
nand U976 (N_976,N_309,N_489);
nor U977 (N_977,In_2335,N_241);
or U978 (N_978,N_442,In_2277);
nand U979 (N_979,N_61,N_378);
nor U980 (N_980,In_2439,N_111);
nor U981 (N_981,In_341,In_1572);
nand U982 (N_982,In_1313,In_909);
nand U983 (N_983,N_166,In_1163);
nand U984 (N_984,N_67,In_1994);
or U985 (N_985,In_2204,In_178);
nand U986 (N_986,N_225,N_454);
or U987 (N_987,In_2468,In_2147);
nor U988 (N_988,In_597,In_1076);
and U989 (N_989,N_124,N_559);
xor U990 (N_990,In_421,N_93);
and U991 (N_991,In_1793,In_1664);
and U992 (N_992,In_2217,N_45);
nor U993 (N_993,N_202,N_344);
nand U994 (N_994,In_956,N_117);
nor U995 (N_995,N_539,In_932);
nand U996 (N_996,In_1041,N_306);
xor U997 (N_997,In_469,In_258);
xnor U998 (N_998,N_556,In_942);
nor U999 (N_999,In_1487,In_133);
or U1000 (N_1000,In_1732,N_521);
and U1001 (N_1001,In_1303,In_2106);
nand U1002 (N_1002,In_1069,In_2340);
nor U1003 (N_1003,In_1626,In_1167);
or U1004 (N_1004,N_311,In_1331);
nor U1005 (N_1005,In_2158,In_1844);
xnor U1006 (N_1006,In_1395,N_592);
nand U1007 (N_1007,In_1297,In_2367);
and U1008 (N_1008,N_298,In_1858);
nor U1009 (N_1009,In_2304,In_2137);
nor U1010 (N_1010,N_468,In_2139);
xnor U1011 (N_1011,In_2103,In_898);
nor U1012 (N_1012,N_517,N_363);
xnor U1013 (N_1013,In_2477,In_1629);
nand U1014 (N_1014,In_2421,In_2402);
and U1015 (N_1015,N_471,In_779);
nand U1016 (N_1016,In_1803,In_405);
and U1017 (N_1017,N_563,N_558);
or U1018 (N_1018,In_750,N_423);
or U1019 (N_1019,In_2394,N_412);
or U1020 (N_1020,In_1176,N_498);
xnor U1021 (N_1021,In_590,In_476);
or U1022 (N_1022,N_121,In_163);
and U1023 (N_1023,In_1232,N_438);
nand U1024 (N_1024,In_1091,N_593);
nand U1025 (N_1025,N_95,In_467);
nor U1026 (N_1026,N_134,In_2455);
nor U1027 (N_1027,In_543,In_2408);
nor U1028 (N_1028,In_2160,In_231);
nand U1029 (N_1029,In_1144,In_1921);
nor U1030 (N_1030,N_496,In_2390);
and U1031 (N_1031,N_494,In_1615);
and U1032 (N_1032,In_196,N_444);
nand U1033 (N_1033,In_2142,In_2317);
nand U1034 (N_1034,N_608,In_1188);
xor U1035 (N_1035,In_358,In_2005);
or U1036 (N_1036,In_1545,N_54);
and U1037 (N_1037,In_1937,In_1338);
nor U1038 (N_1038,In_763,In_488);
xnor U1039 (N_1039,In_682,In_283);
xnor U1040 (N_1040,In_1639,N_3);
or U1041 (N_1041,N_89,In_2000);
or U1042 (N_1042,In_1823,In_850);
nor U1043 (N_1043,N_145,In_2215);
nand U1044 (N_1044,In_1386,In_1372);
xnor U1045 (N_1045,In_1415,In_238);
nand U1046 (N_1046,In_483,In_1433);
and U1047 (N_1047,N_51,N_484);
and U1048 (N_1048,In_56,In_2400);
nand U1049 (N_1049,In_1461,N_548);
xnor U1050 (N_1050,In_1538,In_2122);
nor U1051 (N_1051,In_1687,In_1239);
xor U1052 (N_1052,In_1453,In_934);
nand U1053 (N_1053,N_105,N_525);
xor U1054 (N_1054,In_557,In_683);
nand U1055 (N_1055,In_877,In_223);
nor U1056 (N_1056,In_1696,In_1080);
and U1057 (N_1057,In_42,N_457);
nor U1058 (N_1058,In_1869,N_187);
nand U1059 (N_1059,N_106,N_247);
xor U1060 (N_1060,N_293,N_613);
and U1061 (N_1061,N_402,In_1253);
and U1062 (N_1062,N_251,In_400);
nand U1063 (N_1063,N_129,In_1804);
nand U1064 (N_1064,In_677,N_6);
nor U1065 (N_1065,In_1374,In_1174);
nand U1066 (N_1066,N_329,In_1103);
nor U1067 (N_1067,In_2193,In_926);
or U1068 (N_1068,In_1532,N_368);
and U1069 (N_1069,N_44,In_1759);
nor U1070 (N_1070,In_655,In_1197);
or U1071 (N_1071,N_180,In_904);
nand U1072 (N_1072,In_375,N_267);
xnor U1073 (N_1073,N_38,In_441);
and U1074 (N_1074,In_1178,In_1408);
xor U1075 (N_1075,In_1865,N_348);
or U1076 (N_1076,In_836,In_2032);
nand U1077 (N_1077,N_0,In_386);
or U1078 (N_1078,N_340,N_605);
or U1079 (N_1079,N_250,N_154);
nor U1080 (N_1080,N_57,In_1888);
xor U1081 (N_1081,In_506,In_489);
nor U1082 (N_1082,In_1525,N_431);
and U1083 (N_1083,In_213,N_583);
nand U1084 (N_1084,In_212,In_474);
nand U1085 (N_1085,In_1370,In_1563);
xor U1086 (N_1086,In_1537,N_286);
nand U1087 (N_1087,N_46,N_506);
nor U1088 (N_1088,In_1443,In_1794);
and U1089 (N_1089,In_793,N_416);
xnor U1090 (N_1090,In_2244,In_678);
or U1091 (N_1091,In_1423,In_1252);
and U1092 (N_1092,In_177,In_1360);
and U1093 (N_1093,In_2104,In_373);
and U1094 (N_1094,In_1767,N_59);
nor U1095 (N_1095,In_1951,In_1506);
and U1096 (N_1096,In_979,In_1319);
xor U1097 (N_1097,N_64,N_300);
and U1098 (N_1098,In_2035,N_534);
or U1099 (N_1099,In_1043,N_545);
nand U1100 (N_1100,In_1644,N_221);
or U1101 (N_1101,N_502,N_499);
or U1102 (N_1102,In_339,N_328);
and U1103 (N_1103,In_1500,In_2329);
xnor U1104 (N_1104,N_501,In_1265);
nand U1105 (N_1105,In_2478,In_1748);
nand U1106 (N_1106,N_25,In_1673);
or U1107 (N_1107,N_490,In_2274);
nor U1108 (N_1108,N_268,In_1838);
nor U1109 (N_1109,In_240,N_397);
nand U1110 (N_1110,In_2322,N_317);
xor U1111 (N_1111,N_580,In_2332);
nand U1112 (N_1112,In_1884,In_507);
nand U1113 (N_1113,N_263,N_79);
nor U1114 (N_1114,In_1270,In_1548);
xnor U1115 (N_1115,In_284,In_1653);
or U1116 (N_1116,N_275,N_547);
nand U1117 (N_1117,In_427,In_1796);
nand U1118 (N_1118,N_254,N_260);
xnor U1119 (N_1119,N_122,In_224);
or U1120 (N_1120,In_673,N_237);
xnor U1121 (N_1121,In_1881,N_526);
or U1122 (N_1122,N_170,N_601);
nor U1123 (N_1123,N_459,In_2278);
xor U1124 (N_1124,In_1708,In_41);
nand U1125 (N_1125,In_1859,In_1070);
nand U1126 (N_1126,In_1233,In_560);
and U1127 (N_1127,In_388,N_341);
and U1128 (N_1128,In_336,In_2068);
and U1129 (N_1129,In_2375,In_2180);
or U1130 (N_1130,N_234,In_2368);
and U1131 (N_1131,N_590,In_2055);
nor U1132 (N_1132,In_958,In_1410);
and U1133 (N_1133,In_44,In_1645);
xnor U1134 (N_1134,In_15,In_2258);
nand U1135 (N_1135,N_296,In_708);
and U1136 (N_1136,In_1683,N_135);
or U1137 (N_1137,In_844,In_1284);
nand U1138 (N_1138,In_297,In_2062);
or U1139 (N_1139,In_528,In_1271);
nand U1140 (N_1140,In_2090,N_30);
nand U1141 (N_1141,In_996,In_70);
nor U1142 (N_1142,In_1554,In_1470);
xor U1143 (N_1143,In_754,In_335);
nor U1144 (N_1144,N_595,In_75);
and U1145 (N_1145,In_666,In_1774);
or U1146 (N_1146,In_631,In_1121);
xnor U1147 (N_1147,In_1427,In_737);
xnor U1148 (N_1148,N_48,N_615);
nor U1149 (N_1149,N_602,In_309);
or U1150 (N_1150,N_100,In_2054);
nand U1151 (N_1151,In_796,N_359);
nand U1152 (N_1152,In_1206,In_2295);
or U1153 (N_1153,In_152,N_414);
xnor U1154 (N_1154,N_83,N_351);
xnor U1155 (N_1155,N_586,N_244);
and U1156 (N_1156,N_410,In_2262);
or U1157 (N_1157,In_523,In_1483);
nand U1158 (N_1158,In_937,In_176);
xor U1159 (N_1159,In_207,N_345);
nor U1160 (N_1160,In_1099,In_1278);
or U1161 (N_1161,In_553,In_1390);
nand U1162 (N_1162,In_1025,In_449);
nor U1163 (N_1163,In_12,In_1256);
xnor U1164 (N_1164,In_1118,N_464);
and U1165 (N_1165,In_525,In_172);
nor U1166 (N_1166,In_2036,In_452);
and U1167 (N_1167,In_921,In_868);
and U1168 (N_1168,In_1699,N_316);
and U1169 (N_1169,In_910,In_1044);
nor U1170 (N_1170,N_171,In_29);
nor U1171 (N_1171,In_2206,In_58);
or U1172 (N_1172,N_43,N_284);
nor U1173 (N_1173,N_262,N_425);
xnor U1174 (N_1174,N_178,In_64);
and U1175 (N_1175,N_463,In_1294);
or U1176 (N_1176,N_23,N_573);
nand U1177 (N_1177,In_1660,N_568);
nand U1178 (N_1178,In_2308,In_1857);
nand U1179 (N_1179,N_257,In_84);
nor U1180 (N_1180,In_260,In_203);
and U1181 (N_1181,In_1097,In_2316);
and U1182 (N_1182,N_104,N_233);
nor U1183 (N_1183,In_2369,In_259);
and U1184 (N_1184,N_295,N_473);
and U1185 (N_1185,N_14,N_203);
or U1186 (N_1186,In_1790,In_234);
and U1187 (N_1187,In_1250,In_122);
nor U1188 (N_1188,In_338,N_151);
or U1189 (N_1189,In_859,In_2312);
nand U1190 (N_1190,In_2433,In_78);
or U1191 (N_1191,In_1428,In_537);
or U1192 (N_1192,In_2407,In_1522);
nor U1193 (N_1193,In_1277,In_1062);
and U1194 (N_1194,In_1248,In_1576);
xnor U1195 (N_1195,N_549,N_137);
xnor U1196 (N_1196,N_610,In_1783);
xor U1197 (N_1197,N_72,In_1542);
nor U1198 (N_1198,In_491,N_392);
or U1199 (N_1199,N_261,N_26);
nand U1200 (N_1200,In_450,N_290);
xor U1201 (N_1201,In_2251,In_1763);
or U1202 (N_1202,In_980,In_1047);
or U1203 (N_1203,In_2392,In_1493);
and U1204 (N_1204,N_552,In_888);
or U1205 (N_1205,In_2416,In_185);
and U1206 (N_1206,In_1403,In_2017);
nand U1207 (N_1207,N_409,In_348);
and U1208 (N_1208,In_2283,N_219);
nor U1209 (N_1209,N_91,N_513);
and U1210 (N_1210,In_971,In_1189);
and U1211 (N_1211,In_1800,N_575);
xor U1212 (N_1212,In_2325,In_459);
nor U1213 (N_1213,N_492,In_1492);
or U1214 (N_1214,In_1923,In_2079);
xnor U1215 (N_1215,In_61,In_1613);
and U1216 (N_1216,N_56,In_343);
and U1217 (N_1217,In_580,In_1494);
or U1218 (N_1218,N_382,In_72);
nor U1219 (N_1219,In_973,In_134);
or U1220 (N_1220,N_585,N_94);
and U1221 (N_1221,In_1889,N_31);
xor U1222 (N_1222,In_502,In_809);
or U1223 (N_1223,In_1017,N_430);
nand U1224 (N_1224,N_115,N_355);
nor U1225 (N_1225,In_2422,In_1681);
and U1226 (N_1226,N_491,In_748);
nor U1227 (N_1227,In_366,In_1715);
xnor U1228 (N_1228,In_2117,In_1105);
xor U1229 (N_1229,In_292,In_2219);
nand U1230 (N_1230,In_1142,N_159);
and U1231 (N_1231,In_565,In_179);
xnor U1232 (N_1232,In_721,N_441);
nor U1233 (N_1233,In_1367,In_1227);
xnor U1234 (N_1234,N_481,In_323);
or U1235 (N_1235,In_1987,N_113);
nor U1236 (N_1236,In_1426,In_1324);
or U1237 (N_1237,In_555,In_1352);
nand U1238 (N_1238,In_1379,N_196);
or U1239 (N_1239,In_319,In_1381);
nand U1240 (N_1240,In_1887,N_53);
nor U1241 (N_1241,In_475,In_1321);
or U1242 (N_1242,In_933,In_743);
or U1243 (N_1243,N_614,In_20);
xor U1244 (N_1244,In_800,In_511);
xnor U1245 (N_1245,In_982,In_1833);
nand U1246 (N_1246,N_434,In_2230);
and U1247 (N_1247,In_2161,N_456);
or U1248 (N_1248,N_435,In_394);
and U1249 (N_1249,In_2163,N_477);
nor U1250 (N_1250,N_873,In_731);
or U1251 (N_1251,In_2411,N_970);
nand U1252 (N_1252,N_791,N_639);
nand U1253 (N_1253,In_2146,N_532);
xnor U1254 (N_1254,N_16,N_342);
xnor U1255 (N_1255,In_536,N_1152);
xnor U1256 (N_1256,In_149,In_936);
xor U1257 (N_1257,In_899,In_254);
or U1258 (N_1258,In_1733,In_2084);
and U1259 (N_1259,N_188,N_798);
or U1260 (N_1260,In_524,N_1177);
nor U1261 (N_1261,N_944,In_723);
nand U1262 (N_1262,N_1033,N_1233);
nand U1263 (N_1263,In_519,N_1175);
and U1264 (N_1264,N_123,N_1027);
or U1265 (N_1265,N_19,N_966);
nand U1266 (N_1266,N_411,In_2429);
or U1267 (N_1267,In_2336,In_1993);
or U1268 (N_1268,N_938,In_1669);
or U1269 (N_1269,N_1147,In_1919);
xnor U1270 (N_1270,In_1575,N_1002);
nor U1271 (N_1271,In_90,N_1082);
nand U1272 (N_1272,In_1400,N_797);
xnor U1273 (N_1273,N_209,In_2115);
nor U1274 (N_1274,In_1805,In_815);
xor U1275 (N_1275,In_1975,In_1289);
nor U1276 (N_1276,In_2261,N_252);
nor U1277 (N_1277,N_156,In_332);
and U1278 (N_1278,In_814,N_542);
nor U1279 (N_1279,In_2080,N_979);
nor U1280 (N_1280,N_1196,In_1603);
and U1281 (N_1281,In_2222,N_1085);
nand U1282 (N_1282,N_727,In_732);
nand U1283 (N_1283,N_943,N_1054);
or U1284 (N_1284,N_1194,In_1192);
nand U1285 (N_1285,N_1060,N_1218);
and U1286 (N_1286,In_1851,N_836);
nand U1287 (N_1287,N_403,N_1017);
or U1288 (N_1288,N_1045,N_714);
xor U1289 (N_1289,N_623,N_1035);
nor U1290 (N_1290,N_1234,N_1224);
and U1291 (N_1291,N_1216,In_1991);
or U1292 (N_1292,N_928,N_1098);
xnor U1293 (N_1293,N_827,In_23);
or U1294 (N_1294,N_778,N_742);
and U1295 (N_1295,N_269,N_265);
xor U1296 (N_1296,N_854,N_751);
or U1297 (N_1297,N_1068,N_671);
xnor U1298 (N_1298,N_777,N_68);
and U1299 (N_1299,N_388,N_880);
nand U1300 (N_1300,In_2372,In_1724);
nand U1301 (N_1301,N_684,N_1003);
nor U1302 (N_1302,N_1171,N_379);
or U1303 (N_1303,N_1136,In_861);
nand U1304 (N_1304,N_749,N_1110);
or U1305 (N_1305,N_192,In_1810);
nor U1306 (N_1306,In_473,N_1090);
nand U1307 (N_1307,N_384,In_2208);
nor U1308 (N_1308,In_2156,N_164);
or U1309 (N_1309,N_844,In_821);
nor U1310 (N_1310,N_12,N_616);
or U1311 (N_1311,N_439,N_1056);
and U1312 (N_1312,In_1123,In_1512);
xor U1313 (N_1313,In_686,In_1368);
nand U1314 (N_1314,N_693,N_788);
xnor U1315 (N_1315,N_1084,In_2399);
or U1316 (N_1316,N_843,N_1005);
nor U1317 (N_1317,N_76,N_677);
nor U1318 (N_1318,N_903,N_1021);
nand U1319 (N_1319,N_1030,N_461);
nor U1320 (N_1320,N_308,N_1248);
or U1321 (N_1321,N_169,N_361);
nand U1322 (N_1322,In_995,In_437);
xnor U1323 (N_1323,N_1225,In_1775);
or U1324 (N_1324,In_1871,N_238);
nand U1325 (N_1325,N_855,N_1126);
and U1326 (N_1326,In_831,In_1973);
nor U1327 (N_1327,In_2481,N_1059);
nor U1328 (N_1328,In_744,In_579);
or U1329 (N_1329,In_161,In_1059);
xnor U1330 (N_1330,N_959,N_579);
nand U1331 (N_1331,In_458,N_879);
nand U1332 (N_1332,N_913,N_782);
and U1333 (N_1333,N_679,N_1151);
xor U1334 (N_1334,N_1228,In_1413);
or U1335 (N_1335,N_987,N_925);
nand U1336 (N_1336,N_200,N_349);
nor U1337 (N_1337,N_810,In_188);
or U1338 (N_1338,In_780,In_2085);
or U1339 (N_1339,N_274,N_1107);
nand U1340 (N_1340,N_839,In_1053);
xnor U1341 (N_1341,N_857,N_222);
or U1342 (N_1342,N_232,N_794);
or U1343 (N_1343,N_694,N_906);
xor U1344 (N_1344,N_1235,N_760);
nand U1345 (N_1345,N_635,N_980);
or U1346 (N_1346,N_1232,N_754);
or U1347 (N_1347,N_1067,In_1402);
nor U1348 (N_1348,N_1018,N_34);
nor U1349 (N_1349,N_748,In_985);
nand U1350 (N_1350,In_930,N_954);
nor U1351 (N_1351,N_962,In_1723);
nor U1352 (N_1352,N_852,N_1001);
xnor U1353 (N_1353,N_1073,N_362);
xnor U1354 (N_1354,N_1181,In_1597);
and U1355 (N_1355,In_2240,In_1691);
or U1356 (N_1356,N_533,In_1168);
or U1357 (N_1357,N_189,In_2227);
nor U1358 (N_1358,In_756,In_0);
or U1359 (N_1359,N_546,N_755);
xor U1360 (N_1360,N_708,N_815);
nor U1361 (N_1361,N_469,In_1787);
and U1362 (N_1362,N_226,N_960);
xnor U1363 (N_1363,N_1172,N_811);
nand U1364 (N_1364,N_1249,In_1323);
or U1365 (N_1365,N_685,In_1827);
xnor U1366 (N_1366,In_1115,N_942);
or U1367 (N_1367,In_1491,In_471);
and U1368 (N_1368,In_281,N_1133);
nand U1369 (N_1369,N_862,N_1185);
xnor U1370 (N_1370,In_1962,N_932);
nand U1371 (N_1371,In_438,In_108);
xor U1372 (N_1372,In_2291,N_1091);
nand U1373 (N_1373,N_320,N_1074);
nand U1374 (N_1374,In_1037,N_765);
or U1375 (N_1375,In_2428,N_771);
nand U1376 (N_1376,N_207,In_1703);
or U1377 (N_1377,In_944,N_1170);
nor U1378 (N_1378,N_1078,In_2248);
xor U1379 (N_1379,N_374,N_538);
and U1380 (N_1380,N_536,N_1031);
nor U1381 (N_1381,N_861,N_1204);
and U1382 (N_1382,In_635,N_1199);
and U1383 (N_1383,N_689,N_1141);
or U1384 (N_1384,In_1157,In_1758);
and U1385 (N_1385,N_1061,N_972);
xnor U1386 (N_1386,N_1182,N_845);
or U1387 (N_1387,N_194,N_523);
nor U1388 (N_1388,In_1725,In_1543);
nand U1389 (N_1389,N_1162,N_182);
nand U1390 (N_1390,In_1918,In_195);
xnor U1391 (N_1391,In_2452,N_1069);
and U1392 (N_1392,In_623,N_707);
nand U1393 (N_1393,N_377,N_1221);
xor U1394 (N_1394,In_660,N_817);
nor U1395 (N_1395,N_937,In_436);
or U1396 (N_1396,N_720,In_1567);
or U1397 (N_1397,In_665,N_1143);
nor U1398 (N_1398,N_992,In_1299);
and U1399 (N_1399,N_1208,N_1132);
or U1400 (N_1400,In_1219,N_640);
nor U1401 (N_1401,In_1511,N_571);
or U1402 (N_1402,In_2190,N_1097);
xnor U1403 (N_1403,N_768,N_1108);
or U1404 (N_1404,In_2131,N_690);
and U1405 (N_1405,In_2179,N_184);
and U1406 (N_1406,N_333,N_632);
and U1407 (N_1407,N_779,In_1982);
or U1408 (N_1408,N_1120,N_631);
and U1409 (N_1409,N_1047,In_1754);
and U1410 (N_1410,N_947,In_1193);
xor U1411 (N_1411,In_534,N_1019);
or U1412 (N_1412,N_893,In_1964);
and U1413 (N_1413,N_92,N_700);
or U1414 (N_1414,N_1,N_629);
xor U1415 (N_1415,N_759,N_515);
nor U1416 (N_1416,N_850,N_395);
or U1417 (N_1417,N_774,N_884);
nor U1418 (N_1418,N_1014,N_618);
nand U1419 (N_1419,N_952,N_664);
nor U1420 (N_1420,N_661,In_430);
and U1421 (N_1421,In_268,In_2281);
and U1422 (N_1422,In_1489,N_651);
and U1423 (N_1423,N_1135,N_1245);
nand U1424 (N_1424,N_488,In_2380);
and U1425 (N_1425,N_975,N_912);
nand U1426 (N_1426,N_1193,N_385);
and U1427 (N_1427,In_166,N_114);
or U1428 (N_1428,In_1721,In_2445);
xor U1429 (N_1429,In_1585,In_1465);
and U1430 (N_1430,In_1072,In_10);
nor U1431 (N_1431,In_1998,N_853);
or U1432 (N_1432,N_813,N_848);
xnor U1433 (N_1433,In_1096,N_990);
and U1434 (N_1434,N_96,In_1304);
or U1435 (N_1435,N_865,N_1125);
xnor U1436 (N_1436,N_821,N_898);
xor U1437 (N_1437,In_851,In_310);
and U1438 (N_1438,N_235,N_758);
nand U1439 (N_1439,In_613,In_190);
or U1440 (N_1440,N_923,N_1086);
xnor U1441 (N_1441,In_1942,N_902);
xor U1442 (N_1442,In_1662,N_712);
nand U1443 (N_1443,In_714,N_919);
xor U1444 (N_1444,N_939,N_1072);
xor U1445 (N_1445,N_1008,N_1149);
or U1446 (N_1446,In_171,N_653);
nor U1447 (N_1447,N_807,N_846);
xnor U1448 (N_1448,N_1103,N_883);
xnor U1449 (N_1449,N_401,N_405);
nand U1450 (N_1450,N_483,N_564);
nand U1451 (N_1451,N_1244,In_1932);
or U1452 (N_1452,N_1131,N_989);
xnor U1453 (N_1453,N_369,N_911);
and U1454 (N_1454,N_799,In_143);
or U1455 (N_1455,N_740,N_1160);
nand U1456 (N_1456,N_953,In_1257);
nor U1457 (N_1457,In_709,In_1570);
and U1458 (N_1458,N_654,N_620);
nand U1459 (N_1459,N_982,N_736);
xor U1460 (N_1460,N_10,N_645);
and U1461 (N_1461,N_981,In_387);
or U1462 (N_1462,N_1009,N_18);
or U1463 (N_1463,N_901,N_569);
and U1464 (N_1464,N_826,N_847);
and U1465 (N_1465,In_443,In_2096);
or U1466 (N_1466,In_2379,N_783);
xnor U1467 (N_1467,In_1431,In_2462);
or U1468 (N_1468,N_638,N_950);
nand U1469 (N_1469,N_1161,N_1039);
or U1470 (N_1470,N_801,In_1772);
xor U1471 (N_1471,N_681,In_2448);
xor U1472 (N_1472,In_1300,N_633);
nand U1473 (N_1473,N_173,N_1015);
nor U1474 (N_1474,N_1066,N_983);
and U1475 (N_1475,N_891,N_600);
nor U1476 (N_1476,N_1140,N_897);
or U1477 (N_1477,N_1154,In_1139);
nand U1478 (N_1478,In_2238,In_379);
or U1479 (N_1479,N_745,N_1057);
nand U1480 (N_1480,N_1094,In_1214);
nand U1481 (N_1481,In_783,N_761);
and U1482 (N_1482,N_851,N_1064);
or U1483 (N_1483,N_1222,In_1546);
xnor U1484 (N_1484,N_338,N_508);
or U1485 (N_1485,N_781,N_920);
xor U1486 (N_1486,In_970,N_1238);
xor U1487 (N_1487,In_1863,N_780);
nor U1488 (N_1488,N_824,N_1080);
nor U1489 (N_1489,N_746,In_2086);
or U1490 (N_1490,N_699,In_1345);
and U1491 (N_1491,In_1516,N_1006);
xnor U1492 (N_1492,N_453,N_800);
or U1493 (N_1493,N_220,N_686);
nand U1494 (N_1494,N_805,N_665);
xnor U1495 (N_1495,In_1583,N_460);
and U1496 (N_1496,N_396,In_806);
nand U1497 (N_1497,In_1336,N_1079);
xor U1498 (N_1498,In_1276,N_330);
and U1499 (N_1499,N_1237,N_1178);
or U1500 (N_1500,N_994,N_1163);
or U1501 (N_1501,N_136,In_1420);
nor U1502 (N_1502,N_347,N_663);
or U1503 (N_1503,In_1092,N_835);
nand U1504 (N_1504,In_1246,N_1242);
xnor U1505 (N_1505,N_724,N_1124);
nand U1506 (N_1506,N_1158,N_1071);
nor U1507 (N_1507,N_193,N_630);
or U1508 (N_1508,N_822,N_702);
nor U1509 (N_1509,N_1190,In_2121);
or U1510 (N_1510,N_732,N_790);
and U1511 (N_1511,N_78,In_749);
and U1512 (N_1512,N_1029,N_522);
or U1513 (N_1513,N_1145,N_366);
nor U1514 (N_1514,In_256,N_831);
nand U1515 (N_1515,N_33,N_860);
xnor U1516 (N_1516,In_1154,In_1659);
and U1517 (N_1517,In_1156,N_926);
nor U1518 (N_1518,In_987,N_339);
or U1519 (N_1519,N_753,N_577);
and U1520 (N_1520,In_2056,N_1062);
nand U1521 (N_1521,N_721,N_935);
nand U1522 (N_1522,N_1028,In_91);
and U1523 (N_1523,N_866,N_1134);
and U1524 (N_1524,N_598,In_1882);
nor U1525 (N_1525,In_2450,N_882);
nand U1526 (N_1526,N_97,In_572);
and U1527 (N_1527,N_956,In_211);
nand U1528 (N_1528,N_795,N_544);
or U1529 (N_1529,In_607,N_769);
or U1530 (N_1530,In_752,N_1236);
nor U1531 (N_1531,N_1093,In_137);
and U1532 (N_1532,N_264,In_1764);
or U1533 (N_1533,N_969,N_1167);
nand U1534 (N_1534,In_2497,N_945);
nand U1535 (N_1535,N_606,N_24);
or U1536 (N_1536,N_634,In_407);
or U1537 (N_1537,N_687,N_1184);
nor U1538 (N_1538,N_326,N_705);
or U1539 (N_1539,In_1497,N_391);
nor U1540 (N_1540,In_422,In_2181);
xor U1541 (N_1541,In_66,N_1065);
and U1542 (N_1542,N_766,In_1815);
nand U1543 (N_1543,N_1112,N_118);
nand U1544 (N_1544,N_1050,N_868);
nand U1545 (N_1545,N_1042,In_76);
nor U1546 (N_1546,N_1130,N_804);
and U1547 (N_1547,N_1166,In_1114);
nor U1548 (N_1548,N_128,N_881);
and U1549 (N_1549,N_1138,In_1831);
xor U1550 (N_1550,N_259,N_812);
nand U1551 (N_1551,In_1102,In_222);
and U1552 (N_1552,N_668,N_512);
nand U1553 (N_1553,N_1117,N_715);
nand U1554 (N_1554,N_655,In_2363);
nor U1555 (N_1555,N_752,N_967);
or U1556 (N_1556,N_905,N_670);
or U1557 (N_1557,In_2060,In_1880);
and U1558 (N_1558,N_1220,In_22);
xor U1559 (N_1559,N_272,N_212);
nand U1560 (N_1560,N_1115,N_725);
xor U1561 (N_1561,N_1179,N_927);
or U1562 (N_1562,N_666,N_871);
or U1563 (N_1563,N_957,N_675);
xnor U1564 (N_1564,N_214,N_1122);
or U1565 (N_1565,In_27,In_1501);
xnor U1566 (N_1566,In_1275,N_659);
nor U1567 (N_1567,N_730,In_695);
and U1568 (N_1568,N_924,In_521);
xnor U1569 (N_1569,N_1187,N_900);
xnor U1570 (N_1570,N_4,N_168);
nor U1571 (N_1571,In_1956,In_1450);
nor U1572 (N_1572,In_2318,N_1076);
nor U1573 (N_1573,N_776,In_93);
nand U1574 (N_1574,N_1189,N_1075);
xnor U1575 (N_1575,N_825,In_1678);
xor U1576 (N_1576,N_1088,In_662);
nand U1577 (N_1577,N_680,N_398);
or U1578 (N_1578,N_803,N_916);
and U1579 (N_1579,In_2172,N_1229);
nand U1580 (N_1580,N_1127,N_292);
or U1581 (N_1581,N_657,N_215);
nand U1582 (N_1582,N_1206,N_289);
nand U1583 (N_1583,N_818,In_582);
nand U1584 (N_1584,N_142,N_867);
nor U1585 (N_1585,N_1000,N_789);
or U1586 (N_1586,In_2488,N_1188);
nand U1587 (N_1587,N_936,N_747);
nor U1588 (N_1588,N_1038,N_660);
nand U1589 (N_1589,N_672,N_1173);
nand U1590 (N_1590,N_921,In_272);
and U1591 (N_1591,N_722,In_1243);
and U1592 (N_1592,N_896,N_1165);
and U1593 (N_1593,In_717,N_1037);
nand U1594 (N_1594,In_1913,In_470);
nand U1595 (N_1595,N_890,In_1269);
and U1596 (N_1596,In_642,In_2328);
xnor U1597 (N_1597,In_1985,N_1041);
nor U1598 (N_1598,N_870,N_73);
nand U1599 (N_1599,N_888,In_1598);
and U1600 (N_1600,N_206,In_233);
nand U1601 (N_1601,In_1316,In_321);
or U1602 (N_1602,N_849,N_98);
nor U1603 (N_1603,N_1123,N_1150);
or U1604 (N_1604,N_163,N_1155);
or U1605 (N_1605,N_998,In_1457);
nand U1606 (N_1606,In_1317,N_1192);
xor U1607 (N_1607,N_1053,N_334);
xnor U1608 (N_1608,N_647,In_667);
xnor U1609 (N_1609,In_1924,In_767);
and U1610 (N_1610,In_716,In_484);
nand U1611 (N_1611,N_682,In_522);
xnor U1612 (N_1612,N_859,In_1504);
and U1613 (N_1613,N_917,N_356);
or U1614 (N_1614,N_958,N_354);
or U1615 (N_1615,In_1136,N_1052);
and U1616 (N_1616,N_15,N_869);
or U1617 (N_1617,N_1099,In_3);
xor U1618 (N_1618,In_1843,In_981);
nor U1619 (N_1619,N_918,N_649);
xnor U1620 (N_1620,N_673,N_695);
nand U1621 (N_1621,N_863,N_1113);
or U1622 (N_1622,N_718,N_723);
and U1623 (N_1623,In_252,In_54);
and U1624 (N_1624,N_894,N_892);
and U1625 (N_1625,N_271,In_1222);
nand U1626 (N_1626,N_792,N_315);
nand U1627 (N_1627,N_946,N_191);
nor U1628 (N_1628,In_191,In_57);
nor U1629 (N_1629,N_1137,N_172);
or U1630 (N_1630,N_313,N_991);
or U1631 (N_1631,In_1674,N_216);
nor U1632 (N_1632,N_713,In_1333);
xnor U1633 (N_1633,In_2435,In_393);
nor U1634 (N_1634,N_786,N_764);
or U1635 (N_1635,In_295,N_1191);
nand U1636 (N_1636,In_1556,N_1186);
or U1637 (N_1637,In_39,N_703);
and U1638 (N_1638,N_834,N_829);
xor U1639 (N_1639,N_500,N_698);
or U1640 (N_1640,N_931,N_302);
xnor U1641 (N_1641,N_1104,N_1205);
nor U1642 (N_1642,N_662,N_1195);
or U1643 (N_1643,N_988,N_190);
and U1644 (N_1644,N_1247,In_1986);
nand U1645 (N_1645,In_2352,N_1212);
xor U1646 (N_1646,N_299,N_433);
and U1647 (N_1647,N_737,N_955);
or U1648 (N_1648,In_2213,N_929);
and U1649 (N_1649,N_806,N_1209);
or U1650 (N_1650,N_1215,In_9);
xnor U1651 (N_1651,N_584,N_149);
xnor U1652 (N_1652,N_1198,N_637);
and U1653 (N_1653,N_1016,N_733);
nand U1654 (N_1654,In_2438,N_757);
or U1655 (N_1655,N_819,N_504);
nand U1656 (N_1656,N_1011,In_1917);
nor U1657 (N_1657,N_1024,In_1840);
and U1658 (N_1658,N_802,In_2001);
and U1659 (N_1659,N_1231,N_1180);
and U1660 (N_1660,N_1004,In_1255);
or U1661 (N_1661,N_941,N_1121);
nand U1662 (N_1662,N_505,N_785);
nand U1663 (N_1663,N_1020,N_495);
xnor U1664 (N_1664,N_1176,N_1217);
nor U1665 (N_1665,N_678,In_2185);
nand U1666 (N_1666,N_249,In_180);
nor U1667 (N_1667,N_420,N_1164);
nor U1668 (N_1668,N_706,In_340);
nor U1669 (N_1669,N_773,In_685);
nor U1670 (N_1670,N_1223,N_1240);
and U1671 (N_1671,N_1013,In_1056);
xnor U1672 (N_1672,In_867,N_162);
and U1673 (N_1673,In_2220,In_1467);
nand U1674 (N_1674,N_1077,N_674);
and U1675 (N_1675,N_1111,N_1032);
nor U1676 (N_1676,N_1174,N_858);
xnor U1677 (N_1677,In_2223,N_762);
nor U1678 (N_1678,In_2293,N_995);
nand U1679 (N_1679,N_158,N_763);
nand U1680 (N_1680,In_2414,N_17);
nor U1681 (N_1681,N_479,N_371);
nor U1682 (N_1682,N_1202,N_1148);
xnor U1683 (N_1683,In_30,N_205);
or U1684 (N_1684,In_983,N_126);
or U1685 (N_1685,N_1246,N_909);
xnor U1686 (N_1686,N_997,N_731);
nand U1687 (N_1687,N_697,N_132);
or U1688 (N_1688,N_907,N_148);
or U1689 (N_1689,N_529,N_130);
or U1690 (N_1690,In_772,In_43);
xnor U1691 (N_1691,In_1620,N_719);
or U1692 (N_1692,N_287,N_327);
or U1693 (N_1693,In_719,N_726);
nand U1694 (N_1694,In_530,N_1227);
xor U1695 (N_1695,In_1818,N_55);
nor U1696 (N_1696,N_840,N_628);
and U1697 (N_1697,In_648,N_1087);
nand U1698 (N_1698,N_965,N_968);
and U1699 (N_1699,N_832,N_1063);
xor U1700 (N_1700,In_505,N_1051);
nor U1701 (N_1701,In_1588,N_1153);
and U1702 (N_1702,In_1766,N_1239);
nand U1703 (N_1703,N_1095,N_331);
and U1704 (N_1704,N_838,N_1210);
and U1705 (N_1705,In_445,N_451);
or U1706 (N_1706,N_323,N_1214);
and U1707 (N_1707,In_1517,In_1042);
or U1708 (N_1708,N_770,N_218);
and U1709 (N_1709,N_949,N_1169);
xor U1710 (N_1710,N_1114,N_985);
and U1711 (N_1711,In_757,N_1049);
nand U1712 (N_1712,N_82,N_1012);
and U1713 (N_1713,N_1102,N_750);
nor U1714 (N_1714,N_876,N_318);
nor U1715 (N_1715,In_1283,N_1201);
nand U1716 (N_1716,In_1016,N_604);
nand U1717 (N_1717,N_570,N_658);
and U1718 (N_1718,N_1026,N_1144);
xor U1719 (N_1719,N_908,In_2083);
nand U1720 (N_1720,In_704,N_716);
and U1721 (N_1721,In_2129,In_1873);
nand U1722 (N_1722,N_734,N_230);
nand U1723 (N_1723,N_627,N_1100);
nand U1724 (N_1724,N_426,N_743);
xor U1725 (N_1725,N_691,N_710);
and U1726 (N_1726,In_2436,N_1096);
nand U1727 (N_1727,N_165,In_2116);
xnor U1728 (N_1728,N_594,N_842);
and U1729 (N_1729,N_1089,In_1518);
and U1730 (N_1730,In_729,N_41);
nand U1731 (N_1731,N_85,In_294);
and U1732 (N_1732,N_80,N_683);
xnor U1733 (N_1733,In_1145,N_1044);
nand U1734 (N_1734,In_411,In_1460);
or U1735 (N_1735,N_886,N_993);
and U1736 (N_1736,N_877,N_52);
nor U1737 (N_1737,N_1200,N_974);
nand U1738 (N_1738,In_2451,In_1984);
nand U1739 (N_1739,N_621,N_626);
nand U1740 (N_1740,N_139,In_2020);
xor U1741 (N_1741,N_531,N_1106);
and U1742 (N_1742,N_167,In_1302);
nand U1743 (N_1743,N_930,N_977);
or U1744 (N_1744,N_497,N_784);
nand U1745 (N_1745,In_1566,N_641);
or U1746 (N_1746,N_999,N_174);
or U1747 (N_1747,N_964,In_976);
or U1748 (N_1748,N_1036,In_1890);
nand U1749 (N_1749,N_823,N_305);
and U1750 (N_1750,In_621,In_1226);
xnor U1751 (N_1751,N_1207,N_808);
nor U1752 (N_1752,In_1014,N_157);
and U1753 (N_1753,In_1738,In_1915);
or U1754 (N_1754,In_2496,In_939);
nor U1755 (N_1755,In_1811,In_73);
nand U1756 (N_1756,N_787,In_2149);
or U1757 (N_1757,N_312,N_1070);
or U1758 (N_1758,N_528,N_1048);
nor U1759 (N_1759,N_1213,N_2);
or U1760 (N_1760,N_1105,N_904);
or U1761 (N_1761,N_1055,N_984);
or U1762 (N_1762,N_729,In_2355);
nor U1763 (N_1763,N_1046,N_711);
nand U1764 (N_1764,N_837,N_429);
or U1765 (N_1765,In_327,N_146);
nand U1766 (N_1766,N_1119,In_1478);
xor U1767 (N_1767,N_667,N_996);
nand U1768 (N_1768,N_704,N_1109);
nor U1769 (N_1769,N_814,N_437);
and U1770 (N_1770,In_71,In_912);
and U1771 (N_1771,N_646,N_914);
nand U1772 (N_1772,N_1243,N_841);
nand U1773 (N_1773,In_201,N_50);
xor U1774 (N_1774,In_1505,N_971);
nand U1775 (N_1775,In_354,N_301);
and U1776 (N_1776,N_258,N_828);
nor U1777 (N_1777,In_1628,N_709);
or U1778 (N_1778,N_796,N_1142);
nor U1779 (N_1779,N_319,N_131);
or U1780 (N_1780,In_2016,N_217);
xor U1781 (N_1781,N_692,In_1885);
or U1782 (N_1782,N_978,In_402);
or U1783 (N_1783,In_696,N_669);
or U1784 (N_1784,N_566,In_314);
nand U1785 (N_1785,N_622,N_1203);
xnor U1786 (N_1786,In_1172,N_933);
nor U1787 (N_1787,N_1241,N_551);
nand U1788 (N_1788,In_680,In_136);
or U1789 (N_1789,N_1197,In_1421);
nand U1790 (N_1790,N_643,N_688);
and U1791 (N_1791,N_922,In_1152);
and U1792 (N_1792,N_1010,N_322);
nor U1793 (N_1793,N_280,N_910);
or U1794 (N_1794,In_189,N_343);
nand U1795 (N_1795,N_553,N_885);
nand U1796 (N_1796,In_641,N_976);
nand U1797 (N_1797,N_1219,In_855);
nand U1798 (N_1798,In_1038,N_739);
nand U1799 (N_1799,N_138,N_1146);
xnor U1800 (N_1800,In_512,N_332);
nor U1801 (N_1801,N_1023,In_1066);
nand U1802 (N_1802,N_986,In_1961);
and U1803 (N_1803,In_2069,N_1230);
or U1804 (N_1804,In_657,N_387);
xor U1805 (N_1805,In_448,In_395);
nor U1806 (N_1806,In_881,N_574);
nor U1807 (N_1807,In_49,N_948);
xor U1808 (N_1808,N_961,In_351);
and U1809 (N_1809,In_67,In_1574);
and U1810 (N_1810,N_772,N_728);
nand U1811 (N_1811,N_1058,In_935);
and U1812 (N_1812,N_1081,N_1168);
nand U1813 (N_1813,N_8,In_2130);
xnor U1814 (N_1814,N_963,N_636);
nor U1815 (N_1815,In_1671,N_125);
nand U1816 (N_1816,N_1092,In_1285);
nand U1817 (N_1817,N_1139,In_1791);
nor U1818 (N_1818,N_744,N_1156);
and U1819 (N_1819,N_809,N_940);
nor U1820 (N_1820,N_738,N_1043);
xor U1821 (N_1821,In_1322,N_864);
nand U1822 (N_1822,N_887,In_1692);
nor U1823 (N_1823,In_2175,N_1129);
nor U1824 (N_1824,N_650,N_1157);
xor U1825 (N_1825,N_103,In_614);
nand U1826 (N_1826,N_1083,In_355);
nor U1827 (N_1827,N_288,N_1159);
xor U1828 (N_1828,N_1007,N_816);
nand U1829 (N_1829,N_1118,N_1211);
or U1830 (N_1830,In_125,N_1116);
nand U1831 (N_1831,In_508,N_701);
xor U1832 (N_1832,In_999,N_644);
nand U1833 (N_1833,In_992,N_676);
or U1834 (N_1834,In_1706,In_977);
and U1835 (N_1835,N_1128,In_1242);
nor U1836 (N_1836,N_875,N_642);
nor U1837 (N_1837,N_775,In_1716);
nand U1838 (N_1838,N_767,N_889);
xor U1839 (N_1839,In_1655,In_372);
and U1840 (N_1840,In_1676,In_1822);
or U1841 (N_1841,N_895,N_856);
and U1842 (N_1842,N_793,N_872);
xnor U1843 (N_1843,N_270,In_1883);
xor U1844 (N_1844,N_1101,In_2273);
xor U1845 (N_1845,In_1553,In_345);
nand U1846 (N_1846,N_1183,N_27);
or U1847 (N_1847,N_1022,In_1018);
nand U1848 (N_1848,N_364,In_103);
or U1849 (N_1849,N_899,N_1226);
nand U1850 (N_1850,N_915,In_948);
and U1851 (N_1851,N_717,N_147);
nor U1852 (N_1852,In_902,N_625);
xor U1853 (N_1853,N_656,In_1530);
nor U1854 (N_1854,N_652,In_1947);
xor U1855 (N_1855,In_1730,N_874);
xnor U1856 (N_1856,N_833,In_65);
nand U1857 (N_1857,In_208,In_1035);
nor U1858 (N_1858,In_1221,N_756);
nor U1859 (N_1859,In_1362,N_934);
xnor U1860 (N_1860,In_1179,N_951);
xor U1861 (N_1861,N_820,In_1854);
or U1862 (N_1862,N_116,N_830);
and U1863 (N_1863,N_619,N_735);
xnor U1864 (N_1864,N_696,N_155);
xnor U1865 (N_1865,In_504,N_878);
xnor U1866 (N_1866,N_741,N_1034);
nor U1867 (N_1867,N_304,In_2409);
xnor U1868 (N_1868,N_1025,N_1040);
xor U1869 (N_1869,In_705,N_472);
nor U1870 (N_1870,N_256,In_1026);
xor U1871 (N_1871,In_862,N_973);
nand U1872 (N_1872,In_1995,N_183);
nor U1873 (N_1873,In_2487,N_413);
and U1874 (N_1874,N_648,In_1771);
and U1875 (N_1875,N_1521,N_1328);
xor U1876 (N_1876,N_1371,N_1443);
and U1877 (N_1877,N_1586,N_1338);
nor U1878 (N_1878,N_1310,N_1726);
nand U1879 (N_1879,N_1427,N_1531);
and U1880 (N_1880,N_1296,N_1513);
and U1881 (N_1881,N_1672,N_1461);
nor U1882 (N_1882,N_1384,N_1861);
and U1883 (N_1883,N_1783,N_1494);
or U1884 (N_1884,N_1509,N_1421);
or U1885 (N_1885,N_1593,N_1626);
and U1886 (N_1886,N_1800,N_1841);
or U1887 (N_1887,N_1411,N_1763);
nand U1888 (N_1888,N_1614,N_1399);
nor U1889 (N_1889,N_1568,N_1317);
or U1890 (N_1890,N_1265,N_1860);
and U1891 (N_1891,N_1590,N_1862);
xor U1892 (N_1892,N_1511,N_1830);
xor U1893 (N_1893,N_1829,N_1331);
nor U1894 (N_1894,N_1572,N_1629);
or U1895 (N_1895,N_1667,N_1804);
nor U1896 (N_1896,N_1577,N_1368);
nand U1897 (N_1897,N_1423,N_1524);
nand U1898 (N_1898,N_1369,N_1447);
and U1899 (N_1899,N_1698,N_1744);
xor U1900 (N_1900,N_1482,N_1676);
xnor U1901 (N_1901,N_1498,N_1462);
nand U1902 (N_1902,N_1446,N_1848);
nor U1903 (N_1903,N_1458,N_1375);
nor U1904 (N_1904,N_1449,N_1668);
or U1905 (N_1905,N_1859,N_1267);
xor U1906 (N_1906,N_1313,N_1632);
xor U1907 (N_1907,N_1775,N_1566);
or U1908 (N_1908,N_1413,N_1567);
nand U1909 (N_1909,N_1554,N_1319);
nor U1910 (N_1910,N_1451,N_1504);
xnor U1911 (N_1911,N_1683,N_1866);
and U1912 (N_1912,N_1790,N_1682);
or U1913 (N_1913,N_1537,N_1795);
nand U1914 (N_1914,N_1376,N_1630);
nor U1915 (N_1915,N_1681,N_1735);
or U1916 (N_1916,N_1569,N_1496);
nand U1917 (N_1917,N_1424,N_1438);
or U1918 (N_1918,N_1311,N_1801);
nor U1919 (N_1919,N_1769,N_1733);
nand U1920 (N_1920,N_1722,N_1432);
nand U1921 (N_1921,N_1362,N_1575);
or U1922 (N_1922,N_1491,N_1640);
nand U1923 (N_1923,N_1401,N_1826);
or U1924 (N_1924,N_1792,N_1811);
or U1925 (N_1925,N_1659,N_1366);
or U1926 (N_1926,N_1639,N_1767);
nand U1927 (N_1927,N_1470,N_1431);
and U1928 (N_1928,N_1275,N_1784);
xnor U1929 (N_1929,N_1484,N_1869);
nand U1930 (N_1930,N_1605,N_1654);
and U1931 (N_1931,N_1557,N_1836);
or U1932 (N_1932,N_1812,N_1307);
xnor U1933 (N_1933,N_1270,N_1351);
and U1934 (N_1934,N_1625,N_1348);
nor U1935 (N_1935,N_1476,N_1678);
and U1936 (N_1936,N_1430,N_1643);
or U1937 (N_1937,N_1774,N_1293);
and U1938 (N_1938,N_1428,N_1757);
xnor U1939 (N_1939,N_1747,N_1336);
and U1940 (N_1940,N_1392,N_1810);
nand U1941 (N_1941,N_1488,N_1847);
or U1942 (N_1942,N_1713,N_1358);
xnor U1943 (N_1943,N_1578,N_1613);
and U1944 (N_1944,N_1679,N_1731);
or U1945 (N_1945,N_1495,N_1515);
nand U1946 (N_1946,N_1522,N_1409);
xor U1947 (N_1947,N_1356,N_1502);
nor U1948 (N_1948,N_1686,N_1636);
and U1949 (N_1949,N_1279,N_1365);
or U1950 (N_1950,N_1288,N_1696);
nor U1951 (N_1951,N_1634,N_1408);
nor U1952 (N_1952,N_1777,N_1334);
xor U1953 (N_1953,N_1844,N_1762);
and U1954 (N_1954,N_1268,N_1749);
nor U1955 (N_1955,N_1734,N_1393);
xor U1956 (N_1956,N_1283,N_1587);
nand U1957 (N_1957,N_1483,N_1526);
nor U1958 (N_1958,N_1727,N_1426);
and U1959 (N_1959,N_1740,N_1463);
nor U1960 (N_1960,N_1353,N_1623);
xnor U1961 (N_1961,N_1326,N_1490);
and U1962 (N_1962,N_1454,N_1573);
and U1963 (N_1963,N_1519,N_1730);
xor U1964 (N_1964,N_1418,N_1817);
or U1965 (N_1965,N_1304,N_1318);
nor U1966 (N_1966,N_1361,N_1388);
nand U1967 (N_1967,N_1385,N_1746);
xnor U1968 (N_1968,N_1448,N_1555);
nor U1969 (N_1969,N_1489,N_1687);
nor U1970 (N_1970,N_1598,N_1445);
or U1971 (N_1971,N_1729,N_1584);
nand U1972 (N_1972,N_1329,N_1711);
or U1973 (N_1973,N_1666,N_1793);
nand U1974 (N_1974,N_1501,N_1620);
or U1975 (N_1975,N_1335,N_1545);
xnor U1976 (N_1976,N_1758,N_1534);
or U1977 (N_1977,N_1716,N_1802);
nor U1978 (N_1978,N_1583,N_1635);
nor U1979 (N_1979,N_1252,N_1433);
nand U1980 (N_1980,N_1284,N_1548);
nand U1981 (N_1981,N_1437,N_1373);
xnor U1982 (N_1982,N_1292,N_1536);
or U1983 (N_1983,N_1720,N_1680);
xor U1984 (N_1984,N_1417,N_1853);
or U1985 (N_1985,N_1407,N_1723);
xor U1986 (N_1986,N_1434,N_1379);
nor U1987 (N_1987,N_1585,N_1559);
nand U1988 (N_1988,N_1674,N_1602);
xnor U1989 (N_1989,N_1520,N_1833);
xnor U1990 (N_1990,N_1360,N_1425);
and U1991 (N_1991,N_1503,N_1255);
nor U1992 (N_1992,N_1805,N_1717);
nand U1993 (N_1993,N_1277,N_1694);
and U1994 (N_1994,N_1506,N_1764);
nor U1995 (N_1995,N_1685,N_1415);
nor U1996 (N_1996,N_1647,N_1301);
nand U1997 (N_1997,N_1819,N_1761);
and U1998 (N_1998,N_1637,N_1597);
xor U1999 (N_1999,N_1465,N_1325);
and U2000 (N_2000,N_1493,N_1652);
xor U2001 (N_2001,N_1823,N_1760);
or U2002 (N_2002,N_1565,N_1420);
nor U2003 (N_2003,N_1646,N_1551);
nand U2004 (N_2004,N_1851,N_1297);
or U2005 (N_2005,N_1755,N_1294);
xnor U2006 (N_2006,N_1736,N_1701);
or U2007 (N_2007,N_1258,N_1481);
or U2008 (N_2008,N_1603,N_1276);
nor U2009 (N_2009,N_1803,N_1464);
xor U2010 (N_2010,N_1611,N_1570);
nor U2011 (N_2011,N_1825,N_1260);
and U2012 (N_2012,N_1324,N_1299);
and U2013 (N_2013,N_1724,N_1673);
and U2014 (N_2014,N_1344,N_1846);
nor U2015 (N_2015,N_1670,N_1601);
and U2016 (N_2016,N_1486,N_1858);
nor U2017 (N_2017,N_1671,N_1455);
nand U2018 (N_2018,N_1719,N_1771);
xnor U2019 (N_2019,N_1786,N_1395);
nand U2020 (N_2020,N_1269,N_1868);
nor U2021 (N_2021,N_1658,N_1410);
xor U2022 (N_2022,N_1633,N_1403);
or U2023 (N_2023,N_1839,N_1263);
and U2024 (N_2024,N_1814,N_1333);
and U2025 (N_2025,N_1499,N_1391);
xnor U2026 (N_2026,N_1542,N_1660);
and U2027 (N_2027,N_1781,N_1553);
and U2028 (N_2028,N_1316,N_1380);
nand U2029 (N_2029,N_1725,N_1469);
xnor U2030 (N_2030,N_1549,N_1312);
nand U2031 (N_2031,N_1828,N_1827);
or U2032 (N_2032,N_1364,N_1574);
nor U2033 (N_2033,N_1648,N_1303);
nand U2034 (N_2034,N_1842,N_1571);
nand U2035 (N_2035,N_1541,N_1337);
xor U2036 (N_2036,N_1782,N_1436);
nor U2037 (N_2037,N_1352,N_1527);
or U2038 (N_2038,N_1628,N_1840);
and U2039 (N_2039,N_1808,N_1510);
nor U2040 (N_2040,N_1273,N_1552);
nor U2041 (N_2041,N_1765,N_1530);
or U2042 (N_2042,N_1261,N_1645);
or U2043 (N_2043,N_1374,N_1264);
nor U2044 (N_2044,N_1308,N_1608);
nand U2045 (N_2045,N_1435,N_1357);
and U2046 (N_2046,N_1305,N_1271);
or U2047 (N_2047,N_1251,N_1355);
and U2048 (N_2048,N_1295,N_1416);
nand U2049 (N_2049,N_1745,N_1475);
xnor U2050 (N_2050,N_1759,N_1457);
xnor U2051 (N_2051,N_1546,N_1581);
nand U2052 (N_2052,N_1291,N_1831);
nor U2053 (N_2053,N_1865,N_1523);
and U2054 (N_2054,N_1856,N_1773);
nand U2055 (N_2055,N_1768,N_1772);
nor U2056 (N_2056,N_1700,N_1286);
nor U2057 (N_2057,N_1444,N_1327);
and U2058 (N_2058,N_1341,N_1580);
nand U2059 (N_2059,N_1622,N_1532);
xor U2060 (N_2060,N_1383,N_1835);
and U2061 (N_2061,N_1377,N_1330);
or U2062 (N_2062,N_1750,N_1867);
nand U2063 (N_2063,N_1824,N_1439);
and U2064 (N_2064,N_1616,N_1429);
or U2065 (N_2065,N_1266,N_1770);
nand U2066 (N_2066,N_1562,N_1378);
nand U2067 (N_2067,N_1663,N_1564);
nor U2068 (N_2068,N_1738,N_1529);
or U2069 (N_2069,N_1864,N_1650);
nand U2070 (N_2070,N_1543,N_1699);
xor U2071 (N_2071,N_1386,N_1332);
nor U2072 (N_2072,N_1820,N_1797);
or U2073 (N_2073,N_1871,N_1752);
nand U2074 (N_2074,N_1872,N_1815);
xnor U2075 (N_2075,N_1619,N_1540);
nand U2076 (N_2076,N_1776,N_1525);
xor U2077 (N_2077,N_1664,N_1278);
or U2078 (N_2078,N_1422,N_1472);
nand U2079 (N_2079,N_1306,N_1346);
nand U2080 (N_2080,N_1282,N_1606);
xnor U2081 (N_2081,N_1838,N_1561);
or U2082 (N_2082,N_1528,N_1320);
nor U2083 (N_2083,N_1589,N_1692);
or U2084 (N_2084,N_1816,N_1550);
xor U2085 (N_2085,N_1505,N_1691);
or U2086 (N_2086,N_1257,N_1787);
nand U2087 (N_2087,N_1697,N_1788);
or U2088 (N_2088,N_1556,N_1834);
nor U2089 (N_2089,N_1467,N_1742);
or U2090 (N_2090,N_1289,N_1456);
nand U2091 (N_2091,N_1857,N_1706);
xor U2092 (N_2092,N_1404,N_1707);
nor U2093 (N_2093,N_1753,N_1398);
nor U2094 (N_2094,N_1402,N_1539);
and U2095 (N_2095,N_1414,N_1695);
xnor U2096 (N_2096,N_1662,N_1712);
or U2097 (N_2097,N_1615,N_1314);
or U2098 (N_2098,N_1500,N_1843);
and U2099 (N_2099,N_1644,N_1394);
nand U2100 (N_2100,N_1354,N_1302);
or U2101 (N_2101,N_1485,N_1689);
or U2102 (N_2102,N_1617,N_1592);
nand U2103 (N_2103,N_1604,N_1832);
nor U2104 (N_2104,N_1480,N_1280);
xnor U2105 (N_2105,N_1778,N_1518);
and U2106 (N_2106,N_1582,N_1653);
xnor U2107 (N_2107,N_1612,N_1400);
nand U2108 (N_2108,N_1492,N_1850);
nor U2109 (N_2109,N_1642,N_1487);
and U2110 (N_2110,N_1262,N_1821);
and U2111 (N_2111,N_1512,N_1533);
nand U2112 (N_2112,N_1796,N_1818);
or U2113 (N_2113,N_1721,N_1779);
nand U2114 (N_2114,N_1627,N_1798);
xnor U2115 (N_2115,N_1459,N_1323);
nand U2116 (N_2116,N_1870,N_1372);
nand U2117 (N_2117,N_1347,N_1558);
xnor U2118 (N_2118,N_1703,N_1718);
nand U2119 (N_2119,N_1780,N_1466);
xor U2120 (N_2120,N_1340,N_1478);
nor U2121 (N_2121,N_1477,N_1600);
xor U2122 (N_2122,N_1250,N_1799);
nor U2123 (N_2123,N_1785,N_1544);
or U2124 (N_2124,N_1656,N_1382);
and U2125 (N_2125,N_1684,N_1560);
xnor U2126 (N_2126,N_1732,N_1579);
xnor U2127 (N_2127,N_1516,N_1254);
and U2128 (N_2128,N_1507,N_1479);
xor U2129 (N_2129,N_1397,N_1538);
or U2130 (N_2130,N_1594,N_1791);
or U2131 (N_2131,N_1471,N_1290);
and U2132 (N_2132,N_1693,N_1442);
xnor U2133 (N_2133,N_1661,N_1343);
or U2134 (N_2134,N_1708,N_1591);
nor U2135 (N_2135,N_1837,N_1655);
nand U2136 (N_2136,N_1657,N_1794);
or U2137 (N_2137,N_1690,N_1474);
nand U2138 (N_2138,N_1274,N_1563);
or U2139 (N_2139,N_1595,N_1813);
xor U2140 (N_2140,N_1610,N_1754);
nand U2141 (N_2141,N_1321,N_1517);
xor U2142 (N_2142,N_1677,N_1728);
xor U2143 (N_2143,N_1367,N_1345);
nand U2144 (N_2144,N_1272,N_1535);
and U2145 (N_2145,N_1350,N_1396);
nor U2146 (N_2146,N_1705,N_1873);
xnor U2147 (N_2147,N_1370,N_1669);
nand U2148 (N_2148,N_1675,N_1342);
nor U2149 (N_2149,N_1387,N_1460);
and U2150 (N_2150,N_1849,N_1298);
nand U2151 (N_2151,N_1704,N_1756);
nand U2152 (N_2152,N_1389,N_1709);
nor U2153 (N_2153,N_1855,N_1748);
xor U2154 (N_2154,N_1599,N_1822);
and U2155 (N_2155,N_1441,N_1363);
xnor U2156 (N_2156,N_1741,N_1497);
or U2157 (N_2157,N_1309,N_1473);
or U2158 (N_2158,N_1638,N_1300);
nand U2159 (N_2159,N_1285,N_1453);
nand U2160 (N_2160,N_1412,N_1874);
nor U2161 (N_2161,N_1596,N_1649);
nor U2162 (N_2162,N_1508,N_1621);
and U2163 (N_2163,N_1468,N_1406);
nor U2164 (N_2164,N_1766,N_1852);
and U2165 (N_2165,N_1624,N_1806);
nand U2166 (N_2166,N_1514,N_1259);
nand U2167 (N_2167,N_1609,N_1607);
nor U2168 (N_2168,N_1854,N_1381);
or U2169 (N_2169,N_1359,N_1588);
xor U2170 (N_2170,N_1702,N_1440);
or U2171 (N_2171,N_1863,N_1281);
xnor U2172 (N_2172,N_1751,N_1665);
nand U2173 (N_2173,N_1807,N_1743);
xnor U2174 (N_2174,N_1349,N_1287);
nand U2175 (N_2175,N_1631,N_1714);
xor U2176 (N_2176,N_1253,N_1845);
and U2177 (N_2177,N_1450,N_1739);
and U2178 (N_2178,N_1315,N_1715);
nand U2179 (N_2179,N_1688,N_1737);
and U2180 (N_2180,N_1322,N_1419);
xor U2181 (N_2181,N_1618,N_1651);
nor U2182 (N_2182,N_1256,N_1390);
or U2183 (N_2183,N_1339,N_1547);
nand U2184 (N_2184,N_1405,N_1576);
xnor U2185 (N_2185,N_1710,N_1789);
and U2186 (N_2186,N_1452,N_1641);
nand U2187 (N_2187,N_1809,N_1801);
nand U2188 (N_2188,N_1844,N_1611);
xnor U2189 (N_2189,N_1416,N_1502);
nor U2190 (N_2190,N_1794,N_1411);
and U2191 (N_2191,N_1591,N_1395);
nor U2192 (N_2192,N_1866,N_1821);
and U2193 (N_2193,N_1829,N_1459);
nand U2194 (N_2194,N_1695,N_1367);
nor U2195 (N_2195,N_1741,N_1775);
or U2196 (N_2196,N_1428,N_1817);
and U2197 (N_2197,N_1583,N_1483);
nor U2198 (N_2198,N_1282,N_1823);
or U2199 (N_2199,N_1712,N_1579);
and U2200 (N_2200,N_1279,N_1601);
and U2201 (N_2201,N_1254,N_1431);
xor U2202 (N_2202,N_1555,N_1265);
nand U2203 (N_2203,N_1344,N_1811);
or U2204 (N_2204,N_1543,N_1282);
xnor U2205 (N_2205,N_1324,N_1502);
xnor U2206 (N_2206,N_1551,N_1376);
nand U2207 (N_2207,N_1810,N_1633);
and U2208 (N_2208,N_1619,N_1744);
or U2209 (N_2209,N_1667,N_1475);
and U2210 (N_2210,N_1392,N_1818);
or U2211 (N_2211,N_1525,N_1557);
nand U2212 (N_2212,N_1644,N_1716);
or U2213 (N_2213,N_1560,N_1334);
or U2214 (N_2214,N_1258,N_1294);
xnor U2215 (N_2215,N_1293,N_1368);
and U2216 (N_2216,N_1642,N_1399);
nand U2217 (N_2217,N_1799,N_1270);
nand U2218 (N_2218,N_1394,N_1462);
or U2219 (N_2219,N_1745,N_1697);
nand U2220 (N_2220,N_1809,N_1498);
and U2221 (N_2221,N_1392,N_1369);
and U2222 (N_2222,N_1496,N_1358);
nand U2223 (N_2223,N_1419,N_1306);
xnor U2224 (N_2224,N_1687,N_1784);
and U2225 (N_2225,N_1517,N_1818);
nor U2226 (N_2226,N_1345,N_1831);
nand U2227 (N_2227,N_1332,N_1707);
xor U2228 (N_2228,N_1256,N_1813);
nand U2229 (N_2229,N_1430,N_1367);
nand U2230 (N_2230,N_1639,N_1278);
or U2231 (N_2231,N_1327,N_1496);
nor U2232 (N_2232,N_1715,N_1651);
nor U2233 (N_2233,N_1254,N_1851);
xor U2234 (N_2234,N_1658,N_1296);
xor U2235 (N_2235,N_1263,N_1376);
nand U2236 (N_2236,N_1846,N_1662);
or U2237 (N_2237,N_1811,N_1688);
and U2238 (N_2238,N_1568,N_1741);
xnor U2239 (N_2239,N_1405,N_1553);
xnor U2240 (N_2240,N_1626,N_1661);
or U2241 (N_2241,N_1370,N_1255);
nand U2242 (N_2242,N_1718,N_1411);
nor U2243 (N_2243,N_1778,N_1595);
and U2244 (N_2244,N_1418,N_1474);
nand U2245 (N_2245,N_1471,N_1423);
and U2246 (N_2246,N_1614,N_1476);
nor U2247 (N_2247,N_1735,N_1708);
xor U2248 (N_2248,N_1479,N_1733);
nand U2249 (N_2249,N_1339,N_1559);
nand U2250 (N_2250,N_1845,N_1568);
and U2251 (N_2251,N_1624,N_1397);
nand U2252 (N_2252,N_1826,N_1503);
nor U2253 (N_2253,N_1382,N_1310);
xor U2254 (N_2254,N_1711,N_1708);
or U2255 (N_2255,N_1374,N_1661);
and U2256 (N_2256,N_1860,N_1842);
xnor U2257 (N_2257,N_1282,N_1357);
and U2258 (N_2258,N_1694,N_1257);
xnor U2259 (N_2259,N_1431,N_1584);
and U2260 (N_2260,N_1790,N_1414);
or U2261 (N_2261,N_1531,N_1688);
xnor U2262 (N_2262,N_1461,N_1384);
or U2263 (N_2263,N_1472,N_1395);
nand U2264 (N_2264,N_1684,N_1687);
nor U2265 (N_2265,N_1397,N_1818);
xor U2266 (N_2266,N_1259,N_1440);
nand U2267 (N_2267,N_1672,N_1713);
nor U2268 (N_2268,N_1707,N_1271);
and U2269 (N_2269,N_1538,N_1834);
nand U2270 (N_2270,N_1669,N_1399);
nor U2271 (N_2271,N_1477,N_1522);
xor U2272 (N_2272,N_1572,N_1253);
nand U2273 (N_2273,N_1847,N_1734);
and U2274 (N_2274,N_1300,N_1352);
nand U2275 (N_2275,N_1735,N_1543);
xnor U2276 (N_2276,N_1788,N_1368);
nor U2277 (N_2277,N_1364,N_1523);
and U2278 (N_2278,N_1865,N_1795);
or U2279 (N_2279,N_1596,N_1563);
xor U2280 (N_2280,N_1605,N_1404);
nand U2281 (N_2281,N_1393,N_1870);
xnor U2282 (N_2282,N_1275,N_1365);
nor U2283 (N_2283,N_1429,N_1641);
and U2284 (N_2284,N_1730,N_1497);
and U2285 (N_2285,N_1826,N_1469);
or U2286 (N_2286,N_1791,N_1633);
and U2287 (N_2287,N_1331,N_1283);
nor U2288 (N_2288,N_1457,N_1714);
nor U2289 (N_2289,N_1382,N_1567);
nand U2290 (N_2290,N_1766,N_1388);
and U2291 (N_2291,N_1715,N_1366);
nand U2292 (N_2292,N_1699,N_1393);
nand U2293 (N_2293,N_1432,N_1343);
nor U2294 (N_2294,N_1686,N_1632);
nand U2295 (N_2295,N_1691,N_1728);
nand U2296 (N_2296,N_1326,N_1740);
or U2297 (N_2297,N_1495,N_1394);
nor U2298 (N_2298,N_1288,N_1591);
or U2299 (N_2299,N_1681,N_1763);
or U2300 (N_2300,N_1575,N_1597);
nand U2301 (N_2301,N_1686,N_1384);
or U2302 (N_2302,N_1803,N_1772);
nor U2303 (N_2303,N_1479,N_1748);
nand U2304 (N_2304,N_1621,N_1336);
nor U2305 (N_2305,N_1466,N_1327);
xor U2306 (N_2306,N_1330,N_1299);
nand U2307 (N_2307,N_1840,N_1707);
nand U2308 (N_2308,N_1843,N_1825);
or U2309 (N_2309,N_1367,N_1789);
and U2310 (N_2310,N_1532,N_1342);
nand U2311 (N_2311,N_1771,N_1413);
xnor U2312 (N_2312,N_1413,N_1585);
nor U2313 (N_2313,N_1713,N_1685);
or U2314 (N_2314,N_1647,N_1819);
xnor U2315 (N_2315,N_1396,N_1299);
nor U2316 (N_2316,N_1741,N_1364);
or U2317 (N_2317,N_1778,N_1731);
xnor U2318 (N_2318,N_1860,N_1254);
nor U2319 (N_2319,N_1641,N_1462);
nand U2320 (N_2320,N_1279,N_1330);
or U2321 (N_2321,N_1285,N_1793);
nand U2322 (N_2322,N_1609,N_1665);
nand U2323 (N_2323,N_1461,N_1454);
or U2324 (N_2324,N_1476,N_1263);
nor U2325 (N_2325,N_1318,N_1259);
nand U2326 (N_2326,N_1258,N_1270);
nor U2327 (N_2327,N_1338,N_1333);
and U2328 (N_2328,N_1725,N_1317);
and U2329 (N_2329,N_1753,N_1363);
and U2330 (N_2330,N_1819,N_1297);
and U2331 (N_2331,N_1723,N_1550);
xor U2332 (N_2332,N_1758,N_1342);
and U2333 (N_2333,N_1735,N_1775);
nor U2334 (N_2334,N_1643,N_1299);
or U2335 (N_2335,N_1576,N_1538);
or U2336 (N_2336,N_1582,N_1424);
xor U2337 (N_2337,N_1652,N_1475);
nor U2338 (N_2338,N_1292,N_1769);
or U2339 (N_2339,N_1293,N_1743);
nor U2340 (N_2340,N_1840,N_1684);
nor U2341 (N_2341,N_1678,N_1865);
xnor U2342 (N_2342,N_1399,N_1674);
nand U2343 (N_2343,N_1269,N_1818);
and U2344 (N_2344,N_1716,N_1597);
or U2345 (N_2345,N_1452,N_1260);
and U2346 (N_2346,N_1308,N_1854);
or U2347 (N_2347,N_1873,N_1710);
nor U2348 (N_2348,N_1475,N_1654);
or U2349 (N_2349,N_1816,N_1568);
or U2350 (N_2350,N_1284,N_1336);
or U2351 (N_2351,N_1827,N_1723);
nor U2352 (N_2352,N_1379,N_1724);
or U2353 (N_2353,N_1549,N_1758);
nand U2354 (N_2354,N_1831,N_1273);
or U2355 (N_2355,N_1258,N_1420);
and U2356 (N_2356,N_1722,N_1728);
nand U2357 (N_2357,N_1651,N_1632);
or U2358 (N_2358,N_1461,N_1742);
nor U2359 (N_2359,N_1335,N_1408);
nand U2360 (N_2360,N_1725,N_1295);
nand U2361 (N_2361,N_1554,N_1344);
or U2362 (N_2362,N_1699,N_1652);
nand U2363 (N_2363,N_1468,N_1715);
xnor U2364 (N_2364,N_1254,N_1520);
and U2365 (N_2365,N_1433,N_1776);
and U2366 (N_2366,N_1316,N_1577);
nand U2367 (N_2367,N_1301,N_1745);
nand U2368 (N_2368,N_1585,N_1671);
and U2369 (N_2369,N_1807,N_1511);
or U2370 (N_2370,N_1602,N_1619);
and U2371 (N_2371,N_1288,N_1671);
xnor U2372 (N_2372,N_1256,N_1461);
xnor U2373 (N_2373,N_1671,N_1664);
and U2374 (N_2374,N_1714,N_1639);
nor U2375 (N_2375,N_1714,N_1480);
or U2376 (N_2376,N_1857,N_1253);
and U2377 (N_2377,N_1744,N_1700);
nand U2378 (N_2378,N_1445,N_1669);
nor U2379 (N_2379,N_1672,N_1555);
nor U2380 (N_2380,N_1870,N_1601);
xnor U2381 (N_2381,N_1643,N_1302);
or U2382 (N_2382,N_1254,N_1381);
or U2383 (N_2383,N_1803,N_1610);
nor U2384 (N_2384,N_1590,N_1321);
and U2385 (N_2385,N_1728,N_1840);
nand U2386 (N_2386,N_1538,N_1278);
and U2387 (N_2387,N_1373,N_1789);
nor U2388 (N_2388,N_1622,N_1389);
and U2389 (N_2389,N_1703,N_1729);
and U2390 (N_2390,N_1452,N_1632);
nand U2391 (N_2391,N_1347,N_1369);
and U2392 (N_2392,N_1862,N_1624);
nor U2393 (N_2393,N_1326,N_1679);
xnor U2394 (N_2394,N_1502,N_1592);
xor U2395 (N_2395,N_1309,N_1266);
xnor U2396 (N_2396,N_1767,N_1329);
and U2397 (N_2397,N_1307,N_1818);
nand U2398 (N_2398,N_1818,N_1394);
and U2399 (N_2399,N_1792,N_1323);
nor U2400 (N_2400,N_1694,N_1560);
and U2401 (N_2401,N_1271,N_1565);
nand U2402 (N_2402,N_1387,N_1450);
or U2403 (N_2403,N_1567,N_1420);
nand U2404 (N_2404,N_1421,N_1554);
xnor U2405 (N_2405,N_1445,N_1293);
nor U2406 (N_2406,N_1817,N_1574);
and U2407 (N_2407,N_1336,N_1312);
or U2408 (N_2408,N_1297,N_1577);
xor U2409 (N_2409,N_1256,N_1874);
and U2410 (N_2410,N_1693,N_1716);
and U2411 (N_2411,N_1766,N_1452);
or U2412 (N_2412,N_1523,N_1500);
and U2413 (N_2413,N_1447,N_1354);
nand U2414 (N_2414,N_1326,N_1539);
nand U2415 (N_2415,N_1539,N_1690);
xnor U2416 (N_2416,N_1844,N_1719);
xnor U2417 (N_2417,N_1715,N_1487);
nand U2418 (N_2418,N_1497,N_1794);
and U2419 (N_2419,N_1583,N_1822);
nand U2420 (N_2420,N_1685,N_1332);
nor U2421 (N_2421,N_1613,N_1283);
xnor U2422 (N_2422,N_1844,N_1401);
and U2423 (N_2423,N_1831,N_1354);
and U2424 (N_2424,N_1702,N_1318);
nor U2425 (N_2425,N_1555,N_1682);
and U2426 (N_2426,N_1862,N_1335);
or U2427 (N_2427,N_1807,N_1721);
nand U2428 (N_2428,N_1814,N_1498);
xor U2429 (N_2429,N_1492,N_1254);
nand U2430 (N_2430,N_1708,N_1579);
or U2431 (N_2431,N_1805,N_1820);
nand U2432 (N_2432,N_1828,N_1340);
and U2433 (N_2433,N_1384,N_1446);
nand U2434 (N_2434,N_1737,N_1827);
xor U2435 (N_2435,N_1280,N_1573);
or U2436 (N_2436,N_1511,N_1671);
nand U2437 (N_2437,N_1260,N_1387);
or U2438 (N_2438,N_1656,N_1633);
and U2439 (N_2439,N_1871,N_1337);
nand U2440 (N_2440,N_1749,N_1837);
nand U2441 (N_2441,N_1357,N_1584);
and U2442 (N_2442,N_1626,N_1802);
nand U2443 (N_2443,N_1427,N_1571);
xor U2444 (N_2444,N_1666,N_1538);
xnor U2445 (N_2445,N_1458,N_1777);
nand U2446 (N_2446,N_1807,N_1596);
or U2447 (N_2447,N_1356,N_1809);
and U2448 (N_2448,N_1670,N_1599);
nand U2449 (N_2449,N_1471,N_1411);
nand U2450 (N_2450,N_1757,N_1630);
nor U2451 (N_2451,N_1680,N_1372);
nor U2452 (N_2452,N_1798,N_1408);
nor U2453 (N_2453,N_1603,N_1627);
and U2454 (N_2454,N_1541,N_1614);
xnor U2455 (N_2455,N_1442,N_1703);
nor U2456 (N_2456,N_1663,N_1448);
and U2457 (N_2457,N_1350,N_1628);
and U2458 (N_2458,N_1725,N_1447);
nand U2459 (N_2459,N_1689,N_1529);
xnor U2460 (N_2460,N_1792,N_1771);
xor U2461 (N_2461,N_1532,N_1700);
nand U2462 (N_2462,N_1777,N_1742);
or U2463 (N_2463,N_1482,N_1842);
nor U2464 (N_2464,N_1310,N_1321);
or U2465 (N_2465,N_1803,N_1710);
nor U2466 (N_2466,N_1349,N_1784);
nor U2467 (N_2467,N_1773,N_1293);
xnor U2468 (N_2468,N_1825,N_1734);
nand U2469 (N_2469,N_1291,N_1705);
or U2470 (N_2470,N_1304,N_1326);
nor U2471 (N_2471,N_1269,N_1753);
and U2472 (N_2472,N_1352,N_1442);
or U2473 (N_2473,N_1580,N_1828);
xor U2474 (N_2474,N_1787,N_1685);
and U2475 (N_2475,N_1732,N_1314);
nor U2476 (N_2476,N_1553,N_1347);
xor U2477 (N_2477,N_1304,N_1611);
nand U2478 (N_2478,N_1432,N_1582);
and U2479 (N_2479,N_1770,N_1561);
and U2480 (N_2480,N_1444,N_1295);
and U2481 (N_2481,N_1271,N_1710);
and U2482 (N_2482,N_1386,N_1488);
nand U2483 (N_2483,N_1872,N_1259);
and U2484 (N_2484,N_1388,N_1304);
nand U2485 (N_2485,N_1835,N_1828);
nor U2486 (N_2486,N_1848,N_1547);
nor U2487 (N_2487,N_1498,N_1807);
and U2488 (N_2488,N_1526,N_1395);
nor U2489 (N_2489,N_1844,N_1414);
nor U2490 (N_2490,N_1796,N_1790);
and U2491 (N_2491,N_1655,N_1565);
or U2492 (N_2492,N_1610,N_1444);
and U2493 (N_2493,N_1747,N_1768);
or U2494 (N_2494,N_1293,N_1539);
and U2495 (N_2495,N_1530,N_1778);
nor U2496 (N_2496,N_1796,N_1491);
and U2497 (N_2497,N_1707,N_1548);
xnor U2498 (N_2498,N_1381,N_1710);
nor U2499 (N_2499,N_1372,N_1820);
or U2500 (N_2500,N_2033,N_2323);
xor U2501 (N_2501,N_2247,N_2248);
nand U2502 (N_2502,N_2147,N_2173);
or U2503 (N_2503,N_2051,N_2488);
or U2504 (N_2504,N_2151,N_2338);
xnor U2505 (N_2505,N_2220,N_2039);
nand U2506 (N_2506,N_2295,N_2257);
nand U2507 (N_2507,N_2028,N_2397);
or U2508 (N_2508,N_2399,N_2358);
nand U2509 (N_2509,N_1960,N_2268);
and U2510 (N_2510,N_2105,N_1987);
or U2511 (N_2511,N_2064,N_2393);
nor U2512 (N_2512,N_2158,N_2049);
xnor U2513 (N_2513,N_2265,N_1980);
and U2514 (N_2514,N_1941,N_1938);
and U2515 (N_2515,N_2448,N_2102);
and U2516 (N_2516,N_1890,N_2355);
nand U2517 (N_2517,N_2334,N_2450);
or U2518 (N_2518,N_2080,N_2078);
nand U2519 (N_2519,N_2086,N_2280);
nand U2520 (N_2520,N_2189,N_2202);
or U2521 (N_2521,N_2308,N_2255);
and U2522 (N_2522,N_2238,N_2429);
and U2523 (N_2523,N_2228,N_1956);
and U2524 (N_2524,N_2481,N_2412);
or U2525 (N_2525,N_2035,N_2050);
or U2526 (N_2526,N_1933,N_1889);
or U2527 (N_2527,N_2281,N_2328);
nor U2528 (N_2528,N_2146,N_2004);
xnor U2529 (N_2529,N_2266,N_2366);
nand U2530 (N_2530,N_2377,N_1962);
nor U2531 (N_2531,N_1986,N_2071);
xnor U2532 (N_2532,N_2285,N_2075);
and U2533 (N_2533,N_2458,N_2074);
nor U2534 (N_2534,N_2212,N_2394);
or U2535 (N_2535,N_1882,N_2110);
or U2536 (N_2536,N_2474,N_2020);
xnor U2537 (N_2537,N_2201,N_2204);
nor U2538 (N_2538,N_2341,N_2207);
and U2539 (N_2539,N_2083,N_1918);
nand U2540 (N_2540,N_1920,N_2188);
nand U2541 (N_2541,N_2123,N_2109);
nor U2542 (N_2542,N_2104,N_1884);
or U2543 (N_2543,N_1954,N_2421);
nor U2544 (N_2544,N_2413,N_2274);
and U2545 (N_2545,N_2335,N_2000);
and U2546 (N_2546,N_1886,N_1879);
or U2547 (N_2547,N_2427,N_2239);
xor U2548 (N_2548,N_1963,N_2008);
xnor U2549 (N_2549,N_2447,N_1896);
or U2550 (N_2550,N_1924,N_1952);
nor U2551 (N_2551,N_2246,N_2398);
and U2552 (N_2552,N_2015,N_2292);
or U2553 (N_2553,N_2116,N_2057);
xnor U2554 (N_2554,N_2009,N_2137);
xnor U2555 (N_2555,N_1935,N_2289);
xnor U2556 (N_2556,N_2085,N_2478);
nor U2557 (N_2557,N_2061,N_1922);
xnor U2558 (N_2558,N_2479,N_2079);
nand U2559 (N_2559,N_2496,N_2164);
xnor U2560 (N_2560,N_2376,N_2172);
nand U2561 (N_2561,N_2345,N_1950);
and U2562 (N_2562,N_2272,N_1978);
and U2563 (N_2563,N_1985,N_2311);
nand U2564 (N_2564,N_2305,N_2143);
and U2565 (N_2565,N_2245,N_1901);
and U2566 (N_2566,N_2254,N_2475);
nand U2567 (N_2567,N_2237,N_1939);
xnor U2568 (N_2568,N_2203,N_2395);
and U2569 (N_2569,N_1965,N_2271);
nand U2570 (N_2570,N_2495,N_1931);
xnor U2571 (N_2571,N_2416,N_1923);
nand U2572 (N_2572,N_2296,N_2419);
nor U2573 (N_2573,N_2144,N_2310);
and U2574 (N_2574,N_2286,N_2177);
nand U2575 (N_2575,N_2457,N_2312);
or U2576 (N_2576,N_2042,N_2122);
xnor U2577 (N_2577,N_1971,N_2499);
nand U2578 (N_2578,N_2263,N_2026);
nand U2579 (N_2579,N_2170,N_2279);
xnor U2580 (N_2580,N_2152,N_2477);
or U2581 (N_2581,N_2016,N_2317);
or U2582 (N_2582,N_1947,N_2411);
or U2583 (N_2583,N_2396,N_2389);
nand U2584 (N_2584,N_2476,N_2215);
xnor U2585 (N_2585,N_1906,N_2277);
xor U2586 (N_2586,N_2364,N_2169);
nand U2587 (N_2587,N_2002,N_2131);
xor U2588 (N_2588,N_2387,N_1903);
and U2589 (N_2589,N_2340,N_2150);
xnor U2590 (N_2590,N_2187,N_2357);
or U2591 (N_2591,N_2494,N_2430);
or U2592 (N_2592,N_2302,N_2362);
nand U2593 (N_2593,N_1984,N_2480);
xor U2594 (N_2594,N_2270,N_2017);
and U2595 (N_2595,N_1899,N_2040);
or U2596 (N_2596,N_2249,N_2134);
xnor U2597 (N_2597,N_2052,N_2346);
or U2598 (N_2598,N_2185,N_1940);
xor U2599 (N_2599,N_1902,N_2153);
and U2600 (N_2600,N_2044,N_2375);
nor U2601 (N_2601,N_2225,N_2114);
nor U2602 (N_2602,N_2157,N_2120);
xor U2603 (N_2603,N_2350,N_2252);
and U2604 (N_2604,N_2463,N_2130);
and U2605 (N_2605,N_2363,N_2365);
or U2606 (N_2606,N_1898,N_2351);
nor U2607 (N_2607,N_2227,N_1991);
and U2608 (N_2608,N_1885,N_1976);
and U2609 (N_2609,N_1988,N_2337);
nand U2610 (N_2610,N_2330,N_2007);
or U2611 (N_2611,N_2210,N_2234);
xor U2612 (N_2612,N_2165,N_2195);
or U2613 (N_2613,N_2062,N_2233);
nor U2614 (N_2614,N_2031,N_2339);
nor U2615 (N_2615,N_2367,N_2417);
and U2616 (N_2616,N_1911,N_2406);
xor U2617 (N_2617,N_2038,N_2149);
or U2618 (N_2618,N_2344,N_2293);
xnor U2619 (N_2619,N_2409,N_1883);
nand U2620 (N_2620,N_2467,N_2069);
or U2621 (N_2621,N_2382,N_2168);
xor U2622 (N_2622,N_2403,N_2320);
nand U2623 (N_2623,N_1995,N_2163);
nand U2624 (N_2624,N_2091,N_2348);
xnor U2625 (N_2625,N_2063,N_1977);
nand U2626 (N_2626,N_2156,N_2390);
nor U2627 (N_2627,N_1887,N_2036);
nand U2628 (N_2628,N_2118,N_2297);
nor U2629 (N_2629,N_1925,N_1996);
xor U2630 (N_2630,N_2332,N_2258);
xor U2631 (N_2631,N_2283,N_2013);
and U2632 (N_2632,N_1937,N_2298);
or U2633 (N_2633,N_2162,N_2371);
nor U2634 (N_2634,N_2441,N_2360);
or U2635 (N_2635,N_2089,N_2353);
or U2636 (N_2636,N_2464,N_2370);
xnor U2637 (N_2637,N_2384,N_2326);
or U2638 (N_2638,N_2001,N_2456);
nand U2639 (N_2639,N_2461,N_2401);
nor U2640 (N_2640,N_2282,N_2423);
nor U2641 (N_2641,N_2445,N_2094);
or U2642 (N_2642,N_2453,N_2096);
or U2643 (N_2643,N_2253,N_2073);
or U2644 (N_2644,N_2099,N_2192);
xor U2645 (N_2645,N_2030,N_1973);
nor U2646 (N_2646,N_1921,N_1893);
and U2647 (N_2647,N_2113,N_2194);
or U2648 (N_2648,N_1982,N_2490);
nor U2649 (N_2649,N_2327,N_2487);
nand U2650 (N_2650,N_1997,N_2438);
or U2651 (N_2651,N_2489,N_2313);
xor U2652 (N_2652,N_2223,N_2361);
nor U2653 (N_2653,N_2316,N_2444);
nor U2654 (N_2654,N_2299,N_2003);
nand U2655 (N_2655,N_1992,N_2431);
or U2656 (N_2656,N_2442,N_2404);
or U2657 (N_2657,N_1930,N_2267);
nor U2658 (N_2658,N_2161,N_1949);
xnor U2659 (N_2659,N_2133,N_2378);
and U2660 (N_2660,N_2288,N_1964);
or U2661 (N_2661,N_1989,N_1958);
or U2662 (N_2662,N_2325,N_2300);
or U2663 (N_2663,N_2333,N_1934);
and U2664 (N_2664,N_2059,N_2446);
xor U2665 (N_2665,N_2352,N_2392);
or U2666 (N_2666,N_1913,N_2428);
nor U2667 (N_2667,N_2136,N_1929);
or U2668 (N_2668,N_2218,N_1951);
or U2669 (N_2669,N_2386,N_2148);
and U2670 (N_2670,N_2193,N_2180);
and U2671 (N_2671,N_2088,N_2055);
xnor U2672 (N_2672,N_2471,N_2097);
xnor U2673 (N_2673,N_2451,N_2251);
nor U2674 (N_2674,N_2385,N_1888);
or U2675 (N_2675,N_2183,N_2294);
xnor U2676 (N_2676,N_2132,N_1990);
nand U2677 (N_2677,N_2236,N_2243);
nor U2678 (N_2678,N_1919,N_2229);
xnor U2679 (N_2679,N_2287,N_1926);
nand U2680 (N_2680,N_2190,N_2372);
or U2681 (N_2681,N_2273,N_2250);
xnor U2682 (N_2682,N_2410,N_1975);
nand U2683 (N_2683,N_2117,N_2373);
xnor U2684 (N_2684,N_2459,N_2029);
nand U2685 (N_2685,N_1946,N_2437);
nor U2686 (N_2686,N_2124,N_2432);
and U2687 (N_2687,N_2200,N_2082);
nor U2688 (N_2688,N_2244,N_2126);
nor U2689 (N_2689,N_2470,N_2084);
and U2690 (N_2690,N_2206,N_2145);
and U2691 (N_2691,N_2154,N_2402);
or U2692 (N_2692,N_2443,N_2435);
and U2693 (N_2693,N_2240,N_1932);
nor U2694 (N_2694,N_2424,N_1917);
and U2695 (N_2695,N_2066,N_2107);
xnor U2696 (N_2696,N_1944,N_1905);
xor U2697 (N_2697,N_2485,N_2213);
or U2698 (N_2698,N_2418,N_2301);
or U2699 (N_2699,N_2196,N_1936);
or U2700 (N_2700,N_1881,N_2216);
nand U2701 (N_2701,N_2019,N_1910);
nor U2702 (N_2702,N_2482,N_2174);
nand U2703 (N_2703,N_2208,N_2095);
nand U2704 (N_2704,N_2491,N_2127);
nor U2705 (N_2705,N_2129,N_2211);
xnor U2706 (N_2706,N_2226,N_1877);
nor U2707 (N_2707,N_2291,N_2359);
xnor U2708 (N_2708,N_2103,N_2199);
nor U2709 (N_2709,N_2065,N_2436);
and U2710 (N_2710,N_2100,N_1928);
and U2711 (N_2711,N_1892,N_2006);
or U2712 (N_2712,N_1967,N_2497);
and U2713 (N_2713,N_2492,N_2415);
nor U2714 (N_2714,N_2259,N_2224);
or U2715 (N_2715,N_2336,N_2101);
xor U2716 (N_2716,N_2264,N_2381);
or U2717 (N_2717,N_2354,N_2262);
xnor U2718 (N_2718,N_1943,N_2021);
or U2719 (N_2719,N_2242,N_2349);
nor U2720 (N_2720,N_2235,N_2391);
and U2721 (N_2721,N_1957,N_2053);
xor U2722 (N_2722,N_1876,N_2261);
nand U2723 (N_2723,N_2166,N_2139);
xnor U2724 (N_2724,N_2454,N_2462);
nor U2725 (N_2725,N_2369,N_2037);
xnor U2726 (N_2726,N_2452,N_2414);
or U2727 (N_2727,N_2181,N_1959);
or U2728 (N_2728,N_2024,N_1968);
and U2729 (N_2729,N_2388,N_2011);
nand U2730 (N_2730,N_2440,N_2045);
nand U2731 (N_2731,N_2449,N_2425);
xor U2732 (N_2732,N_2290,N_1908);
or U2733 (N_2733,N_2047,N_2138);
nand U2734 (N_2734,N_2275,N_2434);
nor U2735 (N_2735,N_1999,N_2380);
nand U2736 (N_2736,N_2022,N_2058);
nand U2737 (N_2737,N_2217,N_1961);
and U2738 (N_2738,N_2056,N_2422);
xor U2739 (N_2739,N_2314,N_2178);
nand U2740 (N_2740,N_2171,N_2405);
xnor U2741 (N_2741,N_2315,N_2175);
nand U2742 (N_2742,N_2324,N_2232);
nand U2743 (N_2743,N_2407,N_2230);
nor U2744 (N_2744,N_2121,N_2303);
nand U2745 (N_2745,N_2374,N_2018);
xnor U2746 (N_2746,N_2379,N_2486);
and U2747 (N_2747,N_2400,N_1914);
xor U2748 (N_2748,N_2306,N_1875);
xor U2749 (N_2749,N_2222,N_2012);
or U2750 (N_2750,N_2342,N_1948);
nand U2751 (N_2751,N_1904,N_2241);
nand U2752 (N_2752,N_2115,N_2420);
nand U2753 (N_2753,N_2408,N_2276);
or U2754 (N_2754,N_2093,N_2209);
nor U2755 (N_2755,N_2135,N_2319);
xnor U2756 (N_2756,N_1979,N_2460);
nor U2757 (N_2757,N_2119,N_1927);
xor U2758 (N_2758,N_2090,N_2014);
xnor U2759 (N_2759,N_1945,N_2125);
and U2760 (N_2760,N_2067,N_2128);
xor U2761 (N_2761,N_1916,N_1894);
xor U2762 (N_2762,N_2068,N_2112);
nand U2763 (N_2763,N_2005,N_2484);
nor U2764 (N_2764,N_2347,N_2191);
nand U2765 (N_2765,N_2160,N_2010);
or U2766 (N_2766,N_2142,N_2186);
xnor U2767 (N_2767,N_2284,N_2046);
nor U2768 (N_2768,N_2219,N_1983);
xnor U2769 (N_2769,N_2077,N_1880);
and U2770 (N_2770,N_2081,N_2155);
nor U2771 (N_2771,N_2060,N_2214);
nor U2772 (N_2772,N_1895,N_2304);
and U2773 (N_2773,N_2072,N_2309);
and U2774 (N_2774,N_2455,N_1966);
and U2775 (N_2775,N_2034,N_1955);
xnor U2776 (N_2776,N_2111,N_2176);
nor U2777 (N_2777,N_2329,N_2098);
or U2778 (N_2778,N_2269,N_2483);
nand U2779 (N_2779,N_1878,N_1993);
nor U2780 (N_2780,N_2184,N_2179);
xor U2781 (N_2781,N_2473,N_2433);
nor U2782 (N_2782,N_1942,N_1891);
or U2783 (N_2783,N_2322,N_2256);
xor U2784 (N_2784,N_2321,N_2032);
nand U2785 (N_2785,N_2498,N_2043);
nand U2786 (N_2786,N_2159,N_2025);
xnor U2787 (N_2787,N_2469,N_2106);
nor U2788 (N_2788,N_2197,N_2278);
nor U2789 (N_2789,N_2041,N_1969);
xnor U2790 (N_2790,N_1974,N_1912);
xor U2791 (N_2791,N_2054,N_2356);
nor U2792 (N_2792,N_2318,N_1994);
xnor U2793 (N_2793,N_2383,N_2468);
nor U2794 (N_2794,N_2260,N_2472);
nand U2795 (N_2795,N_2466,N_1915);
nand U2796 (N_2796,N_2205,N_1909);
and U2797 (N_2797,N_2141,N_1907);
nand U2798 (N_2798,N_2076,N_2221);
nor U2799 (N_2799,N_2231,N_2331);
nand U2800 (N_2800,N_2198,N_2087);
nand U2801 (N_2801,N_1981,N_2426);
xor U2802 (N_2802,N_2108,N_2368);
or U2803 (N_2803,N_1970,N_2465);
nor U2804 (N_2804,N_2140,N_2182);
nand U2805 (N_2805,N_2307,N_1998);
and U2806 (N_2806,N_2167,N_2493);
nor U2807 (N_2807,N_2023,N_2027);
and U2808 (N_2808,N_2048,N_1897);
nor U2809 (N_2809,N_2092,N_2343);
xor U2810 (N_2810,N_2439,N_1953);
or U2811 (N_2811,N_1972,N_1900);
nor U2812 (N_2812,N_2070,N_2231);
and U2813 (N_2813,N_2335,N_1996);
nor U2814 (N_2814,N_1894,N_2212);
or U2815 (N_2815,N_2269,N_2493);
nand U2816 (N_2816,N_2447,N_2324);
and U2817 (N_2817,N_1899,N_2174);
nor U2818 (N_2818,N_2474,N_2001);
xnor U2819 (N_2819,N_1901,N_2353);
nor U2820 (N_2820,N_2107,N_2480);
nand U2821 (N_2821,N_1961,N_2108);
nor U2822 (N_2822,N_2414,N_1922);
xor U2823 (N_2823,N_2233,N_2482);
or U2824 (N_2824,N_2146,N_2348);
nand U2825 (N_2825,N_1909,N_1971);
xnor U2826 (N_2826,N_1988,N_2249);
nand U2827 (N_2827,N_2428,N_2184);
xor U2828 (N_2828,N_1911,N_2467);
and U2829 (N_2829,N_2179,N_1890);
nor U2830 (N_2830,N_2316,N_1938);
nor U2831 (N_2831,N_2283,N_2082);
nand U2832 (N_2832,N_2084,N_2092);
and U2833 (N_2833,N_2023,N_2164);
nand U2834 (N_2834,N_2161,N_2084);
or U2835 (N_2835,N_2463,N_2333);
nand U2836 (N_2836,N_2397,N_2225);
xnor U2837 (N_2837,N_2495,N_2146);
or U2838 (N_2838,N_2313,N_2225);
nor U2839 (N_2839,N_1978,N_2354);
nand U2840 (N_2840,N_2230,N_2063);
and U2841 (N_2841,N_2151,N_2423);
xnor U2842 (N_2842,N_2278,N_2224);
and U2843 (N_2843,N_2258,N_1929);
nor U2844 (N_2844,N_2157,N_2464);
and U2845 (N_2845,N_1939,N_2370);
nand U2846 (N_2846,N_2333,N_2246);
nand U2847 (N_2847,N_2486,N_2194);
and U2848 (N_2848,N_2202,N_1915);
nor U2849 (N_2849,N_2359,N_2240);
and U2850 (N_2850,N_2283,N_1995);
nor U2851 (N_2851,N_2061,N_2115);
xor U2852 (N_2852,N_2281,N_2312);
nand U2853 (N_2853,N_2071,N_2243);
xnor U2854 (N_2854,N_2099,N_2362);
xnor U2855 (N_2855,N_2444,N_2345);
nor U2856 (N_2856,N_2328,N_2036);
and U2857 (N_2857,N_2108,N_2084);
xnor U2858 (N_2858,N_2261,N_2494);
xor U2859 (N_2859,N_2164,N_1964);
and U2860 (N_2860,N_2230,N_1984);
nand U2861 (N_2861,N_2117,N_2171);
nand U2862 (N_2862,N_2478,N_2258);
nand U2863 (N_2863,N_1986,N_2245);
or U2864 (N_2864,N_2223,N_2115);
nand U2865 (N_2865,N_2136,N_2112);
or U2866 (N_2866,N_2454,N_2333);
xor U2867 (N_2867,N_2059,N_1875);
nor U2868 (N_2868,N_2134,N_1935);
nand U2869 (N_2869,N_2294,N_2251);
nand U2870 (N_2870,N_1960,N_1998);
xor U2871 (N_2871,N_2364,N_1993);
nand U2872 (N_2872,N_2238,N_2071);
and U2873 (N_2873,N_2289,N_1980);
xnor U2874 (N_2874,N_2493,N_2240);
nor U2875 (N_2875,N_2377,N_2418);
nand U2876 (N_2876,N_2230,N_2169);
and U2877 (N_2877,N_2143,N_2442);
or U2878 (N_2878,N_2369,N_2428);
xnor U2879 (N_2879,N_2181,N_2388);
xor U2880 (N_2880,N_1973,N_2431);
or U2881 (N_2881,N_2325,N_1922);
nand U2882 (N_2882,N_2348,N_2499);
or U2883 (N_2883,N_2165,N_2172);
or U2884 (N_2884,N_2006,N_2261);
and U2885 (N_2885,N_2390,N_2471);
and U2886 (N_2886,N_2445,N_2181);
nor U2887 (N_2887,N_2143,N_1996);
nand U2888 (N_2888,N_2453,N_2408);
and U2889 (N_2889,N_2117,N_2330);
nand U2890 (N_2890,N_2220,N_2060);
and U2891 (N_2891,N_2469,N_1923);
xnor U2892 (N_2892,N_2017,N_2313);
or U2893 (N_2893,N_2000,N_1936);
and U2894 (N_2894,N_2156,N_2292);
or U2895 (N_2895,N_2076,N_2147);
and U2896 (N_2896,N_2095,N_2243);
nand U2897 (N_2897,N_2314,N_2138);
or U2898 (N_2898,N_1937,N_2134);
nand U2899 (N_2899,N_2419,N_2082);
xnor U2900 (N_2900,N_2095,N_1919);
xor U2901 (N_2901,N_1881,N_1895);
xor U2902 (N_2902,N_2131,N_2337);
and U2903 (N_2903,N_2495,N_1920);
and U2904 (N_2904,N_1987,N_2273);
nor U2905 (N_2905,N_1948,N_2307);
nor U2906 (N_2906,N_2464,N_1960);
nor U2907 (N_2907,N_2236,N_2297);
and U2908 (N_2908,N_2137,N_1942);
and U2909 (N_2909,N_2065,N_2282);
or U2910 (N_2910,N_2063,N_2409);
or U2911 (N_2911,N_2218,N_1893);
xor U2912 (N_2912,N_2492,N_2071);
and U2913 (N_2913,N_2400,N_2198);
nor U2914 (N_2914,N_1944,N_2239);
or U2915 (N_2915,N_2291,N_1935);
xor U2916 (N_2916,N_1949,N_2317);
nand U2917 (N_2917,N_1907,N_1916);
or U2918 (N_2918,N_2471,N_2201);
xnor U2919 (N_2919,N_1988,N_2305);
and U2920 (N_2920,N_2162,N_2087);
nand U2921 (N_2921,N_2097,N_2095);
xor U2922 (N_2922,N_2313,N_1933);
and U2923 (N_2923,N_2369,N_2032);
nor U2924 (N_2924,N_2144,N_1879);
xor U2925 (N_2925,N_1906,N_2447);
and U2926 (N_2926,N_2422,N_2025);
or U2927 (N_2927,N_2098,N_2357);
nand U2928 (N_2928,N_2356,N_2460);
nand U2929 (N_2929,N_2213,N_1946);
xnor U2930 (N_2930,N_2116,N_1962);
and U2931 (N_2931,N_2282,N_2011);
nand U2932 (N_2932,N_2200,N_2418);
xor U2933 (N_2933,N_2133,N_1995);
and U2934 (N_2934,N_1934,N_2296);
or U2935 (N_2935,N_2324,N_2268);
or U2936 (N_2936,N_2369,N_2186);
and U2937 (N_2937,N_2333,N_2397);
xor U2938 (N_2938,N_2465,N_2067);
nand U2939 (N_2939,N_2437,N_2267);
and U2940 (N_2940,N_2395,N_2420);
xnor U2941 (N_2941,N_2210,N_2196);
or U2942 (N_2942,N_2038,N_2206);
nor U2943 (N_2943,N_2084,N_2273);
and U2944 (N_2944,N_2006,N_2215);
or U2945 (N_2945,N_2449,N_2144);
and U2946 (N_2946,N_2077,N_2181);
nor U2947 (N_2947,N_1879,N_2375);
or U2948 (N_2948,N_2304,N_2205);
or U2949 (N_2949,N_1960,N_2065);
xor U2950 (N_2950,N_2407,N_2457);
nand U2951 (N_2951,N_2290,N_2292);
nand U2952 (N_2952,N_2391,N_1891);
and U2953 (N_2953,N_2377,N_2332);
and U2954 (N_2954,N_2383,N_2437);
nand U2955 (N_2955,N_2154,N_1932);
or U2956 (N_2956,N_2185,N_2003);
nand U2957 (N_2957,N_2339,N_2440);
and U2958 (N_2958,N_1997,N_1877);
xor U2959 (N_2959,N_1977,N_2339);
nand U2960 (N_2960,N_1920,N_2375);
xor U2961 (N_2961,N_2057,N_2218);
xor U2962 (N_2962,N_2411,N_2247);
nor U2963 (N_2963,N_2441,N_2280);
xor U2964 (N_2964,N_2425,N_2457);
nand U2965 (N_2965,N_1926,N_2478);
and U2966 (N_2966,N_1953,N_2312);
nor U2967 (N_2967,N_2149,N_2075);
nand U2968 (N_2968,N_2078,N_2175);
xor U2969 (N_2969,N_2477,N_2408);
or U2970 (N_2970,N_1887,N_2440);
nand U2971 (N_2971,N_2014,N_2013);
nor U2972 (N_2972,N_2053,N_2455);
xnor U2973 (N_2973,N_2196,N_2069);
nor U2974 (N_2974,N_2279,N_2041);
or U2975 (N_2975,N_2352,N_2183);
and U2976 (N_2976,N_1965,N_2156);
nor U2977 (N_2977,N_2151,N_2436);
nand U2978 (N_2978,N_2073,N_1988);
or U2979 (N_2979,N_2370,N_1978);
and U2980 (N_2980,N_2313,N_2298);
nor U2981 (N_2981,N_2052,N_2451);
nand U2982 (N_2982,N_1903,N_2260);
nor U2983 (N_2983,N_2467,N_2266);
and U2984 (N_2984,N_2002,N_2498);
nor U2985 (N_2985,N_2235,N_2071);
or U2986 (N_2986,N_2258,N_1877);
and U2987 (N_2987,N_2447,N_2065);
or U2988 (N_2988,N_1966,N_1993);
nand U2989 (N_2989,N_1901,N_2389);
xnor U2990 (N_2990,N_1898,N_2297);
or U2991 (N_2991,N_2090,N_1920);
or U2992 (N_2992,N_2173,N_2263);
nor U2993 (N_2993,N_2439,N_2280);
xor U2994 (N_2994,N_2268,N_2205);
or U2995 (N_2995,N_2384,N_2327);
nand U2996 (N_2996,N_2493,N_2004);
and U2997 (N_2997,N_1966,N_2467);
nand U2998 (N_2998,N_2329,N_2068);
nor U2999 (N_2999,N_2482,N_2226);
xor U3000 (N_3000,N_2085,N_2032);
xnor U3001 (N_3001,N_1934,N_2201);
nand U3002 (N_3002,N_2282,N_2330);
nor U3003 (N_3003,N_1927,N_1887);
or U3004 (N_3004,N_2088,N_1914);
and U3005 (N_3005,N_1952,N_2046);
xor U3006 (N_3006,N_2279,N_2472);
or U3007 (N_3007,N_2142,N_2403);
xnor U3008 (N_3008,N_2312,N_2163);
xor U3009 (N_3009,N_2420,N_1951);
nor U3010 (N_3010,N_2049,N_2156);
xnor U3011 (N_3011,N_2272,N_2233);
and U3012 (N_3012,N_2349,N_2180);
xor U3013 (N_3013,N_2058,N_2056);
nor U3014 (N_3014,N_2124,N_1902);
and U3015 (N_3015,N_2415,N_2125);
xor U3016 (N_3016,N_2482,N_2328);
and U3017 (N_3017,N_2044,N_2289);
and U3018 (N_3018,N_1894,N_2308);
and U3019 (N_3019,N_2401,N_2163);
nand U3020 (N_3020,N_2229,N_2312);
nor U3021 (N_3021,N_1902,N_2412);
nor U3022 (N_3022,N_2396,N_2484);
or U3023 (N_3023,N_2275,N_2091);
xnor U3024 (N_3024,N_2135,N_2491);
xnor U3025 (N_3025,N_2132,N_2106);
nand U3026 (N_3026,N_2238,N_2325);
xor U3027 (N_3027,N_2174,N_1992);
or U3028 (N_3028,N_2030,N_2408);
xor U3029 (N_3029,N_1932,N_2482);
or U3030 (N_3030,N_2078,N_2230);
nor U3031 (N_3031,N_2123,N_2253);
and U3032 (N_3032,N_2171,N_2005);
xnor U3033 (N_3033,N_2298,N_2305);
and U3034 (N_3034,N_2013,N_2046);
and U3035 (N_3035,N_2481,N_1877);
or U3036 (N_3036,N_2422,N_2420);
nand U3037 (N_3037,N_2067,N_2425);
nand U3038 (N_3038,N_2207,N_2071);
nand U3039 (N_3039,N_2315,N_2255);
and U3040 (N_3040,N_2463,N_1952);
or U3041 (N_3041,N_2227,N_2333);
and U3042 (N_3042,N_2197,N_2087);
and U3043 (N_3043,N_2035,N_2339);
and U3044 (N_3044,N_2015,N_2471);
nor U3045 (N_3045,N_1959,N_2348);
nor U3046 (N_3046,N_2071,N_2387);
or U3047 (N_3047,N_2482,N_2079);
nor U3048 (N_3048,N_2357,N_2102);
or U3049 (N_3049,N_2330,N_2081);
and U3050 (N_3050,N_2220,N_2464);
nand U3051 (N_3051,N_2237,N_2313);
and U3052 (N_3052,N_2190,N_2145);
nand U3053 (N_3053,N_2467,N_2459);
and U3054 (N_3054,N_2122,N_1897);
and U3055 (N_3055,N_2478,N_2076);
or U3056 (N_3056,N_2362,N_2012);
xnor U3057 (N_3057,N_2354,N_1952);
nand U3058 (N_3058,N_2446,N_2448);
nand U3059 (N_3059,N_2490,N_2378);
xnor U3060 (N_3060,N_2479,N_1961);
nor U3061 (N_3061,N_2353,N_2166);
nand U3062 (N_3062,N_1985,N_2035);
nand U3063 (N_3063,N_2330,N_2429);
nand U3064 (N_3064,N_2302,N_2357);
nor U3065 (N_3065,N_2470,N_1954);
nand U3066 (N_3066,N_2143,N_1922);
and U3067 (N_3067,N_2191,N_1885);
nor U3068 (N_3068,N_2317,N_1957);
nand U3069 (N_3069,N_2231,N_2207);
or U3070 (N_3070,N_1948,N_2408);
xor U3071 (N_3071,N_2079,N_1902);
nor U3072 (N_3072,N_2271,N_2196);
and U3073 (N_3073,N_2405,N_1981);
or U3074 (N_3074,N_2406,N_2377);
or U3075 (N_3075,N_2054,N_2498);
or U3076 (N_3076,N_2251,N_2094);
nor U3077 (N_3077,N_1926,N_1923);
xor U3078 (N_3078,N_2323,N_2471);
nor U3079 (N_3079,N_2464,N_1904);
nand U3080 (N_3080,N_2367,N_2038);
nand U3081 (N_3081,N_2229,N_2166);
nand U3082 (N_3082,N_2162,N_2344);
and U3083 (N_3083,N_1979,N_2495);
or U3084 (N_3084,N_1927,N_2474);
or U3085 (N_3085,N_2428,N_1983);
xnor U3086 (N_3086,N_2273,N_2269);
xor U3087 (N_3087,N_2004,N_2065);
nand U3088 (N_3088,N_2071,N_2398);
or U3089 (N_3089,N_1978,N_2379);
and U3090 (N_3090,N_2288,N_2243);
and U3091 (N_3091,N_2012,N_2107);
or U3092 (N_3092,N_2437,N_2300);
xor U3093 (N_3093,N_1948,N_2040);
nand U3094 (N_3094,N_2451,N_2199);
and U3095 (N_3095,N_2352,N_2379);
nand U3096 (N_3096,N_2197,N_1961);
and U3097 (N_3097,N_2146,N_2248);
nand U3098 (N_3098,N_2100,N_2015);
xnor U3099 (N_3099,N_1956,N_2251);
xnor U3100 (N_3100,N_2429,N_1973);
or U3101 (N_3101,N_2022,N_2322);
nand U3102 (N_3102,N_2246,N_2015);
nor U3103 (N_3103,N_2381,N_2162);
nand U3104 (N_3104,N_1910,N_2297);
nand U3105 (N_3105,N_2417,N_2343);
and U3106 (N_3106,N_2379,N_2443);
or U3107 (N_3107,N_2164,N_1991);
and U3108 (N_3108,N_2055,N_2133);
nor U3109 (N_3109,N_2035,N_2384);
xor U3110 (N_3110,N_2020,N_2143);
or U3111 (N_3111,N_2180,N_1936);
nand U3112 (N_3112,N_2283,N_2108);
or U3113 (N_3113,N_2433,N_1945);
xor U3114 (N_3114,N_2055,N_2273);
or U3115 (N_3115,N_2315,N_1912);
or U3116 (N_3116,N_2226,N_2043);
nand U3117 (N_3117,N_2391,N_1964);
and U3118 (N_3118,N_2457,N_2430);
and U3119 (N_3119,N_2197,N_2405);
and U3120 (N_3120,N_2420,N_2030);
xnor U3121 (N_3121,N_2164,N_2315);
nor U3122 (N_3122,N_2426,N_2149);
or U3123 (N_3123,N_2400,N_2080);
or U3124 (N_3124,N_2287,N_2285);
and U3125 (N_3125,N_2733,N_2746);
or U3126 (N_3126,N_2742,N_2951);
nor U3127 (N_3127,N_2639,N_2881);
nor U3128 (N_3128,N_2520,N_2936);
xnor U3129 (N_3129,N_2553,N_2605);
nor U3130 (N_3130,N_3111,N_2863);
nand U3131 (N_3131,N_3079,N_2775);
or U3132 (N_3132,N_2523,N_2714);
nor U3133 (N_3133,N_3121,N_3026);
xnor U3134 (N_3134,N_2508,N_2877);
nor U3135 (N_3135,N_2716,N_2814);
nand U3136 (N_3136,N_2680,N_2654);
nor U3137 (N_3137,N_2817,N_2942);
or U3138 (N_3138,N_3073,N_2768);
nor U3139 (N_3139,N_2686,N_2901);
or U3140 (N_3140,N_2862,N_2671);
xnor U3141 (N_3141,N_2699,N_2771);
nand U3142 (N_3142,N_2601,N_2642);
or U3143 (N_3143,N_2609,N_2801);
nor U3144 (N_3144,N_2596,N_2736);
or U3145 (N_3145,N_2792,N_2777);
or U3146 (N_3146,N_2574,N_2581);
xor U3147 (N_3147,N_2712,N_2667);
nand U3148 (N_3148,N_2916,N_3081);
xor U3149 (N_3149,N_2846,N_2859);
xor U3150 (N_3150,N_2961,N_3066);
nand U3151 (N_3151,N_3008,N_2891);
or U3152 (N_3152,N_3052,N_2614);
nor U3153 (N_3153,N_2977,N_2715);
or U3154 (N_3154,N_2630,N_3041);
xor U3155 (N_3155,N_2578,N_3013);
and U3156 (N_3156,N_2935,N_2782);
xor U3157 (N_3157,N_2602,N_3090);
or U3158 (N_3158,N_3064,N_3037);
xor U3159 (N_3159,N_2845,N_2926);
or U3160 (N_3160,N_2939,N_3012);
xnor U3161 (N_3161,N_2732,N_2534);
or U3162 (N_3162,N_2503,N_3040);
nand U3163 (N_3163,N_2838,N_2887);
and U3164 (N_3164,N_2629,N_2844);
nor U3165 (N_3165,N_2567,N_2541);
nor U3166 (N_3166,N_2949,N_3042);
nor U3167 (N_3167,N_2860,N_2592);
nand U3168 (N_3168,N_2538,N_3108);
nor U3169 (N_3169,N_2624,N_2735);
nand U3170 (N_3170,N_2940,N_3100);
nand U3171 (N_3171,N_2606,N_2710);
and U3172 (N_3172,N_2655,N_2984);
and U3173 (N_3173,N_2644,N_2711);
nand U3174 (N_3174,N_2823,N_2645);
or U3175 (N_3175,N_3092,N_2632);
nand U3176 (N_3176,N_2761,N_3115);
and U3177 (N_3177,N_2666,N_3022);
nand U3178 (N_3178,N_3032,N_2669);
xnor U3179 (N_3179,N_2793,N_2837);
xnor U3180 (N_3180,N_2767,N_3082);
xnor U3181 (N_3181,N_3001,N_2973);
and U3182 (N_3182,N_3056,N_2996);
nor U3183 (N_3183,N_3101,N_2597);
nand U3184 (N_3184,N_2584,N_3007);
nand U3185 (N_3185,N_3099,N_3088);
or U3186 (N_3186,N_2679,N_2618);
nand U3187 (N_3187,N_2565,N_3050);
xor U3188 (N_3188,N_2695,N_3021);
nand U3189 (N_3189,N_2812,N_2910);
and U3190 (N_3190,N_3076,N_2818);
nand U3191 (N_3191,N_2756,N_2590);
xnor U3192 (N_3192,N_2525,N_2617);
nor U3193 (N_3193,N_3048,N_2813);
xor U3194 (N_3194,N_2968,N_3053);
nand U3195 (N_3195,N_3046,N_2506);
nand U3196 (N_3196,N_3093,N_2750);
xnor U3197 (N_3197,N_2964,N_2952);
nor U3198 (N_3198,N_2696,N_2720);
nand U3199 (N_3199,N_2899,N_3067);
or U3200 (N_3200,N_2551,N_2988);
nor U3201 (N_3201,N_2993,N_3085);
nand U3202 (N_3202,N_3004,N_2962);
nor U3203 (N_3203,N_2744,N_3054);
xnor U3204 (N_3204,N_2959,N_2911);
or U3205 (N_3205,N_2886,N_2780);
xor U3206 (N_3206,N_2647,N_2613);
nor U3207 (N_3207,N_2924,N_2890);
nand U3208 (N_3208,N_2950,N_2995);
and U3209 (N_3209,N_3024,N_2878);
nor U3210 (N_3210,N_2955,N_2743);
nor U3211 (N_3211,N_3002,N_2786);
nor U3212 (N_3212,N_3071,N_2542);
nor U3213 (N_3213,N_2562,N_2787);
nand U3214 (N_3214,N_2799,N_3117);
nor U3215 (N_3215,N_2776,N_2824);
xnor U3216 (N_3216,N_3011,N_2688);
nand U3217 (N_3217,N_2789,N_2804);
nand U3218 (N_3218,N_3029,N_3028);
nor U3219 (N_3219,N_2726,N_3044);
or U3220 (N_3220,N_3031,N_2559);
or U3221 (N_3221,N_2634,N_2925);
or U3222 (N_3222,N_2861,N_3094);
or U3223 (N_3223,N_2876,N_2648);
nand U3224 (N_3224,N_2843,N_2727);
nor U3225 (N_3225,N_2785,N_2566);
and U3226 (N_3226,N_2963,N_2848);
nor U3227 (N_3227,N_2980,N_2663);
xor U3228 (N_3228,N_2797,N_2905);
nor U3229 (N_3229,N_2524,N_2858);
nor U3230 (N_3230,N_2957,N_2664);
nand U3231 (N_3231,N_2779,N_2515);
and U3232 (N_3232,N_3009,N_2920);
nor U3233 (N_3233,N_2637,N_3049);
and U3234 (N_3234,N_2909,N_2947);
nand U3235 (N_3235,N_2897,N_2880);
and U3236 (N_3236,N_3106,N_2918);
nand U3237 (N_3237,N_2649,N_3015);
and U3238 (N_3238,N_2852,N_2903);
or U3239 (N_3239,N_2640,N_3060);
or U3240 (N_3240,N_2564,N_2738);
or U3241 (N_3241,N_3045,N_2672);
xnor U3242 (N_3242,N_2941,N_2514);
nor U3243 (N_3243,N_2554,N_2892);
nor U3244 (N_3244,N_2802,N_3095);
nand U3245 (N_3245,N_2999,N_2622);
nor U3246 (N_3246,N_3005,N_2673);
xor U3247 (N_3247,N_2604,N_2573);
and U3248 (N_3248,N_3038,N_2660);
and U3249 (N_3249,N_2557,N_2721);
nor U3250 (N_3250,N_2795,N_2850);
nor U3251 (N_3251,N_2810,N_2815);
nand U3252 (N_3252,N_2504,N_3091);
xor U3253 (N_3253,N_2619,N_2983);
nand U3254 (N_3254,N_2943,N_2770);
nor U3255 (N_3255,N_3020,N_2883);
nor U3256 (N_3256,N_2552,N_3077);
nor U3257 (N_3257,N_2841,N_3113);
and U3258 (N_3258,N_2741,N_2965);
nand U3259 (N_3259,N_2874,N_2987);
nand U3260 (N_3260,N_2616,N_3097);
or U3261 (N_3261,N_2718,N_2946);
nor U3262 (N_3262,N_3000,N_2643);
and U3263 (N_3263,N_2708,N_2893);
or U3264 (N_3264,N_2600,N_2588);
and U3265 (N_3265,N_3080,N_2788);
and U3266 (N_3266,N_2707,N_2774);
nand U3267 (N_3267,N_2539,N_2638);
and U3268 (N_3268,N_3016,N_2889);
nand U3269 (N_3269,N_2835,N_2598);
and U3270 (N_3270,N_2626,N_2826);
nor U3271 (N_3271,N_2998,N_3057);
or U3272 (N_3272,N_2675,N_2937);
xnor U3273 (N_3273,N_2650,N_3074);
xnor U3274 (N_3274,N_2931,N_2513);
nor U3275 (N_3275,N_2807,N_3030);
and U3276 (N_3276,N_2811,N_2627);
or U3277 (N_3277,N_2927,N_2805);
or U3278 (N_3278,N_2612,N_3124);
and U3279 (N_3279,N_3059,N_2682);
and U3280 (N_3280,N_2621,N_2803);
nor U3281 (N_3281,N_2678,N_2966);
or U3282 (N_3282,N_2625,N_2709);
nor U3283 (N_3283,N_2646,N_3036);
and U3284 (N_3284,N_2840,N_2583);
nor U3285 (N_3285,N_2773,N_3025);
nand U3286 (N_3286,N_3075,N_2898);
and U3287 (N_3287,N_2798,N_3096);
nor U3288 (N_3288,N_2651,N_2888);
and U3289 (N_3289,N_3003,N_3065);
and U3290 (N_3290,N_2791,N_2749);
nand U3291 (N_3291,N_2537,N_2923);
or U3292 (N_3292,N_2723,N_2734);
xor U3293 (N_3293,N_2759,N_3118);
xnor U3294 (N_3294,N_2658,N_2533);
and U3295 (N_3295,N_2752,N_2954);
nand U3296 (N_3296,N_2575,N_2623);
nand U3297 (N_3297,N_2670,N_2500);
and U3298 (N_3298,N_2641,N_2908);
nor U3299 (N_3299,N_2800,N_2991);
nor U3300 (N_3300,N_2758,N_2576);
or U3301 (N_3301,N_3058,N_2737);
or U3302 (N_3302,N_2747,N_2972);
nor U3303 (N_3303,N_2507,N_2974);
nor U3304 (N_3304,N_2689,N_3018);
and U3305 (N_3305,N_2687,N_2816);
nor U3306 (N_3306,N_2599,N_2982);
nand U3307 (N_3307,N_2822,N_2528);
xnor U3308 (N_3308,N_2677,N_2906);
xnor U3309 (N_3309,N_2607,N_2577);
xor U3310 (N_3310,N_2847,N_3078);
or U3311 (N_3311,N_2769,N_2833);
and U3312 (N_3312,N_2543,N_2976);
xor U3313 (N_3313,N_2569,N_2697);
nor U3314 (N_3314,N_2512,N_2919);
xor U3315 (N_3315,N_2871,N_2705);
and U3316 (N_3316,N_3107,N_3084);
and U3317 (N_3317,N_2685,N_3047);
nand U3318 (N_3318,N_3116,N_2635);
xor U3319 (N_3319,N_2518,N_2516);
nor U3320 (N_3320,N_2527,N_2560);
xor U3321 (N_3321,N_2684,N_2713);
nor U3322 (N_3322,N_2904,N_2867);
nand U3323 (N_3323,N_2917,N_2875);
or U3324 (N_3324,N_2778,N_2585);
or U3325 (N_3325,N_2879,N_2809);
or U3326 (N_3326,N_2872,N_2511);
nor U3327 (N_3327,N_2820,N_2631);
nor U3328 (N_3328,N_2784,N_2633);
nand U3329 (N_3329,N_2691,N_3120);
nand U3330 (N_3330,N_2970,N_2702);
nand U3331 (N_3331,N_2894,N_2839);
nor U3332 (N_3332,N_2532,N_2692);
xnor U3333 (N_3333,N_3063,N_2945);
nor U3334 (N_3334,N_2882,N_2994);
nor U3335 (N_3335,N_3034,N_2561);
nand U3336 (N_3336,N_2907,N_2763);
or U3337 (N_3337,N_2808,N_3089);
xnor U3338 (N_3338,N_2563,N_2704);
or U3339 (N_3339,N_2851,N_3072);
or U3340 (N_3340,N_2587,N_2796);
nor U3341 (N_3341,N_2580,N_2956);
nand U3342 (N_3342,N_2884,N_2895);
and U3343 (N_3343,N_2544,N_2510);
or U3344 (N_3344,N_3055,N_2849);
nor U3345 (N_3345,N_2558,N_2981);
nor U3346 (N_3346,N_2864,N_3051);
or U3347 (N_3347,N_2975,N_2519);
and U3348 (N_3348,N_3039,N_2522);
nor U3349 (N_3349,N_3069,N_2668);
nand U3350 (N_3350,N_2555,N_2620);
nand U3351 (N_3351,N_2912,N_2665);
or U3352 (N_3352,N_2928,N_3043);
or U3353 (N_3353,N_2757,N_3017);
nand U3354 (N_3354,N_2703,N_2536);
xnor U3355 (N_3355,N_2915,N_2608);
nor U3356 (N_3356,N_2700,N_2591);
and U3357 (N_3357,N_3102,N_3103);
xor U3358 (N_3358,N_2806,N_2535);
and U3359 (N_3359,N_2694,N_2900);
nand U3360 (N_3360,N_2885,N_3014);
and U3361 (N_3361,N_3112,N_2571);
or U3362 (N_3362,N_2821,N_2896);
and U3363 (N_3363,N_2681,N_2971);
or U3364 (N_3364,N_2985,N_2550);
nand U3365 (N_3365,N_2674,N_2960);
nand U3366 (N_3366,N_2701,N_2913);
and U3367 (N_3367,N_2603,N_2857);
nand U3368 (N_3368,N_3098,N_2832);
nor U3369 (N_3369,N_2502,N_3068);
nor U3370 (N_3370,N_3070,N_2717);
xnor U3371 (N_3371,N_2568,N_2921);
nand U3372 (N_3372,N_2611,N_2997);
nor U3373 (N_3373,N_2969,N_3061);
xnor U3374 (N_3374,N_3119,N_2834);
xnor U3375 (N_3375,N_2772,N_2745);
or U3376 (N_3376,N_2783,N_3104);
nor U3377 (N_3377,N_2854,N_2579);
xnor U3378 (N_3378,N_2819,N_2829);
nor U3379 (N_3379,N_2517,N_2760);
or U3380 (N_3380,N_2986,N_3110);
or U3381 (N_3381,N_2556,N_2868);
and U3382 (N_3382,N_3035,N_2728);
nand U3383 (N_3383,N_2661,N_2902);
and U3384 (N_3384,N_2827,N_2676);
nand U3385 (N_3385,N_2546,N_2693);
nand U3386 (N_3386,N_2825,N_2754);
nor U3387 (N_3387,N_2547,N_3109);
or U3388 (N_3388,N_2914,N_2766);
nor U3389 (N_3389,N_2615,N_2549);
nor U3390 (N_3390,N_2948,N_2659);
and U3391 (N_3391,N_2967,N_2724);
and U3392 (N_3392,N_2698,N_2842);
and U3393 (N_3393,N_2540,N_3087);
xnor U3394 (N_3394,N_2958,N_2657);
nand U3395 (N_3395,N_3122,N_2932);
xor U3396 (N_3396,N_2853,N_2683);
or U3397 (N_3397,N_3086,N_2831);
nor U3398 (N_3398,N_2589,N_2866);
nor U3399 (N_3399,N_2953,N_3123);
and U3400 (N_3400,N_2989,N_2929);
and U3401 (N_3401,N_3114,N_2739);
nor U3402 (N_3402,N_2652,N_2530);
or U3403 (N_3403,N_2790,N_2992);
nand U3404 (N_3404,N_3083,N_2731);
and U3405 (N_3405,N_2855,N_2740);
nand U3406 (N_3406,N_2934,N_2990);
xor U3407 (N_3407,N_2836,N_2765);
and U3408 (N_3408,N_2719,N_2922);
nand U3409 (N_3409,N_2869,N_2653);
and U3410 (N_3410,N_2628,N_3006);
xnor U3411 (N_3411,N_2764,N_2762);
and U3412 (N_3412,N_2751,N_2570);
and U3413 (N_3413,N_2870,N_2505);
nand U3414 (N_3414,N_2830,N_2586);
or U3415 (N_3415,N_2978,N_2572);
xnor U3416 (N_3416,N_3105,N_2865);
nor U3417 (N_3417,N_2690,N_2781);
nor U3418 (N_3418,N_2938,N_2610);
xnor U3419 (N_3419,N_2979,N_2593);
and U3420 (N_3420,N_2548,N_3062);
xor U3421 (N_3421,N_2730,N_2656);
nand U3422 (N_3422,N_2662,N_2545);
and U3423 (N_3423,N_2526,N_2529);
nand U3424 (N_3424,N_2828,N_2521);
nor U3425 (N_3425,N_2582,N_3027);
xnor U3426 (N_3426,N_2748,N_2706);
xnor U3427 (N_3427,N_2753,N_2729);
xor U3428 (N_3428,N_2725,N_2856);
nand U3429 (N_3429,N_3033,N_3023);
nand U3430 (N_3430,N_2930,N_2509);
nand U3431 (N_3431,N_3019,N_2594);
nand U3432 (N_3432,N_2595,N_2501);
and U3433 (N_3433,N_2794,N_2722);
nor U3434 (N_3434,N_2873,N_2636);
and U3435 (N_3435,N_3010,N_2944);
nand U3436 (N_3436,N_2531,N_2755);
xor U3437 (N_3437,N_2933,N_3065);
xnor U3438 (N_3438,N_3097,N_2998);
and U3439 (N_3439,N_2557,N_2774);
nor U3440 (N_3440,N_2912,N_3022);
nand U3441 (N_3441,N_2695,N_2932);
and U3442 (N_3442,N_2562,N_2823);
or U3443 (N_3443,N_3065,N_2815);
nor U3444 (N_3444,N_2679,N_3010);
nor U3445 (N_3445,N_2961,N_2651);
and U3446 (N_3446,N_2758,N_2560);
xnor U3447 (N_3447,N_2986,N_2743);
nor U3448 (N_3448,N_2916,N_2652);
xor U3449 (N_3449,N_2605,N_3047);
or U3450 (N_3450,N_2681,N_2626);
nor U3451 (N_3451,N_3065,N_2884);
xor U3452 (N_3452,N_2655,N_2773);
or U3453 (N_3453,N_2837,N_2670);
nand U3454 (N_3454,N_3035,N_2570);
nand U3455 (N_3455,N_2631,N_3122);
nand U3456 (N_3456,N_2582,N_2875);
xor U3457 (N_3457,N_2716,N_3117);
or U3458 (N_3458,N_2961,N_2744);
xor U3459 (N_3459,N_2938,N_2750);
or U3460 (N_3460,N_2808,N_2543);
or U3461 (N_3461,N_2939,N_3005);
nor U3462 (N_3462,N_2911,N_2830);
nor U3463 (N_3463,N_2966,N_2874);
or U3464 (N_3464,N_2539,N_2622);
and U3465 (N_3465,N_3113,N_2852);
or U3466 (N_3466,N_2993,N_2729);
or U3467 (N_3467,N_2905,N_2666);
or U3468 (N_3468,N_2525,N_2513);
and U3469 (N_3469,N_2669,N_2660);
and U3470 (N_3470,N_3038,N_2941);
xnor U3471 (N_3471,N_3100,N_2794);
or U3472 (N_3472,N_2963,N_3034);
xnor U3473 (N_3473,N_3072,N_2843);
or U3474 (N_3474,N_2925,N_3087);
nand U3475 (N_3475,N_2676,N_3026);
and U3476 (N_3476,N_2947,N_2647);
or U3477 (N_3477,N_2793,N_3051);
nand U3478 (N_3478,N_2656,N_2948);
nor U3479 (N_3479,N_2630,N_2654);
and U3480 (N_3480,N_2633,N_3009);
xor U3481 (N_3481,N_2980,N_3096);
nand U3482 (N_3482,N_2530,N_2824);
nor U3483 (N_3483,N_2502,N_2651);
or U3484 (N_3484,N_2775,N_2852);
nor U3485 (N_3485,N_2636,N_2554);
xor U3486 (N_3486,N_3029,N_2995);
or U3487 (N_3487,N_2759,N_3001);
nor U3488 (N_3488,N_2910,N_2783);
nand U3489 (N_3489,N_2958,N_2612);
xnor U3490 (N_3490,N_2573,N_2589);
or U3491 (N_3491,N_2999,N_2790);
or U3492 (N_3492,N_3086,N_2848);
xnor U3493 (N_3493,N_3043,N_2892);
or U3494 (N_3494,N_2810,N_2920);
or U3495 (N_3495,N_3040,N_2557);
and U3496 (N_3496,N_2630,N_3036);
nand U3497 (N_3497,N_2615,N_2964);
xnor U3498 (N_3498,N_2636,N_2878);
nand U3499 (N_3499,N_2721,N_2797);
xor U3500 (N_3500,N_2566,N_2688);
and U3501 (N_3501,N_2887,N_2903);
and U3502 (N_3502,N_2580,N_2700);
xor U3503 (N_3503,N_2539,N_3057);
xor U3504 (N_3504,N_3095,N_2803);
nand U3505 (N_3505,N_2631,N_2988);
and U3506 (N_3506,N_3027,N_2656);
nand U3507 (N_3507,N_2545,N_2915);
xor U3508 (N_3508,N_2820,N_2845);
xnor U3509 (N_3509,N_2940,N_2511);
nand U3510 (N_3510,N_2517,N_2604);
and U3511 (N_3511,N_2965,N_2882);
and U3512 (N_3512,N_2756,N_3074);
or U3513 (N_3513,N_3098,N_2773);
or U3514 (N_3514,N_2775,N_2876);
nor U3515 (N_3515,N_2545,N_2745);
and U3516 (N_3516,N_3118,N_3079);
xor U3517 (N_3517,N_2890,N_2759);
xor U3518 (N_3518,N_2910,N_3053);
or U3519 (N_3519,N_3008,N_2866);
nand U3520 (N_3520,N_2998,N_3029);
or U3521 (N_3521,N_2863,N_2546);
or U3522 (N_3522,N_2924,N_2563);
nor U3523 (N_3523,N_2669,N_2802);
nor U3524 (N_3524,N_2980,N_2899);
nand U3525 (N_3525,N_2933,N_2997);
nor U3526 (N_3526,N_3086,N_2742);
or U3527 (N_3527,N_2663,N_2856);
and U3528 (N_3528,N_3076,N_2902);
xor U3529 (N_3529,N_2934,N_2915);
or U3530 (N_3530,N_2698,N_2558);
xnor U3531 (N_3531,N_3122,N_3019);
or U3532 (N_3532,N_2975,N_2670);
nor U3533 (N_3533,N_3040,N_2852);
and U3534 (N_3534,N_2836,N_2946);
nor U3535 (N_3535,N_2746,N_2705);
and U3536 (N_3536,N_2754,N_2750);
and U3537 (N_3537,N_3068,N_2685);
nand U3538 (N_3538,N_2930,N_3095);
and U3539 (N_3539,N_2957,N_3070);
and U3540 (N_3540,N_2717,N_2705);
xor U3541 (N_3541,N_2584,N_2872);
nor U3542 (N_3542,N_2732,N_2676);
nand U3543 (N_3543,N_2622,N_2703);
nand U3544 (N_3544,N_3044,N_2831);
and U3545 (N_3545,N_2513,N_2657);
and U3546 (N_3546,N_2794,N_2796);
and U3547 (N_3547,N_2704,N_3046);
nand U3548 (N_3548,N_2807,N_2871);
nor U3549 (N_3549,N_2863,N_2784);
nor U3550 (N_3550,N_2877,N_2685);
nand U3551 (N_3551,N_2621,N_2810);
xor U3552 (N_3552,N_2837,N_3082);
or U3553 (N_3553,N_2772,N_3079);
and U3554 (N_3554,N_2831,N_3028);
xnor U3555 (N_3555,N_2546,N_3002);
xor U3556 (N_3556,N_2531,N_2847);
or U3557 (N_3557,N_2689,N_2576);
or U3558 (N_3558,N_3099,N_3012);
xnor U3559 (N_3559,N_3094,N_2954);
xnor U3560 (N_3560,N_2699,N_2858);
xor U3561 (N_3561,N_3117,N_3037);
xor U3562 (N_3562,N_3042,N_2708);
or U3563 (N_3563,N_2501,N_2643);
or U3564 (N_3564,N_3077,N_3117);
nor U3565 (N_3565,N_3014,N_3115);
or U3566 (N_3566,N_2607,N_2667);
or U3567 (N_3567,N_3047,N_2690);
xor U3568 (N_3568,N_2909,N_3034);
nand U3569 (N_3569,N_2914,N_3030);
and U3570 (N_3570,N_2639,N_2744);
nor U3571 (N_3571,N_2570,N_3023);
or U3572 (N_3572,N_3061,N_2944);
and U3573 (N_3573,N_3038,N_2825);
and U3574 (N_3574,N_2555,N_2744);
xnor U3575 (N_3575,N_2666,N_2766);
and U3576 (N_3576,N_2703,N_3041);
nor U3577 (N_3577,N_3014,N_3104);
and U3578 (N_3578,N_2955,N_2624);
nand U3579 (N_3579,N_2678,N_3041);
and U3580 (N_3580,N_2924,N_2538);
nor U3581 (N_3581,N_2850,N_2984);
or U3582 (N_3582,N_3068,N_3042);
nand U3583 (N_3583,N_2931,N_2821);
or U3584 (N_3584,N_2882,N_2748);
nand U3585 (N_3585,N_3040,N_3059);
nand U3586 (N_3586,N_2785,N_2904);
and U3587 (N_3587,N_3010,N_2583);
nand U3588 (N_3588,N_2597,N_2808);
xnor U3589 (N_3589,N_2589,N_3049);
nor U3590 (N_3590,N_3028,N_2686);
and U3591 (N_3591,N_3045,N_2574);
or U3592 (N_3592,N_3002,N_3028);
nor U3593 (N_3593,N_2875,N_2821);
xor U3594 (N_3594,N_2795,N_3001);
xnor U3595 (N_3595,N_2723,N_2977);
and U3596 (N_3596,N_2782,N_2830);
nand U3597 (N_3597,N_2991,N_2688);
or U3598 (N_3598,N_2931,N_3076);
nor U3599 (N_3599,N_2515,N_2865);
and U3600 (N_3600,N_2956,N_2679);
xnor U3601 (N_3601,N_2651,N_2686);
nor U3602 (N_3602,N_2634,N_2659);
nand U3603 (N_3603,N_2830,N_2992);
and U3604 (N_3604,N_2580,N_2780);
and U3605 (N_3605,N_2589,N_2511);
or U3606 (N_3606,N_2725,N_3074);
nor U3607 (N_3607,N_2999,N_2913);
or U3608 (N_3608,N_2527,N_2528);
xor U3609 (N_3609,N_2776,N_2952);
xor U3610 (N_3610,N_2835,N_2937);
or U3611 (N_3611,N_3101,N_2785);
and U3612 (N_3612,N_2638,N_2688);
nand U3613 (N_3613,N_3121,N_3066);
nand U3614 (N_3614,N_3093,N_2663);
and U3615 (N_3615,N_2730,N_3043);
and U3616 (N_3616,N_2986,N_2990);
nor U3617 (N_3617,N_2703,N_3049);
or U3618 (N_3618,N_2592,N_2750);
and U3619 (N_3619,N_2740,N_2991);
xnor U3620 (N_3620,N_2827,N_2559);
or U3621 (N_3621,N_2536,N_3062);
or U3622 (N_3622,N_2754,N_2510);
nor U3623 (N_3623,N_2632,N_2737);
nor U3624 (N_3624,N_2586,N_3009);
xor U3625 (N_3625,N_2977,N_2676);
and U3626 (N_3626,N_2976,N_2973);
and U3627 (N_3627,N_2742,N_2647);
and U3628 (N_3628,N_2629,N_2679);
or U3629 (N_3629,N_2650,N_2802);
and U3630 (N_3630,N_2677,N_3034);
or U3631 (N_3631,N_2854,N_2765);
xor U3632 (N_3632,N_2897,N_2586);
nand U3633 (N_3633,N_2769,N_2819);
xnor U3634 (N_3634,N_2670,N_2696);
nor U3635 (N_3635,N_2851,N_2698);
xor U3636 (N_3636,N_2905,N_2549);
or U3637 (N_3637,N_2602,N_2832);
nor U3638 (N_3638,N_3086,N_2717);
xnor U3639 (N_3639,N_2588,N_2555);
or U3640 (N_3640,N_3096,N_2711);
nand U3641 (N_3641,N_2891,N_3119);
or U3642 (N_3642,N_2540,N_3107);
nand U3643 (N_3643,N_2603,N_2955);
and U3644 (N_3644,N_2709,N_2802);
or U3645 (N_3645,N_2557,N_3026);
and U3646 (N_3646,N_2582,N_2836);
or U3647 (N_3647,N_3039,N_2890);
or U3648 (N_3648,N_3066,N_2769);
or U3649 (N_3649,N_2926,N_3016);
or U3650 (N_3650,N_2932,N_3021);
and U3651 (N_3651,N_2691,N_3017);
nand U3652 (N_3652,N_2818,N_2677);
and U3653 (N_3653,N_2526,N_2813);
nor U3654 (N_3654,N_2717,N_2788);
nor U3655 (N_3655,N_2863,N_3009);
nor U3656 (N_3656,N_2692,N_2744);
xor U3657 (N_3657,N_2517,N_2740);
or U3658 (N_3658,N_2858,N_2964);
nand U3659 (N_3659,N_2770,N_2624);
xor U3660 (N_3660,N_3018,N_3080);
and U3661 (N_3661,N_2593,N_2653);
nand U3662 (N_3662,N_3022,N_2819);
nand U3663 (N_3663,N_3049,N_2705);
nor U3664 (N_3664,N_3121,N_2793);
xnor U3665 (N_3665,N_2807,N_2760);
or U3666 (N_3666,N_3071,N_3123);
or U3667 (N_3667,N_2876,N_2510);
nand U3668 (N_3668,N_2733,N_2604);
nor U3669 (N_3669,N_2736,N_2609);
or U3670 (N_3670,N_2556,N_2871);
xor U3671 (N_3671,N_2986,N_2559);
or U3672 (N_3672,N_2823,N_2686);
and U3673 (N_3673,N_2563,N_3070);
xor U3674 (N_3674,N_2769,N_2881);
xnor U3675 (N_3675,N_2838,N_2991);
or U3676 (N_3676,N_3121,N_3067);
nand U3677 (N_3677,N_2638,N_2640);
nand U3678 (N_3678,N_2540,N_2606);
nand U3679 (N_3679,N_2527,N_2620);
xor U3680 (N_3680,N_2735,N_2669);
xor U3681 (N_3681,N_2507,N_2613);
xor U3682 (N_3682,N_2645,N_2842);
and U3683 (N_3683,N_2670,N_2982);
xor U3684 (N_3684,N_2921,N_2581);
or U3685 (N_3685,N_2822,N_2525);
nand U3686 (N_3686,N_2892,N_2678);
or U3687 (N_3687,N_2735,N_2671);
nand U3688 (N_3688,N_2606,N_2559);
nor U3689 (N_3689,N_3030,N_2924);
xnor U3690 (N_3690,N_2938,N_2524);
or U3691 (N_3691,N_2724,N_2558);
nor U3692 (N_3692,N_2979,N_2840);
nand U3693 (N_3693,N_2731,N_2889);
and U3694 (N_3694,N_2712,N_2945);
nand U3695 (N_3695,N_2611,N_2715);
and U3696 (N_3696,N_2971,N_3119);
xnor U3697 (N_3697,N_2554,N_3111);
nand U3698 (N_3698,N_2516,N_2878);
and U3699 (N_3699,N_2612,N_2756);
nor U3700 (N_3700,N_2677,N_2860);
or U3701 (N_3701,N_2662,N_2847);
xnor U3702 (N_3702,N_2722,N_3080);
nand U3703 (N_3703,N_2733,N_2835);
nor U3704 (N_3704,N_2768,N_2817);
nor U3705 (N_3705,N_2864,N_2836);
and U3706 (N_3706,N_2761,N_2962);
nor U3707 (N_3707,N_2840,N_2723);
xnor U3708 (N_3708,N_2732,N_2992);
xor U3709 (N_3709,N_2596,N_3065);
and U3710 (N_3710,N_2616,N_2505);
or U3711 (N_3711,N_2893,N_2771);
xor U3712 (N_3712,N_2509,N_2770);
and U3713 (N_3713,N_2883,N_2529);
nand U3714 (N_3714,N_2788,N_2903);
and U3715 (N_3715,N_2682,N_2927);
and U3716 (N_3716,N_2619,N_2956);
xor U3717 (N_3717,N_3122,N_2925);
xor U3718 (N_3718,N_2573,N_2525);
xnor U3719 (N_3719,N_2730,N_2761);
nand U3720 (N_3720,N_3084,N_2960);
and U3721 (N_3721,N_2914,N_2693);
and U3722 (N_3722,N_2975,N_2952);
or U3723 (N_3723,N_2803,N_2851);
nand U3724 (N_3724,N_2942,N_3102);
xor U3725 (N_3725,N_2518,N_2870);
xnor U3726 (N_3726,N_3011,N_3019);
nor U3727 (N_3727,N_2710,N_2510);
nand U3728 (N_3728,N_2632,N_2647);
nand U3729 (N_3729,N_2572,N_2812);
nand U3730 (N_3730,N_2915,N_2798);
nor U3731 (N_3731,N_2725,N_2807);
nand U3732 (N_3732,N_3095,N_3092);
or U3733 (N_3733,N_2859,N_3101);
and U3734 (N_3734,N_2940,N_2734);
or U3735 (N_3735,N_2563,N_2761);
or U3736 (N_3736,N_2541,N_2889);
nand U3737 (N_3737,N_2770,N_3057);
nand U3738 (N_3738,N_2641,N_2828);
xnor U3739 (N_3739,N_2901,N_2852);
nor U3740 (N_3740,N_2738,N_2705);
nor U3741 (N_3741,N_2775,N_3000);
and U3742 (N_3742,N_2999,N_3035);
nand U3743 (N_3743,N_2750,N_2812);
xnor U3744 (N_3744,N_2922,N_2720);
or U3745 (N_3745,N_2699,N_3124);
and U3746 (N_3746,N_3056,N_2734);
nand U3747 (N_3747,N_3026,N_2867);
nand U3748 (N_3748,N_2911,N_2760);
xnor U3749 (N_3749,N_2852,N_2659);
nand U3750 (N_3750,N_3466,N_3738);
or U3751 (N_3751,N_3746,N_3335);
or U3752 (N_3752,N_3640,N_3730);
xnor U3753 (N_3753,N_3623,N_3423);
xor U3754 (N_3754,N_3439,N_3127);
and U3755 (N_3755,N_3362,N_3317);
nand U3756 (N_3756,N_3564,N_3229);
and U3757 (N_3757,N_3269,N_3566);
and U3758 (N_3758,N_3342,N_3310);
or U3759 (N_3759,N_3479,N_3489);
and U3760 (N_3760,N_3484,N_3225);
and U3761 (N_3761,N_3363,N_3185);
or U3762 (N_3762,N_3646,N_3560);
and U3763 (N_3763,N_3700,N_3556);
xor U3764 (N_3764,N_3542,N_3731);
xnor U3765 (N_3765,N_3638,N_3268);
xnor U3766 (N_3766,N_3681,N_3178);
or U3767 (N_3767,N_3683,N_3382);
xor U3768 (N_3768,N_3380,N_3415);
or U3769 (N_3769,N_3475,N_3161);
xor U3770 (N_3770,N_3308,N_3534);
or U3771 (N_3771,N_3678,N_3387);
xor U3772 (N_3772,N_3287,N_3451);
or U3773 (N_3773,N_3265,N_3421);
nor U3774 (N_3774,N_3435,N_3684);
xor U3775 (N_3775,N_3369,N_3692);
nand U3776 (N_3776,N_3548,N_3272);
nor U3777 (N_3777,N_3199,N_3192);
or U3778 (N_3778,N_3256,N_3729);
or U3779 (N_3779,N_3339,N_3652);
nand U3780 (N_3780,N_3430,N_3142);
nor U3781 (N_3781,N_3516,N_3708);
nor U3782 (N_3782,N_3695,N_3513);
or U3783 (N_3783,N_3530,N_3266);
nor U3784 (N_3784,N_3605,N_3591);
xnor U3785 (N_3785,N_3667,N_3609);
or U3786 (N_3786,N_3747,N_3514);
and U3787 (N_3787,N_3223,N_3410);
nand U3788 (N_3788,N_3467,N_3303);
nand U3789 (N_3789,N_3414,N_3138);
and U3790 (N_3790,N_3541,N_3179);
or U3791 (N_3791,N_3334,N_3570);
and U3792 (N_3792,N_3180,N_3291);
and U3793 (N_3793,N_3422,N_3386);
and U3794 (N_3794,N_3726,N_3299);
or U3795 (N_3795,N_3601,N_3505);
xor U3796 (N_3796,N_3704,N_3455);
xor U3797 (N_3797,N_3206,N_3690);
and U3798 (N_3798,N_3599,N_3733);
or U3799 (N_3799,N_3366,N_3580);
nand U3800 (N_3800,N_3420,N_3491);
xor U3801 (N_3801,N_3281,N_3452);
nor U3802 (N_3802,N_3359,N_3527);
xnor U3803 (N_3803,N_3216,N_3249);
nand U3804 (N_3804,N_3594,N_3186);
xor U3805 (N_3805,N_3578,N_3252);
or U3806 (N_3806,N_3551,N_3177);
xor U3807 (N_3807,N_3523,N_3368);
and U3808 (N_3808,N_3728,N_3176);
or U3809 (N_3809,N_3436,N_3137);
or U3810 (N_3810,N_3665,N_3231);
or U3811 (N_3811,N_3468,N_3337);
nor U3812 (N_3812,N_3535,N_3627);
nand U3813 (N_3813,N_3321,N_3714);
and U3814 (N_3814,N_3583,N_3183);
and U3815 (N_3815,N_3156,N_3151);
xor U3816 (N_3816,N_3628,N_3538);
and U3817 (N_3817,N_3712,N_3220);
nand U3818 (N_3818,N_3477,N_3128);
xnor U3819 (N_3819,N_3447,N_3540);
nor U3820 (N_3820,N_3260,N_3394);
nor U3821 (N_3821,N_3145,N_3649);
or U3822 (N_3822,N_3597,N_3413);
or U3823 (N_3823,N_3552,N_3641);
nand U3824 (N_3824,N_3383,N_3515);
and U3825 (N_3825,N_3693,N_3585);
nor U3826 (N_3826,N_3230,N_3647);
and U3827 (N_3827,N_3642,N_3353);
and U3828 (N_3828,N_3531,N_3444);
xnor U3829 (N_3829,N_3718,N_3679);
nor U3830 (N_3830,N_3318,N_3717);
xnor U3831 (N_3831,N_3471,N_3191);
nand U3832 (N_3832,N_3289,N_3358);
nor U3833 (N_3833,N_3481,N_3407);
nor U3834 (N_3834,N_3493,N_3418);
and U3835 (N_3835,N_3309,N_3711);
xnor U3836 (N_3836,N_3685,N_3559);
nand U3837 (N_3837,N_3456,N_3241);
xnor U3838 (N_3838,N_3221,N_3297);
or U3839 (N_3839,N_3307,N_3565);
or U3840 (N_3840,N_3153,N_3217);
nand U3841 (N_3841,N_3461,N_3533);
nand U3842 (N_3842,N_3416,N_3190);
xnor U3843 (N_3843,N_3319,N_3469);
xnor U3844 (N_3844,N_3248,N_3125);
and U3845 (N_3845,N_3553,N_3616);
or U3846 (N_3846,N_3748,N_3227);
and U3847 (N_3847,N_3460,N_3412);
nor U3848 (N_3848,N_3454,N_3348);
or U3849 (N_3849,N_3499,N_3724);
xor U3850 (N_3850,N_3236,N_3244);
nand U3851 (N_3851,N_3170,N_3441);
or U3852 (N_3852,N_3429,N_3402);
nor U3853 (N_3853,N_3376,N_3129);
and U3854 (N_3854,N_3618,N_3650);
or U3855 (N_3855,N_3694,N_3581);
nand U3856 (N_3856,N_3582,N_3670);
nor U3857 (N_3857,N_3340,N_3482);
nor U3858 (N_3858,N_3546,N_3437);
nand U3859 (N_3859,N_3575,N_3240);
nand U3860 (N_3860,N_3209,N_3476);
nor U3861 (N_3861,N_3238,N_3443);
and U3862 (N_3862,N_3164,N_3433);
and U3863 (N_3863,N_3235,N_3653);
or U3864 (N_3864,N_3740,N_3390);
nor U3865 (N_3865,N_3403,N_3341);
nor U3866 (N_3866,N_3497,N_3356);
or U3867 (N_3867,N_3350,N_3345);
or U3868 (N_3868,N_3725,N_3417);
nor U3869 (N_3869,N_3522,N_3160);
or U3870 (N_3870,N_3676,N_3432);
nor U3871 (N_3871,N_3263,N_3374);
and U3872 (N_3872,N_3181,N_3346);
or U3873 (N_3873,N_3709,N_3696);
nand U3874 (N_3874,N_3517,N_3504);
nand U3875 (N_3875,N_3325,N_3526);
and U3876 (N_3876,N_3478,N_3408);
and U3877 (N_3877,N_3198,N_3354);
nand U3878 (N_3878,N_3329,N_3463);
xor U3879 (N_3879,N_3537,N_3296);
nand U3880 (N_3880,N_3657,N_3702);
xnor U3881 (N_3881,N_3590,N_3384);
or U3882 (N_3882,N_3361,N_3487);
xnor U3883 (N_3883,N_3637,N_3301);
or U3884 (N_3884,N_3302,N_3473);
and U3885 (N_3885,N_3434,N_3648);
xor U3886 (N_3886,N_3598,N_3674);
nor U3887 (N_3887,N_3154,N_3490);
nand U3888 (N_3888,N_3257,N_3411);
or U3889 (N_3889,N_3425,N_3157);
xor U3890 (N_3890,N_3624,N_3389);
or U3891 (N_3891,N_3131,N_3519);
xnor U3892 (N_3892,N_3520,N_3464);
xor U3893 (N_3893,N_3328,N_3502);
nand U3894 (N_3894,N_3659,N_3713);
xnor U3895 (N_3895,N_3501,N_3237);
nor U3896 (N_3896,N_3682,N_3529);
xnor U3897 (N_3897,N_3656,N_3633);
nor U3898 (N_3898,N_3214,N_3330);
nor U3899 (N_3899,N_3351,N_3458);
nand U3900 (N_3900,N_3453,N_3506);
and U3901 (N_3901,N_3737,N_3370);
nand U3902 (N_3902,N_3210,N_3169);
or U3903 (N_3903,N_3654,N_3593);
xnor U3904 (N_3904,N_3586,N_3596);
nor U3905 (N_3905,N_3595,N_3568);
nor U3906 (N_3906,N_3399,N_3222);
nand U3907 (N_3907,N_3528,N_3132);
or U3908 (N_3908,N_3349,N_3270);
or U3909 (N_3909,N_3562,N_3572);
nor U3910 (N_3910,N_3701,N_3735);
or U3911 (N_3911,N_3732,N_3508);
nand U3912 (N_3912,N_3187,N_3669);
xor U3913 (N_3913,N_3472,N_3344);
or U3914 (N_3914,N_3364,N_3294);
nand U3915 (N_3915,N_3691,N_3126);
nor U3916 (N_3916,N_3152,N_3459);
or U3917 (N_3917,N_3201,N_3391);
or U3918 (N_3918,N_3234,N_3193);
and U3919 (N_3919,N_3720,N_3293);
and U3920 (N_3920,N_3574,N_3215);
xor U3921 (N_3921,N_3280,N_3278);
nor U3922 (N_3922,N_3621,N_3147);
and U3923 (N_3923,N_3474,N_3555);
and U3924 (N_3924,N_3203,N_3604);
nor U3925 (N_3925,N_3189,N_3273);
or U3926 (N_3926,N_3277,N_3242);
or U3927 (N_3927,N_3224,N_3144);
nor U3928 (N_3928,N_3705,N_3134);
nand U3929 (N_3929,N_3488,N_3322);
or U3930 (N_3930,N_3372,N_3419);
or U3931 (N_3931,N_3155,N_3606);
or U3932 (N_3932,N_3158,N_3603);
nand U3933 (N_3933,N_3584,N_3228);
or U3934 (N_3934,N_3393,N_3442);
nor U3935 (N_3935,N_3173,N_3557);
and U3936 (N_3936,N_3140,N_3205);
nor U3937 (N_3937,N_3392,N_3483);
and U3938 (N_3938,N_3449,N_3744);
and U3939 (N_3939,N_3500,N_3743);
nand U3940 (N_3940,N_3741,N_3554);
nand U3941 (N_3941,N_3233,N_3511);
nand U3942 (N_3942,N_3405,N_3680);
or U3943 (N_3943,N_3465,N_3749);
xor U3944 (N_3944,N_3381,N_3660);
and U3945 (N_3945,N_3261,N_3645);
nand U3946 (N_3946,N_3635,N_3607);
xnor U3947 (N_3947,N_3611,N_3589);
nor U3948 (N_3948,N_3327,N_3347);
and U3949 (N_3949,N_3194,N_3247);
xnor U3950 (N_3950,N_3632,N_3576);
nor U3951 (N_3951,N_3719,N_3258);
xnor U3952 (N_3952,N_3355,N_3614);
nand U3953 (N_3953,N_3510,N_3672);
xor U3954 (N_3954,N_3426,N_3323);
nor U3955 (N_3955,N_3612,N_3406);
nand U3956 (N_3956,N_3274,N_3245);
xnor U3957 (N_3957,N_3569,N_3636);
xor U3958 (N_3958,N_3166,N_3699);
or U3959 (N_3959,N_3630,N_3561);
nor U3960 (N_3960,N_3480,N_3503);
xor U3961 (N_3961,N_3388,N_3305);
nand U3962 (N_3962,N_3404,N_3644);
nor U3963 (N_3963,N_3365,N_3375);
nor U3964 (N_3964,N_3279,N_3525);
nor U3965 (N_3965,N_3314,N_3723);
or U3966 (N_3966,N_3254,N_3655);
xor U3967 (N_3967,N_3663,N_3697);
xnor U3968 (N_3968,N_3378,N_3698);
xor U3969 (N_3969,N_3651,N_3243);
nand U3970 (N_3970,N_3333,N_3250);
nor U3971 (N_3971,N_3620,N_3136);
or U3972 (N_3972,N_3662,N_3558);
nand U3973 (N_3973,N_3664,N_3445);
or U3974 (N_3974,N_3440,N_3218);
xor U3975 (N_3975,N_3495,N_3130);
and U3976 (N_3976,N_3271,N_3331);
nor U3977 (N_3977,N_3188,N_3195);
nand U3978 (N_3978,N_3457,N_3686);
nor U3979 (N_3979,N_3300,N_3689);
or U3980 (N_3980,N_3431,N_3608);
and U3981 (N_3981,N_3715,N_3587);
or U3982 (N_3982,N_3615,N_3485);
and U3983 (N_3983,N_3518,N_3316);
nor U3984 (N_3984,N_3172,N_3211);
xnor U3985 (N_3985,N_3239,N_3543);
or U3986 (N_3986,N_3545,N_3196);
nor U3987 (N_3987,N_3496,N_3338);
nor U3988 (N_3988,N_3610,N_3171);
nand U3989 (N_3989,N_3286,N_3143);
xor U3990 (N_3990,N_3688,N_3311);
nand U3991 (N_3991,N_3470,N_3722);
nand U3992 (N_3992,N_3671,N_3424);
xnor U3993 (N_3993,N_3745,N_3326);
and U3994 (N_3994,N_3204,N_3285);
nor U3995 (N_3995,N_3275,N_3661);
xnor U3996 (N_3996,N_3133,N_3446);
xor U3997 (N_3997,N_3313,N_3532);
xnor U3998 (N_3998,N_3288,N_3282);
and U3999 (N_3999,N_3295,N_3577);
nor U4000 (N_4000,N_3159,N_3600);
or U4001 (N_4001,N_3219,N_3739);
or U4002 (N_4002,N_3324,N_3197);
nand U4003 (N_4003,N_3687,N_3284);
and U4004 (N_4004,N_3675,N_3563);
nand U4005 (N_4005,N_3148,N_3397);
nor U4006 (N_4006,N_3677,N_3658);
nand U4007 (N_4007,N_3734,N_3264);
or U4008 (N_4008,N_3592,N_3312);
nor U4009 (N_4009,N_3213,N_3544);
nor U4010 (N_4010,N_3706,N_3336);
and U4011 (N_4011,N_3276,N_3507);
xnor U4012 (N_4012,N_3617,N_3146);
nor U4013 (N_4013,N_3385,N_3255);
nor U4014 (N_4014,N_3267,N_3571);
nor U4015 (N_4015,N_3721,N_3486);
nand U4016 (N_4016,N_3668,N_3549);
nand U4017 (N_4017,N_3304,N_3212);
nand U4018 (N_4018,N_3742,N_3707);
xnor U4019 (N_4019,N_3139,N_3165);
xor U4020 (N_4020,N_3547,N_3184);
or U4021 (N_4021,N_3631,N_3207);
or U4022 (N_4022,N_3494,N_3232);
nand U4023 (N_4023,N_3251,N_3629);
nand U4024 (N_4024,N_3371,N_3539);
nand U4025 (N_4025,N_3373,N_3283);
and U4026 (N_4026,N_3710,N_3567);
and U4027 (N_4027,N_3167,N_3666);
and U4028 (N_4028,N_3262,N_3200);
nand U4029 (N_4029,N_3332,N_3428);
xnor U4030 (N_4030,N_3360,N_3352);
and U4031 (N_4031,N_3448,N_3579);
xor U4032 (N_4032,N_3524,N_3320);
and U4033 (N_4033,N_3673,N_3492);
nand U4034 (N_4034,N_3409,N_3202);
xor U4035 (N_4035,N_3550,N_3259);
xor U4036 (N_4036,N_3639,N_3377);
nand U4037 (N_4037,N_3149,N_3298);
and U4038 (N_4038,N_3401,N_3306);
or U4039 (N_4039,N_3253,N_3246);
or U4040 (N_4040,N_3162,N_3626);
nor U4041 (N_4041,N_3703,N_3357);
or U4042 (N_4042,N_3498,N_3588);
and U4043 (N_4043,N_3175,N_3622);
and U4044 (N_4044,N_3625,N_3602);
xor U4045 (N_4045,N_3716,N_3141);
or U4046 (N_4046,N_3135,N_3509);
or U4047 (N_4047,N_3226,N_3438);
nand U4048 (N_4048,N_3292,N_3643);
or U4049 (N_4049,N_3395,N_3573);
nor U4050 (N_4050,N_3343,N_3613);
xor U4051 (N_4051,N_3462,N_3367);
xor U4052 (N_4052,N_3174,N_3536);
xor U4053 (N_4053,N_3521,N_3379);
and U4054 (N_4054,N_3396,N_3727);
nor U4055 (N_4055,N_3619,N_3427);
nor U4056 (N_4056,N_3450,N_3400);
or U4057 (N_4057,N_3208,N_3634);
and U4058 (N_4058,N_3512,N_3736);
nor U4059 (N_4059,N_3163,N_3398);
or U4060 (N_4060,N_3150,N_3315);
and U4061 (N_4061,N_3290,N_3168);
and U4062 (N_4062,N_3182,N_3130);
and U4063 (N_4063,N_3645,N_3205);
nor U4064 (N_4064,N_3234,N_3307);
or U4065 (N_4065,N_3596,N_3315);
and U4066 (N_4066,N_3294,N_3212);
or U4067 (N_4067,N_3564,N_3194);
nor U4068 (N_4068,N_3267,N_3590);
nand U4069 (N_4069,N_3569,N_3606);
or U4070 (N_4070,N_3550,N_3682);
nand U4071 (N_4071,N_3569,N_3129);
nor U4072 (N_4072,N_3675,N_3548);
nor U4073 (N_4073,N_3711,N_3244);
and U4074 (N_4074,N_3573,N_3702);
or U4075 (N_4075,N_3604,N_3581);
or U4076 (N_4076,N_3132,N_3488);
nand U4077 (N_4077,N_3383,N_3459);
nand U4078 (N_4078,N_3289,N_3230);
or U4079 (N_4079,N_3481,N_3203);
nor U4080 (N_4080,N_3684,N_3525);
nor U4081 (N_4081,N_3492,N_3713);
nor U4082 (N_4082,N_3742,N_3593);
xor U4083 (N_4083,N_3218,N_3717);
nand U4084 (N_4084,N_3599,N_3655);
nand U4085 (N_4085,N_3279,N_3493);
nor U4086 (N_4086,N_3282,N_3419);
and U4087 (N_4087,N_3297,N_3285);
nand U4088 (N_4088,N_3453,N_3508);
nor U4089 (N_4089,N_3675,N_3326);
or U4090 (N_4090,N_3224,N_3521);
nor U4091 (N_4091,N_3458,N_3159);
nor U4092 (N_4092,N_3147,N_3262);
nor U4093 (N_4093,N_3642,N_3339);
and U4094 (N_4094,N_3267,N_3238);
nor U4095 (N_4095,N_3599,N_3610);
or U4096 (N_4096,N_3445,N_3748);
nor U4097 (N_4097,N_3466,N_3355);
xor U4098 (N_4098,N_3385,N_3260);
nor U4099 (N_4099,N_3430,N_3584);
nand U4100 (N_4100,N_3334,N_3158);
and U4101 (N_4101,N_3201,N_3681);
nor U4102 (N_4102,N_3534,N_3655);
and U4103 (N_4103,N_3468,N_3471);
or U4104 (N_4104,N_3315,N_3284);
nor U4105 (N_4105,N_3327,N_3593);
and U4106 (N_4106,N_3683,N_3519);
and U4107 (N_4107,N_3468,N_3408);
nor U4108 (N_4108,N_3232,N_3648);
nor U4109 (N_4109,N_3724,N_3424);
xnor U4110 (N_4110,N_3622,N_3623);
nand U4111 (N_4111,N_3162,N_3376);
nor U4112 (N_4112,N_3328,N_3699);
and U4113 (N_4113,N_3337,N_3166);
xnor U4114 (N_4114,N_3254,N_3202);
xor U4115 (N_4115,N_3244,N_3556);
nor U4116 (N_4116,N_3545,N_3633);
or U4117 (N_4117,N_3198,N_3262);
or U4118 (N_4118,N_3232,N_3362);
nand U4119 (N_4119,N_3547,N_3317);
nor U4120 (N_4120,N_3390,N_3270);
or U4121 (N_4121,N_3382,N_3455);
nor U4122 (N_4122,N_3267,N_3331);
xnor U4123 (N_4123,N_3722,N_3581);
xor U4124 (N_4124,N_3241,N_3228);
nor U4125 (N_4125,N_3689,N_3291);
xnor U4126 (N_4126,N_3497,N_3746);
nand U4127 (N_4127,N_3436,N_3723);
or U4128 (N_4128,N_3233,N_3714);
and U4129 (N_4129,N_3719,N_3674);
nand U4130 (N_4130,N_3511,N_3307);
nor U4131 (N_4131,N_3610,N_3133);
and U4132 (N_4132,N_3625,N_3512);
and U4133 (N_4133,N_3667,N_3705);
or U4134 (N_4134,N_3304,N_3454);
and U4135 (N_4135,N_3196,N_3414);
and U4136 (N_4136,N_3463,N_3747);
and U4137 (N_4137,N_3599,N_3145);
nand U4138 (N_4138,N_3606,N_3680);
xor U4139 (N_4139,N_3157,N_3572);
nor U4140 (N_4140,N_3395,N_3495);
and U4141 (N_4141,N_3659,N_3359);
xnor U4142 (N_4142,N_3158,N_3377);
nand U4143 (N_4143,N_3159,N_3269);
nand U4144 (N_4144,N_3707,N_3642);
and U4145 (N_4145,N_3264,N_3705);
and U4146 (N_4146,N_3713,N_3516);
xnor U4147 (N_4147,N_3581,N_3224);
xor U4148 (N_4148,N_3261,N_3240);
or U4149 (N_4149,N_3537,N_3631);
nor U4150 (N_4150,N_3383,N_3674);
xnor U4151 (N_4151,N_3528,N_3468);
and U4152 (N_4152,N_3592,N_3390);
nor U4153 (N_4153,N_3457,N_3478);
and U4154 (N_4154,N_3683,N_3686);
nand U4155 (N_4155,N_3436,N_3231);
xnor U4156 (N_4156,N_3446,N_3730);
and U4157 (N_4157,N_3461,N_3321);
and U4158 (N_4158,N_3722,N_3413);
or U4159 (N_4159,N_3239,N_3559);
or U4160 (N_4160,N_3224,N_3353);
and U4161 (N_4161,N_3189,N_3504);
xnor U4162 (N_4162,N_3604,N_3531);
nor U4163 (N_4163,N_3408,N_3608);
nor U4164 (N_4164,N_3369,N_3419);
nand U4165 (N_4165,N_3281,N_3674);
xor U4166 (N_4166,N_3337,N_3377);
or U4167 (N_4167,N_3644,N_3465);
nor U4168 (N_4168,N_3395,N_3674);
or U4169 (N_4169,N_3529,N_3695);
and U4170 (N_4170,N_3522,N_3279);
xor U4171 (N_4171,N_3608,N_3602);
and U4172 (N_4172,N_3488,N_3196);
nand U4173 (N_4173,N_3341,N_3412);
nor U4174 (N_4174,N_3691,N_3589);
nor U4175 (N_4175,N_3355,N_3233);
or U4176 (N_4176,N_3660,N_3711);
and U4177 (N_4177,N_3371,N_3522);
nor U4178 (N_4178,N_3562,N_3244);
and U4179 (N_4179,N_3240,N_3503);
nand U4180 (N_4180,N_3423,N_3413);
nand U4181 (N_4181,N_3563,N_3539);
nand U4182 (N_4182,N_3310,N_3285);
xnor U4183 (N_4183,N_3159,N_3387);
and U4184 (N_4184,N_3475,N_3714);
xor U4185 (N_4185,N_3315,N_3318);
and U4186 (N_4186,N_3626,N_3731);
xnor U4187 (N_4187,N_3262,N_3562);
and U4188 (N_4188,N_3736,N_3738);
xor U4189 (N_4189,N_3548,N_3274);
nor U4190 (N_4190,N_3190,N_3216);
nor U4191 (N_4191,N_3391,N_3411);
and U4192 (N_4192,N_3178,N_3242);
or U4193 (N_4193,N_3699,N_3665);
or U4194 (N_4194,N_3415,N_3318);
nand U4195 (N_4195,N_3140,N_3529);
or U4196 (N_4196,N_3660,N_3252);
nor U4197 (N_4197,N_3218,N_3427);
xnor U4198 (N_4198,N_3243,N_3324);
nor U4199 (N_4199,N_3611,N_3255);
xnor U4200 (N_4200,N_3684,N_3605);
and U4201 (N_4201,N_3150,N_3397);
and U4202 (N_4202,N_3640,N_3738);
xnor U4203 (N_4203,N_3482,N_3317);
nor U4204 (N_4204,N_3622,N_3522);
nand U4205 (N_4205,N_3675,N_3496);
and U4206 (N_4206,N_3175,N_3460);
nor U4207 (N_4207,N_3317,N_3158);
xor U4208 (N_4208,N_3377,N_3524);
or U4209 (N_4209,N_3393,N_3294);
nor U4210 (N_4210,N_3506,N_3202);
xnor U4211 (N_4211,N_3514,N_3681);
nand U4212 (N_4212,N_3299,N_3185);
nor U4213 (N_4213,N_3270,N_3161);
nor U4214 (N_4214,N_3177,N_3431);
or U4215 (N_4215,N_3148,N_3439);
nand U4216 (N_4216,N_3312,N_3722);
nand U4217 (N_4217,N_3285,N_3663);
xnor U4218 (N_4218,N_3545,N_3254);
or U4219 (N_4219,N_3592,N_3586);
nor U4220 (N_4220,N_3438,N_3544);
nor U4221 (N_4221,N_3463,N_3362);
nor U4222 (N_4222,N_3349,N_3512);
nor U4223 (N_4223,N_3214,N_3461);
nor U4224 (N_4224,N_3518,N_3222);
xor U4225 (N_4225,N_3621,N_3157);
and U4226 (N_4226,N_3323,N_3140);
nor U4227 (N_4227,N_3364,N_3637);
xor U4228 (N_4228,N_3157,N_3564);
or U4229 (N_4229,N_3314,N_3304);
xor U4230 (N_4230,N_3266,N_3672);
nor U4231 (N_4231,N_3201,N_3283);
nor U4232 (N_4232,N_3428,N_3183);
nor U4233 (N_4233,N_3493,N_3171);
nor U4234 (N_4234,N_3688,N_3690);
nor U4235 (N_4235,N_3251,N_3712);
xnor U4236 (N_4236,N_3368,N_3130);
and U4237 (N_4237,N_3589,N_3453);
nand U4238 (N_4238,N_3223,N_3154);
nand U4239 (N_4239,N_3172,N_3140);
or U4240 (N_4240,N_3499,N_3393);
nand U4241 (N_4241,N_3477,N_3209);
nand U4242 (N_4242,N_3178,N_3510);
xnor U4243 (N_4243,N_3592,N_3467);
nor U4244 (N_4244,N_3492,N_3365);
and U4245 (N_4245,N_3472,N_3229);
nand U4246 (N_4246,N_3367,N_3401);
xor U4247 (N_4247,N_3354,N_3154);
or U4248 (N_4248,N_3600,N_3403);
xnor U4249 (N_4249,N_3658,N_3376);
nor U4250 (N_4250,N_3184,N_3160);
nor U4251 (N_4251,N_3429,N_3361);
nand U4252 (N_4252,N_3587,N_3382);
nand U4253 (N_4253,N_3619,N_3140);
nor U4254 (N_4254,N_3623,N_3159);
nand U4255 (N_4255,N_3489,N_3256);
and U4256 (N_4256,N_3380,N_3621);
nand U4257 (N_4257,N_3622,N_3128);
or U4258 (N_4258,N_3160,N_3645);
and U4259 (N_4259,N_3232,N_3409);
and U4260 (N_4260,N_3647,N_3418);
nand U4261 (N_4261,N_3553,N_3497);
or U4262 (N_4262,N_3476,N_3685);
or U4263 (N_4263,N_3652,N_3579);
nand U4264 (N_4264,N_3402,N_3477);
nor U4265 (N_4265,N_3725,N_3419);
nand U4266 (N_4266,N_3650,N_3666);
and U4267 (N_4267,N_3654,N_3740);
and U4268 (N_4268,N_3429,N_3492);
and U4269 (N_4269,N_3419,N_3651);
nand U4270 (N_4270,N_3325,N_3674);
or U4271 (N_4271,N_3635,N_3189);
nand U4272 (N_4272,N_3715,N_3689);
or U4273 (N_4273,N_3363,N_3142);
nand U4274 (N_4274,N_3697,N_3170);
and U4275 (N_4275,N_3258,N_3138);
nand U4276 (N_4276,N_3401,N_3288);
and U4277 (N_4277,N_3471,N_3731);
nor U4278 (N_4278,N_3147,N_3604);
or U4279 (N_4279,N_3479,N_3656);
or U4280 (N_4280,N_3670,N_3533);
and U4281 (N_4281,N_3662,N_3748);
nor U4282 (N_4282,N_3270,N_3735);
xnor U4283 (N_4283,N_3698,N_3746);
nor U4284 (N_4284,N_3509,N_3571);
or U4285 (N_4285,N_3562,N_3439);
xnor U4286 (N_4286,N_3682,N_3159);
or U4287 (N_4287,N_3259,N_3434);
and U4288 (N_4288,N_3691,N_3326);
and U4289 (N_4289,N_3606,N_3678);
nand U4290 (N_4290,N_3172,N_3728);
and U4291 (N_4291,N_3591,N_3648);
or U4292 (N_4292,N_3151,N_3587);
or U4293 (N_4293,N_3286,N_3413);
nand U4294 (N_4294,N_3415,N_3423);
or U4295 (N_4295,N_3441,N_3626);
and U4296 (N_4296,N_3155,N_3272);
nand U4297 (N_4297,N_3433,N_3498);
nor U4298 (N_4298,N_3704,N_3190);
nand U4299 (N_4299,N_3171,N_3416);
nand U4300 (N_4300,N_3414,N_3360);
nand U4301 (N_4301,N_3236,N_3716);
nor U4302 (N_4302,N_3265,N_3718);
or U4303 (N_4303,N_3295,N_3589);
nand U4304 (N_4304,N_3385,N_3696);
nor U4305 (N_4305,N_3283,N_3644);
nand U4306 (N_4306,N_3170,N_3727);
xnor U4307 (N_4307,N_3516,N_3319);
nand U4308 (N_4308,N_3360,N_3278);
xnor U4309 (N_4309,N_3272,N_3214);
nand U4310 (N_4310,N_3256,N_3467);
nand U4311 (N_4311,N_3268,N_3667);
nor U4312 (N_4312,N_3492,N_3688);
nand U4313 (N_4313,N_3465,N_3395);
nand U4314 (N_4314,N_3243,N_3362);
xnor U4315 (N_4315,N_3572,N_3252);
nand U4316 (N_4316,N_3148,N_3400);
and U4317 (N_4317,N_3338,N_3718);
and U4318 (N_4318,N_3227,N_3396);
nand U4319 (N_4319,N_3223,N_3743);
nand U4320 (N_4320,N_3127,N_3684);
and U4321 (N_4321,N_3347,N_3597);
and U4322 (N_4322,N_3470,N_3368);
nor U4323 (N_4323,N_3322,N_3249);
nor U4324 (N_4324,N_3641,N_3311);
xnor U4325 (N_4325,N_3704,N_3467);
xnor U4326 (N_4326,N_3676,N_3257);
nor U4327 (N_4327,N_3255,N_3125);
or U4328 (N_4328,N_3201,N_3487);
or U4329 (N_4329,N_3548,N_3263);
xnor U4330 (N_4330,N_3143,N_3317);
and U4331 (N_4331,N_3559,N_3714);
nand U4332 (N_4332,N_3428,N_3463);
or U4333 (N_4333,N_3506,N_3635);
nand U4334 (N_4334,N_3164,N_3449);
nand U4335 (N_4335,N_3520,N_3274);
nand U4336 (N_4336,N_3511,N_3415);
and U4337 (N_4337,N_3368,N_3631);
nor U4338 (N_4338,N_3140,N_3174);
nand U4339 (N_4339,N_3484,N_3551);
and U4340 (N_4340,N_3308,N_3492);
xnor U4341 (N_4341,N_3746,N_3526);
or U4342 (N_4342,N_3281,N_3525);
and U4343 (N_4343,N_3177,N_3307);
or U4344 (N_4344,N_3593,N_3441);
and U4345 (N_4345,N_3318,N_3320);
nor U4346 (N_4346,N_3324,N_3694);
or U4347 (N_4347,N_3435,N_3725);
nand U4348 (N_4348,N_3388,N_3686);
nor U4349 (N_4349,N_3430,N_3609);
xor U4350 (N_4350,N_3290,N_3712);
nor U4351 (N_4351,N_3699,N_3656);
nand U4352 (N_4352,N_3336,N_3702);
xor U4353 (N_4353,N_3671,N_3615);
and U4354 (N_4354,N_3331,N_3716);
nor U4355 (N_4355,N_3379,N_3497);
nor U4356 (N_4356,N_3223,N_3373);
or U4357 (N_4357,N_3587,N_3284);
and U4358 (N_4358,N_3679,N_3262);
nor U4359 (N_4359,N_3688,N_3684);
nor U4360 (N_4360,N_3548,N_3584);
or U4361 (N_4361,N_3434,N_3182);
xnor U4362 (N_4362,N_3519,N_3460);
nor U4363 (N_4363,N_3195,N_3208);
xor U4364 (N_4364,N_3539,N_3687);
or U4365 (N_4365,N_3520,N_3356);
xnor U4366 (N_4366,N_3378,N_3164);
nand U4367 (N_4367,N_3175,N_3744);
xor U4368 (N_4368,N_3274,N_3594);
or U4369 (N_4369,N_3186,N_3506);
nor U4370 (N_4370,N_3684,N_3281);
and U4371 (N_4371,N_3611,N_3741);
nor U4372 (N_4372,N_3197,N_3415);
and U4373 (N_4373,N_3214,N_3247);
xnor U4374 (N_4374,N_3635,N_3533);
nand U4375 (N_4375,N_4262,N_4177);
or U4376 (N_4376,N_4315,N_3817);
or U4377 (N_4377,N_4123,N_4280);
and U4378 (N_4378,N_4001,N_3798);
nand U4379 (N_4379,N_4149,N_3826);
xnor U4380 (N_4380,N_4034,N_4341);
nand U4381 (N_4381,N_4121,N_4006);
xnor U4382 (N_4382,N_3775,N_4270);
nor U4383 (N_4383,N_4061,N_3875);
xor U4384 (N_4384,N_3959,N_3838);
xnor U4385 (N_4385,N_4134,N_4287);
nor U4386 (N_4386,N_4297,N_3890);
or U4387 (N_4387,N_4348,N_4035);
or U4388 (N_4388,N_4225,N_4019);
and U4389 (N_4389,N_4150,N_3753);
or U4390 (N_4390,N_3870,N_3984);
nor U4391 (N_4391,N_4336,N_3951);
and U4392 (N_4392,N_4263,N_3778);
and U4393 (N_4393,N_4255,N_3789);
nand U4394 (N_4394,N_4283,N_3972);
xor U4395 (N_4395,N_4248,N_4357);
and U4396 (N_4396,N_4093,N_4139);
xnor U4397 (N_4397,N_3835,N_4127);
nor U4398 (N_4398,N_3812,N_3954);
and U4399 (N_4399,N_3962,N_4200);
nor U4400 (N_4400,N_4013,N_3828);
nand U4401 (N_4401,N_4038,N_4004);
and U4402 (N_4402,N_4236,N_3925);
nor U4403 (N_4403,N_4055,N_4037);
and U4404 (N_4404,N_4163,N_4084);
xor U4405 (N_4405,N_4296,N_3821);
or U4406 (N_4406,N_4189,N_4063);
nand U4407 (N_4407,N_4036,N_4166);
nand U4408 (N_4408,N_4126,N_3788);
or U4409 (N_4409,N_3783,N_3806);
and U4410 (N_4410,N_4021,N_3889);
or U4411 (N_4411,N_4107,N_4042);
xor U4412 (N_4412,N_4095,N_4087);
xnor U4413 (N_4413,N_4051,N_4098);
or U4414 (N_4414,N_3764,N_4347);
nand U4415 (N_4415,N_4114,N_3865);
or U4416 (N_4416,N_4143,N_4085);
and U4417 (N_4417,N_3781,N_3937);
or U4418 (N_4418,N_3825,N_4302);
xor U4419 (N_4419,N_3864,N_4322);
xnor U4420 (N_4420,N_4254,N_4246);
nor U4421 (N_4421,N_3866,N_4062);
and U4422 (N_4422,N_4147,N_4181);
nor U4423 (N_4423,N_4113,N_4244);
xnor U4424 (N_4424,N_3832,N_4237);
or U4425 (N_4425,N_3861,N_4268);
and U4426 (N_4426,N_4281,N_4235);
or U4427 (N_4427,N_4140,N_4288);
and U4428 (N_4428,N_4015,N_3762);
or U4429 (N_4429,N_4202,N_4229);
or U4430 (N_4430,N_3916,N_3948);
or U4431 (N_4431,N_4290,N_4124);
or U4432 (N_4432,N_3772,N_3961);
xor U4433 (N_4433,N_3779,N_4151);
xor U4434 (N_4434,N_3852,N_4203);
and U4435 (N_4435,N_3897,N_4245);
xor U4436 (N_4436,N_4058,N_4090);
or U4437 (N_4437,N_4240,N_3769);
or U4438 (N_4438,N_4041,N_4313);
nor U4439 (N_4439,N_3845,N_4369);
or U4440 (N_4440,N_3914,N_3922);
nor U4441 (N_4441,N_4308,N_3928);
and U4442 (N_4442,N_3955,N_3807);
xor U4443 (N_4443,N_4223,N_3879);
nand U4444 (N_4444,N_3982,N_4108);
xor U4445 (N_4445,N_4269,N_3911);
xor U4446 (N_4446,N_4072,N_4299);
nor U4447 (N_4447,N_3985,N_3987);
or U4448 (N_4448,N_4188,N_4125);
nand U4449 (N_4449,N_4067,N_4106);
xnor U4450 (N_4450,N_3882,N_4137);
xor U4451 (N_4451,N_3795,N_4096);
nand U4452 (N_4452,N_4148,N_3856);
xnor U4453 (N_4453,N_4231,N_4184);
nand U4454 (N_4454,N_3824,N_3813);
nand U4455 (N_4455,N_3834,N_4243);
nor U4456 (N_4456,N_3917,N_4079);
nand U4457 (N_4457,N_4054,N_4094);
and U4458 (N_4458,N_3857,N_4170);
or U4459 (N_4459,N_4208,N_4216);
or U4460 (N_4460,N_4284,N_3858);
and U4461 (N_4461,N_3844,N_3968);
nor U4462 (N_4462,N_4352,N_4256);
and U4463 (N_4463,N_3923,N_3965);
or U4464 (N_4464,N_4122,N_3763);
or U4465 (N_4465,N_3767,N_4092);
nand U4466 (N_4466,N_3770,N_4179);
nand U4467 (N_4467,N_3973,N_4048);
or U4468 (N_4468,N_4100,N_4360);
nand U4469 (N_4469,N_4301,N_4345);
nor U4470 (N_4470,N_3886,N_4209);
nand U4471 (N_4471,N_4350,N_4278);
or U4472 (N_4472,N_3918,N_4167);
xnor U4473 (N_4473,N_3932,N_3904);
and U4474 (N_4474,N_4372,N_3888);
and U4475 (N_4475,N_3799,N_4059);
or U4476 (N_4476,N_3878,N_3940);
xnor U4477 (N_4477,N_4277,N_4312);
or U4478 (N_4478,N_4158,N_4339);
or U4479 (N_4479,N_3766,N_3883);
xnor U4480 (N_4480,N_4355,N_3797);
nand U4481 (N_4481,N_4213,N_4201);
and U4482 (N_4482,N_3862,N_3787);
xnor U4483 (N_4483,N_4053,N_4349);
xor U4484 (N_4484,N_3945,N_4191);
or U4485 (N_4485,N_4196,N_4309);
nor U4486 (N_4486,N_4195,N_3790);
nand U4487 (N_4487,N_4340,N_4138);
or U4488 (N_4488,N_4070,N_4161);
xnor U4489 (N_4489,N_4091,N_3823);
and U4490 (N_4490,N_4132,N_3809);
nor U4491 (N_4491,N_3872,N_3816);
or U4492 (N_4492,N_4077,N_4180);
nor U4493 (N_4493,N_4217,N_3854);
or U4494 (N_4494,N_4317,N_4344);
nand U4495 (N_4495,N_4076,N_4222);
and U4496 (N_4496,N_3998,N_4117);
nand U4497 (N_4497,N_4265,N_4071);
nor U4498 (N_4498,N_3771,N_4030);
or U4499 (N_4499,N_4185,N_4361);
or U4500 (N_4500,N_3943,N_4156);
and U4501 (N_4501,N_4286,N_3814);
nand U4502 (N_4502,N_4105,N_4174);
nand U4503 (N_4503,N_3805,N_4104);
or U4504 (N_4504,N_4324,N_3808);
nand U4505 (N_4505,N_4332,N_3927);
and U4506 (N_4506,N_4314,N_3876);
and U4507 (N_4507,N_3792,N_4016);
and U4508 (N_4508,N_4274,N_3933);
nand U4509 (N_4509,N_3877,N_3949);
nand U4510 (N_4510,N_4101,N_3830);
and U4511 (N_4511,N_4111,N_4227);
nand U4512 (N_4512,N_4285,N_3979);
and U4513 (N_4513,N_3907,N_3754);
xor U4514 (N_4514,N_3993,N_4261);
nand U4515 (N_4515,N_4320,N_3896);
xnor U4516 (N_4516,N_4289,N_4011);
xnor U4517 (N_4517,N_4178,N_4075);
xor U4518 (N_4518,N_3869,N_4146);
and U4519 (N_4519,N_3793,N_3990);
nand U4520 (N_4520,N_3853,N_4359);
and U4521 (N_4521,N_3751,N_3855);
nor U4522 (N_4522,N_4168,N_3801);
nand U4523 (N_4523,N_4258,N_3846);
or U4524 (N_4524,N_4321,N_3991);
and U4525 (N_4525,N_3784,N_3867);
and U4526 (N_4526,N_4131,N_3761);
or U4527 (N_4527,N_3837,N_3818);
and U4528 (N_4528,N_3782,N_4337);
or U4529 (N_4529,N_3803,N_4207);
nand U4530 (N_4530,N_4211,N_3836);
and U4531 (N_4531,N_3831,N_4120);
nand U4532 (N_4532,N_3786,N_3820);
nor U4533 (N_4533,N_4044,N_4017);
xor U4534 (N_4534,N_3941,N_3868);
nand U4535 (N_4535,N_4330,N_4102);
or U4536 (N_4536,N_4215,N_3765);
nor U4537 (N_4537,N_4366,N_4198);
xor U4538 (N_4538,N_3760,N_4026);
and U4539 (N_4539,N_4214,N_4218);
nand U4540 (N_4540,N_4129,N_4190);
nor U4541 (N_4541,N_3777,N_4230);
and U4542 (N_4542,N_3822,N_4005);
or U4543 (N_4543,N_3947,N_3924);
nor U4544 (N_4544,N_4292,N_3980);
xor U4545 (N_4545,N_4024,N_4039);
nor U4546 (N_4546,N_3859,N_4193);
xnor U4547 (N_4547,N_4353,N_3946);
and U4548 (N_4548,N_4014,N_4370);
nor U4549 (N_4549,N_4128,N_4069);
or U4550 (N_4550,N_3921,N_4160);
and U4551 (N_4551,N_3848,N_3910);
nand U4552 (N_4552,N_3989,N_4367);
xnor U4553 (N_4553,N_4241,N_3893);
or U4554 (N_4554,N_4298,N_4046);
nand U4555 (N_4555,N_3915,N_3986);
nor U4556 (N_4556,N_3935,N_4338);
nand U4557 (N_4557,N_4220,N_4354);
or U4558 (N_4558,N_4264,N_3847);
or U4559 (N_4559,N_4175,N_3849);
xnor U4560 (N_4560,N_4266,N_4010);
nor U4561 (N_4561,N_4343,N_4346);
xor U4562 (N_4562,N_3776,N_3981);
nor U4563 (N_4563,N_3895,N_3988);
xor U4564 (N_4564,N_4043,N_3898);
xnor U4565 (N_4565,N_4282,N_4373);
nand U4566 (N_4566,N_4194,N_3758);
nand U4567 (N_4567,N_4003,N_4169);
xnor U4568 (N_4568,N_4173,N_4275);
nand U4569 (N_4569,N_4257,N_4159);
xnor U4570 (N_4570,N_4239,N_3936);
nor U4571 (N_4571,N_4306,N_3887);
nor U4572 (N_4572,N_4116,N_4212);
and U4573 (N_4573,N_4089,N_3956);
and U4574 (N_4574,N_3796,N_4234);
nand U4575 (N_4575,N_4182,N_3755);
xor U4576 (N_4576,N_4119,N_3950);
nor U4577 (N_4577,N_4192,N_4144);
or U4578 (N_4578,N_4267,N_4065);
nand U4579 (N_4579,N_3995,N_4115);
nor U4580 (N_4580,N_3756,N_4233);
nand U4581 (N_4581,N_3811,N_4327);
and U4582 (N_4582,N_4103,N_4145);
xnor U4583 (N_4583,N_3912,N_3819);
nand U4584 (N_4584,N_4060,N_4365);
nand U4585 (N_4585,N_4002,N_4351);
nand U4586 (N_4586,N_4009,N_4221);
nor U4587 (N_4587,N_4056,N_4078);
and U4588 (N_4588,N_3942,N_3977);
or U4589 (N_4589,N_4097,N_3833);
nand U4590 (N_4590,N_4112,N_4291);
or U4591 (N_4591,N_3905,N_4165);
and U4592 (N_4592,N_3964,N_4325);
xor U4593 (N_4593,N_3920,N_4186);
nor U4594 (N_4594,N_3885,N_3841);
or U4595 (N_4595,N_3996,N_3850);
and U4596 (N_4596,N_4210,N_3815);
xnor U4597 (N_4597,N_4049,N_4323);
and U4598 (N_4598,N_3874,N_4300);
xnor U4599 (N_4599,N_3900,N_3960);
xor U4600 (N_4600,N_4232,N_4368);
xor U4601 (N_4601,N_3906,N_3938);
and U4602 (N_4602,N_4074,N_4066);
xnor U4603 (N_4603,N_3842,N_3967);
and U4604 (N_4604,N_4133,N_3759);
xnor U4605 (N_4605,N_4303,N_3902);
or U4606 (N_4606,N_4206,N_4154);
xor U4607 (N_4607,N_3903,N_3901);
nor U4608 (N_4608,N_4247,N_4228);
nand U4609 (N_4609,N_3880,N_4199);
or U4610 (N_4610,N_3939,N_4276);
nand U4611 (N_4611,N_4294,N_4226);
or U4612 (N_4612,N_4205,N_4068);
nand U4613 (N_4613,N_4335,N_4334);
nor U4614 (N_4614,N_3774,N_4025);
and U4615 (N_4615,N_3944,N_4007);
and U4616 (N_4616,N_3891,N_4157);
nand U4617 (N_4617,N_4374,N_3768);
xnor U4618 (N_4618,N_4242,N_4171);
nor U4619 (N_4619,N_4172,N_3800);
or U4620 (N_4620,N_3963,N_3791);
nor U4621 (N_4621,N_3999,N_4272);
nor U4622 (N_4622,N_4328,N_3931);
or U4623 (N_4623,N_4251,N_3802);
or U4624 (N_4624,N_4086,N_4135);
and U4625 (N_4625,N_4057,N_3804);
nand U4626 (N_4626,N_3952,N_4316);
nand U4627 (N_4627,N_3975,N_3953);
nor U4628 (N_4628,N_4176,N_3970);
or U4629 (N_4629,N_3863,N_4142);
xor U4630 (N_4630,N_3934,N_4155);
and U4631 (N_4631,N_3827,N_3884);
nand U4632 (N_4632,N_4141,N_4304);
nand U4633 (N_4633,N_4153,N_3757);
or U4634 (N_4634,N_4183,N_3908);
nand U4635 (N_4635,N_4136,N_4083);
nand U4636 (N_4636,N_3810,N_4080);
and U4637 (N_4637,N_3785,N_4187);
nand U4638 (N_4638,N_3873,N_4318);
or U4639 (N_4639,N_4082,N_4204);
nor U4640 (N_4640,N_4333,N_3958);
nor U4641 (N_4641,N_4273,N_3974);
nor U4642 (N_4642,N_3752,N_4259);
xnor U4643 (N_4643,N_4000,N_3930);
nand U4644 (N_4644,N_4088,N_3871);
nand U4645 (N_4645,N_4029,N_3892);
nor U4646 (N_4646,N_3978,N_4028);
or U4647 (N_4647,N_4224,N_4032);
xor U4648 (N_4648,N_4364,N_3881);
and U4649 (N_4649,N_4064,N_4356);
nand U4650 (N_4650,N_4073,N_4047);
and U4651 (N_4651,N_4307,N_3983);
nand U4652 (N_4652,N_4219,N_4031);
and U4653 (N_4653,N_4164,N_3997);
nor U4654 (N_4654,N_4279,N_3957);
xor U4655 (N_4655,N_4371,N_4293);
or U4656 (N_4656,N_4081,N_4099);
xor U4657 (N_4657,N_3829,N_4052);
xor U4658 (N_4658,N_4250,N_4109);
nand U4659 (N_4659,N_4331,N_3773);
or U4660 (N_4660,N_3750,N_4022);
or U4661 (N_4661,N_3919,N_3976);
and U4662 (N_4662,N_4249,N_3860);
and U4663 (N_4663,N_3851,N_3971);
xnor U4664 (N_4664,N_4152,N_3994);
and U4665 (N_4665,N_4362,N_3926);
nor U4666 (N_4666,N_4252,N_4018);
and U4667 (N_4667,N_4045,N_4342);
nor U4668 (N_4668,N_4358,N_4050);
nand U4669 (N_4669,N_3794,N_4027);
xnor U4670 (N_4670,N_4008,N_3839);
nor U4671 (N_4671,N_4130,N_3780);
nand U4672 (N_4672,N_4253,N_3913);
and U4673 (N_4673,N_4305,N_3969);
or U4674 (N_4674,N_4110,N_4260);
xnor U4675 (N_4675,N_3929,N_4326);
xor U4676 (N_4676,N_4319,N_3909);
or U4677 (N_4677,N_4197,N_4363);
or U4678 (N_4678,N_4033,N_3843);
nor U4679 (N_4679,N_3840,N_4023);
and U4680 (N_4680,N_4329,N_4012);
xor U4681 (N_4681,N_4311,N_4162);
and U4682 (N_4682,N_4310,N_3992);
xor U4683 (N_4683,N_3966,N_3899);
xnor U4684 (N_4684,N_4020,N_4295);
or U4685 (N_4685,N_3894,N_4118);
or U4686 (N_4686,N_4238,N_4040);
xor U4687 (N_4687,N_4271,N_3763);
and U4688 (N_4688,N_4358,N_3819);
nand U4689 (N_4689,N_4006,N_4139);
or U4690 (N_4690,N_4327,N_4088);
nand U4691 (N_4691,N_3889,N_3885);
nor U4692 (N_4692,N_4149,N_3865);
nand U4693 (N_4693,N_4275,N_4189);
nor U4694 (N_4694,N_4261,N_4312);
and U4695 (N_4695,N_3873,N_4090);
and U4696 (N_4696,N_4329,N_3930);
nand U4697 (N_4697,N_3905,N_3903);
xor U4698 (N_4698,N_4034,N_4291);
xor U4699 (N_4699,N_3910,N_4357);
and U4700 (N_4700,N_3757,N_3769);
or U4701 (N_4701,N_4090,N_3931);
nand U4702 (N_4702,N_3786,N_3776);
nor U4703 (N_4703,N_3762,N_3834);
xnor U4704 (N_4704,N_3915,N_4185);
and U4705 (N_4705,N_4285,N_3958);
xor U4706 (N_4706,N_4034,N_4233);
nand U4707 (N_4707,N_4153,N_4122);
nor U4708 (N_4708,N_4142,N_4100);
or U4709 (N_4709,N_3932,N_4114);
nor U4710 (N_4710,N_4175,N_3869);
or U4711 (N_4711,N_4172,N_3830);
and U4712 (N_4712,N_4024,N_3932);
nor U4713 (N_4713,N_4084,N_4344);
nor U4714 (N_4714,N_3783,N_3916);
and U4715 (N_4715,N_4030,N_4195);
or U4716 (N_4716,N_3768,N_4290);
or U4717 (N_4717,N_4145,N_4051);
xor U4718 (N_4718,N_3931,N_3981);
nand U4719 (N_4719,N_3975,N_4314);
nor U4720 (N_4720,N_3965,N_4118);
nor U4721 (N_4721,N_3898,N_4035);
and U4722 (N_4722,N_4216,N_3773);
nor U4723 (N_4723,N_3925,N_3980);
nand U4724 (N_4724,N_4122,N_4100);
nor U4725 (N_4725,N_3800,N_3986);
xor U4726 (N_4726,N_3779,N_4099);
or U4727 (N_4727,N_4073,N_3982);
and U4728 (N_4728,N_4136,N_4081);
or U4729 (N_4729,N_4271,N_3802);
nor U4730 (N_4730,N_4272,N_3980);
xnor U4731 (N_4731,N_4095,N_4225);
nor U4732 (N_4732,N_3839,N_3832);
nand U4733 (N_4733,N_4265,N_4343);
nor U4734 (N_4734,N_3778,N_3849);
or U4735 (N_4735,N_4142,N_3968);
and U4736 (N_4736,N_4015,N_3966);
or U4737 (N_4737,N_4043,N_4348);
nand U4738 (N_4738,N_4351,N_4343);
nand U4739 (N_4739,N_4054,N_3913);
or U4740 (N_4740,N_3977,N_4315);
nand U4741 (N_4741,N_3898,N_4001);
or U4742 (N_4742,N_3983,N_4371);
or U4743 (N_4743,N_4196,N_4217);
and U4744 (N_4744,N_4080,N_4239);
nor U4745 (N_4745,N_4296,N_3991);
and U4746 (N_4746,N_3912,N_4140);
xnor U4747 (N_4747,N_3789,N_3968);
xor U4748 (N_4748,N_4363,N_4058);
xnor U4749 (N_4749,N_3876,N_3777);
and U4750 (N_4750,N_4149,N_3968);
xnor U4751 (N_4751,N_3822,N_4342);
nand U4752 (N_4752,N_4094,N_4186);
or U4753 (N_4753,N_3795,N_3948);
nor U4754 (N_4754,N_4246,N_3751);
xnor U4755 (N_4755,N_4001,N_4029);
nand U4756 (N_4756,N_4303,N_4304);
xor U4757 (N_4757,N_4272,N_4209);
nand U4758 (N_4758,N_4363,N_4215);
nor U4759 (N_4759,N_4040,N_4341);
xnor U4760 (N_4760,N_3775,N_3859);
xor U4761 (N_4761,N_3750,N_3852);
nand U4762 (N_4762,N_3827,N_3985);
or U4763 (N_4763,N_4112,N_4212);
nand U4764 (N_4764,N_4003,N_4181);
xnor U4765 (N_4765,N_4206,N_3988);
nor U4766 (N_4766,N_4267,N_4269);
or U4767 (N_4767,N_4221,N_4036);
nor U4768 (N_4768,N_4230,N_4290);
xnor U4769 (N_4769,N_4083,N_4147);
nand U4770 (N_4770,N_3867,N_4198);
nand U4771 (N_4771,N_4317,N_3942);
and U4772 (N_4772,N_4188,N_4320);
or U4773 (N_4773,N_4050,N_4054);
nand U4774 (N_4774,N_4242,N_4238);
xnor U4775 (N_4775,N_4368,N_4353);
or U4776 (N_4776,N_4054,N_4329);
and U4777 (N_4777,N_4176,N_4155);
xnor U4778 (N_4778,N_4177,N_4141);
nor U4779 (N_4779,N_3947,N_4318);
nor U4780 (N_4780,N_3808,N_4049);
and U4781 (N_4781,N_4003,N_4253);
xor U4782 (N_4782,N_3840,N_3802);
xnor U4783 (N_4783,N_4178,N_4203);
nor U4784 (N_4784,N_4012,N_4005);
and U4785 (N_4785,N_4031,N_4310);
and U4786 (N_4786,N_4306,N_4256);
and U4787 (N_4787,N_3807,N_4309);
or U4788 (N_4788,N_4372,N_4225);
and U4789 (N_4789,N_3768,N_4100);
or U4790 (N_4790,N_4208,N_3947);
nor U4791 (N_4791,N_3755,N_4171);
nand U4792 (N_4792,N_3842,N_4344);
nor U4793 (N_4793,N_4014,N_3863);
nand U4794 (N_4794,N_4017,N_4320);
xnor U4795 (N_4795,N_4072,N_3754);
and U4796 (N_4796,N_3858,N_3908);
nand U4797 (N_4797,N_4145,N_4059);
nor U4798 (N_4798,N_3932,N_4203);
or U4799 (N_4799,N_4103,N_3975);
nand U4800 (N_4800,N_4146,N_4008);
or U4801 (N_4801,N_4201,N_3814);
or U4802 (N_4802,N_4079,N_3939);
nand U4803 (N_4803,N_3846,N_4168);
nand U4804 (N_4804,N_4172,N_4347);
and U4805 (N_4805,N_3995,N_3943);
and U4806 (N_4806,N_3752,N_4128);
or U4807 (N_4807,N_4318,N_4173);
or U4808 (N_4808,N_4255,N_4208);
nor U4809 (N_4809,N_3967,N_4232);
xnor U4810 (N_4810,N_4360,N_3853);
and U4811 (N_4811,N_4040,N_3889);
xnor U4812 (N_4812,N_4128,N_4083);
and U4813 (N_4813,N_4004,N_3967);
xor U4814 (N_4814,N_4253,N_4147);
xor U4815 (N_4815,N_4253,N_4239);
or U4816 (N_4816,N_3973,N_4284);
xnor U4817 (N_4817,N_4163,N_3987);
or U4818 (N_4818,N_3956,N_3914);
xor U4819 (N_4819,N_4307,N_4075);
xnor U4820 (N_4820,N_4016,N_4113);
xor U4821 (N_4821,N_3819,N_4090);
and U4822 (N_4822,N_3806,N_4208);
nand U4823 (N_4823,N_4269,N_4237);
and U4824 (N_4824,N_4037,N_4118);
nand U4825 (N_4825,N_4108,N_4092);
or U4826 (N_4826,N_4359,N_3761);
nand U4827 (N_4827,N_3869,N_4152);
and U4828 (N_4828,N_4172,N_3805);
nor U4829 (N_4829,N_4286,N_3913);
or U4830 (N_4830,N_3895,N_4298);
and U4831 (N_4831,N_3841,N_4232);
and U4832 (N_4832,N_3885,N_3947);
nor U4833 (N_4833,N_3954,N_3936);
or U4834 (N_4834,N_3976,N_4148);
nor U4835 (N_4835,N_4070,N_3770);
nand U4836 (N_4836,N_4254,N_3752);
xnor U4837 (N_4837,N_4154,N_4106);
xor U4838 (N_4838,N_3909,N_3867);
and U4839 (N_4839,N_4162,N_3830);
xnor U4840 (N_4840,N_4222,N_4303);
xor U4841 (N_4841,N_4274,N_4162);
xnor U4842 (N_4842,N_3901,N_4246);
xnor U4843 (N_4843,N_3785,N_3830);
xnor U4844 (N_4844,N_4201,N_4090);
nor U4845 (N_4845,N_3927,N_4055);
or U4846 (N_4846,N_4009,N_4081);
and U4847 (N_4847,N_4192,N_4059);
or U4848 (N_4848,N_4293,N_4159);
xnor U4849 (N_4849,N_4124,N_4012);
and U4850 (N_4850,N_4038,N_4315);
xnor U4851 (N_4851,N_4014,N_4068);
xor U4852 (N_4852,N_3894,N_3882);
and U4853 (N_4853,N_3854,N_3964);
xnor U4854 (N_4854,N_3848,N_4329);
and U4855 (N_4855,N_3782,N_4289);
xor U4856 (N_4856,N_4170,N_4227);
and U4857 (N_4857,N_4101,N_3779);
or U4858 (N_4858,N_4299,N_4108);
nand U4859 (N_4859,N_3848,N_4243);
nand U4860 (N_4860,N_4274,N_3751);
and U4861 (N_4861,N_4036,N_4259);
nor U4862 (N_4862,N_3897,N_4033);
nand U4863 (N_4863,N_3928,N_4070);
nand U4864 (N_4864,N_4322,N_4197);
and U4865 (N_4865,N_3774,N_3927);
nor U4866 (N_4866,N_4011,N_4068);
or U4867 (N_4867,N_4060,N_3778);
and U4868 (N_4868,N_3874,N_3884);
nor U4869 (N_4869,N_4326,N_4011);
or U4870 (N_4870,N_4362,N_3917);
nand U4871 (N_4871,N_4226,N_4290);
and U4872 (N_4872,N_4326,N_4169);
xor U4873 (N_4873,N_4213,N_4365);
or U4874 (N_4874,N_4214,N_3923);
or U4875 (N_4875,N_4149,N_4228);
and U4876 (N_4876,N_3963,N_3930);
nand U4877 (N_4877,N_4233,N_4025);
or U4878 (N_4878,N_4208,N_4263);
nor U4879 (N_4879,N_4020,N_4148);
xor U4880 (N_4880,N_3898,N_3756);
nand U4881 (N_4881,N_4232,N_3966);
xnor U4882 (N_4882,N_3896,N_4173);
nand U4883 (N_4883,N_4008,N_4304);
xnor U4884 (N_4884,N_4122,N_3988);
or U4885 (N_4885,N_3834,N_4303);
and U4886 (N_4886,N_4012,N_3888);
or U4887 (N_4887,N_4070,N_4047);
or U4888 (N_4888,N_3805,N_3755);
nand U4889 (N_4889,N_4144,N_3913);
or U4890 (N_4890,N_3982,N_4080);
nor U4891 (N_4891,N_4325,N_3818);
nor U4892 (N_4892,N_4321,N_3820);
xor U4893 (N_4893,N_3938,N_3819);
or U4894 (N_4894,N_3944,N_3881);
or U4895 (N_4895,N_4053,N_3880);
xnor U4896 (N_4896,N_3951,N_4181);
xnor U4897 (N_4897,N_3910,N_4095);
or U4898 (N_4898,N_4186,N_4029);
and U4899 (N_4899,N_4370,N_3934);
nand U4900 (N_4900,N_4302,N_3964);
nor U4901 (N_4901,N_4340,N_4314);
and U4902 (N_4902,N_4363,N_3759);
xor U4903 (N_4903,N_4343,N_4060);
or U4904 (N_4904,N_4039,N_4028);
nor U4905 (N_4905,N_3838,N_4031);
or U4906 (N_4906,N_3805,N_3917);
xnor U4907 (N_4907,N_4203,N_4262);
nand U4908 (N_4908,N_4085,N_4014);
nand U4909 (N_4909,N_4133,N_4057);
xor U4910 (N_4910,N_4198,N_3773);
nand U4911 (N_4911,N_4358,N_4270);
xor U4912 (N_4912,N_4172,N_4056);
nand U4913 (N_4913,N_4250,N_4029);
and U4914 (N_4914,N_4024,N_3785);
and U4915 (N_4915,N_4075,N_4276);
and U4916 (N_4916,N_3751,N_3903);
or U4917 (N_4917,N_4103,N_4017);
xnor U4918 (N_4918,N_3996,N_3908);
nand U4919 (N_4919,N_4122,N_3977);
xnor U4920 (N_4920,N_3783,N_4261);
or U4921 (N_4921,N_4225,N_4068);
nand U4922 (N_4922,N_4328,N_4368);
or U4923 (N_4923,N_4069,N_3940);
and U4924 (N_4924,N_4171,N_4326);
nor U4925 (N_4925,N_4082,N_3908);
and U4926 (N_4926,N_3794,N_3861);
nor U4927 (N_4927,N_4067,N_3794);
or U4928 (N_4928,N_4132,N_4250);
xnor U4929 (N_4929,N_3873,N_4259);
or U4930 (N_4930,N_4262,N_3769);
nand U4931 (N_4931,N_3977,N_3907);
nor U4932 (N_4932,N_4015,N_4269);
nand U4933 (N_4933,N_4298,N_4295);
nor U4934 (N_4934,N_4161,N_4126);
and U4935 (N_4935,N_4366,N_4159);
and U4936 (N_4936,N_4368,N_3936);
xor U4937 (N_4937,N_4336,N_4188);
xor U4938 (N_4938,N_4361,N_4113);
nor U4939 (N_4939,N_3916,N_4370);
nand U4940 (N_4940,N_4009,N_3968);
nor U4941 (N_4941,N_4124,N_3893);
nor U4942 (N_4942,N_4075,N_4069);
nand U4943 (N_4943,N_4058,N_4123);
nand U4944 (N_4944,N_3757,N_3761);
xnor U4945 (N_4945,N_4176,N_4255);
and U4946 (N_4946,N_4307,N_4351);
nor U4947 (N_4947,N_4302,N_4339);
nand U4948 (N_4948,N_4152,N_3948);
or U4949 (N_4949,N_3885,N_4203);
and U4950 (N_4950,N_4162,N_3956);
nor U4951 (N_4951,N_3927,N_4290);
nand U4952 (N_4952,N_4352,N_3896);
nand U4953 (N_4953,N_3866,N_4330);
or U4954 (N_4954,N_4285,N_4055);
xor U4955 (N_4955,N_4181,N_4081);
nand U4956 (N_4956,N_3998,N_4262);
nand U4957 (N_4957,N_4117,N_4015);
or U4958 (N_4958,N_4307,N_3865);
and U4959 (N_4959,N_4139,N_3812);
and U4960 (N_4960,N_4201,N_3826);
and U4961 (N_4961,N_4049,N_4106);
or U4962 (N_4962,N_4092,N_3843);
nor U4963 (N_4963,N_3811,N_4219);
and U4964 (N_4964,N_4246,N_3863);
xor U4965 (N_4965,N_4240,N_3991);
nor U4966 (N_4966,N_3990,N_3839);
nor U4967 (N_4967,N_4132,N_4272);
xnor U4968 (N_4968,N_3984,N_3882);
nand U4969 (N_4969,N_3853,N_4143);
or U4970 (N_4970,N_4108,N_3914);
or U4971 (N_4971,N_3864,N_4047);
nand U4972 (N_4972,N_4120,N_3918);
nand U4973 (N_4973,N_3832,N_4162);
nor U4974 (N_4974,N_3789,N_3811);
and U4975 (N_4975,N_4027,N_3815);
xnor U4976 (N_4976,N_3847,N_4175);
or U4977 (N_4977,N_3967,N_3867);
nor U4978 (N_4978,N_3891,N_4080);
xnor U4979 (N_4979,N_3762,N_4264);
or U4980 (N_4980,N_4099,N_4317);
nand U4981 (N_4981,N_3906,N_3967);
nand U4982 (N_4982,N_4250,N_3771);
or U4983 (N_4983,N_4147,N_4351);
nor U4984 (N_4984,N_3928,N_4347);
nor U4985 (N_4985,N_4026,N_4100);
nand U4986 (N_4986,N_3985,N_3964);
nand U4987 (N_4987,N_3790,N_4274);
nor U4988 (N_4988,N_4114,N_4341);
xor U4989 (N_4989,N_3946,N_4257);
xnor U4990 (N_4990,N_4314,N_3939);
nor U4991 (N_4991,N_3926,N_4127);
xor U4992 (N_4992,N_3884,N_3761);
xor U4993 (N_4993,N_4324,N_3917);
nand U4994 (N_4994,N_3928,N_4176);
or U4995 (N_4995,N_3983,N_4278);
nand U4996 (N_4996,N_3902,N_4284);
or U4997 (N_4997,N_4195,N_4070);
nor U4998 (N_4998,N_4262,N_4095);
and U4999 (N_4999,N_3777,N_3857);
nor U5000 (N_5000,N_4573,N_4670);
xor U5001 (N_5001,N_4383,N_4871);
or U5002 (N_5002,N_4745,N_4813);
nand U5003 (N_5003,N_4420,N_4946);
or U5004 (N_5004,N_4993,N_4534);
or U5005 (N_5005,N_4977,N_4866);
or U5006 (N_5006,N_4679,N_4740);
or U5007 (N_5007,N_4390,N_4429);
or U5008 (N_5008,N_4956,N_4439);
xnor U5009 (N_5009,N_4730,N_4673);
nor U5010 (N_5010,N_4845,N_4792);
xnor U5011 (N_5011,N_4947,N_4450);
xnor U5012 (N_5012,N_4413,N_4958);
xnor U5013 (N_5013,N_4680,N_4566);
xor U5014 (N_5014,N_4384,N_4378);
or U5015 (N_5015,N_4481,N_4614);
or U5016 (N_5016,N_4987,N_4437);
and U5017 (N_5017,N_4391,N_4684);
xor U5018 (N_5018,N_4436,N_4662);
nor U5019 (N_5019,N_4504,N_4830);
or U5020 (N_5020,N_4715,N_4774);
xnor U5021 (N_5021,N_4948,N_4550);
and U5022 (N_5022,N_4982,N_4878);
nor U5023 (N_5023,N_4756,N_4454);
and U5024 (N_5024,N_4653,N_4621);
nand U5025 (N_5025,N_4505,N_4885);
and U5026 (N_5026,N_4508,N_4905);
xor U5027 (N_5027,N_4640,N_4913);
or U5028 (N_5028,N_4605,N_4512);
or U5029 (N_5029,N_4906,N_4953);
and U5030 (N_5030,N_4582,N_4775);
xor U5031 (N_5031,N_4585,N_4691);
and U5032 (N_5032,N_4502,N_4549);
and U5033 (N_5033,N_4951,N_4942);
nor U5034 (N_5034,N_4786,N_4731);
nand U5035 (N_5035,N_4506,N_4648);
nand U5036 (N_5036,N_4674,N_4675);
nand U5037 (N_5037,N_4726,N_4791);
nand U5038 (N_5038,N_4503,N_4753);
and U5039 (N_5039,N_4625,N_4750);
xnor U5040 (N_5040,N_4485,N_4552);
or U5041 (N_5041,N_4794,N_4613);
nand U5042 (N_5042,N_4989,N_4421);
and U5043 (N_5043,N_4583,N_4759);
xor U5044 (N_5044,N_4842,N_4941);
xor U5045 (N_5045,N_4976,N_4603);
nand U5046 (N_5046,N_4397,N_4382);
xor U5047 (N_5047,N_4782,N_4672);
nand U5048 (N_5048,N_4797,N_4570);
nor U5049 (N_5049,N_4881,N_4516);
nand U5050 (N_5050,N_4839,N_4994);
and U5051 (N_5051,N_4960,N_4571);
nand U5052 (N_5052,N_4376,N_4379);
and U5053 (N_5053,N_4617,N_4739);
xnor U5054 (N_5054,N_4712,N_4800);
and U5055 (N_5055,N_4575,N_4627);
xor U5056 (N_5056,N_4579,N_4785);
or U5057 (N_5057,N_4464,N_4381);
nor U5058 (N_5058,N_4581,N_4689);
nor U5059 (N_5059,N_4387,N_4499);
or U5060 (N_5060,N_4696,N_4978);
xor U5061 (N_5061,N_4523,N_4686);
or U5062 (N_5062,N_4752,N_4854);
xnor U5063 (N_5063,N_4798,N_4496);
nor U5064 (N_5064,N_4713,N_4404);
nor U5065 (N_5065,N_4709,N_4911);
xor U5066 (N_5066,N_4644,N_4665);
nor U5067 (N_5067,N_4377,N_4862);
or U5068 (N_5068,N_4923,N_4576);
nor U5069 (N_5069,N_4417,N_4443);
nand U5070 (N_5070,N_4940,N_4449);
or U5071 (N_5071,N_4388,N_4755);
xor U5072 (N_5072,N_4671,N_4721);
xnor U5073 (N_5073,N_4760,N_4749);
xor U5074 (N_5074,N_4385,N_4761);
or U5075 (N_5075,N_4668,N_4427);
nor U5076 (N_5076,N_4807,N_4804);
xnor U5077 (N_5077,N_4663,N_4495);
or U5078 (N_5078,N_4514,N_4560);
or U5079 (N_5079,N_4771,N_4902);
nand U5080 (N_5080,N_4536,N_4773);
xor U5081 (N_5081,N_4546,N_4667);
xnor U5082 (N_5082,N_4971,N_4848);
nor U5083 (N_5083,N_4861,N_4984);
and U5084 (N_5084,N_4895,N_4612);
and U5085 (N_5085,N_4720,N_4635);
or U5086 (N_5086,N_4875,N_4609);
nor U5087 (N_5087,N_4727,N_4400);
and U5088 (N_5088,N_4882,N_4451);
nand U5089 (N_5089,N_4944,N_4651);
xor U5090 (N_5090,N_4970,N_4735);
or U5091 (N_5091,N_4434,N_4584);
or U5092 (N_5092,N_4828,N_4950);
or U5093 (N_5093,N_4685,N_4746);
or U5094 (N_5094,N_4949,N_4452);
and U5095 (N_5095,N_4530,N_4867);
xor U5096 (N_5096,N_4559,N_4593);
nor U5097 (N_5097,N_4743,N_4849);
nor U5098 (N_5098,N_4961,N_4986);
and U5099 (N_5099,N_4545,N_4393);
and U5100 (N_5100,N_4482,N_4541);
nor U5101 (N_5101,N_4469,N_4654);
xor U5102 (N_5102,N_4925,N_4580);
xnor U5103 (N_5103,N_4988,N_4677);
xnor U5104 (N_5104,N_4995,N_4922);
or U5105 (N_5105,N_4710,N_4729);
xnor U5106 (N_5106,N_4836,N_4733);
and U5107 (N_5107,N_4399,N_4569);
nor U5108 (N_5108,N_4870,N_4493);
xor U5109 (N_5109,N_4829,N_4463);
nor U5110 (N_5110,N_4738,N_4600);
or U5111 (N_5111,N_4456,N_4490);
nor U5112 (N_5112,N_4525,N_4630);
and U5113 (N_5113,N_4426,N_4998);
nor U5114 (N_5114,N_4847,N_4466);
or U5115 (N_5115,N_4598,N_4823);
nor U5116 (N_5116,N_4835,N_4962);
xnor U5117 (N_5117,N_4589,N_4532);
nand U5118 (N_5118,N_4938,N_4824);
nand U5119 (N_5119,N_4412,N_4681);
nor U5120 (N_5120,N_4687,N_4623);
xnor U5121 (N_5121,N_4954,N_4487);
and U5122 (N_5122,N_4535,N_4943);
nand U5123 (N_5123,N_4860,N_4915);
nor U5124 (N_5124,N_4781,N_4544);
or U5125 (N_5125,N_4747,N_4457);
nand U5126 (N_5126,N_4821,N_4921);
nand U5127 (N_5127,N_4784,N_4478);
xor U5128 (N_5128,N_4832,N_4779);
or U5129 (N_5129,N_4834,N_4825);
nor U5130 (N_5130,N_4893,N_4539);
and U5131 (N_5131,N_4442,N_4997);
nor U5132 (N_5132,N_4594,N_4879);
nor U5133 (N_5133,N_4669,N_4891);
nor U5134 (N_5134,N_4856,N_4886);
and U5135 (N_5135,N_4957,N_4959);
nor U5136 (N_5136,N_4857,N_4725);
nand U5137 (N_5137,N_4864,N_4742);
nand U5138 (N_5138,N_4990,N_4551);
or U5139 (N_5139,N_4701,N_4751);
xnor U5140 (N_5140,N_4587,N_4386);
and U5141 (N_5141,N_4766,N_4658);
nand U5142 (N_5142,N_4980,N_4409);
or U5143 (N_5143,N_4458,N_4432);
or U5144 (N_5144,N_4966,N_4477);
xor U5145 (N_5145,N_4897,N_4642);
xnor U5146 (N_5146,N_4690,N_4435);
xor U5147 (N_5147,N_4611,N_4963);
and U5148 (N_5148,N_4419,N_4732);
or U5149 (N_5149,N_4765,N_4935);
nor U5150 (N_5150,N_4931,N_4633);
and U5151 (N_5151,N_4933,N_4380);
or U5152 (N_5152,N_4416,N_4641);
nand U5153 (N_5153,N_4634,N_4799);
and U5154 (N_5154,N_4637,N_4407);
xor U5155 (N_5155,N_4453,N_4850);
nor U5156 (N_5156,N_4812,N_4707);
nor U5157 (N_5157,N_4736,N_4903);
or U5158 (N_5158,N_4652,N_4822);
nand U5159 (N_5159,N_4700,N_4405);
nand U5160 (N_5160,N_4441,N_4428);
nand U5161 (N_5161,N_4607,N_4618);
xor U5162 (N_5162,N_4410,N_4790);
or U5163 (N_5163,N_4659,N_4509);
nand U5164 (N_5164,N_4447,N_4928);
nor U5165 (N_5165,N_4554,N_4926);
and U5166 (N_5166,N_4664,N_4425);
xor U5167 (N_5167,N_4719,N_4969);
nand U5168 (N_5168,N_4558,N_4704);
xnor U5169 (N_5169,N_4567,N_4770);
nor U5170 (N_5170,N_4661,N_4624);
xor U5171 (N_5171,N_4778,N_4757);
nor U5172 (N_5172,N_4952,N_4531);
nand U5173 (N_5173,N_4924,N_4810);
xor U5174 (N_5174,N_4660,N_4401);
xor U5175 (N_5175,N_4929,N_4446);
nand U5176 (N_5176,N_4803,N_4939);
nand U5177 (N_5177,N_4484,N_4565);
nor U5178 (N_5178,N_4787,N_4595);
xor U5179 (N_5179,N_4843,N_4471);
or U5180 (N_5180,N_4838,N_4392);
xnor U5181 (N_5181,N_4932,N_4455);
nand U5182 (N_5182,N_4851,N_4480);
xnor U5183 (N_5183,N_4894,N_4936);
nor U5184 (N_5184,N_4876,N_4744);
or U5185 (N_5185,N_4795,N_4826);
xor U5186 (N_5186,N_4398,N_4394);
or U5187 (N_5187,N_4459,N_4622);
nor U5188 (N_5188,N_4853,N_4763);
or U5189 (N_5189,N_4568,N_4473);
and U5190 (N_5190,N_4937,N_4748);
nor U5191 (N_5191,N_4793,N_4811);
nand U5192 (N_5192,N_4991,N_4780);
xnor U5193 (N_5193,N_4467,N_4840);
and U5194 (N_5194,N_4896,N_4688);
or U5195 (N_5195,N_4912,N_4403);
or U5196 (N_5196,N_4494,N_4777);
or U5197 (N_5197,N_4528,N_4515);
and U5198 (N_5198,N_4483,N_4796);
or U5199 (N_5199,N_4734,N_4979);
nor U5200 (N_5200,N_4917,N_4999);
nor U5201 (N_5201,N_4975,N_4527);
nand U5202 (N_5202,N_4533,N_4817);
nand U5203 (N_5203,N_4629,N_4815);
xor U5204 (N_5204,N_4764,N_4522);
nor U5205 (N_5205,N_4448,N_4521);
xnor U5206 (N_5206,N_4908,N_4722);
nand U5207 (N_5207,N_4555,N_4406);
or U5208 (N_5208,N_4683,N_4865);
nand U5209 (N_5209,N_4604,N_4626);
or U5210 (N_5210,N_4694,N_4818);
nand U5211 (N_5211,N_4474,N_4968);
and U5212 (N_5212,N_4837,N_4819);
or U5213 (N_5213,N_4616,N_4714);
nor U5214 (N_5214,N_4945,N_4649);
and U5215 (N_5215,N_4880,N_4577);
and U5216 (N_5216,N_4646,N_4596);
nand U5217 (N_5217,N_4591,N_4476);
nor U5218 (N_5218,N_4619,N_4547);
and U5219 (N_5219,N_4833,N_4820);
and U5220 (N_5220,N_4754,N_4898);
xnor U5221 (N_5221,N_4762,N_4656);
xor U5222 (N_5222,N_4973,N_4491);
nor U5223 (N_5223,N_4827,N_4708);
and U5224 (N_5224,N_4615,N_4444);
and U5225 (N_5225,N_4438,N_4996);
and U5226 (N_5226,N_4479,N_4666);
or U5227 (N_5227,N_4588,N_4553);
nand U5228 (N_5228,N_4507,N_4657);
nor U5229 (N_5229,N_4647,N_4572);
xor U5230 (N_5230,N_4841,N_4716);
nor U5231 (N_5231,N_4855,N_4529);
or U5232 (N_5232,N_4610,N_4518);
and U5233 (N_5233,N_4538,N_4557);
and U5234 (N_5234,N_4498,N_4769);
and U5235 (N_5235,N_4678,N_4934);
and U5236 (N_5236,N_4914,N_4389);
nor U5237 (N_5237,N_4645,N_4741);
nor U5238 (N_5238,N_4564,N_4758);
or U5239 (N_5239,N_4517,N_4431);
or U5240 (N_5240,N_4693,N_4816);
or U5241 (N_5241,N_4433,N_4983);
and U5242 (N_5242,N_4526,N_4711);
xnor U5243 (N_5243,N_4972,N_4702);
nand U5244 (N_5244,N_4461,N_4703);
or U5245 (N_5245,N_4814,N_4873);
or U5246 (N_5246,N_4422,N_4974);
or U5247 (N_5247,N_4801,N_4904);
nand U5248 (N_5248,N_4632,N_4465);
nor U5249 (N_5249,N_4501,N_4520);
nor U5250 (N_5250,N_4601,N_4964);
and U5251 (N_5251,N_4806,N_4631);
nand U5252 (N_5252,N_4486,N_4430);
nand U5253 (N_5253,N_4643,N_4985);
xnor U5254 (N_5254,N_4682,N_4537);
xnor U5255 (N_5255,N_4883,N_4788);
and U5256 (N_5256,N_4863,N_4440);
and U5257 (N_5257,N_4650,N_4424);
and U5258 (N_5258,N_4699,N_4415);
nand U5259 (N_5259,N_4488,N_4590);
xnor U5260 (N_5260,N_4918,N_4890);
nor U5261 (N_5261,N_4916,N_4723);
and U5262 (N_5262,N_4561,N_4414);
nand U5263 (N_5263,N_4697,N_4805);
or U5264 (N_5264,N_4556,N_4638);
nand U5265 (N_5265,N_4869,N_4844);
xor U5266 (N_5266,N_4767,N_4639);
nand U5267 (N_5267,N_4563,N_4472);
xor U5268 (N_5268,N_4602,N_4909);
xnor U5269 (N_5269,N_4955,N_4606);
nand U5270 (N_5270,N_4592,N_4899);
nand U5271 (N_5271,N_4408,N_4511);
and U5272 (N_5272,N_4724,N_4868);
xnor U5273 (N_5273,N_4872,N_4470);
nor U5274 (N_5274,N_4900,N_4468);
nor U5275 (N_5275,N_4620,N_4887);
or U5276 (N_5276,N_4846,N_4578);
and U5277 (N_5277,N_4831,N_4396);
nand U5278 (N_5278,N_4965,N_4423);
nor U5279 (N_5279,N_4809,N_4475);
xnor U5280 (N_5280,N_4717,N_4608);
xnor U5281 (N_5281,N_4889,N_4852);
and U5282 (N_5282,N_4884,N_4728);
and U5283 (N_5283,N_4574,N_4586);
xor U5284 (N_5284,N_4992,N_4930);
or U5285 (N_5285,N_4519,N_4901);
nor U5286 (N_5286,N_4920,N_4789);
nand U5287 (N_5287,N_4411,N_4698);
nor U5288 (N_5288,N_4737,N_4597);
nor U5289 (N_5289,N_4636,N_4892);
or U5290 (N_5290,N_4874,N_4858);
xor U5291 (N_5291,N_4500,N_4776);
xor U5292 (N_5292,N_4460,N_4445);
nand U5293 (N_5293,N_4543,N_4497);
nor U5294 (N_5294,N_4513,N_4705);
nor U5295 (N_5295,N_4375,N_4462);
nand U5296 (N_5296,N_4562,N_4524);
and U5297 (N_5297,N_4695,N_4888);
nor U5298 (N_5298,N_4542,N_4967);
and U5299 (N_5299,N_4927,N_4540);
xnor U5300 (N_5300,N_4628,N_4418);
nor U5301 (N_5301,N_4706,N_4808);
and U5302 (N_5302,N_4859,N_4910);
nor U5303 (N_5303,N_4877,N_4599);
or U5304 (N_5304,N_4489,N_4402);
xor U5305 (N_5305,N_4919,N_4676);
nand U5306 (N_5306,N_4510,N_4772);
nand U5307 (N_5307,N_4548,N_4655);
nand U5308 (N_5308,N_4692,N_4783);
and U5309 (N_5309,N_4718,N_4802);
nand U5310 (N_5310,N_4981,N_4907);
nor U5311 (N_5311,N_4492,N_4768);
or U5312 (N_5312,N_4395,N_4984);
nand U5313 (N_5313,N_4395,N_4756);
nand U5314 (N_5314,N_4653,N_4396);
nor U5315 (N_5315,N_4403,N_4829);
or U5316 (N_5316,N_4724,N_4558);
nand U5317 (N_5317,N_4678,N_4595);
and U5318 (N_5318,N_4594,N_4501);
or U5319 (N_5319,N_4738,N_4848);
and U5320 (N_5320,N_4732,N_4911);
nor U5321 (N_5321,N_4558,N_4442);
nand U5322 (N_5322,N_4976,N_4906);
nand U5323 (N_5323,N_4816,N_4795);
nor U5324 (N_5324,N_4637,N_4396);
nand U5325 (N_5325,N_4536,N_4758);
nor U5326 (N_5326,N_4722,N_4949);
or U5327 (N_5327,N_4732,N_4885);
or U5328 (N_5328,N_4992,N_4714);
or U5329 (N_5329,N_4848,N_4577);
nor U5330 (N_5330,N_4658,N_4945);
xor U5331 (N_5331,N_4540,N_4778);
and U5332 (N_5332,N_4416,N_4677);
or U5333 (N_5333,N_4588,N_4658);
and U5334 (N_5334,N_4521,N_4578);
xnor U5335 (N_5335,N_4376,N_4469);
xnor U5336 (N_5336,N_4473,N_4604);
and U5337 (N_5337,N_4472,N_4794);
or U5338 (N_5338,N_4939,N_4888);
or U5339 (N_5339,N_4763,N_4533);
nand U5340 (N_5340,N_4817,N_4519);
or U5341 (N_5341,N_4529,N_4593);
nor U5342 (N_5342,N_4776,N_4470);
nand U5343 (N_5343,N_4793,N_4481);
xnor U5344 (N_5344,N_4533,N_4431);
nor U5345 (N_5345,N_4593,N_4509);
and U5346 (N_5346,N_4844,N_4589);
and U5347 (N_5347,N_4904,N_4600);
xnor U5348 (N_5348,N_4538,N_4523);
xor U5349 (N_5349,N_4392,N_4916);
and U5350 (N_5350,N_4467,N_4961);
or U5351 (N_5351,N_4835,N_4636);
or U5352 (N_5352,N_4897,N_4422);
nor U5353 (N_5353,N_4533,N_4590);
and U5354 (N_5354,N_4400,N_4630);
nor U5355 (N_5355,N_4614,N_4881);
nand U5356 (N_5356,N_4846,N_4732);
nand U5357 (N_5357,N_4853,N_4581);
or U5358 (N_5358,N_4764,N_4763);
nor U5359 (N_5359,N_4725,N_4995);
nor U5360 (N_5360,N_4964,N_4639);
or U5361 (N_5361,N_4843,N_4807);
nor U5362 (N_5362,N_4773,N_4431);
nor U5363 (N_5363,N_4772,N_4624);
xor U5364 (N_5364,N_4933,N_4981);
nor U5365 (N_5365,N_4830,N_4896);
and U5366 (N_5366,N_4606,N_4895);
xnor U5367 (N_5367,N_4619,N_4469);
nor U5368 (N_5368,N_4730,N_4826);
nand U5369 (N_5369,N_4604,N_4435);
nand U5370 (N_5370,N_4513,N_4557);
xnor U5371 (N_5371,N_4442,N_4779);
xnor U5372 (N_5372,N_4703,N_4793);
and U5373 (N_5373,N_4523,N_4681);
nand U5374 (N_5374,N_4725,N_4867);
xor U5375 (N_5375,N_4751,N_4755);
and U5376 (N_5376,N_4937,N_4892);
or U5377 (N_5377,N_4513,N_4910);
nand U5378 (N_5378,N_4386,N_4487);
and U5379 (N_5379,N_4466,N_4741);
nor U5380 (N_5380,N_4876,N_4616);
and U5381 (N_5381,N_4910,N_4839);
nor U5382 (N_5382,N_4851,N_4960);
nor U5383 (N_5383,N_4659,N_4847);
or U5384 (N_5384,N_4699,N_4965);
or U5385 (N_5385,N_4832,N_4602);
and U5386 (N_5386,N_4649,N_4506);
nor U5387 (N_5387,N_4621,N_4847);
nand U5388 (N_5388,N_4816,N_4645);
nor U5389 (N_5389,N_4410,N_4571);
and U5390 (N_5390,N_4615,N_4724);
nand U5391 (N_5391,N_4836,N_4942);
and U5392 (N_5392,N_4731,N_4735);
nor U5393 (N_5393,N_4835,N_4477);
nand U5394 (N_5394,N_4565,N_4923);
or U5395 (N_5395,N_4598,N_4520);
and U5396 (N_5396,N_4935,N_4929);
and U5397 (N_5397,N_4489,N_4728);
nor U5398 (N_5398,N_4502,N_4962);
or U5399 (N_5399,N_4630,N_4759);
xnor U5400 (N_5400,N_4784,N_4686);
xnor U5401 (N_5401,N_4609,N_4944);
or U5402 (N_5402,N_4636,N_4597);
and U5403 (N_5403,N_4975,N_4428);
nand U5404 (N_5404,N_4633,N_4912);
xnor U5405 (N_5405,N_4802,N_4553);
nor U5406 (N_5406,N_4787,N_4857);
nand U5407 (N_5407,N_4737,N_4913);
xor U5408 (N_5408,N_4481,N_4889);
or U5409 (N_5409,N_4707,N_4934);
nand U5410 (N_5410,N_4451,N_4732);
nor U5411 (N_5411,N_4709,N_4646);
nor U5412 (N_5412,N_4556,N_4398);
nor U5413 (N_5413,N_4816,N_4640);
and U5414 (N_5414,N_4918,N_4944);
or U5415 (N_5415,N_4473,N_4597);
and U5416 (N_5416,N_4402,N_4905);
and U5417 (N_5417,N_4383,N_4658);
and U5418 (N_5418,N_4648,N_4959);
nor U5419 (N_5419,N_4977,N_4610);
nor U5420 (N_5420,N_4953,N_4619);
or U5421 (N_5421,N_4527,N_4720);
nor U5422 (N_5422,N_4603,N_4521);
and U5423 (N_5423,N_4954,N_4738);
nor U5424 (N_5424,N_4627,N_4535);
or U5425 (N_5425,N_4383,N_4890);
nand U5426 (N_5426,N_4488,N_4582);
and U5427 (N_5427,N_4440,N_4773);
or U5428 (N_5428,N_4643,N_4838);
and U5429 (N_5429,N_4376,N_4860);
or U5430 (N_5430,N_4552,N_4604);
or U5431 (N_5431,N_4684,N_4545);
or U5432 (N_5432,N_4869,N_4409);
nand U5433 (N_5433,N_4899,N_4402);
xnor U5434 (N_5434,N_4932,N_4740);
and U5435 (N_5435,N_4718,N_4900);
and U5436 (N_5436,N_4593,N_4803);
nor U5437 (N_5437,N_4568,N_4930);
xor U5438 (N_5438,N_4848,N_4979);
xnor U5439 (N_5439,N_4554,N_4653);
nor U5440 (N_5440,N_4417,N_4952);
or U5441 (N_5441,N_4942,N_4861);
nand U5442 (N_5442,N_4860,N_4961);
xnor U5443 (N_5443,N_4462,N_4515);
nand U5444 (N_5444,N_4868,N_4880);
or U5445 (N_5445,N_4730,N_4629);
or U5446 (N_5446,N_4858,N_4565);
nor U5447 (N_5447,N_4641,N_4919);
xnor U5448 (N_5448,N_4852,N_4839);
or U5449 (N_5449,N_4662,N_4677);
or U5450 (N_5450,N_4952,N_4985);
nor U5451 (N_5451,N_4632,N_4455);
nor U5452 (N_5452,N_4589,N_4974);
and U5453 (N_5453,N_4813,N_4650);
nor U5454 (N_5454,N_4865,N_4442);
or U5455 (N_5455,N_4533,N_4883);
nor U5456 (N_5456,N_4970,N_4875);
and U5457 (N_5457,N_4523,N_4916);
and U5458 (N_5458,N_4587,N_4721);
nor U5459 (N_5459,N_4981,N_4384);
or U5460 (N_5460,N_4643,N_4809);
or U5461 (N_5461,N_4462,N_4680);
and U5462 (N_5462,N_4780,N_4478);
xor U5463 (N_5463,N_4421,N_4621);
xor U5464 (N_5464,N_4480,N_4791);
nor U5465 (N_5465,N_4841,N_4785);
xnor U5466 (N_5466,N_4439,N_4935);
xor U5467 (N_5467,N_4922,N_4561);
or U5468 (N_5468,N_4662,N_4426);
or U5469 (N_5469,N_4660,N_4697);
nor U5470 (N_5470,N_4753,N_4898);
and U5471 (N_5471,N_4555,N_4762);
nand U5472 (N_5472,N_4714,N_4850);
nand U5473 (N_5473,N_4942,N_4822);
nand U5474 (N_5474,N_4959,N_4718);
nand U5475 (N_5475,N_4593,N_4886);
or U5476 (N_5476,N_4969,N_4502);
xor U5477 (N_5477,N_4728,N_4532);
and U5478 (N_5478,N_4539,N_4960);
and U5479 (N_5479,N_4729,N_4968);
nand U5480 (N_5480,N_4413,N_4866);
nor U5481 (N_5481,N_4684,N_4939);
xnor U5482 (N_5482,N_4620,N_4415);
and U5483 (N_5483,N_4427,N_4426);
nand U5484 (N_5484,N_4829,N_4642);
xor U5485 (N_5485,N_4866,N_4895);
xor U5486 (N_5486,N_4654,N_4413);
and U5487 (N_5487,N_4537,N_4946);
nand U5488 (N_5488,N_4823,N_4581);
nor U5489 (N_5489,N_4703,N_4789);
nor U5490 (N_5490,N_4731,N_4661);
xnor U5491 (N_5491,N_4773,N_4937);
or U5492 (N_5492,N_4637,N_4586);
nor U5493 (N_5493,N_4665,N_4730);
and U5494 (N_5494,N_4503,N_4487);
xnor U5495 (N_5495,N_4440,N_4464);
and U5496 (N_5496,N_4755,N_4868);
and U5497 (N_5497,N_4816,N_4755);
xor U5498 (N_5498,N_4486,N_4928);
nand U5499 (N_5499,N_4514,N_4594);
and U5500 (N_5500,N_4519,N_4812);
and U5501 (N_5501,N_4656,N_4651);
or U5502 (N_5502,N_4381,N_4909);
and U5503 (N_5503,N_4915,N_4986);
nor U5504 (N_5504,N_4483,N_4815);
xor U5505 (N_5505,N_4916,N_4825);
and U5506 (N_5506,N_4631,N_4933);
nand U5507 (N_5507,N_4964,N_4514);
or U5508 (N_5508,N_4727,N_4766);
nand U5509 (N_5509,N_4589,N_4742);
nand U5510 (N_5510,N_4862,N_4574);
nand U5511 (N_5511,N_4925,N_4728);
xnor U5512 (N_5512,N_4528,N_4973);
xnor U5513 (N_5513,N_4862,N_4915);
or U5514 (N_5514,N_4709,N_4912);
nor U5515 (N_5515,N_4879,N_4666);
xnor U5516 (N_5516,N_4860,N_4858);
and U5517 (N_5517,N_4794,N_4762);
xnor U5518 (N_5518,N_4949,N_4761);
or U5519 (N_5519,N_4490,N_4939);
or U5520 (N_5520,N_4523,N_4800);
nor U5521 (N_5521,N_4906,N_4872);
or U5522 (N_5522,N_4490,N_4520);
or U5523 (N_5523,N_4975,N_4642);
nor U5524 (N_5524,N_4976,N_4932);
or U5525 (N_5525,N_4899,N_4428);
nor U5526 (N_5526,N_4536,N_4422);
nor U5527 (N_5527,N_4454,N_4410);
or U5528 (N_5528,N_4675,N_4773);
nor U5529 (N_5529,N_4717,N_4687);
and U5530 (N_5530,N_4982,N_4993);
nor U5531 (N_5531,N_4384,N_4885);
nor U5532 (N_5532,N_4703,N_4653);
nor U5533 (N_5533,N_4752,N_4563);
nand U5534 (N_5534,N_4483,N_4873);
nor U5535 (N_5535,N_4686,N_4677);
nor U5536 (N_5536,N_4715,N_4999);
nand U5537 (N_5537,N_4671,N_4719);
and U5538 (N_5538,N_4782,N_4622);
nor U5539 (N_5539,N_4817,N_4772);
nand U5540 (N_5540,N_4457,N_4706);
and U5541 (N_5541,N_4679,N_4654);
nand U5542 (N_5542,N_4479,N_4834);
xor U5543 (N_5543,N_4441,N_4781);
nor U5544 (N_5544,N_4627,N_4552);
and U5545 (N_5545,N_4678,N_4553);
nor U5546 (N_5546,N_4419,N_4792);
or U5547 (N_5547,N_4690,N_4686);
xor U5548 (N_5548,N_4745,N_4690);
nand U5549 (N_5549,N_4389,N_4408);
or U5550 (N_5550,N_4642,N_4836);
or U5551 (N_5551,N_4627,N_4613);
and U5552 (N_5552,N_4567,N_4995);
xor U5553 (N_5553,N_4764,N_4779);
xor U5554 (N_5554,N_4671,N_4805);
and U5555 (N_5555,N_4766,N_4816);
nor U5556 (N_5556,N_4385,N_4763);
nor U5557 (N_5557,N_4403,N_4827);
nand U5558 (N_5558,N_4495,N_4941);
nor U5559 (N_5559,N_4694,N_4912);
nand U5560 (N_5560,N_4497,N_4894);
xor U5561 (N_5561,N_4786,N_4956);
and U5562 (N_5562,N_4673,N_4852);
or U5563 (N_5563,N_4734,N_4569);
xor U5564 (N_5564,N_4693,N_4830);
nand U5565 (N_5565,N_4436,N_4432);
nand U5566 (N_5566,N_4977,N_4976);
nand U5567 (N_5567,N_4515,N_4437);
nand U5568 (N_5568,N_4603,N_4838);
and U5569 (N_5569,N_4527,N_4684);
nand U5570 (N_5570,N_4867,N_4724);
or U5571 (N_5571,N_4837,N_4533);
nor U5572 (N_5572,N_4712,N_4450);
and U5573 (N_5573,N_4779,N_4399);
and U5574 (N_5574,N_4579,N_4866);
nor U5575 (N_5575,N_4853,N_4786);
xnor U5576 (N_5576,N_4463,N_4460);
nor U5577 (N_5577,N_4500,N_4969);
nor U5578 (N_5578,N_4432,N_4924);
or U5579 (N_5579,N_4436,N_4659);
xnor U5580 (N_5580,N_4707,N_4599);
and U5581 (N_5581,N_4403,N_4837);
and U5582 (N_5582,N_4765,N_4563);
nand U5583 (N_5583,N_4456,N_4982);
or U5584 (N_5584,N_4564,N_4478);
and U5585 (N_5585,N_4433,N_4551);
and U5586 (N_5586,N_4959,N_4724);
or U5587 (N_5587,N_4778,N_4869);
nor U5588 (N_5588,N_4814,N_4557);
nand U5589 (N_5589,N_4816,N_4474);
nand U5590 (N_5590,N_4673,N_4472);
and U5591 (N_5591,N_4816,N_4527);
or U5592 (N_5592,N_4624,N_4561);
or U5593 (N_5593,N_4464,N_4693);
nor U5594 (N_5594,N_4681,N_4414);
nand U5595 (N_5595,N_4649,N_4395);
and U5596 (N_5596,N_4555,N_4631);
or U5597 (N_5597,N_4397,N_4743);
nor U5598 (N_5598,N_4942,N_4793);
or U5599 (N_5599,N_4406,N_4725);
or U5600 (N_5600,N_4430,N_4573);
or U5601 (N_5601,N_4840,N_4750);
and U5602 (N_5602,N_4509,N_4697);
nand U5603 (N_5603,N_4734,N_4962);
or U5604 (N_5604,N_4537,N_4906);
and U5605 (N_5605,N_4723,N_4491);
nor U5606 (N_5606,N_4879,N_4890);
nand U5607 (N_5607,N_4734,N_4807);
nor U5608 (N_5608,N_4866,N_4709);
nand U5609 (N_5609,N_4964,N_4795);
or U5610 (N_5610,N_4726,N_4951);
or U5611 (N_5611,N_4679,N_4665);
nand U5612 (N_5612,N_4964,N_4892);
xor U5613 (N_5613,N_4598,N_4897);
nand U5614 (N_5614,N_4637,N_4400);
nor U5615 (N_5615,N_4383,N_4932);
nand U5616 (N_5616,N_4505,N_4601);
or U5617 (N_5617,N_4806,N_4998);
nand U5618 (N_5618,N_4429,N_4391);
or U5619 (N_5619,N_4465,N_4611);
and U5620 (N_5620,N_4779,N_4927);
and U5621 (N_5621,N_4548,N_4479);
nand U5622 (N_5622,N_4807,N_4849);
or U5623 (N_5623,N_4590,N_4950);
or U5624 (N_5624,N_4880,N_4390);
xnor U5625 (N_5625,N_5016,N_5056);
nand U5626 (N_5626,N_5276,N_5359);
nand U5627 (N_5627,N_5408,N_5450);
and U5628 (N_5628,N_5343,N_5103);
or U5629 (N_5629,N_5458,N_5085);
nor U5630 (N_5630,N_5368,N_5165);
nor U5631 (N_5631,N_5378,N_5415);
nor U5632 (N_5632,N_5088,N_5568);
nand U5633 (N_5633,N_5502,N_5204);
nor U5634 (N_5634,N_5000,N_5309);
or U5635 (N_5635,N_5434,N_5025);
nor U5636 (N_5636,N_5589,N_5208);
nand U5637 (N_5637,N_5100,N_5459);
or U5638 (N_5638,N_5023,N_5325);
and U5639 (N_5639,N_5521,N_5440);
and U5640 (N_5640,N_5512,N_5477);
or U5641 (N_5641,N_5139,N_5209);
or U5642 (N_5642,N_5247,N_5092);
and U5643 (N_5643,N_5038,N_5246);
xnor U5644 (N_5644,N_5101,N_5072);
nand U5645 (N_5645,N_5363,N_5607);
nand U5646 (N_5646,N_5515,N_5431);
or U5647 (N_5647,N_5281,N_5506);
and U5648 (N_5648,N_5347,N_5429);
or U5649 (N_5649,N_5416,N_5127);
xor U5650 (N_5650,N_5511,N_5467);
or U5651 (N_5651,N_5211,N_5134);
or U5652 (N_5652,N_5575,N_5004);
nand U5653 (N_5653,N_5465,N_5540);
nor U5654 (N_5654,N_5417,N_5572);
or U5655 (N_5655,N_5194,N_5484);
and U5656 (N_5656,N_5037,N_5482);
or U5657 (N_5657,N_5151,N_5448);
nor U5658 (N_5658,N_5195,N_5220);
nand U5659 (N_5659,N_5530,N_5495);
xor U5660 (N_5660,N_5449,N_5093);
nand U5661 (N_5661,N_5558,N_5140);
or U5662 (N_5662,N_5393,N_5435);
xnor U5663 (N_5663,N_5132,N_5469);
or U5664 (N_5664,N_5376,N_5602);
and U5665 (N_5665,N_5517,N_5245);
and U5666 (N_5666,N_5544,N_5051);
nand U5667 (N_5667,N_5239,N_5345);
xor U5668 (N_5668,N_5294,N_5096);
xnor U5669 (N_5669,N_5503,N_5609);
and U5670 (N_5670,N_5562,N_5284);
or U5671 (N_5671,N_5375,N_5003);
nand U5672 (N_5672,N_5362,N_5041);
nand U5673 (N_5673,N_5260,N_5184);
or U5674 (N_5674,N_5039,N_5066);
nor U5675 (N_5675,N_5462,N_5222);
and U5676 (N_5676,N_5249,N_5201);
or U5677 (N_5677,N_5352,N_5547);
xor U5678 (N_5678,N_5070,N_5313);
nand U5679 (N_5679,N_5310,N_5028);
nand U5680 (N_5680,N_5116,N_5399);
nor U5681 (N_5681,N_5040,N_5586);
and U5682 (N_5682,N_5299,N_5414);
and U5683 (N_5683,N_5120,N_5427);
or U5684 (N_5684,N_5109,N_5391);
xnor U5685 (N_5685,N_5419,N_5373);
and U5686 (N_5686,N_5206,N_5150);
nand U5687 (N_5687,N_5269,N_5090);
nor U5688 (N_5688,N_5240,N_5546);
nor U5689 (N_5689,N_5557,N_5332);
or U5690 (N_5690,N_5102,N_5580);
xor U5691 (N_5691,N_5185,N_5318);
or U5692 (N_5692,N_5122,N_5069);
or U5693 (N_5693,N_5125,N_5560);
and U5694 (N_5694,N_5623,N_5168);
xnor U5695 (N_5695,N_5190,N_5279);
or U5696 (N_5696,N_5339,N_5006);
nor U5697 (N_5697,N_5288,N_5036);
or U5698 (N_5698,N_5254,N_5573);
nor U5699 (N_5699,N_5175,N_5329);
nand U5700 (N_5700,N_5397,N_5364);
nor U5701 (N_5701,N_5272,N_5112);
or U5702 (N_5702,N_5044,N_5019);
and U5703 (N_5703,N_5026,N_5191);
xnor U5704 (N_5704,N_5271,N_5403);
nand U5705 (N_5705,N_5218,N_5149);
or U5706 (N_5706,N_5119,N_5105);
or U5707 (N_5707,N_5014,N_5320);
or U5708 (N_5708,N_5154,N_5554);
and U5709 (N_5709,N_5323,N_5241);
and U5710 (N_5710,N_5307,N_5242);
nand U5711 (N_5711,N_5361,N_5505);
xor U5712 (N_5712,N_5387,N_5395);
nand U5713 (N_5713,N_5174,N_5483);
or U5714 (N_5714,N_5567,N_5366);
nor U5715 (N_5715,N_5214,N_5486);
and U5716 (N_5716,N_5328,N_5301);
xnor U5717 (N_5717,N_5166,N_5113);
or U5718 (N_5718,N_5596,N_5570);
nor U5719 (N_5719,N_5489,N_5581);
nand U5720 (N_5720,N_5330,N_5182);
and U5721 (N_5721,N_5423,N_5615);
nor U5722 (N_5722,N_5461,N_5509);
nor U5723 (N_5723,N_5578,N_5020);
xor U5724 (N_5724,N_5525,N_5262);
xnor U5725 (N_5725,N_5009,N_5107);
xnor U5726 (N_5726,N_5608,N_5087);
or U5727 (N_5727,N_5147,N_5532);
or U5728 (N_5728,N_5582,N_5253);
nand U5729 (N_5729,N_5292,N_5111);
xor U5730 (N_5730,N_5453,N_5454);
and U5731 (N_5731,N_5543,N_5338);
nor U5732 (N_5732,N_5114,N_5372);
xor U5733 (N_5733,N_5264,N_5229);
nand U5734 (N_5734,N_5073,N_5142);
nand U5735 (N_5735,N_5110,N_5189);
xnor U5736 (N_5736,N_5106,N_5232);
or U5737 (N_5737,N_5157,N_5621);
xnor U5738 (N_5738,N_5564,N_5042);
nor U5739 (N_5739,N_5425,N_5277);
and U5740 (N_5740,N_5289,N_5050);
nand U5741 (N_5741,N_5563,N_5624);
and U5742 (N_5742,N_5534,N_5349);
or U5743 (N_5743,N_5612,N_5494);
xor U5744 (N_5744,N_5555,N_5183);
nor U5745 (N_5745,N_5351,N_5048);
and U5746 (N_5746,N_5296,N_5407);
nand U5747 (N_5747,N_5333,N_5371);
or U5748 (N_5748,N_5398,N_5198);
nand U5749 (N_5749,N_5322,N_5237);
and U5750 (N_5750,N_5479,N_5238);
or U5751 (N_5751,N_5455,N_5584);
nor U5752 (N_5752,N_5305,N_5381);
xnor U5753 (N_5753,N_5585,N_5457);
or U5754 (N_5754,N_5045,N_5569);
nand U5755 (N_5755,N_5619,N_5541);
or U5756 (N_5756,N_5452,N_5614);
nor U5757 (N_5757,N_5031,N_5071);
xnor U5758 (N_5758,N_5551,N_5062);
and U5759 (N_5759,N_5146,N_5021);
and U5760 (N_5760,N_5576,N_5143);
xor U5761 (N_5761,N_5059,N_5410);
nor U5762 (N_5762,N_5057,N_5148);
or U5763 (N_5763,N_5034,N_5430);
xor U5764 (N_5764,N_5266,N_5601);
or U5765 (N_5765,N_5524,N_5317);
and U5766 (N_5766,N_5196,N_5136);
nor U5767 (N_5767,N_5225,N_5497);
xnor U5768 (N_5768,N_5357,N_5163);
nor U5769 (N_5769,N_5426,N_5518);
and U5770 (N_5770,N_5538,N_5137);
and U5771 (N_5771,N_5478,N_5268);
or U5772 (N_5772,N_5155,N_5013);
nor U5773 (N_5773,N_5243,N_5011);
nor U5774 (N_5774,N_5265,N_5123);
xor U5775 (N_5775,N_5049,N_5267);
or U5776 (N_5776,N_5421,N_5303);
and U5777 (N_5777,N_5565,N_5300);
nand U5778 (N_5778,N_5500,N_5287);
nor U5779 (N_5779,N_5533,N_5445);
nor U5780 (N_5780,N_5583,N_5474);
nand U5781 (N_5781,N_5015,N_5598);
xnor U5782 (N_5782,N_5354,N_5248);
nor U5783 (N_5783,N_5600,N_5064);
nand U5784 (N_5784,N_5144,N_5231);
and U5785 (N_5785,N_5358,N_5290);
nand U5786 (N_5786,N_5176,N_5178);
or U5787 (N_5787,N_5438,N_5161);
and U5788 (N_5788,N_5224,N_5274);
xnor U5789 (N_5789,N_5389,N_5033);
or U5790 (N_5790,N_5523,N_5162);
xor U5791 (N_5791,N_5418,N_5032);
or U5792 (N_5792,N_5388,N_5047);
xor U5793 (N_5793,N_5250,N_5251);
nor U5794 (N_5794,N_5367,N_5542);
nand U5795 (N_5795,N_5193,N_5436);
nor U5796 (N_5796,N_5210,N_5086);
xor U5797 (N_5797,N_5216,N_5094);
nand U5798 (N_5798,N_5587,N_5304);
nor U5799 (N_5799,N_5063,N_5017);
nand U5800 (N_5800,N_5377,N_5291);
and U5801 (N_5801,N_5188,N_5475);
xnor U5802 (N_5802,N_5441,N_5259);
nor U5803 (N_5803,N_5537,N_5622);
xor U5804 (N_5804,N_5030,N_5295);
and U5805 (N_5805,N_5091,N_5571);
nor U5806 (N_5806,N_5539,N_5470);
and U5807 (N_5807,N_5215,N_5255);
xnor U5808 (N_5808,N_5058,N_5553);
nor U5809 (N_5809,N_5485,N_5012);
nand U5810 (N_5810,N_5024,N_5256);
xor U5811 (N_5811,N_5171,N_5187);
xor U5812 (N_5812,N_5007,N_5331);
nor U5813 (N_5813,N_5529,N_5404);
nor U5814 (N_5814,N_5592,N_5080);
nand U5815 (N_5815,N_5074,N_5337);
and U5816 (N_5816,N_5460,N_5067);
or U5817 (N_5817,N_5442,N_5535);
nand U5818 (N_5818,N_5411,N_5052);
xnor U5819 (N_5819,N_5356,N_5008);
nor U5820 (N_5820,N_5492,N_5095);
or U5821 (N_5821,N_5129,N_5374);
xnor U5822 (N_5822,N_5488,N_5599);
xnor U5823 (N_5823,N_5212,N_5043);
and U5824 (N_5824,N_5590,N_5531);
nor U5825 (N_5825,N_5466,N_5481);
and U5826 (N_5826,N_5022,N_5227);
nand U5827 (N_5827,N_5468,N_5130);
and U5828 (N_5828,N_5406,N_5396);
and U5829 (N_5829,N_5158,N_5226);
xor U5830 (N_5830,N_5593,N_5412);
and U5831 (N_5831,N_5350,N_5117);
nand U5832 (N_5832,N_5611,N_5223);
nor U5833 (N_5833,N_5556,N_5451);
and U5834 (N_5834,N_5499,N_5496);
or U5835 (N_5835,N_5464,N_5258);
xnor U5836 (N_5836,N_5420,N_5360);
or U5837 (N_5837,N_5319,N_5604);
xor U5838 (N_5838,N_5054,N_5365);
and U5839 (N_5839,N_5081,N_5579);
nand U5840 (N_5840,N_5205,N_5405);
nand U5841 (N_5841,N_5446,N_5536);
and U5842 (N_5842,N_5186,N_5340);
nand U5843 (N_5843,N_5380,N_5180);
xor U5844 (N_5844,N_5386,N_5079);
and U5845 (N_5845,N_5055,N_5392);
and U5846 (N_5846,N_5574,N_5172);
or U5847 (N_5847,N_5336,N_5083);
xor U5848 (N_5848,N_5257,N_5527);
nand U5849 (N_5849,N_5471,N_5552);
nand U5850 (N_5850,N_5278,N_5275);
nor U5851 (N_5851,N_5545,N_5202);
and U5852 (N_5852,N_5520,N_5487);
nor U5853 (N_5853,N_5522,N_5402);
and U5854 (N_5854,N_5594,N_5618);
nand U5855 (N_5855,N_5385,N_5498);
nor U5856 (N_5856,N_5181,N_5472);
nand U5857 (N_5857,N_5595,N_5480);
or U5858 (N_5858,N_5312,N_5315);
and U5859 (N_5859,N_5233,N_5409);
and U5860 (N_5860,N_5270,N_5613);
xor U5861 (N_5861,N_5610,N_5507);
or U5862 (N_5862,N_5170,N_5010);
xor U5863 (N_5863,N_5179,N_5566);
or U5864 (N_5864,N_5065,N_5353);
and U5865 (N_5865,N_5316,N_5514);
or U5866 (N_5866,N_5207,N_5124);
or U5867 (N_5867,N_5035,N_5422);
nor U5868 (N_5868,N_5327,N_5559);
nor U5869 (N_5869,N_5005,N_5456);
xnor U5870 (N_5870,N_5550,N_5128);
nand U5871 (N_5871,N_5235,N_5145);
or U5872 (N_5872,N_5463,N_5027);
nor U5873 (N_5873,N_5261,N_5342);
and U5874 (N_5874,N_5597,N_5297);
xnor U5875 (N_5875,N_5561,N_5493);
or U5876 (N_5876,N_5219,N_5159);
nor U5877 (N_5877,N_5306,N_5401);
nand U5878 (N_5878,N_5283,N_5141);
or U5879 (N_5879,N_5603,N_5591);
nor U5880 (N_5880,N_5280,N_5549);
nor U5881 (N_5881,N_5302,N_5002);
and U5882 (N_5882,N_5138,N_5428);
or U5883 (N_5883,N_5199,N_5606);
nor U5884 (N_5884,N_5348,N_5516);
xor U5885 (N_5885,N_5588,N_5234);
nor U5886 (N_5886,N_5617,N_5053);
nand U5887 (N_5887,N_5383,N_5286);
nor U5888 (N_5888,N_5321,N_5164);
and U5889 (N_5889,N_5018,N_5504);
or U5890 (N_5890,N_5616,N_5273);
or U5891 (N_5891,N_5473,N_5156);
nand U5892 (N_5892,N_5135,N_5513);
and U5893 (N_5893,N_5217,N_5098);
nand U5894 (N_5894,N_5326,N_5282);
and U5895 (N_5895,N_5252,N_5061);
nand U5896 (N_5896,N_5221,N_5424);
nor U5897 (N_5897,N_5153,N_5335);
nand U5898 (N_5898,N_5001,N_5519);
or U5899 (N_5899,N_5447,N_5528);
xor U5900 (N_5900,N_5308,N_5177);
and U5901 (N_5901,N_5060,N_5548);
xor U5902 (N_5902,N_5046,N_5476);
nor U5903 (N_5903,N_5501,N_5230);
nor U5904 (N_5904,N_5334,N_5344);
and U5905 (N_5905,N_5213,N_5413);
xnor U5906 (N_5906,N_5169,N_5443);
xnor U5907 (N_5907,N_5394,N_5369);
or U5908 (N_5908,N_5075,N_5076);
xor U5909 (N_5909,N_5197,N_5167);
or U5910 (N_5910,N_5311,N_5131);
nand U5911 (N_5911,N_5605,N_5510);
xor U5912 (N_5912,N_5384,N_5341);
nor U5913 (N_5913,N_5444,N_5078);
nand U5914 (N_5914,N_5084,N_5160);
xnor U5915 (N_5915,N_5491,N_5432);
nand U5916 (N_5916,N_5200,N_5508);
nand U5917 (N_5917,N_5192,N_5433);
or U5918 (N_5918,N_5029,N_5314);
and U5919 (N_5919,N_5173,N_5382);
nor U5920 (N_5920,N_5121,N_5379);
xnor U5921 (N_5921,N_5104,N_5133);
xor U5922 (N_5922,N_5346,N_5244);
or U5923 (N_5923,N_5355,N_5228);
nand U5924 (N_5924,N_5370,N_5068);
nand U5925 (N_5925,N_5400,N_5115);
and U5926 (N_5926,N_5298,N_5077);
xnor U5927 (N_5927,N_5437,N_5118);
nand U5928 (N_5928,N_5293,N_5108);
and U5929 (N_5929,N_5490,N_5089);
nand U5930 (N_5930,N_5097,N_5285);
and U5931 (N_5931,N_5324,N_5620);
nor U5932 (N_5932,N_5126,N_5439);
nor U5933 (N_5933,N_5526,N_5236);
xnor U5934 (N_5934,N_5577,N_5099);
or U5935 (N_5935,N_5082,N_5390);
or U5936 (N_5936,N_5263,N_5152);
xor U5937 (N_5937,N_5203,N_5558);
xnor U5938 (N_5938,N_5485,N_5253);
nand U5939 (N_5939,N_5318,N_5506);
xor U5940 (N_5940,N_5417,N_5211);
nand U5941 (N_5941,N_5399,N_5553);
nand U5942 (N_5942,N_5043,N_5591);
nor U5943 (N_5943,N_5108,N_5259);
nor U5944 (N_5944,N_5508,N_5073);
nand U5945 (N_5945,N_5559,N_5348);
and U5946 (N_5946,N_5499,N_5163);
and U5947 (N_5947,N_5487,N_5342);
and U5948 (N_5948,N_5572,N_5544);
nand U5949 (N_5949,N_5311,N_5340);
nand U5950 (N_5950,N_5585,N_5549);
nand U5951 (N_5951,N_5263,N_5019);
and U5952 (N_5952,N_5561,N_5349);
xnor U5953 (N_5953,N_5172,N_5307);
nor U5954 (N_5954,N_5161,N_5064);
nor U5955 (N_5955,N_5304,N_5316);
xor U5956 (N_5956,N_5400,N_5363);
and U5957 (N_5957,N_5611,N_5030);
or U5958 (N_5958,N_5046,N_5246);
or U5959 (N_5959,N_5030,N_5209);
nand U5960 (N_5960,N_5158,N_5243);
nand U5961 (N_5961,N_5153,N_5308);
nor U5962 (N_5962,N_5420,N_5530);
nand U5963 (N_5963,N_5589,N_5405);
nand U5964 (N_5964,N_5464,N_5167);
and U5965 (N_5965,N_5065,N_5603);
nand U5966 (N_5966,N_5130,N_5255);
and U5967 (N_5967,N_5239,N_5604);
nand U5968 (N_5968,N_5497,N_5146);
nand U5969 (N_5969,N_5127,N_5564);
nand U5970 (N_5970,N_5116,N_5165);
xnor U5971 (N_5971,N_5281,N_5370);
nor U5972 (N_5972,N_5497,N_5569);
and U5973 (N_5973,N_5583,N_5529);
xnor U5974 (N_5974,N_5008,N_5222);
and U5975 (N_5975,N_5300,N_5550);
nor U5976 (N_5976,N_5395,N_5457);
or U5977 (N_5977,N_5082,N_5484);
nand U5978 (N_5978,N_5033,N_5003);
xnor U5979 (N_5979,N_5249,N_5054);
or U5980 (N_5980,N_5307,N_5186);
or U5981 (N_5981,N_5530,N_5423);
xnor U5982 (N_5982,N_5293,N_5232);
nand U5983 (N_5983,N_5176,N_5350);
and U5984 (N_5984,N_5401,N_5201);
nor U5985 (N_5985,N_5328,N_5109);
and U5986 (N_5986,N_5025,N_5404);
or U5987 (N_5987,N_5026,N_5185);
nor U5988 (N_5988,N_5117,N_5260);
or U5989 (N_5989,N_5225,N_5410);
or U5990 (N_5990,N_5035,N_5330);
xor U5991 (N_5991,N_5002,N_5393);
nor U5992 (N_5992,N_5272,N_5085);
xor U5993 (N_5993,N_5272,N_5309);
xor U5994 (N_5994,N_5143,N_5365);
or U5995 (N_5995,N_5135,N_5493);
nor U5996 (N_5996,N_5353,N_5426);
nor U5997 (N_5997,N_5468,N_5049);
and U5998 (N_5998,N_5163,N_5455);
or U5999 (N_5999,N_5448,N_5223);
nand U6000 (N_6000,N_5189,N_5494);
xnor U6001 (N_6001,N_5470,N_5521);
xor U6002 (N_6002,N_5555,N_5245);
xor U6003 (N_6003,N_5402,N_5241);
and U6004 (N_6004,N_5039,N_5185);
or U6005 (N_6005,N_5291,N_5351);
and U6006 (N_6006,N_5140,N_5472);
and U6007 (N_6007,N_5153,N_5045);
or U6008 (N_6008,N_5050,N_5013);
nand U6009 (N_6009,N_5266,N_5147);
nor U6010 (N_6010,N_5302,N_5429);
nand U6011 (N_6011,N_5369,N_5461);
xor U6012 (N_6012,N_5511,N_5125);
or U6013 (N_6013,N_5494,N_5153);
or U6014 (N_6014,N_5185,N_5571);
nand U6015 (N_6015,N_5395,N_5604);
xnor U6016 (N_6016,N_5446,N_5257);
nand U6017 (N_6017,N_5528,N_5042);
xnor U6018 (N_6018,N_5422,N_5090);
and U6019 (N_6019,N_5070,N_5188);
nand U6020 (N_6020,N_5213,N_5478);
nor U6021 (N_6021,N_5041,N_5333);
or U6022 (N_6022,N_5554,N_5517);
xnor U6023 (N_6023,N_5381,N_5184);
xnor U6024 (N_6024,N_5441,N_5498);
nor U6025 (N_6025,N_5544,N_5497);
nand U6026 (N_6026,N_5194,N_5374);
xnor U6027 (N_6027,N_5423,N_5178);
and U6028 (N_6028,N_5290,N_5182);
or U6029 (N_6029,N_5580,N_5437);
or U6030 (N_6030,N_5121,N_5294);
and U6031 (N_6031,N_5222,N_5571);
xor U6032 (N_6032,N_5497,N_5292);
nand U6033 (N_6033,N_5155,N_5056);
xor U6034 (N_6034,N_5239,N_5331);
xor U6035 (N_6035,N_5511,N_5403);
or U6036 (N_6036,N_5589,N_5118);
xor U6037 (N_6037,N_5606,N_5175);
or U6038 (N_6038,N_5082,N_5414);
or U6039 (N_6039,N_5307,N_5541);
and U6040 (N_6040,N_5348,N_5142);
xor U6041 (N_6041,N_5051,N_5217);
nor U6042 (N_6042,N_5120,N_5124);
and U6043 (N_6043,N_5448,N_5515);
nor U6044 (N_6044,N_5002,N_5080);
xor U6045 (N_6045,N_5070,N_5068);
nand U6046 (N_6046,N_5380,N_5601);
nor U6047 (N_6047,N_5235,N_5053);
nand U6048 (N_6048,N_5422,N_5078);
xor U6049 (N_6049,N_5481,N_5242);
and U6050 (N_6050,N_5139,N_5008);
or U6051 (N_6051,N_5352,N_5157);
or U6052 (N_6052,N_5424,N_5554);
or U6053 (N_6053,N_5466,N_5293);
nand U6054 (N_6054,N_5160,N_5554);
nor U6055 (N_6055,N_5087,N_5238);
nor U6056 (N_6056,N_5002,N_5597);
xor U6057 (N_6057,N_5026,N_5508);
and U6058 (N_6058,N_5400,N_5125);
and U6059 (N_6059,N_5454,N_5518);
or U6060 (N_6060,N_5219,N_5324);
and U6061 (N_6061,N_5232,N_5534);
nor U6062 (N_6062,N_5473,N_5386);
nand U6063 (N_6063,N_5360,N_5461);
nor U6064 (N_6064,N_5523,N_5267);
xor U6065 (N_6065,N_5516,N_5415);
or U6066 (N_6066,N_5181,N_5493);
and U6067 (N_6067,N_5374,N_5277);
xnor U6068 (N_6068,N_5209,N_5536);
nand U6069 (N_6069,N_5472,N_5231);
nor U6070 (N_6070,N_5282,N_5435);
nand U6071 (N_6071,N_5046,N_5329);
nor U6072 (N_6072,N_5280,N_5537);
nand U6073 (N_6073,N_5227,N_5362);
and U6074 (N_6074,N_5250,N_5293);
and U6075 (N_6075,N_5448,N_5388);
xor U6076 (N_6076,N_5480,N_5579);
or U6077 (N_6077,N_5415,N_5032);
nor U6078 (N_6078,N_5275,N_5345);
nor U6079 (N_6079,N_5433,N_5237);
nor U6080 (N_6080,N_5068,N_5537);
nor U6081 (N_6081,N_5045,N_5080);
and U6082 (N_6082,N_5370,N_5064);
xnor U6083 (N_6083,N_5241,N_5005);
nor U6084 (N_6084,N_5166,N_5583);
xor U6085 (N_6085,N_5272,N_5585);
nand U6086 (N_6086,N_5418,N_5269);
nand U6087 (N_6087,N_5199,N_5605);
xor U6088 (N_6088,N_5517,N_5010);
or U6089 (N_6089,N_5341,N_5126);
or U6090 (N_6090,N_5441,N_5604);
xnor U6091 (N_6091,N_5296,N_5490);
nand U6092 (N_6092,N_5567,N_5010);
xnor U6093 (N_6093,N_5405,N_5069);
xor U6094 (N_6094,N_5029,N_5606);
xnor U6095 (N_6095,N_5093,N_5013);
and U6096 (N_6096,N_5321,N_5134);
nor U6097 (N_6097,N_5176,N_5016);
and U6098 (N_6098,N_5194,N_5271);
and U6099 (N_6099,N_5045,N_5467);
nor U6100 (N_6100,N_5271,N_5099);
nor U6101 (N_6101,N_5304,N_5615);
nand U6102 (N_6102,N_5578,N_5307);
xnor U6103 (N_6103,N_5489,N_5350);
and U6104 (N_6104,N_5388,N_5242);
xor U6105 (N_6105,N_5009,N_5412);
or U6106 (N_6106,N_5430,N_5343);
nor U6107 (N_6107,N_5380,N_5478);
xnor U6108 (N_6108,N_5271,N_5279);
or U6109 (N_6109,N_5448,N_5031);
and U6110 (N_6110,N_5624,N_5171);
and U6111 (N_6111,N_5310,N_5015);
nor U6112 (N_6112,N_5409,N_5038);
or U6113 (N_6113,N_5304,N_5170);
nand U6114 (N_6114,N_5090,N_5223);
nand U6115 (N_6115,N_5082,N_5106);
nor U6116 (N_6116,N_5430,N_5365);
nand U6117 (N_6117,N_5278,N_5377);
nor U6118 (N_6118,N_5034,N_5593);
or U6119 (N_6119,N_5600,N_5167);
and U6120 (N_6120,N_5413,N_5589);
nand U6121 (N_6121,N_5127,N_5484);
or U6122 (N_6122,N_5351,N_5608);
nand U6123 (N_6123,N_5025,N_5135);
xor U6124 (N_6124,N_5092,N_5136);
and U6125 (N_6125,N_5195,N_5455);
nand U6126 (N_6126,N_5366,N_5560);
and U6127 (N_6127,N_5223,N_5089);
nor U6128 (N_6128,N_5373,N_5099);
xor U6129 (N_6129,N_5620,N_5167);
nor U6130 (N_6130,N_5508,N_5583);
nor U6131 (N_6131,N_5584,N_5112);
nand U6132 (N_6132,N_5367,N_5124);
xnor U6133 (N_6133,N_5191,N_5530);
xor U6134 (N_6134,N_5101,N_5541);
or U6135 (N_6135,N_5306,N_5390);
xnor U6136 (N_6136,N_5288,N_5392);
or U6137 (N_6137,N_5538,N_5056);
and U6138 (N_6138,N_5022,N_5318);
nor U6139 (N_6139,N_5037,N_5071);
xor U6140 (N_6140,N_5624,N_5013);
and U6141 (N_6141,N_5085,N_5561);
nand U6142 (N_6142,N_5557,N_5499);
and U6143 (N_6143,N_5135,N_5440);
nand U6144 (N_6144,N_5089,N_5238);
and U6145 (N_6145,N_5608,N_5494);
or U6146 (N_6146,N_5161,N_5394);
and U6147 (N_6147,N_5259,N_5042);
xor U6148 (N_6148,N_5193,N_5351);
nand U6149 (N_6149,N_5333,N_5036);
or U6150 (N_6150,N_5128,N_5171);
xor U6151 (N_6151,N_5465,N_5284);
nor U6152 (N_6152,N_5389,N_5056);
xor U6153 (N_6153,N_5161,N_5005);
nand U6154 (N_6154,N_5589,N_5314);
or U6155 (N_6155,N_5028,N_5149);
nor U6156 (N_6156,N_5108,N_5526);
nand U6157 (N_6157,N_5435,N_5568);
xnor U6158 (N_6158,N_5068,N_5612);
nand U6159 (N_6159,N_5604,N_5536);
or U6160 (N_6160,N_5459,N_5586);
nand U6161 (N_6161,N_5387,N_5186);
or U6162 (N_6162,N_5215,N_5247);
or U6163 (N_6163,N_5427,N_5148);
nor U6164 (N_6164,N_5193,N_5186);
nor U6165 (N_6165,N_5148,N_5478);
or U6166 (N_6166,N_5450,N_5079);
and U6167 (N_6167,N_5258,N_5220);
nand U6168 (N_6168,N_5093,N_5525);
or U6169 (N_6169,N_5243,N_5111);
nor U6170 (N_6170,N_5399,N_5277);
nand U6171 (N_6171,N_5361,N_5457);
nor U6172 (N_6172,N_5074,N_5183);
nor U6173 (N_6173,N_5347,N_5339);
nor U6174 (N_6174,N_5307,N_5606);
or U6175 (N_6175,N_5413,N_5190);
nand U6176 (N_6176,N_5094,N_5387);
or U6177 (N_6177,N_5058,N_5422);
xor U6178 (N_6178,N_5155,N_5257);
nor U6179 (N_6179,N_5284,N_5174);
nand U6180 (N_6180,N_5472,N_5428);
or U6181 (N_6181,N_5111,N_5540);
or U6182 (N_6182,N_5225,N_5298);
and U6183 (N_6183,N_5575,N_5510);
nand U6184 (N_6184,N_5010,N_5571);
and U6185 (N_6185,N_5549,N_5255);
xnor U6186 (N_6186,N_5574,N_5003);
and U6187 (N_6187,N_5062,N_5348);
or U6188 (N_6188,N_5602,N_5473);
and U6189 (N_6189,N_5034,N_5318);
xnor U6190 (N_6190,N_5464,N_5239);
nand U6191 (N_6191,N_5022,N_5475);
or U6192 (N_6192,N_5414,N_5062);
and U6193 (N_6193,N_5436,N_5004);
nor U6194 (N_6194,N_5290,N_5000);
or U6195 (N_6195,N_5497,N_5558);
or U6196 (N_6196,N_5375,N_5229);
xor U6197 (N_6197,N_5172,N_5570);
or U6198 (N_6198,N_5590,N_5272);
nor U6199 (N_6199,N_5215,N_5035);
and U6200 (N_6200,N_5448,N_5356);
nor U6201 (N_6201,N_5107,N_5470);
nand U6202 (N_6202,N_5002,N_5258);
or U6203 (N_6203,N_5389,N_5582);
and U6204 (N_6204,N_5077,N_5201);
and U6205 (N_6205,N_5166,N_5050);
nand U6206 (N_6206,N_5156,N_5390);
and U6207 (N_6207,N_5229,N_5052);
xnor U6208 (N_6208,N_5138,N_5351);
xnor U6209 (N_6209,N_5543,N_5036);
or U6210 (N_6210,N_5115,N_5168);
xnor U6211 (N_6211,N_5110,N_5087);
nor U6212 (N_6212,N_5113,N_5455);
and U6213 (N_6213,N_5294,N_5017);
nand U6214 (N_6214,N_5252,N_5402);
nand U6215 (N_6215,N_5159,N_5460);
and U6216 (N_6216,N_5474,N_5436);
nand U6217 (N_6217,N_5016,N_5009);
and U6218 (N_6218,N_5110,N_5185);
or U6219 (N_6219,N_5038,N_5606);
nand U6220 (N_6220,N_5141,N_5406);
or U6221 (N_6221,N_5387,N_5065);
xor U6222 (N_6222,N_5624,N_5272);
nor U6223 (N_6223,N_5523,N_5618);
and U6224 (N_6224,N_5588,N_5433);
xnor U6225 (N_6225,N_5193,N_5467);
or U6226 (N_6226,N_5112,N_5120);
or U6227 (N_6227,N_5567,N_5012);
nor U6228 (N_6228,N_5345,N_5556);
nor U6229 (N_6229,N_5444,N_5042);
or U6230 (N_6230,N_5478,N_5329);
or U6231 (N_6231,N_5346,N_5023);
xor U6232 (N_6232,N_5007,N_5218);
xnor U6233 (N_6233,N_5168,N_5245);
nand U6234 (N_6234,N_5605,N_5594);
and U6235 (N_6235,N_5422,N_5485);
nand U6236 (N_6236,N_5405,N_5116);
xnor U6237 (N_6237,N_5104,N_5556);
and U6238 (N_6238,N_5123,N_5348);
nand U6239 (N_6239,N_5117,N_5409);
and U6240 (N_6240,N_5441,N_5284);
xor U6241 (N_6241,N_5444,N_5127);
nand U6242 (N_6242,N_5562,N_5157);
nand U6243 (N_6243,N_5508,N_5260);
nor U6244 (N_6244,N_5264,N_5327);
xnor U6245 (N_6245,N_5145,N_5147);
and U6246 (N_6246,N_5478,N_5585);
xor U6247 (N_6247,N_5575,N_5476);
and U6248 (N_6248,N_5115,N_5104);
and U6249 (N_6249,N_5258,N_5589);
or U6250 (N_6250,N_6070,N_5763);
xor U6251 (N_6251,N_5738,N_5630);
or U6252 (N_6252,N_5917,N_5821);
and U6253 (N_6253,N_6158,N_5842);
nor U6254 (N_6254,N_5829,N_5818);
and U6255 (N_6255,N_6025,N_6105);
nor U6256 (N_6256,N_5911,N_6142);
and U6257 (N_6257,N_6176,N_5946);
nand U6258 (N_6258,N_5708,N_6093);
nand U6259 (N_6259,N_5741,N_6069);
and U6260 (N_6260,N_5972,N_5921);
nand U6261 (N_6261,N_5985,N_5631);
or U6262 (N_6262,N_5843,N_6004);
or U6263 (N_6263,N_6067,N_5922);
nand U6264 (N_6264,N_5745,N_6084);
nor U6265 (N_6265,N_5787,N_5670);
nand U6266 (N_6266,N_5797,N_6037);
or U6267 (N_6267,N_6124,N_5712);
or U6268 (N_6268,N_5800,N_6042);
or U6269 (N_6269,N_5662,N_5848);
nor U6270 (N_6270,N_5694,N_6117);
xor U6271 (N_6271,N_5875,N_5638);
nand U6272 (N_6272,N_5807,N_5908);
or U6273 (N_6273,N_6022,N_6178);
and U6274 (N_6274,N_5919,N_5751);
nor U6275 (N_6275,N_5863,N_5758);
xnor U6276 (N_6276,N_6190,N_5831);
nand U6277 (N_6277,N_5846,N_5854);
and U6278 (N_6278,N_6170,N_6019);
and U6279 (N_6279,N_5715,N_5663);
and U6280 (N_6280,N_6165,N_5968);
and U6281 (N_6281,N_6104,N_6131);
or U6282 (N_6282,N_5722,N_5929);
and U6283 (N_6283,N_6210,N_5647);
nor U6284 (N_6284,N_6232,N_5872);
nor U6285 (N_6285,N_5732,N_5949);
xnor U6286 (N_6286,N_5739,N_5635);
xnor U6287 (N_6287,N_6059,N_6229);
or U6288 (N_6288,N_6226,N_6066);
or U6289 (N_6289,N_6000,N_6096);
and U6290 (N_6290,N_5685,N_5626);
and U6291 (N_6291,N_6152,N_5979);
nand U6292 (N_6292,N_5888,N_5884);
xor U6293 (N_6293,N_5999,N_5934);
xor U6294 (N_6294,N_6076,N_5839);
xor U6295 (N_6295,N_5727,N_6218);
and U6296 (N_6296,N_5869,N_6102);
xor U6297 (N_6297,N_5891,N_6144);
xnor U6298 (N_6298,N_5883,N_5943);
and U6299 (N_6299,N_6023,N_6172);
nand U6300 (N_6300,N_5645,N_5696);
or U6301 (N_6301,N_5878,N_6139);
xor U6302 (N_6302,N_6200,N_5826);
nor U6303 (N_6303,N_6249,N_5933);
nand U6304 (N_6304,N_6083,N_5983);
nand U6305 (N_6305,N_6118,N_5802);
xnor U6306 (N_6306,N_5951,N_5958);
nor U6307 (N_6307,N_5918,N_6110);
nor U6308 (N_6308,N_6106,N_5810);
nor U6309 (N_6309,N_5952,N_6143);
or U6310 (N_6310,N_6174,N_6031);
xor U6311 (N_6311,N_6173,N_5734);
xnor U6312 (N_6312,N_6087,N_5967);
or U6313 (N_6313,N_5901,N_6214);
and U6314 (N_6314,N_5729,N_6061);
nor U6315 (N_6315,N_5743,N_5691);
xor U6316 (N_6316,N_5785,N_6114);
xor U6317 (N_6317,N_5666,N_5956);
xnor U6318 (N_6318,N_5844,N_6125);
nand U6319 (N_6319,N_5811,N_5866);
or U6320 (N_6320,N_5966,N_6092);
and U6321 (N_6321,N_5778,N_6021);
nor U6322 (N_6322,N_5927,N_5784);
or U6323 (N_6323,N_5996,N_5757);
or U6324 (N_6324,N_5819,N_5675);
xnor U6325 (N_6325,N_5882,N_6213);
nor U6326 (N_6326,N_6184,N_5948);
and U6327 (N_6327,N_5658,N_5642);
or U6328 (N_6328,N_6147,N_6121);
nand U6329 (N_6329,N_5671,N_5669);
xor U6330 (N_6330,N_6177,N_5782);
and U6331 (N_6331,N_6065,N_5689);
xnor U6332 (N_6332,N_5900,N_5770);
and U6333 (N_6333,N_5865,N_6028);
nand U6334 (N_6334,N_5858,N_5777);
or U6335 (N_6335,N_6048,N_5747);
and U6336 (N_6336,N_5902,N_6133);
and U6337 (N_6337,N_5674,N_5706);
nor U6338 (N_6338,N_5974,N_6217);
nand U6339 (N_6339,N_5648,N_6163);
xnor U6340 (N_6340,N_5700,N_6130);
and U6341 (N_6341,N_6236,N_5938);
or U6342 (N_6342,N_6215,N_6010);
xnor U6343 (N_6343,N_5634,N_5717);
or U6344 (N_6344,N_5841,N_5981);
xor U6345 (N_6345,N_5633,N_5781);
or U6346 (N_6346,N_6049,N_6132);
nor U6347 (N_6347,N_5939,N_5772);
and U6348 (N_6348,N_5737,N_5657);
or U6349 (N_6349,N_6185,N_5711);
nand U6350 (N_6350,N_6242,N_6162);
nor U6351 (N_6351,N_5885,N_6091);
or U6352 (N_6352,N_6113,N_5847);
nand U6353 (N_6353,N_5698,N_5978);
xor U6354 (N_6354,N_5655,N_6088);
and U6355 (N_6355,N_5636,N_6161);
and U6356 (N_6356,N_5969,N_5880);
nand U6357 (N_6357,N_5861,N_6208);
xnor U6358 (N_6358,N_6036,N_5765);
and U6359 (N_6359,N_5879,N_6020);
and U6360 (N_6360,N_6052,N_5906);
xor U6361 (N_6361,N_6013,N_5721);
or U6362 (N_6362,N_6099,N_6224);
or U6363 (N_6363,N_6026,N_5834);
and U6364 (N_6364,N_5980,N_5805);
or U6365 (N_6365,N_5894,N_5795);
and U6366 (N_6366,N_5926,N_6071);
nand U6367 (N_6367,N_5720,N_5783);
nand U6368 (N_6368,N_5724,N_5923);
and U6369 (N_6369,N_6189,N_5740);
nand U6370 (N_6370,N_5965,N_5828);
or U6371 (N_6371,N_6009,N_5870);
or U6372 (N_6372,N_5759,N_6204);
nand U6373 (N_6373,N_5836,N_5849);
or U6374 (N_6374,N_6055,N_6058);
nor U6375 (N_6375,N_5775,N_5650);
or U6376 (N_6376,N_5886,N_6064);
nor U6377 (N_6377,N_5876,N_6078);
or U6378 (N_6378,N_6196,N_5915);
xnor U6379 (N_6379,N_5824,N_5684);
or U6380 (N_6380,N_6129,N_6201);
nand U6381 (N_6381,N_5859,N_6231);
nand U6382 (N_6382,N_6157,N_5726);
or U6383 (N_6383,N_5661,N_5803);
nand U6384 (N_6384,N_5827,N_6018);
and U6385 (N_6385,N_6225,N_5629);
and U6386 (N_6386,N_6047,N_6120);
or U6387 (N_6387,N_6097,N_6151);
and U6388 (N_6388,N_5680,N_6167);
and U6389 (N_6389,N_5823,N_6193);
or U6390 (N_6390,N_5990,N_5731);
and U6391 (N_6391,N_6050,N_6123);
and U6392 (N_6392,N_5699,N_6206);
xnor U6393 (N_6393,N_5768,N_5916);
and U6394 (N_6394,N_5748,N_5769);
nor U6395 (N_6395,N_6075,N_5761);
or U6396 (N_6396,N_6112,N_6111);
and U6397 (N_6397,N_6191,N_5851);
nand U6398 (N_6398,N_6073,N_5753);
nand U6399 (N_6399,N_5840,N_6197);
nand U6400 (N_6400,N_5975,N_5817);
xnor U6401 (N_6401,N_6209,N_5833);
and U6402 (N_6402,N_5871,N_5822);
or U6403 (N_6403,N_5754,N_6238);
and U6404 (N_6404,N_6192,N_6035);
nor U6405 (N_6405,N_5774,N_5905);
nand U6406 (N_6406,N_6101,N_5742);
nor U6407 (N_6407,N_6155,N_6027);
xnor U6408 (N_6408,N_5896,N_6227);
nor U6409 (N_6409,N_5723,N_5936);
nor U6410 (N_6410,N_5677,N_5752);
or U6411 (N_6411,N_6098,N_6199);
or U6412 (N_6412,N_5762,N_6100);
nand U6413 (N_6413,N_5798,N_5925);
nor U6414 (N_6414,N_5835,N_6126);
nor U6415 (N_6415,N_5714,N_6150);
nor U6416 (N_6416,N_6248,N_5730);
and U6417 (N_6417,N_5982,N_5688);
nand U6418 (N_6418,N_5809,N_6103);
xor U6419 (N_6419,N_5856,N_5853);
xnor U6420 (N_6420,N_6243,N_6222);
nand U6421 (N_6421,N_6219,N_5637);
or U6422 (N_6422,N_5707,N_5673);
and U6423 (N_6423,N_5977,N_5660);
nand U6424 (N_6424,N_6221,N_5703);
nand U6425 (N_6425,N_6005,N_6039);
and U6426 (N_6426,N_6082,N_6034);
nor U6427 (N_6427,N_6235,N_5756);
and U6428 (N_6428,N_6085,N_5646);
or U6429 (N_6429,N_5892,N_5656);
or U6430 (N_6430,N_5991,N_5764);
xor U6431 (N_6431,N_5744,N_5945);
nand U6432 (N_6432,N_5643,N_5801);
nor U6433 (N_6433,N_5668,N_5683);
or U6434 (N_6434,N_6171,N_5667);
and U6435 (N_6435,N_5710,N_6179);
and U6436 (N_6436,N_5984,N_5713);
or U6437 (N_6437,N_6068,N_5718);
or U6438 (N_6438,N_5808,N_6134);
nor U6439 (N_6439,N_6038,N_6119);
nand U6440 (N_6440,N_5697,N_6205);
nand U6441 (N_6441,N_6011,N_5640);
nor U6442 (N_6442,N_6175,N_6153);
xor U6443 (N_6443,N_6116,N_6182);
nand U6444 (N_6444,N_6212,N_6079);
or U6445 (N_6445,N_6247,N_6024);
or U6446 (N_6446,N_6045,N_6051);
xnor U6447 (N_6447,N_6223,N_5820);
nor U6448 (N_6448,N_6053,N_5852);
nor U6449 (N_6449,N_6041,N_6080);
xor U6450 (N_6450,N_6240,N_5860);
or U6451 (N_6451,N_6186,N_6046);
xor U6452 (N_6452,N_6183,N_5997);
nor U6453 (N_6453,N_5804,N_5628);
and U6454 (N_6454,N_5962,N_6239);
nand U6455 (N_6455,N_6156,N_5794);
and U6456 (N_6456,N_6115,N_6014);
xnor U6457 (N_6457,N_5904,N_6145);
nor U6458 (N_6458,N_6154,N_6195);
xor U6459 (N_6459,N_5995,N_5789);
or U6460 (N_6460,N_6057,N_6198);
and U6461 (N_6461,N_5625,N_5961);
nand U6462 (N_6462,N_5897,N_6169);
and U6463 (N_6463,N_5989,N_5653);
or U6464 (N_6464,N_5998,N_5947);
or U6465 (N_6465,N_6017,N_5976);
or U6466 (N_6466,N_5899,N_6008);
xor U6467 (N_6467,N_5716,N_6089);
nand U6468 (N_6468,N_5931,N_5725);
or U6469 (N_6469,N_5701,N_6107);
nand U6470 (N_6470,N_5750,N_6246);
and U6471 (N_6471,N_5790,N_6072);
nand U6472 (N_6472,N_5857,N_6140);
xnor U6473 (N_6473,N_5887,N_5672);
nor U6474 (N_6474,N_6180,N_5749);
and U6475 (N_6475,N_6244,N_5719);
and U6476 (N_6476,N_5914,N_5733);
xnor U6477 (N_6477,N_5890,N_5994);
nand U6478 (N_6478,N_6220,N_6245);
xor U6479 (N_6479,N_5986,N_5881);
nand U6480 (N_6480,N_6074,N_6233);
xor U6481 (N_6481,N_5862,N_6166);
nor U6482 (N_6482,N_5903,N_5920);
and U6483 (N_6483,N_5873,N_6043);
and U6484 (N_6484,N_5644,N_6237);
nand U6485 (N_6485,N_5627,N_5813);
or U6486 (N_6486,N_5932,N_6044);
or U6487 (N_6487,N_6188,N_6040);
or U6488 (N_6488,N_6109,N_5867);
xnor U6489 (N_6489,N_6095,N_5639);
or U6490 (N_6490,N_5773,N_5924);
nand U6491 (N_6491,N_5953,N_5755);
nand U6492 (N_6492,N_5678,N_5993);
xnor U6493 (N_6493,N_6203,N_5690);
xnor U6494 (N_6494,N_5850,N_5806);
nor U6495 (N_6495,N_5941,N_5659);
or U6496 (N_6496,N_5907,N_5973);
xor U6497 (N_6497,N_5776,N_6054);
nor U6498 (N_6498,N_6160,N_6230);
xor U6499 (N_6499,N_5791,N_5912);
or U6500 (N_6500,N_5709,N_6187);
or U6501 (N_6501,N_5641,N_6001);
and U6502 (N_6502,N_5735,N_6234);
xor U6503 (N_6503,N_6003,N_6007);
nand U6504 (N_6504,N_5971,N_6033);
nor U6505 (N_6505,N_5970,N_6194);
nor U6506 (N_6506,N_5935,N_5992);
and U6507 (N_6507,N_5954,N_5877);
or U6508 (N_6508,N_5874,N_6168);
or U6509 (N_6509,N_6006,N_5746);
and U6510 (N_6510,N_5788,N_6081);
xnor U6511 (N_6511,N_5959,N_5832);
nor U6512 (N_6512,N_5780,N_5987);
xnor U6513 (N_6513,N_5909,N_5930);
and U6514 (N_6514,N_6228,N_5687);
or U6515 (N_6515,N_6137,N_5942);
xor U6516 (N_6516,N_5695,N_6086);
or U6517 (N_6517,N_6164,N_5898);
nor U6518 (N_6518,N_5893,N_5960);
nand U6519 (N_6519,N_5705,N_5676);
xor U6520 (N_6520,N_6211,N_5704);
xnor U6521 (N_6521,N_5816,N_5937);
and U6522 (N_6522,N_5940,N_5793);
and U6523 (N_6523,N_5928,N_6135);
nor U6524 (N_6524,N_5964,N_5814);
nand U6525 (N_6525,N_5760,N_5812);
xor U6526 (N_6526,N_6056,N_6127);
nor U6527 (N_6527,N_5649,N_6012);
or U6528 (N_6528,N_5910,N_5988);
and U6529 (N_6529,N_5728,N_6148);
nand U6530 (N_6530,N_6136,N_5895);
nand U6531 (N_6531,N_5736,N_5664);
or U6532 (N_6532,N_5963,N_6063);
and U6533 (N_6533,N_5792,N_5838);
and U6534 (N_6534,N_6015,N_6149);
nor U6535 (N_6535,N_6060,N_6159);
nand U6536 (N_6536,N_6029,N_5632);
xor U6537 (N_6537,N_6202,N_6002);
xor U6538 (N_6538,N_5799,N_5830);
xnor U6539 (N_6539,N_5654,N_6090);
and U6540 (N_6540,N_5665,N_5693);
nand U6541 (N_6541,N_5652,N_5913);
nand U6542 (N_6542,N_5855,N_5681);
nand U6543 (N_6543,N_5779,N_5682);
or U6544 (N_6544,N_5766,N_6146);
nor U6545 (N_6545,N_6077,N_5651);
xnor U6546 (N_6546,N_5957,N_5950);
or U6547 (N_6547,N_6032,N_6108);
nand U6548 (N_6548,N_5944,N_6016);
and U6549 (N_6549,N_6241,N_6216);
nand U6550 (N_6550,N_6207,N_6181);
or U6551 (N_6551,N_5868,N_6094);
xnor U6552 (N_6552,N_6138,N_5864);
nand U6553 (N_6553,N_5825,N_5889);
nor U6554 (N_6554,N_5786,N_5955);
xnor U6555 (N_6555,N_6062,N_5837);
nand U6556 (N_6556,N_5815,N_6141);
nand U6557 (N_6557,N_5845,N_5767);
xor U6558 (N_6558,N_5796,N_5679);
nand U6559 (N_6559,N_5692,N_5771);
nand U6560 (N_6560,N_5686,N_6030);
and U6561 (N_6561,N_6128,N_5702);
nand U6562 (N_6562,N_6122,N_5664);
nand U6563 (N_6563,N_6108,N_5886);
nand U6564 (N_6564,N_6137,N_5822);
and U6565 (N_6565,N_6181,N_6110);
or U6566 (N_6566,N_5829,N_5976);
and U6567 (N_6567,N_5765,N_5707);
nand U6568 (N_6568,N_6067,N_5764);
nor U6569 (N_6569,N_5947,N_6143);
or U6570 (N_6570,N_5812,N_6093);
xor U6571 (N_6571,N_5927,N_5706);
and U6572 (N_6572,N_5714,N_6029);
nor U6573 (N_6573,N_5830,N_5724);
and U6574 (N_6574,N_6075,N_6104);
and U6575 (N_6575,N_6039,N_5807);
nand U6576 (N_6576,N_5830,N_5930);
xnor U6577 (N_6577,N_5664,N_5757);
and U6578 (N_6578,N_5941,N_5939);
nand U6579 (N_6579,N_6198,N_6032);
nand U6580 (N_6580,N_6209,N_6065);
xnor U6581 (N_6581,N_5747,N_5659);
and U6582 (N_6582,N_6206,N_5940);
or U6583 (N_6583,N_6094,N_5935);
and U6584 (N_6584,N_6052,N_5897);
nor U6585 (N_6585,N_6144,N_6154);
nand U6586 (N_6586,N_6243,N_5714);
or U6587 (N_6587,N_5694,N_5912);
xor U6588 (N_6588,N_5838,N_5920);
and U6589 (N_6589,N_6012,N_5847);
and U6590 (N_6590,N_6083,N_6131);
nor U6591 (N_6591,N_6098,N_6206);
and U6592 (N_6592,N_6158,N_5997);
and U6593 (N_6593,N_5972,N_6040);
and U6594 (N_6594,N_5692,N_5997);
nand U6595 (N_6595,N_5731,N_6211);
and U6596 (N_6596,N_5748,N_5972);
and U6597 (N_6597,N_5770,N_6016);
nor U6598 (N_6598,N_6221,N_5788);
or U6599 (N_6599,N_5936,N_5853);
or U6600 (N_6600,N_6095,N_5729);
nor U6601 (N_6601,N_6212,N_6061);
or U6602 (N_6602,N_5711,N_6160);
and U6603 (N_6603,N_5985,N_5945);
and U6604 (N_6604,N_6076,N_6146);
or U6605 (N_6605,N_5698,N_5930);
and U6606 (N_6606,N_6047,N_6075);
nor U6607 (N_6607,N_5666,N_5780);
nand U6608 (N_6608,N_6241,N_5711);
or U6609 (N_6609,N_5681,N_6120);
xnor U6610 (N_6610,N_5712,N_5945);
nand U6611 (N_6611,N_5823,N_6203);
xor U6612 (N_6612,N_6196,N_5991);
xor U6613 (N_6613,N_5684,N_5891);
xnor U6614 (N_6614,N_5841,N_5917);
or U6615 (N_6615,N_5977,N_5813);
nor U6616 (N_6616,N_5679,N_6196);
nor U6617 (N_6617,N_5743,N_5703);
xnor U6618 (N_6618,N_6189,N_5716);
xnor U6619 (N_6619,N_6152,N_5872);
xnor U6620 (N_6620,N_6113,N_6015);
and U6621 (N_6621,N_5789,N_5798);
nor U6622 (N_6622,N_5979,N_5882);
nand U6623 (N_6623,N_5860,N_5772);
xnor U6624 (N_6624,N_5873,N_6059);
nand U6625 (N_6625,N_5663,N_5926);
nor U6626 (N_6626,N_5929,N_6118);
xnor U6627 (N_6627,N_6004,N_5852);
and U6628 (N_6628,N_5802,N_5847);
xor U6629 (N_6629,N_6217,N_5976);
or U6630 (N_6630,N_5997,N_5850);
nand U6631 (N_6631,N_5675,N_6114);
nand U6632 (N_6632,N_5879,N_6023);
xor U6633 (N_6633,N_5985,N_6011);
nand U6634 (N_6634,N_6095,N_6119);
or U6635 (N_6635,N_6125,N_5654);
and U6636 (N_6636,N_5866,N_5657);
or U6637 (N_6637,N_5980,N_6073);
or U6638 (N_6638,N_5777,N_5842);
nor U6639 (N_6639,N_5952,N_6194);
or U6640 (N_6640,N_5783,N_5759);
and U6641 (N_6641,N_5889,N_6104);
nand U6642 (N_6642,N_5722,N_5909);
and U6643 (N_6643,N_6049,N_6147);
and U6644 (N_6644,N_5679,N_6222);
nor U6645 (N_6645,N_5863,N_5824);
and U6646 (N_6646,N_6012,N_6122);
nor U6647 (N_6647,N_5946,N_5764);
xor U6648 (N_6648,N_5704,N_6191);
and U6649 (N_6649,N_6223,N_6184);
xor U6650 (N_6650,N_5868,N_5636);
nor U6651 (N_6651,N_6162,N_5890);
nand U6652 (N_6652,N_5762,N_5849);
or U6653 (N_6653,N_6128,N_6217);
or U6654 (N_6654,N_5805,N_6091);
xor U6655 (N_6655,N_6245,N_5894);
xor U6656 (N_6656,N_6023,N_5847);
or U6657 (N_6657,N_6026,N_6065);
xnor U6658 (N_6658,N_5808,N_5880);
xor U6659 (N_6659,N_5721,N_6230);
and U6660 (N_6660,N_5832,N_6056);
and U6661 (N_6661,N_6034,N_6063);
or U6662 (N_6662,N_5814,N_5708);
nand U6663 (N_6663,N_5967,N_5919);
nor U6664 (N_6664,N_5727,N_6053);
nor U6665 (N_6665,N_6219,N_5970);
xor U6666 (N_6666,N_6148,N_6113);
and U6667 (N_6667,N_6005,N_6012);
and U6668 (N_6668,N_5666,N_5896);
xor U6669 (N_6669,N_5868,N_5960);
nor U6670 (N_6670,N_5664,N_6130);
or U6671 (N_6671,N_5770,N_5826);
or U6672 (N_6672,N_5844,N_5656);
xor U6673 (N_6673,N_5695,N_5790);
xnor U6674 (N_6674,N_6172,N_5799);
xor U6675 (N_6675,N_6008,N_5757);
or U6676 (N_6676,N_5726,N_6204);
nand U6677 (N_6677,N_6150,N_5926);
xnor U6678 (N_6678,N_5773,N_6204);
nand U6679 (N_6679,N_6240,N_5937);
nor U6680 (N_6680,N_5690,N_6123);
nor U6681 (N_6681,N_6104,N_6201);
and U6682 (N_6682,N_5856,N_5785);
and U6683 (N_6683,N_6060,N_6059);
xor U6684 (N_6684,N_6202,N_5836);
or U6685 (N_6685,N_6149,N_6067);
nor U6686 (N_6686,N_6151,N_5652);
and U6687 (N_6687,N_5724,N_5949);
nand U6688 (N_6688,N_5666,N_5813);
xor U6689 (N_6689,N_5862,N_5662);
nor U6690 (N_6690,N_5967,N_5631);
xor U6691 (N_6691,N_5865,N_5812);
and U6692 (N_6692,N_5749,N_6083);
and U6693 (N_6693,N_6103,N_6003);
nor U6694 (N_6694,N_5659,N_6176);
nor U6695 (N_6695,N_6002,N_6194);
xor U6696 (N_6696,N_6098,N_6126);
nor U6697 (N_6697,N_6030,N_5862);
nand U6698 (N_6698,N_6171,N_5832);
and U6699 (N_6699,N_6186,N_5625);
or U6700 (N_6700,N_5853,N_6039);
nor U6701 (N_6701,N_6214,N_5639);
and U6702 (N_6702,N_5681,N_5914);
xor U6703 (N_6703,N_5782,N_5851);
nor U6704 (N_6704,N_5732,N_5627);
nand U6705 (N_6705,N_5868,N_5713);
nor U6706 (N_6706,N_5715,N_5887);
nor U6707 (N_6707,N_5984,N_5722);
nand U6708 (N_6708,N_6211,N_6117);
nand U6709 (N_6709,N_6234,N_5955);
or U6710 (N_6710,N_5877,N_5907);
nand U6711 (N_6711,N_6014,N_6040);
nor U6712 (N_6712,N_6022,N_5799);
or U6713 (N_6713,N_5798,N_6229);
nand U6714 (N_6714,N_5807,N_5662);
or U6715 (N_6715,N_6230,N_6121);
xor U6716 (N_6716,N_6005,N_5876);
or U6717 (N_6717,N_5627,N_5838);
or U6718 (N_6718,N_5837,N_5909);
nand U6719 (N_6719,N_6004,N_6030);
and U6720 (N_6720,N_5996,N_5970);
and U6721 (N_6721,N_5675,N_5975);
and U6722 (N_6722,N_6211,N_5947);
and U6723 (N_6723,N_5736,N_6073);
nor U6724 (N_6724,N_6087,N_5646);
xnor U6725 (N_6725,N_6031,N_5708);
xor U6726 (N_6726,N_5684,N_6158);
xor U6727 (N_6727,N_6032,N_5728);
or U6728 (N_6728,N_5909,N_6143);
nor U6729 (N_6729,N_6212,N_5880);
xnor U6730 (N_6730,N_5767,N_5755);
and U6731 (N_6731,N_5746,N_6121);
nor U6732 (N_6732,N_6154,N_6224);
nand U6733 (N_6733,N_5789,N_5654);
or U6734 (N_6734,N_5751,N_6035);
xnor U6735 (N_6735,N_5851,N_5849);
or U6736 (N_6736,N_5885,N_5775);
and U6737 (N_6737,N_6170,N_6107);
nor U6738 (N_6738,N_5694,N_5867);
xor U6739 (N_6739,N_5880,N_6112);
or U6740 (N_6740,N_5687,N_6102);
nor U6741 (N_6741,N_6109,N_5849);
and U6742 (N_6742,N_6153,N_5942);
nand U6743 (N_6743,N_6116,N_5746);
and U6744 (N_6744,N_5790,N_5673);
nand U6745 (N_6745,N_5877,N_5915);
nor U6746 (N_6746,N_6020,N_5805);
nor U6747 (N_6747,N_5734,N_6084);
nand U6748 (N_6748,N_6237,N_5649);
or U6749 (N_6749,N_6019,N_5968);
or U6750 (N_6750,N_5902,N_5932);
and U6751 (N_6751,N_6008,N_5799);
nor U6752 (N_6752,N_6021,N_6199);
nor U6753 (N_6753,N_6190,N_6106);
xnor U6754 (N_6754,N_5656,N_5707);
xnor U6755 (N_6755,N_5694,N_5740);
or U6756 (N_6756,N_5832,N_5874);
or U6757 (N_6757,N_6102,N_6246);
and U6758 (N_6758,N_5871,N_5636);
xnor U6759 (N_6759,N_6208,N_5644);
nand U6760 (N_6760,N_6153,N_6202);
nor U6761 (N_6761,N_5763,N_5758);
nand U6762 (N_6762,N_6126,N_6232);
xor U6763 (N_6763,N_6168,N_6241);
and U6764 (N_6764,N_6021,N_5764);
or U6765 (N_6765,N_6184,N_6109);
nand U6766 (N_6766,N_5716,N_6220);
nor U6767 (N_6767,N_5695,N_5743);
or U6768 (N_6768,N_5751,N_6036);
xor U6769 (N_6769,N_5999,N_5656);
xnor U6770 (N_6770,N_6101,N_5782);
or U6771 (N_6771,N_5734,N_5681);
and U6772 (N_6772,N_5976,N_5734);
and U6773 (N_6773,N_6117,N_5916);
nand U6774 (N_6774,N_5854,N_5809);
xnor U6775 (N_6775,N_5657,N_6013);
nor U6776 (N_6776,N_6115,N_6145);
nor U6777 (N_6777,N_6233,N_6102);
xnor U6778 (N_6778,N_5852,N_6055);
nor U6779 (N_6779,N_6152,N_5705);
or U6780 (N_6780,N_5889,N_5993);
nor U6781 (N_6781,N_5819,N_5981);
xor U6782 (N_6782,N_5934,N_6192);
and U6783 (N_6783,N_5960,N_6183);
xor U6784 (N_6784,N_5648,N_6088);
nand U6785 (N_6785,N_5803,N_6242);
nor U6786 (N_6786,N_6115,N_6111);
xnor U6787 (N_6787,N_5945,N_5967);
xnor U6788 (N_6788,N_5791,N_5965);
nor U6789 (N_6789,N_5918,N_6013);
and U6790 (N_6790,N_5674,N_6056);
xnor U6791 (N_6791,N_5866,N_6092);
xnor U6792 (N_6792,N_5675,N_5955);
or U6793 (N_6793,N_6066,N_5642);
xnor U6794 (N_6794,N_5751,N_6117);
or U6795 (N_6795,N_6115,N_5671);
and U6796 (N_6796,N_6056,N_5852);
nor U6797 (N_6797,N_5942,N_6087);
nand U6798 (N_6798,N_6089,N_5878);
and U6799 (N_6799,N_6041,N_6127);
or U6800 (N_6800,N_6161,N_5971);
xor U6801 (N_6801,N_5750,N_5877);
nand U6802 (N_6802,N_6222,N_6185);
nor U6803 (N_6803,N_5749,N_6165);
nand U6804 (N_6804,N_5841,N_6147);
nand U6805 (N_6805,N_5769,N_6143);
and U6806 (N_6806,N_6071,N_6249);
nor U6807 (N_6807,N_6155,N_6182);
xnor U6808 (N_6808,N_5965,N_5919);
and U6809 (N_6809,N_5714,N_5845);
xnor U6810 (N_6810,N_5817,N_5852);
nand U6811 (N_6811,N_5680,N_5948);
xor U6812 (N_6812,N_6193,N_5975);
or U6813 (N_6813,N_6235,N_5899);
nor U6814 (N_6814,N_6180,N_6048);
nor U6815 (N_6815,N_5991,N_6000);
or U6816 (N_6816,N_5955,N_6215);
nor U6817 (N_6817,N_5697,N_5934);
nand U6818 (N_6818,N_5713,N_5708);
nand U6819 (N_6819,N_5803,N_5840);
and U6820 (N_6820,N_5953,N_5797);
or U6821 (N_6821,N_5752,N_6224);
or U6822 (N_6822,N_5699,N_6058);
nor U6823 (N_6823,N_6021,N_6054);
nor U6824 (N_6824,N_6202,N_6040);
xnor U6825 (N_6825,N_5720,N_5742);
nor U6826 (N_6826,N_5974,N_6154);
nand U6827 (N_6827,N_6215,N_5850);
nand U6828 (N_6828,N_5744,N_5708);
nor U6829 (N_6829,N_5790,N_6033);
xor U6830 (N_6830,N_6239,N_5879);
or U6831 (N_6831,N_6137,N_5974);
nor U6832 (N_6832,N_5948,N_5954);
nand U6833 (N_6833,N_5994,N_6107);
nand U6834 (N_6834,N_5927,N_5729);
or U6835 (N_6835,N_6120,N_5683);
nand U6836 (N_6836,N_5816,N_5745);
or U6837 (N_6837,N_5849,N_5856);
nand U6838 (N_6838,N_6000,N_6244);
nand U6839 (N_6839,N_5935,N_5878);
and U6840 (N_6840,N_5847,N_6231);
nand U6841 (N_6841,N_5726,N_5858);
and U6842 (N_6842,N_5729,N_5626);
nand U6843 (N_6843,N_5954,N_5829);
nor U6844 (N_6844,N_6071,N_5689);
or U6845 (N_6845,N_6128,N_5820);
nor U6846 (N_6846,N_6108,N_5914);
xor U6847 (N_6847,N_6207,N_6244);
xnor U6848 (N_6848,N_5817,N_5943);
xnor U6849 (N_6849,N_6149,N_5668);
nand U6850 (N_6850,N_6113,N_5909);
xnor U6851 (N_6851,N_5946,N_5641);
or U6852 (N_6852,N_5634,N_6006);
nand U6853 (N_6853,N_6077,N_6170);
nor U6854 (N_6854,N_6120,N_6168);
nor U6855 (N_6855,N_5893,N_6175);
or U6856 (N_6856,N_6128,N_5736);
nor U6857 (N_6857,N_5810,N_6096);
nor U6858 (N_6858,N_6121,N_6123);
nand U6859 (N_6859,N_6012,N_5739);
nand U6860 (N_6860,N_5813,N_5925);
and U6861 (N_6861,N_5790,N_5816);
nand U6862 (N_6862,N_6156,N_5665);
nand U6863 (N_6863,N_5853,N_5868);
nand U6864 (N_6864,N_6142,N_5801);
xor U6865 (N_6865,N_5852,N_5978);
xor U6866 (N_6866,N_5903,N_5811);
or U6867 (N_6867,N_6037,N_5686);
nand U6868 (N_6868,N_6043,N_6089);
nor U6869 (N_6869,N_5775,N_6245);
and U6870 (N_6870,N_6133,N_6067);
nand U6871 (N_6871,N_6053,N_6068);
xnor U6872 (N_6872,N_5642,N_6083);
or U6873 (N_6873,N_5665,N_5831);
and U6874 (N_6874,N_5704,N_6026);
and U6875 (N_6875,N_6575,N_6484);
or U6876 (N_6876,N_6828,N_6726);
nor U6877 (N_6877,N_6747,N_6792);
or U6878 (N_6878,N_6387,N_6369);
nand U6879 (N_6879,N_6839,N_6349);
and U6880 (N_6880,N_6346,N_6371);
and U6881 (N_6881,N_6717,N_6427);
and U6882 (N_6882,N_6831,N_6347);
or U6883 (N_6883,N_6825,N_6262);
nand U6884 (N_6884,N_6592,N_6801);
xor U6885 (N_6885,N_6525,N_6664);
nor U6886 (N_6886,N_6284,N_6742);
and U6887 (N_6887,N_6620,N_6848);
xor U6888 (N_6888,N_6844,N_6463);
nand U6889 (N_6889,N_6430,N_6336);
or U6890 (N_6890,N_6351,N_6305);
nand U6891 (N_6891,N_6641,N_6368);
nor U6892 (N_6892,N_6542,N_6373);
or U6893 (N_6893,N_6447,N_6609);
or U6894 (N_6894,N_6297,N_6377);
or U6895 (N_6895,N_6398,N_6335);
nand U6896 (N_6896,N_6822,N_6674);
xor U6897 (N_6897,N_6680,N_6687);
nor U6898 (N_6898,N_6867,N_6590);
nor U6899 (N_6899,N_6526,N_6514);
nor U6900 (N_6900,N_6438,N_6709);
or U6901 (N_6901,N_6589,N_6282);
nor U6902 (N_6902,N_6711,N_6396);
or U6903 (N_6903,N_6385,N_6344);
xor U6904 (N_6904,N_6550,N_6661);
or U6905 (N_6905,N_6751,N_6401);
or U6906 (N_6906,N_6557,N_6395);
nand U6907 (N_6907,N_6653,N_6611);
nor U6908 (N_6908,N_6363,N_6724);
or U6909 (N_6909,N_6291,N_6745);
and U6910 (N_6910,N_6636,N_6800);
and U6911 (N_6911,N_6374,N_6562);
nor U6912 (N_6912,N_6389,N_6418);
and U6913 (N_6913,N_6443,N_6585);
and U6914 (N_6914,N_6362,N_6261);
nor U6915 (N_6915,N_6416,N_6692);
nand U6916 (N_6916,N_6712,N_6422);
or U6917 (N_6917,N_6666,N_6415);
nor U6918 (N_6918,N_6440,N_6569);
xor U6919 (N_6919,N_6798,N_6582);
nand U6920 (N_6920,N_6728,N_6588);
and U6921 (N_6921,N_6504,N_6543);
nor U6922 (N_6922,N_6468,N_6672);
and U6923 (N_6923,N_6546,N_6830);
or U6924 (N_6924,N_6425,N_6823);
xnor U6925 (N_6925,N_6773,N_6849);
and U6926 (N_6926,N_6423,N_6301);
nand U6927 (N_6927,N_6325,N_6675);
nor U6928 (N_6928,N_6690,N_6860);
nand U6929 (N_6929,N_6518,N_6639);
or U6930 (N_6930,N_6775,N_6436);
and U6931 (N_6931,N_6413,N_6458);
or U6932 (N_6932,N_6870,N_6857);
xnor U6933 (N_6933,N_6571,N_6784);
nor U6934 (N_6934,N_6730,N_6670);
xnor U6935 (N_6935,N_6621,N_6497);
nor U6936 (N_6936,N_6281,N_6782);
nor U6937 (N_6937,N_6303,N_6622);
nor U6938 (N_6938,N_6506,N_6854);
xor U6939 (N_6939,N_6759,N_6272);
nand U6940 (N_6940,N_6265,N_6277);
or U6941 (N_6941,N_6250,N_6383);
xnor U6942 (N_6942,N_6379,N_6523);
xor U6943 (N_6943,N_6693,N_6629);
nand U6944 (N_6944,N_6599,N_6421);
or U6945 (N_6945,N_6407,N_6763);
and U6946 (N_6946,N_6818,N_6684);
and U6947 (N_6947,N_6453,N_6428);
nand U6948 (N_6948,N_6686,N_6476);
and U6949 (N_6949,N_6833,N_6827);
nand U6950 (N_6950,N_6604,N_6280);
nor U6951 (N_6951,N_6299,N_6273);
xnor U6952 (N_6952,N_6851,N_6475);
xnor U6953 (N_6953,N_6859,N_6276);
or U6954 (N_6954,N_6507,N_6719);
and U6955 (N_6955,N_6433,N_6834);
nand U6956 (N_6956,N_6545,N_6378);
nor U6957 (N_6957,N_6722,N_6847);
or U6958 (N_6958,N_6419,N_6259);
nand U6959 (N_6959,N_6360,N_6862);
nor U6960 (N_6960,N_6274,N_6630);
and U6961 (N_6961,N_6873,N_6489);
nand U6962 (N_6962,N_6841,N_6323);
xor U6963 (N_6963,N_6471,N_6723);
and U6964 (N_6964,N_6382,N_6289);
nand U6965 (N_6965,N_6766,N_6771);
or U6966 (N_6966,N_6739,N_6527);
xnor U6967 (N_6967,N_6811,N_6406);
and U6968 (N_6968,N_6757,N_6326);
xor U6969 (N_6969,N_6804,N_6375);
or U6970 (N_6970,N_6561,N_6482);
nor U6971 (N_6971,N_6574,N_6705);
or U6972 (N_6972,N_6499,N_6603);
nand U6973 (N_6973,N_6720,N_6531);
xnor U6974 (N_6974,N_6478,N_6270);
xnor U6975 (N_6975,N_6442,N_6338);
nor U6976 (N_6976,N_6738,N_6402);
xnor U6977 (N_6977,N_6740,N_6777);
nand U6978 (N_6978,N_6713,N_6296);
and U6979 (N_6979,N_6364,N_6549);
nor U6980 (N_6980,N_6601,N_6566);
nor U6981 (N_6981,N_6665,N_6736);
and U6982 (N_6982,N_6460,N_6725);
or U6983 (N_6983,N_6619,N_6455);
nor U6984 (N_6984,N_6807,N_6330);
and U6985 (N_6985,N_6733,N_6864);
xnor U6986 (N_6986,N_6477,N_6308);
nor U6987 (N_6987,N_6521,N_6488);
nor U6988 (N_6988,N_6753,N_6492);
nor U6989 (N_6989,N_6858,N_6676);
nor U6990 (N_6990,N_6394,N_6457);
nor U6991 (N_6991,N_6780,N_6474);
and U6992 (N_6992,N_6532,N_6626);
and U6993 (N_6993,N_6449,N_6644);
and U6994 (N_6994,N_6324,N_6637);
nor U6995 (N_6995,N_6699,N_6439);
or U6996 (N_6996,N_6361,N_6555);
or U6997 (N_6997,N_6567,N_6617);
nor U6998 (N_6998,N_6600,N_6372);
xnor U6999 (N_6999,N_6348,N_6317);
or U7000 (N_7000,N_6863,N_6649);
xnor U7001 (N_7001,N_6537,N_6624);
nor U7002 (N_7002,N_6703,N_6657);
and U7003 (N_7003,N_6577,N_6431);
nor U7004 (N_7004,N_6695,N_6528);
or U7005 (N_7005,N_6251,N_6522);
nand U7006 (N_7006,N_6467,N_6683);
and U7007 (N_7007,N_6496,N_6586);
nand U7008 (N_7008,N_6852,N_6832);
and U7009 (N_7009,N_6640,N_6500);
and U7010 (N_7010,N_6815,N_6380);
nand U7011 (N_7011,N_6635,N_6819);
and U7012 (N_7012,N_6610,N_6405);
nand U7013 (N_7013,N_6633,N_6519);
nor U7014 (N_7014,N_6420,N_6721);
and U7015 (N_7015,N_6448,N_6734);
or U7016 (N_7016,N_6573,N_6329);
and U7017 (N_7017,N_6794,N_6316);
nor U7018 (N_7018,N_6286,N_6432);
and U7019 (N_7019,N_6732,N_6283);
nor U7020 (N_7020,N_6824,N_6645);
or U7021 (N_7021,N_6341,N_6466);
nor U7022 (N_7022,N_6812,N_6288);
xor U7023 (N_7023,N_6799,N_6838);
xnor U7024 (N_7024,N_6552,N_6835);
nor U7025 (N_7025,N_6400,N_6746);
xnor U7026 (N_7026,N_6810,N_6454);
nand U7027 (N_7027,N_6483,N_6598);
and U7028 (N_7028,N_6558,N_6581);
nand U7029 (N_7029,N_6874,N_6779);
or U7030 (N_7030,N_6802,N_6370);
or U7031 (N_7031,N_6638,N_6597);
nand U7032 (N_7032,N_6594,N_6365);
nand U7033 (N_7033,N_6718,N_6451);
nand U7034 (N_7034,N_6702,N_6390);
nand U7035 (N_7035,N_6789,N_6342);
or U7036 (N_7036,N_6480,N_6772);
nor U7037 (N_7037,N_6805,N_6333);
or U7038 (N_7038,N_6481,N_6269);
xnor U7039 (N_7039,N_6701,N_6761);
nand U7040 (N_7040,N_6384,N_6691);
nand U7041 (N_7041,N_6788,N_6660);
nand U7042 (N_7042,N_6632,N_6707);
and U7043 (N_7043,N_6503,N_6495);
and U7044 (N_7044,N_6271,N_6354);
xor U7045 (N_7045,N_6461,N_6334);
and U7046 (N_7046,N_6446,N_6696);
nand U7047 (N_7047,N_6541,N_6826);
and U7048 (N_7048,N_6498,N_6714);
or U7049 (N_7049,N_6658,N_6300);
nand U7050 (N_7050,N_6646,N_6345);
nor U7051 (N_7051,N_6313,N_6318);
xor U7052 (N_7052,N_6426,N_6716);
nand U7053 (N_7053,N_6572,N_6790);
nand U7054 (N_7054,N_6530,N_6462);
and U7055 (N_7055,N_6515,N_6791);
and U7056 (N_7056,N_6651,N_6520);
xor U7057 (N_7057,N_6253,N_6294);
nand U7058 (N_7058,N_6627,N_6302);
nand U7059 (N_7059,N_6869,N_6583);
nand U7060 (N_7060,N_6769,N_6606);
nor U7061 (N_7061,N_6605,N_6381);
or U7062 (N_7062,N_6814,N_6536);
and U7063 (N_7063,N_6386,N_6648);
and U7064 (N_7064,N_6358,N_6698);
xnor U7065 (N_7065,N_6332,N_6564);
and U7066 (N_7066,N_6749,N_6285);
xnor U7067 (N_7067,N_6704,N_6319);
xnor U7068 (N_7068,N_6634,N_6808);
and U7069 (N_7069,N_6845,N_6310);
nand U7070 (N_7070,N_6548,N_6786);
and U7071 (N_7071,N_6655,N_6741);
xnor U7072 (N_7072,N_6856,N_6796);
xnor U7073 (N_7073,N_6356,N_6486);
or U7074 (N_7074,N_6544,N_6434);
xor U7075 (N_7075,N_6309,N_6292);
nor U7076 (N_7076,N_6625,N_6682);
and U7077 (N_7077,N_6866,N_6366);
nor U7078 (N_7078,N_6669,N_6776);
nand U7079 (N_7079,N_6256,N_6491);
xnor U7080 (N_7080,N_6524,N_6565);
or U7081 (N_7081,N_6613,N_6450);
nand U7082 (N_7082,N_6821,N_6469);
nand U7083 (N_7083,N_6293,N_6706);
nand U7084 (N_7084,N_6403,N_6560);
xor U7085 (N_7085,N_6459,N_6744);
or U7086 (N_7086,N_6279,N_6511);
nand U7087 (N_7087,N_6809,N_6708);
nor U7088 (N_7088,N_6593,N_6554);
nor U7089 (N_7089,N_6568,N_6659);
nor U7090 (N_7090,N_6322,N_6643);
xnor U7091 (N_7091,N_6367,N_6729);
and U7092 (N_7092,N_6517,N_6410);
xor U7093 (N_7093,N_6836,N_6353);
nand U7094 (N_7094,N_6295,N_6806);
nand U7095 (N_7095,N_6615,N_6429);
nand U7096 (N_7096,N_6260,N_6840);
and U7097 (N_7097,N_6399,N_6444);
or U7098 (N_7098,N_6388,N_6376);
nor U7099 (N_7099,N_6679,N_6578);
or U7100 (N_7100,N_6412,N_6591);
nand U7101 (N_7101,N_6631,N_6414);
and U7102 (N_7102,N_6513,N_6816);
or U7103 (N_7103,N_6352,N_6337);
or U7104 (N_7104,N_6472,N_6465);
nand U7105 (N_7105,N_6464,N_6662);
and U7106 (N_7106,N_6508,N_6781);
or U7107 (N_7107,N_6797,N_6393);
nand U7108 (N_7108,N_6871,N_6311);
nand U7109 (N_7109,N_6538,N_6678);
xor U7110 (N_7110,N_6770,N_6689);
or U7111 (N_7111,N_6473,N_6748);
xnor U7112 (N_7112,N_6268,N_6505);
nor U7113 (N_7113,N_6570,N_6754);
nor U7114 (N_7114,N_6307,N_6304);
nor U7115 (N_7115,N_6512,N_6357);
or U7116 (N_7116,N_6865,N_6737);
nand U7117 (N_7117,N_6793,N_6616);
and U7118 (N_7118,N_6647,N_6339);
and U7119 (N_7119,N_6768,N_6327);
or U7120 (N_7120,N_6846,N_6618);
xor U7121 (N_7121,N_6535,N_6861);
or U7122 (N_7122,N_6563,N_6266);
nor U7123 (N_7123,N_6487,N_6803);
nand U7124 (N_7124,N_6540,N_6392);
nand U7125 (N_7125,N_6391,N_6710);
nor U7126 (N_7126,N_6654,N_6490);
nor U7127 (N_7127,N_6829,N_6758);
or U7128 (N_7128,N_6263,N_6501);
xnor U7129 (N_7129,N_6547,N_6715);
or U7130 (N_7130,N_6756,N_6778);
xor U7131 (N_7131,N_6252,N_6694);
nand U7132 (N_7132,N_6602,N_6350);
xnor U7133 (N_7133,N_6509,N_6556);
and U7134 (N_7134,N_6437,N_6275);
or U7135 (N_7135,N_6853,N_6502);
nand U7136 (N_7136,N_6534,N_6764);
nor U7137 (N_7137,N_6850,N_6516);
xor U7138 (N_7138,N_6494,N_6843);
and U7139 (N_7139,N_6855,N_6559);
xnor U7140 (N_7140,N_6623,N_6652);
and U7141 (N_7141,N_6290,N_6320);
nand U7142 (N_7142,N_6397,N_6355);
nand U7143 (N_7143,N_6668,N_6435);
nor U7144 (N_7144,N_6820,N_6727);
or U7145 (N_7145,N_6842,N_6533);
or U7146 (N_7146,N_6755,N_6743);
nand U7147 (N_7147,N_6872,N_6767);
xnor U7148 (N_7148,N_6612,N_6584);
or U7149 (N_7149,N_6697,N_6596);
nor U7150 (N_7150,N_6783,N_6614);
and U7151 (N_7151,N_6667,N_6331);
or U7152 (N_7152,N_6576,N_6267);
nand U7153 (N_7153,N_6470,N_6595);
or U7154 (N_7154,N_6663,N_6587);
and U7155 (N_7155,N_6813,N_6762);
or U7156 (N_7156,N_6321,N_6411);
or U7157 (N_7157,N_6445,N_6328);
nor U7158 (N_7158,N_6795,N_6343);
nor U7159 (N_7159,N_6314,N_6688);
nor U7160 (N_7160,N_6264,N_6298);
nor U7161 (N_7161,N_6671,N_6685);
nand U7162 (N_7162,N_6485,N_6315);
xnor U7163 (N_7163,N_6539,N_6752);
or U7164 (N_7164,N_6817,N_6765);
or U7165 (N_7165,N_6287,N_6650);
nand U7166 (N_7166,N_6787,N_6456);
or U7167 (N_7167,N_6785,N_6700);
nor U7168 (N_7168,N_6551,N_6579);
nand U7169 (N_7169,N_6404,N_6731);
xnor U7170 (N_7170,N_6750,N_6642);
nor U7171 (N_7171,N_6278,N_6441);
xor U7172 (N_7172,N_6493,N_6673);
or U7173 (N_7173,N_6306,N_6628);
xnor U7174 (N_7174,N_6479,N_6510);
or U7175 (N_7175,N_6258,N_6359);
or U7176 (N_7176,N_6312,N_6340);
xnor U7177 (N_7177,N_6656,N_6607);
nand U7178 (N_7178,N_6580,N_6257);
xor U7179 (N_7179,N_6553,N_6255);
xnor U7180 (N_7180,N_6677,N_6424);
nand U7181 (N_7181,N_6735,N_6837);
nor U7182 (N_7182,N_6774,N_6254);
nor U7183 (N_7183,N_6408,N_6409);
nand U7184 (N_7184,N_6452,N_6868);
nor U7185 (N_7185,N_6681,N_6529);
or U7186 (N_7186,N_6760,N_6608);
nor U7187 (N_7187,N_6417,N_6279);
xor U7188 (N_7188,N_6477,N_6796);
xor U7189 (N_7189,N_6499,N_6419);
and U7190 (N_7190,N_6834,N_6639);
or U7191 (N_7191,N_6560,N_6872);
or U7192 (N_7192,N_6453,N_6789);
or U7193 (N_7193,N_6551,N_6565);
and U7194 (N_7194,N_6469,N_6612);
xnor U7195 (N_7195,N_6574,N_6541);
nor U7196 (N_7196,N_6755,N_6426);
nor U7197 (N_7197,N_6392,N_6631);
or U7198 (N_7198,N_6740,N_6579);
nand U7199 (N_7199,N_6693,N_6442);
or U7200 (N_7200,N_6441,N_6741);
xnor U7201 (N_7201,N_6789,N_6611);
nor U7202 (N_7202,N_6813,N_6810);
nand U7203 (N_7203,N_6477,N_6407);
nor U7204 (N_7204,N_6503,N_6438);
nor U7205 (N_7205,N_6281,N_6523);
nor U7206 (N_7206,N_6822,N_6638);
nand U7207 (N_7207,N_6351,N_6530);
and U7208 (N_7208,N_6623,N_6472);
or U7209 (N_7209,N_6358,N_6830);
or U7210 (N_7210,N_6475,N_6365);
nand U7211 (N_7211,N_6485,N_6694);
xor U7212 (N_7212,N_6584,N_6823);
or U7213 (N_7213,N_6348,N_6851);
or U7214 (N_7214,N_6721,N_6834);
or U7215 (N_7215,N_6711,N_6418);
xnor U7216 (N_7216,N_6264,N_6670);
xor U7217 (N_7217,N_6304,N_6739);
nand U7218 (N_7218,N_6508,N_6544);
xnor U7219 (N_7219,N_6306,N_6329);
or U7220 (N_7220,N_6774,N_6294);
xnor U7221 (N_7221,N_6814,N_6624);
xor U7222 (N_7222,N_6731,N_6342);
or U7223 (N_7223,N_6685,N_6405);
xor U7224 (N_7224,N_6831,N_6796);
and U7225 (N_7225,N_6442,N_6268);
or U7226 (N_7226,N_6540,N_6817);
xnor U7227 (N_7227,N_6681,N_6497);
or U7228 (N_7228,N_6520,N_6828);
and U7229 (N_7229,N_6686,N_6351);
and U7230 (N_7230,N_6400,N_6485);
nor U7231 (N_7231,N_6844,N_6421);
and U7232 (N_7232,N_6596,N_6538);
xnor U7233 (N_7233,N_6762,N_6391);
nand U7234 (N_7234,N_6494,N_6400);
or U7235 (N_7235,N_6574,N_6638);
xnor U7236 (N_7236,N_6530,N_6639);
or U7237 (N_7237,N_6678,N_6613);
and U7238 (N_7238,N_6357,N_6579);
xor U7239 (N_7239,N_6808,N_6681);
nor U7240 (N_7240,N_6497,N_6462);
and U7241 (N_7241,N_6332,N_6615);
or U7242 (N_7242,N_6677,N_6571);
and U7243 (N_7243,N_6522,N_6261);
xor U7244 (N_7244,N_6429,N_6836);
or U7245 (N_7245,N_6695,N_6551);
and U7246 (N_7246,N_6392,N_6469);
or U7247 (N_7247,N_6701,N_6544);
nor U7248 (N_7248,N_6395,N_6465);
nor U7249 (N_7249,N_6322,N_6811);
nor U7250 (N_7250,N_6370,N_6589);
and U7251 (N_7251,N_6807,N_6397);
nor U7252 (N_7252,N_6346,N_6744);
and U7253 (N_7253,N_6439,N_6732);
nor U7254 (N_7254,N_6572,N_6570);
nor U7255 (N_7255,N_6252,N_6397);
xnor U7256 (N_7256,N_6367,N_6739);
nor U7257 (N_7257,N_6854,N_6644);
nand U7258 (N_7258,N_6850,N_6661);
and U7259 (N_7259,N_6436,N_6547);
or U7260 (N_7260,N_6853,N_6441);
xnor U7261 (N_7261,N_6251,N_6585);
nor U7262 (N_7262,N_6623,N_6424);
and U7263 (N_7263,N_6824,N_6805);
xor U7264 (N_7264,N_6698,N_6474);
and U7265 (N_7265,N_6638,N_6730);
xnor U7266 (N_7266,N_6840,N_6709);
nand U7267 (N_7267,N_6361,N_6348);
or U7268 (N_7268,N_6765,N_6850);
nor U7269 (N_7269,N_6688,N_6297);
nand U7270 (N_7270,N_6577,N_6849);
nor U7271 (N_7271,N_6479,N_6467);
nand U7272 (N_7272,N_6320,N_6481);
nand U7273 (N_7273,N_6684,N_6651);
xor U7274 (N_7274,N_6558,N_6519);
nand U7275 (N_7275,N_6561,N_6579);
nand U7276 (N_7276,N_6550,N_6825);
or U7277 (N_7277,N_6523,N_6624);
or U7278 (N_7278,N_6297,N_6787);
or U7279 (N_7279,N_6501,N_6617);
and U7280 (N_7280,N_6345,N_6528);
nor U7281 (N_7281,N_6702,N_6731);
nor U7282 (N_7282,N_6565,N_6340);
nand U7283 (N_7283,N_6478,N_6512);
nor U7284 (N_7284,N_6492,N_6559);
nand U7285 (N_7285,N_6345,N_6687);
or U7286 (N_7286,N_6483,N_6437);
xor U7287 (N_7287,N_6564,N_6528);
and U7288 (N_7288,N_6801,N_6624);
nor U7289 (N_7289,N_6399,N_6501);
nor U7290 (N_7290,N_6343,N_6624);
nor U7291 (N_7291,N_6645,N_6421);
nor U7292 (N_7292,N_6816,N_6324);
nand U7293 (N_7293,N_6498,N_6519);
nor U7294 (N_7294,N_6564,N_6677);
nand U7295 (N_7295,N_6866,N_6826);
xnor U7296 (N_7296,N_6710,N_6614);
or U7297 (N_7297,N_6396,N_6364);
nor U7298 (N_7298,N_6767,N_6637);
or U7299 (N_7299,N_6793,N_6295);
and U7300 (N_7300,N_6788,N_6775);
nor U7301 (N_7301,N_6710,N_6396);
and U7302 (N_7302,N_6574,N_6380);
xnor U7303 (N_7303,N_6374,N_6864);
xnor U7304 (N_7304,N_6309,N_6320);
nor U7305 (N_7305,N_6814,N_6807);
xor U7306 (N_7306,N_6809,N_6354);
or U7307 (N_7307,N_6429,N_6755);
or U7308 (N_7308,N_6424,N_6463);
and U7309 (N_7309,N_6647,N_6273);
nand U7310 (N_7310,N_6466,N_6258);
xor U7311 (N_7311,N_6807,N_6655);
xnor U7312 (N_7312,N_6252,N_6510);
nor U7313 (N_7313,N_6361,N_6778);
nor U7314 (N_7314,N_6715,N_6410);
or U7315 (N_7315,N_6759,N_6251);
xnor U7316 (N_7316,N_6269,N_6304);
and U7317 (N_7317,N_6822,N_6797);
xor U7318 (N_7318,N_6728,N_6322);
xor U7319 (N_7319,N_6414,N_6640);
nor U7320 (N_7320,N_6254,N_6380);
nor U7321 (N_7321,N_6256,N_6375);
and U7322 (N_7322,N_6790,N_6306);
nand U7323 (N_7323,N_6314,N_6363);
and U7324 (N_7324,N_6490,N_6568);
and U7325 (N_7325,N_6301,N_6631);
xor U7326 (N_7326,N_6407,N_6440);
nand U7327 (N_7327,N_6573,N_6686);
nor U7328 (N_7328,N_6527,N_6744);
nor U7329 (N_7329,N_6830,N_6847);
nand U7330 (N_7330,N_6854,N_6250);
nand U7331 (N_7331,N_6460,N_6549);
nor U7332 (N_7332,N_6799,N_6277);
and U7333 (N_7333,N_6787,N_6428);
and U7334 (N_7334,N_6667,N_6571);
or U7335 (N_7335,N_6833,N_6596);
nand U7336 (N_7336,N_6757,N_6786);
and U7337 (N_7337,N_6265,N_6504);
xor U7338 (N_7338,N_6809,N_6335);
and U7339 (N_7339,N_6312,N_6588);
xor U7340 (N_7340,N_6528,N_6701);
nor U7341 (N_7341,N_6610,N_6372);
or U7342 (N_7342,N_6529,N_6469);
xnor U7343 (N_7343,N_6685,N_6494);
and U7344 (N_7344,N_6575,N_6453);
xor U7345 (N_7345,N_6709,N_6809);
xor U7346 (N_7346,N_6408,N_6623);
or U7347 (N_7347,N_6740,N_6480);
nand U7348 (N_7348,N_6416,N_6828);
xor U7349 (N_7349,N_6461,N_6761);
or U7350 (N_7350,N_6357,N_6767);
and U7351 (N_7351,N_6434,N_6750);
and U7352 (N_7352,N_6351,N_6264);
or U7353 (N_7353,N_6724,N_6433);
xor U7354 (N_7354,N_6705,N_6753);
or U7355 (N_7355,N_6376,N_6458);
nand U7356 (N_7356,N_6450,N_6725);
xnor U7357 (N_7357,N_6566,N_6472);
or U7358 (N_7358,N_6648,N_6368);
xor U7359 (N_7359,N_6378,N_6751);
or U7360 (N_7360,N_6614,N_6670);
nand U7361 (N_7361,N_6720,N_6820);
nor U7362 (N_7362,N_6827,N_6385);
nor U7363 (N_7363,N_6760,N_6793);
xnor U7364 (N_7364,N_6527,N_6314);
nor U7365 (N_7365,N_6289,N_6739);
xor U7366 (N_7366,N_6712,N_6606);
nand U7367 (N_7367,N_6252,N_6540);
and U7368 (N_7368,N_6713,N_6668);
or U7369 (N_7369,N_6526,N_6734);
xor U7370 (N_7370,N_6314,N_6698);
nand U7371 (N_7371,N_6590,N_6309);
or U7372 (N_7372,N_6252,N_6261);
xor U7373 (N_7373,N_6806,N_6416);
nor U7374 (N_7374,N_6262,N_6594);
nor U7375 (N_7375,N_6355,N_6802);
or U7376 (N_7376,N_6480,N_6446);
or U7377 (N_7377,N_6798,N_6630);
nor U7378 (N_7378,N_6568,N_6772);
nor U7379 (N_7379,N_6304,N_6648);
or U7380 (N_7380,N_6517,N_6761);
nor U7381 (N_7381,N_6339,N_6299);
nor U7382 (N_7382,N_6419,N_6257);
xor U7383 (N_7383,N_6707,N_6797);
xnor U7384 (N_7384,N_6415,N_6610);
and U7385 (N_7385,N_6570,N_6712);
nand U7386 (N_7386,N_6440,N_6664);
nor U7387 (N_7387,N_6624,N_6492);
nand U7388 (N_7388,N_6332,N_6605);
xor U7389 (N_7389,N_6463,N_6655);
and U7390 (N_7390,N_6547,N_6712);
nand U7391 (N_7391,N_6286,N_6617);
nand U7392 (N_7392,N_6355,N_6323);
nor U7393 (N_7393,N_6312,N_6305);
or U7394 (N_7394,N_6824,N_6267);
nor U7395 (N_7395,N_6343,N_6687);
or U7396 (N_7396,N_6285,N_6358);
and U7397 (N_7397,N_6600,N_6264);
or U7398 (N_7398,N_6369,N_6774);
xnor U7399 (N_7399,N_6369,N_6286);
nor U7400 (N_7400,N_6687,N_6396);
nor U7401 (N_7401,N_6666,N_6559);
nor U7402 (N_7402,N_6727,N_6655);
xnor U7403 (N_7403,N_6579,N_6560);
or U7404 (N_7404,N_6710,N_6828);
or U7405 (N_7405,N_6756,N_6254);
or U7406 (N_7406,N_6494,N_6865);
and U7407 (N_7407,N_6610,N_6516);
nand U7408 (N_7408,N_6836,N_6388);
xnor U7409 (N_7409,N_6701,N_6646);
nand U7410 (N_7410,N_6633,N_6501);
or U7411 (N_7411,N_6369,N_6289);
or U7412 (N_7412,N_6676,N_6527);
or U7413 (N_7413,N_6791,N_6508);
nand U7414 (N_7414,N_6301,N_6291);
xor U7415 (N_7415,N_6737,N_6590);
or U7416 (N_7416,N_6847,N_6631);
nor U7417 (N_7417,N_6414,N_6622);
xnor U7418 (N_7418,N_6722,N_6719);
nand U7419 (N_7419,N_6521,N_6760);
or U7420 (N_7420,N_6505,N_6533);
nand U7421 (N_7421,N_6719,N_6467);
nor U7422 (N_7422,N_6525,N_6306);
nor U7423 (N_7423,N_6462,N_6528);
and U7424 (N_7424,N_6401,N_6763);
or U7425 (N_7425,N_6690,N_6327);
or U7426 (N_7426,N_6544,N_6717);
and U7427 (N_7427,N_6256,N_6857);
or U7428 (N_7428,N_6800,N_6567);
and U7429 (N_7429,N_6722,N_6818);
or U7430 (N_7430,N_6304,N_6396);
nor U7431 (N_7431,N_6431,N_6364);
nor U7432 (N_7432,N_6605,N_6497);
nor U7433 (N_7433,N_6441,N_6386);
nand U7434 (N_7434,N_6331,N_6308);
nor U7435 (N_7435,N_6522,N_6351);
and U7436 (N_7436,N_6381,N_6821);
and U7437 (N_7437,N_6762,N_6561);
xor U7438 (N_7438,N_6853,N_6808);
nand U7439 (N_7439,N_6761,N_6269);
nor U7440 (N_7440,N_6442,N_6260);
nor U7441 (N_7441,N_6694,N_6760);
or U7442 (N_7442,N_6485,N_6280);
xnor U7443 (N_7443,N_6650,N_6519);
xnor U7444 (N_7444,N_6806,N_6442);
and U7445 (N_7445,N_6284,N_6383);
nor U7446 (N_7446,N_6482,N_6331);
and U7447 (N_7447,N_6292,N_6744);
xor U7448 (N_7448,N_6655,N_6413);
xor U7449 (N_7449,N_6724,N_6858);
or U7450 (N_7450,N_6259,N_6795);
nand U7451 (N_7451,N_6619,N_6372);
nor U7452 (N_7452,N_6754,N_6678);
xor U7453 (N_7453,N_6655,N_6561);
xnor U7454 (N_7454,N_6425,N_6660);
nor U7455 (N_7455,N_6670,N_6517);
or U7456 (N_7456,N_6763,N_6833);
or U7457 (N_7457,N_6717,N_6344);
and U7458 (N_7458,N_6837,N_6514);
xor U7459 (N_7459,N_6534,N_6438);
xor U7460 (N_7460,N_6843,N_6372);
nor U7461 (N_7461,N_6432,N_6716);
nor U7462 (N_7462,N_6331,N_6442);
nor U7463 (N_7463,N_6601,N_6402);
nand U7464 (N_7464,N_6820,N_6652);
and U7465 (N_7465,N_6787,N_6597);
and U7466 (N_7466,N_6490,N_6445);
nand U7467 (N_7467,N_6421,N_6667);
nor U7468 (N_7468,N_6843,N_6381);
nand U7469 (N_7469,N_6666,N_6645);
xor U7470 (N_7470,N_6407,N_6430);
or U7471 (N_7471,N_6469,N_6633);
nand U7472 (N_7472,N_6792,N_6341);
or U7473 (N_7473,N_6286,N_6364);
or U7474 (N_7474,N_6814,N_6676);
or U7475 (N_7475,N_6816,N_6464);
nor U7476 (N_7476,N_6269,N_6858);
nor U7477 (N_7477,N_6362,N_6702);
xor U7478 (N_7478,N_6336,N_6293);
xnor U7479 (N_7479,N_6390,N_6430);
or U7480 (N_7480,N_6435,N_6268);
xor U7481 (N_7481,N_6843,N_6493);
xnor U7482 (N_7482,N_6454,N_6538);
nand U7483 (N_7483,N_6347,N_6384);
and U7484 (N_7484,N_6669,N_6754);
or U7485 (N_7485,N_6385,N_6594);
xnor U7486 (N_7486,N_6469,N_6756);
and U7487 (N_7487,N_6390,N_6442);
nand U7488 (N_7488,N_6489,N_6595);
or U7489 (N_7489,N_6625,N_6670);
nor U7490 (N_7490,N_6847,N_6602);
and U7491 (N_7491,N_6844,N_6793);
nor U7492 (N_7492,N_6830,N_6862);
nand U7493 (N_7493,N_6565,N_6373);
and U7494 (N_7494,N_6294,N_6751);
and U7495 (N_7495,N_6654,N_6528);
or U7496 (N_7496,N_6501,N_6553);
xnor U7497 (N_7497,N_6549,N_6588);
xnor U7498 (N_7498,N_6390,N_6306);
nand U7499 (N_7499,N_6583,N_6468);
and U7500 (N_7500,N_6958,N_6964);
and U7501 (N_7501,N_7125,N_6931);
or U7502 (N_7502,N_7313,N_7263);
and U7503 (N_7503,N_7484,N_7452);
nand U7504 (N_7504,N_7179,N_6970);
nor U7505 (N_7505,N_7436,N_6993);
and U7506 (N_7506,N_7060,N_7044);
or U7507 (N_7507,N_6979,N_7265);
nand U7508 (N_7508,N_7302,N_7098);
nand U7509 (N_7509,N_7339,N_7262);
and U7510 (N_7510,N_7204,N_7165);
nand U7511 (N_7511,N_6951,N_6942);
xor U7512 (N_7512,N_7326,N_7232);
and U7513 (N_7513,N_7161,N_7199);
nand U7514 (N_7514,N_7453,N_7107);
and U7515 (N_7515,N_6994,N_7249);
and U7516 (N_7516,N_7282,N_7402);
xor U7517 (N_7517,N_7206,N_7428);
or U7518 (N_7518,N_7145,N_7432);
or U7519 (N_7519,N_7186,N_7413);
and U7520 (N_7520,N_7260,N_7062);
or U7521 (N_7521,N_7029,N_6936);
nand U7522 (N_7522,N_6915,N_7219);
or U7523 (N_7523,N_7016,N_6880);
nand U7524 (N_7524,N_6896,N_7052);
nor U7525 (N_7525,N_6918,N_6925);
xor U7526 (N_7526,N_7374,N_7449);
nor U7527 (N_7527,N_7149,N_7036);
xnor U7528 (N_7528,N_7465,N_7459);
or U7529 (N_7529,N_7497,N_7009);
or U7530 (N_7530,N_6982,N_7401);
nor U7531 (N_7531,N_6984,N_7496);
or U7532 (N_7532,N_7142,N_7133);
xor U7533 (N_7533,N_7338,N_7247);
or U7534 (N_7534,N_7285,N_7064);
or U7535 (N_7535,N_7443,N_7456);
nand U7536 (N_7536,N_6893,N_7154);
and U7537 (N_7537,N_7377,N_7363);
nor U7538 (N_7538,N_7222,N_7234);
and U7539 (N_7539,N_7021,N_7121);
and U7540 (N_7540,N_7385,N_7430);
xor U7541 (N_7541,N_7201,N_7422);
xnor U7542 (N_7542,N_7472,N_7461);
xor U7543 (N_7543,N_7439,N_6988);
nor U7544 (N_7544,N_7137,N_6987);
nand U7545 (N_7545,N_7076,N_6971);
or U7546 (N_7546,N_7487,N_7254);
xnor U7547 (N_7547,N_7235,N_7323);
nand U7548 (N_7548,N_7210,N_6897);
and U7549 (N_7549,N_7274,N_6905);
and U7550 (N_7550,N_7304,N_6885);
nor U7551 (N_7551,N_7404,N_7388);
xnor U7552 (N_7552,N_7096,N_6883);
or U7553 (N_7553,N_7280,N_7160);
or U7554 (N_7554,N_7362,N_7191);
and U7555 (N_7555,N_7291,N_7094);
and U7556 (N_7556,N_7031,N_7354);
and U7557 (N_7557,N_6928,N_7015);
nor U7558 (N_7558,N_7104,N_7348);
or U7559 (N_7559,N_7175,N_7310);
nand U7560 (N_7560,N_6957,N_7469);
xnor U7561 (N_7561,N_7463,N_7039);
nor U7562 (N_7562,N_7103,N_7403);
nand U7563 (N_7563,N_7182,N_7256);
and U7564 (N_7564,N_7226,N_7306);
and U7565 (N_7565,N_6932,N_7297);
or U7566 (N_7566,N_6956,N_7307);
nand U7567 (N_7567,N_7337,N_7314);
nand U7568 (N_7568,N_7088,N_7146);
xor U7569 (N_7569,N_7067,N_6974);
xnor U7570 (N_7570,N_7136,N_7195);
nor U7571 (N_7571,N_7335,N_7084);
and U7572 (N_7572,N_7281,N_7118);
and U7573 (N_7573,N_7267,N_7395);
xnor U7574 (N_7574,N_7290,N_7305);
nand U7575 (N_7575,N_7066,N_7458);
xor U7576 (N_7576,N_7004,N_7320);
or U7577 (N_7577,N_7123,N_7375);
or U7578 (N_7578,N_7228,N_7457);
nand U7579 (N_7579,N_7030,N_7003);
and U7580 (N_7580,N_7147,N_7365);
and U7581 (N_7581,N_7358,N_7419);
nand U7582 (N_7582,N_7209,N_6935);
xor U7583 (N_7583,N_7196,N_7038);
and U7584 (N_7584,N_7057,N_7397);
or U7585 (N_7585,N_7392,N_7382);
xor U7586 (N_7586,N_7427,N_7440);
nand U7587 (N_7587,N_7387,N_6898);
and U7588 (N_7588,N_7061,N_7068);
nand U7589 (N_7589,N_7495,N_6913);
and U7590 (N_7590,N_7250,N_7026);
xor U7591 (N_7591,N_7370,N_7474);
xnor U7592 (N_7592,N_7217,N_7115);
or U7593 (N_7593,N_7318,N_7129);
or U7594 (N_7594,N_7001,N_7278);
nand U7595 (N_7595,N_7312,N_7159);
or U7596 (N_7596,N_7499,N_7489);
xor U7597 (N_7597,N_7223,N_7283);
or U7598 (N_7598,N_6947,N_7156);
and U7599 (N_7599,N_6991,N_6914);
nand U7600 (N_7600,N_7266,N_7086);
and U7601 (N_7601,N_6933,N_7135);
nor U7602 (N_7602,N_7153,N_6944);
nand U7603 (N_7603,N_7194,N_7355);
nor U7604 (N_7604,N_7212,N_7367);
nor U7605 (N_7605,N_7000,N_6976);
or U7606 (N_7606,N_6921,N_7255);
and U7607 (N_7607,N_7032,N_7272);
xor U7608 (N_7608,N_7188,N_7424);
and U7609 (N_7609,N_7231,N_6978);
xnor U7610 (N_7610,N_7099,N_7421);
nor U7611 (N_7611,N_7303,N_7378);
and U7612 (N_7612,N_6955,N_7239);
and U7613 (N_7613,N_7046,N_7479);
xor U7614 (N_7614,N_7264,N_6882);
nor U7615 (N_7615,N_7012,N_7193);
or U7616 (N_7616,N_7298,N_6980);
nand U7617 (N_7617,N_7414,N_7246);
or U7618 (N_7618,N_7309,N_7376);
xor U7619 (N_7619,N_7024,N_7043);
and U7620 (N_7620,N_7293,N_7328);
nand U7621 (N_7621,N_6878,N_7185);
nand U7622 (N_7622,N_6875,N_6884);
nand U7623 (N_7623,N_7073,N_7330);
or U7624 (N_7624,N_7221,N_7059);
nor U7625 (N_7625,N_7475,N_7399);
or U7626 (N_7626,N_7243,N_7183);
nor U7627 (N_7627,N_7360,N_7184);
xor U7628 (N_7628,N_7220,N_6940);
nand U7629 (N_7629,N_7148,N_7359);
nor U7630 (N_7630,N_6906,N_7117);
nand U7631 (N_7631,N_6975,N_7412);
and U7632 (N_7632,N_7049,N_7486);
xnor U7633 (N_7633,N_7132,N_7027);
nand U7634 (N_7634,N_7109,N_7070);
nor U7635 (N_7635,N_7242,N_7394);
xnor U7636 (N_7636,N_6895,N_7420);
xor U7637 (N_7637,N_6894,N_7287);
or U7638 (N_7638,N_7202,N_7130);
xor U7639 (N_7639,N_7172,N_6888);
nand U7640 (N_7640,N_7106,N_6946);
and U7641 (N_7641,N_7433,N_6900);
and U7642 (N_7642,N_7451,N_7295);
nand U7643 (N_7643,N_7013,N_7341);
and U7644 (N_7644,N_7299,N_6962);
nor U7645 (N_7645,N_7467,N_7416);
xor U7646 (N_7646,N_7418,N_7442);
nor U7647 (N_7647,N_6989,N_7319);
xnor U7648 (N_7648,N_6889,N_7390);
and U7649 (N_7649,N_7425,N_7331);
or U7650 (N_7650,N_7100,N_7380);
or U7651 (N_7651,N_7005,N_7462);
and U7652 (N_7652,N_7493,N_7482);
and U7653 (N_7653,N_7491,N_7108);
nand U7654 (N_7654,N_7476,N_7327);
nand U7655 (N_7655,N_7151,N_6903);
and U7656 (N_7656,N_6899,N_7460);
and U7657 (N_7657,N_7152,N_7090);
or U7658 (N_7658,N_7478,N_6972);
or U7659 (N_7659,N_6939,N_7273);
or U7660 (N_7660,N_7240,N_6967);
nor U7661 (N_7661,N_7011,N_6959);
xor U7662 (N_7662,N_6919,N_7321);
and U7663 (N_7663,N_7350,N_7227);
nand U7664 (N_7664,N_7138,N_6920);
nand U7665 (N_7665,N_7400,N_7468);
xor U7666 (N_7666,N_7325,N_7054);
nor U7667 (N_7667,N_7238,N_7368);
nor U7668 (N_7668,N_7237,N_7028);
nor U7669 (N_7669,N_7444,N_6965);
nor U7670 (N_7670,N_7371,N_7033);
xor U7671 (N_7671,N_7271,N_6999);
nand U7672 (N_7672,N_7494,N_7177);
nor U7673 (N_7673,N_7055,N_7174);
nand U7674 (N_7674,N_6886,N_7448);
or U7675 (N_7675,N_7200,N_7351);
nor U7676 (N_7676,N_7071,N_7480);
and U7677 (N_7677,N_7216,N_7346);
nand U7678 (N_7678,N_7379,N_7253);
nor U7679 (N_7679,N_7155,N_7065);
nand U7680 (N_7680,N_7035,N_6943);
xor U7681 (N_7681,N_7329,N_7268);
nor U7682 (N_7682,N_7447,N_7381);
xor U7683 (N_7683,N_7431,N_6937);
nand U7684 (N_7684,N_7292,N_7023);
nor U7685 (N_7685,N_7257,N_6997);
or U7686 (N_7686,N_7372,N_7214);
and U7687 (N_7687,N_6952,N_7356);
xor U7688 (N_7688,N_7483,N_7006);
xor U7689 (N_7689,N_6910,N_7207);
or U7690 (N_7690,N_6983,N_7466);
xor U7691 (N_7691,N_6926,N_7112);
or U7692 (N_7692,N_7241,N_7008);
or U7693 (N_7693,N_7485,N_7294);
or U7694 (N_7694,N_7042,N_6968);
or U7695 (N_7695,N_7077,N_7208);
nand U7696 (N_7696,N_7127,N_7258);
or U7697 (N_7697,N_6995,N_7124);
or U7698 (N_7698,N_7316,N_7353);
and U7699 (N_7699,N_7007,N_7270);
nor U7700 (N_7700,N_7276,N_7284);
xnor U7701 (N_7701,N_7091,N_7162);
xnor U7702 (N_7702,N_7446,N_7308);
nor U7703 (N_7703,N_6901,N_7245);
xnor U7704 (N_7704,N_7192,N_7322);
or U7705 (N_7705,N_7079,N_6960);
nand U7706 (N_7706,N_7190,N_7010);
nor U7707 (N_7707,N_7187,N_7141);
nand U7708 (N_7708,N_7301,N_6927);
xnor U7709 (N_7709,N_7063,N_7464);
and U7710 (N_7710,N_7315,N_7383);
and U7711 (N_7711,N_7047,N_6973);
nor U7712 (N_7712,N_7170,N_7289);
nand U7713 (N_7713,N_6923,N_7101);
xor U7714 (N_7714,N_7014,N_6966);
nor U7715 (N_7715,N_7020,N_7134);
nand U7716 (N_7716,N_7423,N_7164);
and U7717 (N_7717,N_7143,N_7334);
and U7718 (N_7718,N_7120,N_7211);
and U7719 (N_7719,N_7229,N_7150);
and U7720 (N_7720,N_6981,N_7048);
xnor U7721 (N_7721,N_6887,N_6953);
xor U7722 (N_7722,N_7342,N_7252);
nor U7723 (N_7723,N_7105,N_6916);
xor U7724 (N_7724,N_6924,N_7018);
nand U7725 (N_7725,N_7345,N_6890);
or U7726 (N_7726,N_7083,N_7311);
xor U7727 (N_7727,N_7089,N_7167);
and U7728 (N_7728,N_6961,N_7261);
or U7729 (N_7729,N_7198,N_7369);
or U7730 (N_7730,N_7408,N_7471);
and U7731 (N_7731,N_7169,N_6881);
nand U7732 (N_7732,N_7181,N_7116);
xnor U7733 (N_7733,N_7441,N_7366);
or U7734 (N_7734,N_6990,N_7340);
xor U7735 (N_7735,N_6908,N_7128);
xnor U7736 (N_7736,N_7095,N_7407);
xnor U7737 (N_7737,N_7352,N_7473);
nor U7738 (N_7738,N_7236,N_7180);
and U7739 (N_7739,N_7417,N_7126);
xnor U7740 (N_7740,N_7275,N_6929);
nor U7741 (N_7741,N_7470,N_7178);
xor U7742 (N_7742,N_7102,N_6912);
nand U7743 (N_7743,N_7435,N_7317);
or U7744 (N_7744,N_7455,N_7288);
nand U7745 (N_7745,N_7157,N_7454);
or U7746 (N_7746,N_6998,N_7398);
and U7747 (N_7747,N_7437,N_7045);
or U7748 (N_7748,N_7140,N_7093);
nand U7749 (N_7749,N_7041,N_7173);
nand U7750 (N_7750,N_7230,N_7080);
xnor U7751 (N_7751,N_7110,N_7279);
and U7752 (N_7752,N_7072,N_7384);
nor U7753 (N_7753,N_7171,N_7078);
nor U7754 (N_7754,N_6877,N_7324);
nor U7755 (N_7755,N_7373,N_7344);
xnor U7756 (N_7756,N_7248,N_6909);
xor U7757 (N_7757,N_7176,N_6902);
xor U7758 (N_7758,N_6934,N_7224);
and U7759 (N_7759,N_7144,N_7019);
and U7760 (N_7760,N_7445,N_6904);
nand U7761 (N_7761,N_7111,N_7034);
nand U7762 (N_7762,N_7166,N_7051);
or U7763 (N_7763,N_6891,N_7197);
and U7764 (N_7764,N_7058,N_7336);
nand U7765 (N_7765,N_7244,N_7259);
and U7766 (N_7766,N_7410,N_7218);
xor U7767 (N_7767,N_7251,N_7347);
and U7768 (N_7768,N_7233,N_7409);
or U7769 (N_7769,N_7277,N_7332);
and U7770 (N_7770,N_6911,N_7393);
xnor U7771 (N_7771,N_6969,N_7488);
nor U7772 (N_7772,N_6985,N_6876);
or U7773 (N_7773,N_6892,N_7406);
nand U7774 (N_7774,N_6879,N_7364);
and U7775 (N_7775,N_7429,N_7343);
xnor U7776 (N_7776,N_7037,N_7203);
or U7777 (N_7777,N_7411,N_7396);
xnor U7778 (N_7778,N_7349,N_7168);
and U7779 (N_7779,N_7492,N_7300);
or U7780 (N_7780,N_7391,N_7056);
or U7781 (N_7781,N_7481,N_7426);
xnor U7782 (N_7782,N_7002,N_7163);
xor U7783 (N_7783,N_7017,N_7040);
nand U7784 (N_7784,N_7081,N_6954);
and U7785 (N_7785,N_7205,N_6996);
nor U7786 (N_7786,N_7069,N_7082);
xor U7787 (N_7787,N_7092,N_7415);
or U7788 (N_7788,N_6963,N_6930);
nor U7789 (N_7789,N_7333,N_6950);
and U7790 (N_7790,N_7286,N_6949);
or U7791 (N_7791,N_7074,N_7097);
and U7792 (N_7792,N_7022,N_7386);
xor U7793 (N_7793,N_7269,N_6917);
xnor U7794 (N_7794,N_6945,N_7477);
or U7795 (N_7795,N_7296,N_7119);
or U7796 (N_7796,N_7113,N_7053);
or U7797 (N_7797,N_7498,N_7139);
or U7798 (N_7798,N_7189,N_7434);
xnor U7799 (N_7799,N_6922,N_7025);
nor U7800 (N_7800,N_7225,N_7122);
xnor U7801 (N_7801,N_7389,N_7075);
nor U7802 (N_7802,N_7450,N_7361);
or U7803 (N_7803,N_7490,N_6941);
and U7804 (N_7804,N_7357,N_7213);
nand U7805 (N_7805,N_7114,N_6977);
nand U7806 (N_7806,N_7050,N_6938);
or U7807 (N_7807,N_6948,N_7087);
nand U7808 (N_7808,N_6907,N_7158);
nor U7809 (N_7809,N_7085,N_6986);
xnor U7810 (N_7810,N_7215,N_7438);
nand U7811 (N_7811,N_7131,N_6992);
nor U7812 (N_7812,N_7405,N_7191);
xor U7813 (N_7813,N_7001,N_7437);
and U7814 (N_7814,N_7406,N_6921);
and U7815 (N_7815,N_7456,N_7375);
nor U7816 (N_7816,N_7484,N_7256);
xor U7817 (N_7817,N_7043,N_7285);
xor U7818 (N_7818,N_7000,N_7243);
and U7819 (N_7819,N_6876,N_7083);
nor U7820 (N_7820,N_7387,N_7010);
xor U7821 (N_7821,N_7159,N_7414);
or U7822 (N_7822,N_6886,N_7089);
nor U7823 (N_7823,N_6876,N_7448);
xor U7824 (N_7824,N_7217,N_7423);
nor U7825 (N_7825,N_7319,N_7343);
xnor U7826 (N_7826,N_6894,N_7368);
xor U7827 (N_7827,N_6998,N_7061);
or U7828 (N_7828,N_7414,N_7207);
and U7829 (N_7829,N_7460,N_7215);
xnor U7830 (N_7830,N_7400,N_6950);
xor U7831 (N_7831,N_7184,N_7172);
nand U7832 (N_7832,N_7236,N_7270);
xor U7833 (N_7833,N_7214,N_7101);
xor U7834 (N_7834,N_7379,N_6999);
or U7835 (N_7835,N_7232,N_6985);
and U7836 (N_7836,N_7118,N_7141);
xor U7837 (N_7837,N_6965,N_7127);
or U7838 (N_7838,N_7050,N_6916);
nand U7839 (N_7839,N_7055,N_7129);
nand U7840 (N_7840,N_6974,N_7296);
or U7841 (N_7841,N_7148,N_7020);
nand U7842 (N_7842,N_7038,N_6909);
nand U7843 (N_7843,N_6949,N_7238);
nor U7844 (N_7844,N_7493,N_7012);
nor U7845 (N_7845,N_7416,N_7076);
nand U7846 (N_7846,N_7153,N_7305);
nor U7847 (N_7847,N_6938,N_7245);
nor U7848 (N_7848,N_6967,N_6905);
xor U7849 (N_7849,N_7072,N_6980);
or U7850 (N_7850,N_7104,N_7014);
or U7851 (N_7851,N_7009,N_7294);
xor U7852 (N_7852,N_7246,N_7424);
xnor U7853 (N_7853,N_7475,N_7079);
nor U7854 (N_7854,N_7489,N_6927);
and U7855 (N_7855,N_7107,N_7387);
and U7856 (N_7856,N_7059,N_7143);
xor U7857 (N_7857,N_7220,N_7239);
and U7858 (N_7858,N_7141,N_7168);
xor U7859 (N_7859,N_6937,N_7241);
nand U7860 (N_7860,N_7437,N_7428);
nor U7861 (N_7861,N_7142,N_7087);
or U7862 (N_7862,N_7209,N_7353);
xor U7863 (N_7863,N_7319,N_6902);
xor U7864 (N_7864,N_6916,N_7418);
nand U7865 (N_7865,N_7485,N_7256);
nand U7866 (N_7866,N_6938,N_7308);
nand U7867 (N_7867,N_6958,N_7081);
and U7868 (N_7868,N_7004,N_7131);
or U7869 (N_7869,N_7438,N_6953);
and U7870 (N_7870,N_7325,N_6949);
or U7871 (N_7871,N_6987,N_7252);
nand U7872 (N_7872,N_6993,N_7292);
nor U7873 (N_7873,N_7494,N_7469);
or U7874 (N_7874,N_7388,N_7044);
and U7875 (N_7875,N_7202,N_7149);
nor U7876 (N_7876,N_7264,N_6904);
nand U7877 (N_7877,N_7205,N_7480);
xor U7878 (N_7878,N_7086,N_7226);
xnor U7879 (N_7879,N_7169,N_7052);
nand U7880 (N_7880,N_7426,N_7205);
or U7881 (N_7881,N_7302,N_7365);
and U7882 (N_7882,N_7092,N_7485);
nor U7883 (N_7883,N_7261,N_7398);
nand U7884 (N_7884,N_7333,N_7105);
nand U7885 (N_7885,N_6951,N_7414);
nand U7886 (N_7886,N_6934,N_7235);
nor U7887 (N_7887,N_7026,N_7459);
and U7888 (N_7888,N_7400,N_7173);
and U7889 (N_7889,N_6930,N_7482);
and U7890 (N_7890,N_7495,N_6932);
nor U7891 (N_7891,N_7068,N_7283);
xor U7892 (N_7892,N_7035,N_6997);
nor U7893 (N_7893,N_7052,N_7441);
nand U7894 (N_7894,N_7135,N_7270);
nand U7895 (N_7895,N_7124,N_7095);
or U7896 (N_7896,N_6883,N_7451);
or U7897 (N_7897,N_7034,N_6919);
nor U7898 (N_7898,N_7420,N_6964);
or U7899 (N_7899,N_7163,N_7032);
or U7900 (N_7900,N_7065,N_7425);
nor U7901 (N_7901,N_6928,N_7428);
or U7902 (N_7902,N_7468,N_7481);
nand U7903 (N_7903,N_7417,N_7117);
or U7904 (N_7904,N_7394,N_7431);
nand U7905 (N_7905,N_7125,N_6941);
nor U7906 (N_7906,N_7339,N_7395);
xor U7907 (N_7907,N_7258,N_7181);
xnor U7908 (N_7908,N_7297,N_7244);
nand U7909 (N_7909,N_7137,N_7242);
and U7910 (N_7910,N_7465,N_7385);
nand U7911 (N_7911,N_7489,N_7032);
nor U7912 (N_7912,N_7223,N_7060);
or U7913 (N_7913,N_7437,N_7144);
xor U7914 (N_7914,N_6953,N_7471);
or U7915 (N_7915,N_7407,N_7159);
or U7916 (N_7916,N_6899,N_7009);
and U7917 (N_7917,N_7145,N_7487);
or U7918 (N_7918,N_6961,N_7493);
nand U7919 (N_7919,N_7467,N_7076);
nand U7920 (N_7920,N_7443,N_7464);
nor U7921 (N_7921,N_7487,N_7341);
nor U7922 (N_7922,N_7000,N_7018);
xnor U7923 (N_7923,N_7226,N_7450);
nor U7924 (N_7924,N_7129,N_7436);
or U7925 (N_7925,N_6943,N_6907);
nand U7926 (N_7926,N_7462,N_6900);
nand U7927 (N_7927,N_6973,N_7234);
and U7928 (N_7928,N_7086,N_7280);
xnor U7929 (N_7929,N_6971,N_7133);
nand U7930 (N_7930,N_7454,N_7160);
and U7931 (N_7931,N_7382,N_6993);
and U7932 (N_7932,N_6911,N_7050);
and U7933 (N_7933,N_7134,N_7236);
nand U7934 (N_7934,N_7105,N_6881);
or U7935 (N_7935,N_7033,N_7423);
nor U7936 (N_7936,N_6950,N_6903);
xnor U7937 (N_7937,N_6940,N_7094);
and U7938 (N_7938,N_7131,N_7438);
and U7939 (N_7939,N_7237,N_7033);
xnor U7940 (N_7940,N_7408,N_7135);
and U7941 (N_7941,N_6922,N_7460);
nand U7942 (N_7942,N_7021,N_7145);
or U7943 (N_7943,N_6983,N_7050);
and U7944 (N_7944,N_6982,N_6956);
xor U7945 (N_7945,N_7023,N_7249);
xnor U7946 (N_7946,N_7050,N_7439);
nor U7947 (N_7947,N_7033,N_6898);
nand U7948 (N_7948,N_7362,N_7456);
or U7949 (N_7949,N_7233,N_7068);
nor U7950 (N_7950,N_7474,N_7074);
nor U7951 (N_7951,N_7108,N_6988);
nand U7952 (N_7952,N_6945,N_6973);
and U7953 (N_7953,N_7215,N_7146);
nand U7954 (N_7954,N_7088,N_7262);
and U7955 (N_7955,N_7085,N_7320);
and U7956 (N_7956,N_7052,N_6966);
nand U7957 (N_7957,N_7308,N_7173);
nor U7958 (N_7958,N_6888,N_6928);
xor U7959 (N_7959,N_7305,N_6940);
and U7960 (N_7960,N_6896,N_7425);
nand U7961 (N_7961,N_7240,N_7494);
xnor U7962 (N_7962,N_7475,N_7396);
nand U7963 (N_7963,N_7485,N_7352);
nor U7964 (N_7964,N_7016,N_7236);
nand U7965 (N_7965,N_6941,N_7264);
xor U7966 (N_7966,N_7117,N_7013);
or U7967 (N_7967,N_7437,N_7132);
nor U7968 (N_7968,N_7061,N_7110);
and U7969 (N_7969,N_7490,N_7337);
xor U7970 (N_7970,N_6947,N_7358);
and U7971 (N_7971,N_7046,N_7424);
or U7972 (N_7972,N_7486,N_6946);
or U7973 (N_7973,N_7001,N_7075);
or U7974 (N_7974,N_7254,N_7441);
nor U7975 (N_7975,N_7074,N_6921);
and U7976 (N_7976,N_7142,N_7453);
or U7977 (N_7977,N_7316,N_7012);
nand U7978 (N_7978,N_6948,N_7459);
xnor U7979 (N_7979,N_7451,N_6947);
and U7980 (N_7980,N_6901,N_7276);
or U7981 (N_7981,N_7464,N_6914);
xnor U7982 (N_7982,N_6878,N_6875);
and U7983 (N_7983,N_6945,N_7389);
xnor U7984 (N_7984,N_7496,N_6919);
or U7985 (N_7985,N_7456,N_7312);
xor U7986 (N_7986,N_7329,N_7001);
xor U7987 (N_7987,N_7276,N_7440);
and U7988 (N_7988,N_6936,N_7062);
nand U7989 (N_7989,N_6937,N_7323);
and U7990 (N_7990,N_6877,N_7291);
nand U7991 (N_7991,N_7065,N_6960);
xnor U7992 (N_7992,N_6934,N_7272);
or U7993 (N_7993,N_7013,N_6988);
nor U7994 (N_7994,N_7099,N_7370);
or U7995 (N_7995,N_6932,N_7461);
nor U7996 (N_7996,N_7120,N_7311);
nor U7997 (N_7997,N_7190,N_7464);
nand U7998 (N_7998,N_7084,N_7183);
nand U7999 (N_7999,N_7295,N_6885);
nand U8000 (N_8000,N_6971,N_7273);
xor U8001 (N_8001,N_7475,N_7124);
or U8002 (N_8002,N_7002,N_7280);
nand U8003 (N_8003,N_7289,N_7032);
and U8004 (N_8004,N_7449,N_7360);
xnor U8005 (N_8005,N_7107,N_7390);
nor U8006 (N_8006,N_6938,N_7253);
and U8007 (N_8007,N_7168,N_7468);
or U8008 (N_8008,N_7480,N_7350);
nand U8009 (N_8009,N_7312,N_7332);
xnor U8010 (N_8010,N_7309,N_6913);
nor U8011 (N_8011,N_7005,N_6938);
or U8012 (N_8012,N_7079,N_7033);
nor U8013 (N_8013,N_7307,N_7463);
nand U8014 (N_8014,N_7477,N_6985);
xnor U8015 (N_8015,N_7479,N_7066);
nor U8016 (N_8016,N_7411,N_7471);
xor U8017 (N_8017,N_7444,N_7427);
xnor U8018 (N_8018,N_6992,N_7332);
or U8019 (N_8019,N_7305,N_7390);
or U8020 (N_8020,N_7402,N_6913);
or U8021 (N_8021,N_7121,N_6902);
xor U8022 (N_8022,N_7262,N_7031);
or U8023 (N_8023,N_7400,N_7089);
and U8024 (N_8024,N_6997,N_7092);
or U8025 (N_8025,N_7365,N_7497);
or U8026 (N_8026,N_7180,N_7082);
xor U8027 (N_8027,N_6897,N_7080);
nand U8028 (N_8028,N_7017,N_7182);
xnor U8029 (N_8029,N_6883,N_7469);
or U8030 (N_8030,N_7492,N_6998);
nand U8031 (N_8031,N_7484,N_7215);
and U8032 (N_8032,N_6911,N_6884);
nor U8033 (N_8033,N_7131,N_7228);
nand U8034 (N_8034,N_7143,N_7254);
xor U8035 (N_8035,N_7421,N_7353);
nor U8036 (N_8036,N_7051,N_6973);
or U8037 (N_8037,N_7493,N_6983);
or U8038 (N_8038,N_6942,N_7022);
or U8039 (N_8039,N_7112,N_7424);
nand U8040 (N_8040,N_7319,N_6908);
xor U8041 (N_8041,N_7223,N_7192);
or U8042 (N_8042,N_6950,N_7274);
and U8043 (N_8043,N_7456,N_7143);
or U8044 (N_8044,N_7453,N_6952);
nor U8045 (N_8045,N_7338,N_7224);
nand U8046 (N_8046,N_7010,N_6924);
nand U8047 (N_8047,N_7097,N_7481);
nor U8048 (N_8048,N_7154,N_7426);
xor U8049 (N_8049,N_7197,N_6992);
nand U8050 (N_8050,N_7463,N_6908);
and U8051 (N_8051,N_7246,N_7147);
xor U8052 (N_8052,N_7221,N_7110);
or U8053 (N_8053,N_6991,N_6961);
or U8054 (N_8054,N_7490,N_7371);
or U8055 (N_8055,N_7060,N_6994);
nor U8056 (N_8056,N_7044,N_6893);
xor U8057 (N_8057,N_7144,N_7301);
and U8058 (N_8058,N_7284,N_7044);
xor U8059 (N_8059,N_7143,N_7273);
nor U8060 (N_8060,N_7158,N_7392);
nand U8061 (N_8061,N_6894,N_6899);
or U8062 (N_8062,N_7499,N_7098);
or U8063 (N_8063,N_7216,N_7291);
or U8064 (N_8064,N_6943,N_7196);
nor U8065 (N_8065,N_7137,N_7176);
and U8066 (N_8066,N_7300,N_7189);
and U8067 (N_8067,N_7129,N_7120);
and U8068 (N_8068,N_7162,N_6953);
nor U8069 (N_8069,N_7456,N_7289);
nand U8070 (N_8070,N_7185,N_7318);
or U8071 (N_8071,N_7030,N_7255);
nand U8072 (N_8072,N_7135,N_7205);
nor U8073 (N_8073,N_7447,N_6875);
nand U8074 (N_8074,N_7063,N_7243);
nor U8075 (N_8075,N_6917,N_7233);
and U8076 (N_8076,N_7259,N_7058);
nand U8077 (N_8077,N_7166,N_7014);
xnor U8078 (N_8078,N_7152,N_6880);
xnor U8079 (N_8079,N_6944,N_6978);
xnor U8080 (N_8080,N_7472,N_7013);
xnor U8081 (N_8081,N_7270,N_7011);
nand U8082 (N_8082,N_7473,N_7150);
nor U8083 (N_8083,N_7060,N_7390);
or U8084 (N_8084,N_7274,N_7114);
nand U8085 (N_8085,N_7076,N_7256);
nor U8086 (N_8086,N_7465,N_7112);
and U8087 (N_8087,N_7112,N_7422);
nand U8088 (N_8088,N_7002,N_6940);
nor U8089 (N_8089,N_6925,N_7333);
nor U8090 (N_8090,N_7272,N_7300);
xor U8091 (N_8091,N_7442,N_6967);
and U8092 (N_8092,N_7447,N_7264);
nor U8093 (N_8093,N_7366,N_7205);
nor U8094 (N_8094,N_7151,N_6935);
xnor U8095 (N_8095,N_7477,N_7370);
and U8096 (N_8096,N_6936,N_7279);
xor U8097 (N_8097,N_7045,N_6962);
or U8098 (N_8098,N_7357,N_7008);
or U8099 (N_8099,N_7028,N_7264);
nor U8100 (N_8100,N_7302,N_7121);
xnor U8101 (N_8101,N_6988,N_7014);
xnor U8102 (N_8102,N_7408,N_7036);
or U8103 (N_8103,N_6933,N_7144);
nand U8104 (N_8104,N_6909,N_7429);
or U8105 (N_8105,N_7360,N_7125);
and U8106 (N_8106,N_6998,N_7128);
nor U8107 (N_8107,N_7053,N_7047);
nand U8108 (N_8108,N_7113,N_6911);
or U8109 (N_8109,N_7420,N_7244);
and U8110 (N_8110,N_7104,N_6950);
nor U8111 (N_8111,N_7100,N_6989);
and U8112 (N_8112,N_7061,N_6992);
nand U8113 (N_8113,N_7091,N_7380);
or U8114 (N_8114,N_7208,N_6902);
and U8115 (N_8115,N_7295,N_7072);
nor U8116 (N_8116,N_6963,N_6958);
nor U8117 (N_8117,N_7084,N_7359);
or U8118 (N_8118,N_7091,N_7370);
nor U8119 (N_8119,N_7429,N_7098);
or U8120 (N_8120,N_7234,N_6920);
and U8121 (N_8121,N_6956,N_7393);
or U8122 (N_8122,N_7164,N_7354);
nand U8123 (N_8123,N_7158,N_7141);
nand U8124 (N_8124,N_7204,N_7390);
or U8125 (N_8125,N_7958,N_7579);
or U8126 (N_8126,N_7697,N_7738);
nor U8127 (N_8127,N_7560,N_7720);
xnor U8128 (N_8128,N_7822,N_8011);
nand U8129 (N_8129,N_7522,N_7835);
nor U8130 (N_8130,N_7557,N_7563);
nand U8131 (N_8131,N_7675,N_7889);
and U8132 (N_8132,N_8034,N_7705);
nand U8133 (N_8133,N_7943,N_8001);
xor U8134 (N_8134,N_7649,N_8055);
or U8135 (N_8135,N_7722,N_7816);
xnor U8136 (N_8136,N_7575,N_7715);
xnor U8137 (N_8137,N_8060,N_7747);
and U8138 (N_8138,N_7809,N_7952);
nor U8139 (N_8139,N_7772,N_8020);
or U8140 (N_8140,N_7602,N_8022);
xnor U8141 (N_8141,N_7505,N_7581);
and U8142 (N_8142,N_7966,N_7696);
xnor U8143 (N_8143,N_7584,N_7815);
or U8144 (N_8144,N_8052,N_7867);
or U8145 (N_8145,N_7698,N_7871);
nand U8146 (N_8146,N_7704,N_7657);
nor U8147 (N_8147,N_7702,N_7920);
nand U8148 (N_8148,N_7725,N_7717);
and U8149 (N_8149,N_7700,N_8047);
or U8150 (N_8150,N_7787,N_7578);
nor U8151 (N_8151,N_7987,N_7903);
xnor U8152 (N_8152,N_7909,N_8117);
nand U8153 (N_8153,N_7979,N_8062);
nand U8154 (N_8154,N_7542,N_7617);
xnor U8155 (N_8155,N_7729,N_7518);
xor U8156 (N_8156,N_8100,N_7691);
or U8157 (N_8157,N_7667,N_7709);
and U8158 (N_8158,N_8096,N_7508);
nand U8159 (N_8159,N_7842,N_7912);
nand U8160 (N_8160,N_7841,N_7942);
or U8161 (N_8161,N_7670,N_7745);
nor U8162 (N_8162,N_8065,N_7976);
and U8163 (N_8163,N_7821,N_7862);
nor U8164 (N_8164,N_7733,N_7888);
xnor U8165 (N_8165,N_7727,N_7883);
and U8166 (N_8166,N_7805,N_7866);
nand U8167 (N_8167,N_7783,N_8012);
nand U8168 (N_8168,N_7760,N_7592);
nand U8169 (N_8169,N_7806,N_7568);
or U8170 (N_8170,N_7956,N_7734);
or U8171 (N_8171,N_7586,N_7895);
and U8172 (N_8172,N_8085,N_7807);
nand U8173 (N_8173,N_7984,N_7907);
or U8174 (N_8174,N_7863,N_7712);
and U8175 (N_8175,N_7758,N_7910);
nand U8176 (N_8176,N_7716,N_7762);
nor U8177 (N_8177,N_7925,N_7756);
nor U8178 (N_8178,N_7699,N_7547);
nand U8179 (N_8179,N_7701,N_7792);
nor U8180 (N_8180,N_7975,N_7678);
or U8181 (N_8181,N_8005,N_7711);
and U8182 (N_8182,N_7780,N_7744);
nand U8183 (N_8183,N_8109,N_7899);
xor U8184 (N_8184,N_7999,N_8120);
nor U8185 (N_8185,N_7961,N_7662);
xor U8186 (N_8186,N_7650,N_8045);
nand U8187 (N_8187,N_7605,N_7577);
nor U8188 (N_8188,N_7681,N_7730);
xor U8189 (N_8189,N_8110,N_7922);
xor U8190 (N_8190,N_8101,N_7726);
nand U8191 (N_8191,N_7924,N_8018);
and U8192 (N_8192,N_7601,N_7753);
or U8193 (N_8193,N_7990,N_7599);
or U8194 (N_8194,N_7520,N_7562);
xor U8195 (N_8195,N_7865,N_8030);
and U8196 (N_8196,N_7801,N_7763);
and U8197 (N_8197,N_8092,N_7752);
nand U8198 (N_8198,N_7668,N_7981);
xnor U8199 (N_8199,N_7860,N_7527);
nor U8200 (N_8200,N_7960,N_7974);
nand U8201 (N_8201,N_8032,N_7768);
nor U8202 (N_8202,N_7637,N_7513);
nor U8203 (N_8203,N_8112,N_7703);
nand U8204 (N_8204,N_7604,N_7555);
or U8205 (N_8205,N_7764,N_7582);
nand U8206 (N_8206,N_7838,N_7970);
xnor U8207 (N_8207,N_8048,N_8021);
and U8208 (N_8208,N_7785,N_7775);
xor U8209 (N_8209,N_7881,N_7595);
nand U8210 (N_8210,N_7916,N_8063);
or U8211 (N_8211,N_7629,N_8082);
nand U8212 (N_8212,N_8039,N_7671);
and U8213 (N_8213,N_7846,N_7968);
nand U8214 (N_8214,N_7507,N_7872);
xnor U8215 (N_8215,N_7625,N_7569);
nor U8216 (N_8216,N_7992,N_7635);
nand U8217 (N_8217,N_7985,N_7932);
nand U8218 (N_8218,N_7953,N_7611);
nand U8219 (N_8219,N_7906,N_7998);
xor U8220 (N_8220,N_8078,N_8114);
nor U8221 (N_8221,N_7831,N_8106);
and U8222 (N_8222,N_7535,N_8098);
nand U8223 (N_8223,N_7996,N_7844);
nor U8224 (N_8224,N_7501,N_7509);
and U8225 (N_8225,N_7918,N_7880);
and U8226 (N_8226,N_7882,N_7767);
or U8227 (N_8227,N_7761,N_7931);
and U8228 (N_8228,N_8076,N_7536);
or U8229 (N_8229,N_7944,N_7594);
nor U8230 (N_8230,N_7908,N_7828);
nor U8231 (N_8231,N_7973,N_7620);
nor U8232 (N_8232,N_7556,N_7718);
nand U8233 (N_8233,N_7825,N_8027);
and U8234 (N_8234,N_7759,N_8079);
or U8235 (N_8235,N_8091,N_8069);
and U8236 (N_8236,N_7870,N_7945);
nand U8237 (N_8237,N_8102,N_7837);
nor U8238 (N_8238,N_7660,N_7896);
nor U8239 (N_8239,N_7694,N_7814);
nor U8240 (N_8240,N_7724,N_7706);
nand U8241 (N_8241,N_8004,N_7829);
nor U8242 (N_8242,N_8040,N_8046);
nor U8243 (N_8243,N_8073,N_7754);
xnor U8244 (N_8244,N_8086,N_7797);
and U8245 (N_8245,N_7927,N_7651);
and U8246 (N_8246,N_7677,N_7731);
nor U8247 (N_8247,N_7827,N_7962);
nand U8248 (N_8248,N_7955,N_7877);
and U8249 (N_8249,N_7641,N_7665);
and U8250 (N_8250,N_7644,N_8015);
nand U8251 (N_8251,N_7591,N_7868);
and U8252 (N_8252,N_7504,N_7969);
xor U8253 (N_8253,N_7566,N_7808);
nand U8254 (N_8254,N_7776,N_8084);
nand U8255 (N_8255,N_7603,N_7614);
nand U8256 (N_8256,N_7991,N_7989);
or U8257 (N_8257,N_7892,N_8075);
nand U8258 (N_8258,N_7978,N_7533);
xor U8259 (N_8259,N_7551,N_7583);
nor U8260 (N_8260,N_8000,N_7786);
xor U8261 (N_8261,N_7771,N_7800);
nor U8262 (N_8262,N_8122,N_8087);
xnor U8263 (N_8263,N_8119,N_8095);
and U8264 (N_8264,N_7676,N_7654);
nand U8265 (N_8265,N_7859,N_8042);
nor U8266 (N_8266,N_7986,N_7755);
or U8267 (N_8267,N_8103,N_8029);
nor U8268 (N_8268,N_7830,N_7500);
xor U8269 (N_8269,N_7930,N_7549);
and U8270 (N_8270,N_7663,N_7933);
nor U8271 (N_8271,N_7820,N_7684);
xor U8272 (N_8272,N_8017,N_7541);
xor U8273 (N_8273,N_7512,N_7710);
nor U8274 (N_8274,N_7794,N_7689);
or U8275 (N_8275,N_8080,N_7803);
nand U8276 (N_8276,N_7652,N_7915);
and U8277 (N_8277,N_8024,N_7923);
or U8278 (N_8278,N_7648,N_8067);
or U8279 (N_8279,N_7534,N_8051);
nand U8280 (N_8280,N_7928,N_7564);
nor U8281 (N_8281,N_7964,N_8077);
nor U8282 (N_8282,N_7735,N_7610);
xor U8283 (N_8283,N_7972,N_7525);
and U8284 (N_8284,N_7799,N_7836);
or U8285 (N_8285,N_7897,N_8081);
nor U8286 (N_8286,N_7572,N_7538);
xnor U8287 (N_8287,N_7561,N_7823);
xnor U8288 (N_8288,N_7714,N_8070);
xor U8289 (N_8289,N_7951,N_7517);
nor U8290 (N_8290,N_7521,N_7887);
xor U8291 (N_8291,N_7587,N_7963);
nand U8292 (N_8292,N_7921,N_7749);
nand U8293 (N_8293,N_7732,N_7606);
nand U8294 (N_8294,N_8044,N_7742);
or U8295 (N_8295,N_8111,N_7570);
and U8296 (N_8296,N_7971,N_7664);
nor U8297 (N_8297,N_7626,N_7708);
nor U8298 (N_8298,N_7612,N_7632);
nand U8299 (N_8299,N_7545,N_7813);
nand U8300 (N_8300,N_7516,N_7719);
nor U8301 (N_8301,N_7798,N_8071);
nand U8302 (N_8302,N_7861,N_7739);
nor U8303 (N_8303,N_7589,N_7847);
xnor U8304 (N_8304,N_7674,N_7552);
xor U8305 (N_8305,N_8007,N_7543);
and U8306 (N_8306,N_7523,N_7598);
xnor U8307 (N_8307,N_7864,N_7938);
nor U8308 (N_8308,N_7936,N_8115);
and U8309 (N_8309,N_7893,N_7793);
nor U8310 (N_8310,N_7983,N_7688);
and U8311 (N_8311,N_7804,N_8053);
nand U8312 (N_8312,N_7519,N_7854);
and U8313 (N_8313,N_7687,N_8002);
and U8314 (N_8314,N_8033,N_7669);
or U8315 (N_8315,N_7642,N_7993);
and U8316 (N_8316,N_7879,N_7633);
xnor U8317 (N_8317,N_8118,N_7679);
or U8318 (N_8318,N_7634,N_7661);
xor U8319 (N_8319,N_7939,N_7843);
nand U8320 (N_8320,N_7950,N_8066);
and U8321 (N_8321,N_7567,N_7682);
nand U8322 (N_8322,N_7618,N_7796);
nor U8323 (N_8323,N_7802,N_8089);
or U8324 (N_8324,N_7834,N_7766);
and U8325 (N_8325,N_7548,N_7919);
nand U8326 (N_8326,N_7673,N_7851);
or U8327 (N_8327,N_7713,N_7997);
nor U8328 (N_8328,N_7672,N_8028);
xor U8329 (N_8329,N_8010,N_7636);
nor U8330 (N_8330,N_8061,N_8031);
xor U8331 (N_8331,N_7982,N_7839);
and U8332 (N_8332,N_7977,N_8038);
and U8333 (N_8333,N_7576,N_7593);
xor U8334 (N_8334,N_7511,N_7746);
xor U8335 (N_8335,N_7884,N_7631);
and U8336 (N_8336,N_7778,N_7779);
or U8337 (N_8337,N_8064,N_7741);
and U8338 (N_8338,N_7723,N_7869);
xor U8339 (N_8339,N_8019,N_7683);
or U8340 (N_8340,N_7905,N_7937);
xnor U8341 (N_8341,N_7740,N_7515);
xnor U8342 (N_8342,N_8088,N_8043);
and U8343 (N_8343,N_7911,N_7790);
nand U8344 (N_8344,N_8023,N_7812);
xnor U8345 (N_8345,N_8107,N_7935);
nor U8346 (N_8346,N_7934,N_7526);
nand U8347 (N_8347,N_7619,N_7539);
nor U8348 (N_8348,N_8108,N_7900);
xnor U8349 (N_8349,N_7693,N_7622);
xnor U8350 (N_8350,N_7954,N_7967);
nor U8351 (N_8351,N_7613,N_8083);
nor U8352 (N_8352,N_7597,N_7926);
nor U8353 (N_8353,N_7774,N_7600);
nor U8354 (N_8354,N_7546,N_8013);
and U8355 (N_8355,N_8003,N_8006);
nand U8356 (N_8356,N_7885,N_7558);
xor U8357 (N_8357,N_7524,N_8036);
xnor U8358 (N_8358,N_7947,N_7647);
and U8359 (N_8359,N_7994,N_7638);
and U8360 (N_8360,N_8054,N_8093);
or U8361 (N_8361,N_8099,N_7728);
xor U8362 (N_8362,N_7607,N_7721);
nor U8363 (N_8363,N_7686,N_7878);
or U8364 (N_8364,N_7643,N_8104);
nand U8365 (N_8365,N_7949,N_7856);
xnor U8366 (N_8366,N_8049,N_7503);
and U8367 (N_8367,N_8057,N_8008);
nand U8368 (N_8368,N_7781,N_7789);
nor U8369 (N_8369,N_7585,N_7750);
xnor U8370 (N_8370,N_7782,N_7890);
and U8371 (N_8371,N_7874,N_7628);
or U8372 (N_8372,N_8123,N_7692);
nand U8373 (N_8373,N_7737,N_7506);
nand U8374 (N_8374,N_7645,N_7659);
xnor U8375 (N_8375,N_7941,N_7588);
or U8376 (N_8376,N_7510,N_7914);
nand U8377 (N_8377,N_8116,N_7528);
xor U8378 (N_8378,N_7630,N_7819);
and U8379 (N_8379,N_7550,N_8035);
and U8380 (N_8380,N_8058,N_7876);
and U8381 (N_8381,N_7627,N_7609);
xor U8382 (N_8382,N_8113,N_7656);
or U8383 (N_8383,N_7574,N_7748);
xor U8384 (N_8384,N_7788,N_7653);
and U8385 (N_8385,N_7621,N_7743);
nor U8386 (N_8386,N_7777,N_7658);
or U8387 (N_8387,N_7769,N_7917);
and U8388 (N_8388,N_7615,N_7855);
nor U8389 (N_8389,N_8009,N_7554);
xor U8390 (N_8390,N_7810,N_8068);
nand U8391 (N_8391,N_8074,N_8026);
nand U8392 (N_8392,N_7655,N_8041);
xor U8393 (N_8393,N_7833,N_7573);
and U8394 (N_8394,N_8059,N_7824);
nor U8395 (N_8395,N_7646,N_7640);
nand U8396 (N_8396,N_7901,N_7832);
or U8397 (N_8397,N_8016,N_7680);
nand U8398 (N_8398,N_7571,N_7690);
and U8399 (N_8399,N_7580,N_8056);
xnor U8400 (N_8400,N_7530,N_8105);
nor U8401 (N_8401,N_8050,N_7529);
nor U8402 (N_8402,N_8072,N_7770);
and U8403 (N_8403,N_7590,N_7894);
xor U8404 (N_8404,N_7639,N_7565);
nor U8405 (N_8405,N_7898,N_7929);
xnor U8406 (N_8406,N_7904,N_7608);
xor U8407 (N_8407,N_7826,N_7791);
nand U8408 (N_8408,N_7988,N_7559);
nand U8409 (N_8409,N_7886,N_8014);
or U8410 (N_8410,N_7995,N_7616);
or U8411 (N_8411,N_7537,N_8094);
or U8412 (N_8412,N_7858,N_7959);
nand U8413 (N_8413,N_7624,N_7736);
and U8414 (N_8414,N_8090,N_7811);
and U8415 (N_8415,N_7623,N_7853);
or U8416 (N_8416,N_7875,N_7913);
or U8417 (N_8417,N_7852,N_8124);
nor U8418 (N_8418,N_7685,N_8121);
and U8419 (N_8419,N_7795,N_7818);
and U8420 (N_8420,N_7840,N_7845);
nor U8421 (N_8421,N_7502,N_7757);
and U8422 (N_8422,N_8037,N_7784);
and U8423 (N_8423,N_7817,N_7666);
xnor U8424 (N_8424,N_7531,N_7553);
and U8425 (N_8425,N_7540,N_7751);
nor U8426 (N_8426,N_8097,N_7848);
nor U8427 (N_8427,N_7946,N_7857);
and U8428 (N_8428,N_7957,N_7980);
nor U8429 (N_8429,N_7695,N_7544);
and U8430 (N_8430,N_7707,N_7765);
xor U8431 (N_8431,N_7940,N_7596);
or U8432 (N_8432,N_7891,N_8025);
nor U8433 (N_8433,N_7850,N_7965);
xor U8434 (N_8434,N_7514,N_7532);
and U8435 (N_8435,N_7948,N_7773);
nand U8436 (N_8436,N_7849,N_7902);
nand U8437 (N_8437,N_7873,N_7930);
nand U8438 (N_8438,N_7544,N_7806);
or U8439 (N_8439,N_7763,N_8018);
nand U8440 (N_8440,N_7795,N_7759);
nand U8441 (N_8441,N_8108,N_7681);
nor U8442 (N_8442,N_8115,N_7715);
nand U8443 (N_8443,N_7804,N_7658);
nand U8444 (N_8444,N_7770,N_7713);
or U8445 (N_8445,N_7827,N_7568);
nor U8446 (N_8446,N_7821,N_8075);
nand U8447 (N_8447,N_7940,N_7561);
or U8448 (N_8448,N_7796,N_8030);
nor U8449 (N_8449,N_7946,N_7549);
nand U8450 (N_8450,N_7873,N_7653);
and U8451 (N_8451,N_8102,N_7939);
nand U8452 (N_8452,N_8094,N_7959);
nand U8453 (N_8453,N_7576,N_7908);
and U8454 (N_8454,N_8050,N_7822);
or U8455 (N_8455,N_8084,N_7681);
nor U8456 (N_8456,N_7636,N_8072);
xnor U8457 (N_8457,N_7768,N_8080);
xor U8458 (N_8458,N_7780,N_7700);
and U8459 (N_8459,N_7551,N_7612);
xnor U8460 (N_8460,N_7879,N_7962);
and U8461 (N_8461,N_7514,N_7966);
and U8462 (N_8462,N_7625,N_7568);
and U8463 (N_8463,N_7861,N_8101);
nand U8464 (N_8464,N_7566,N_7853);
nor U8465 (N_8465,N_7531,N_8033);
or U8466 (N_8466,N_7541,N_7738);
nor U8467 (N_8467,N_7631,N_7680);
nor U8468 (N_8468,N_7765,N_7604);
and U8469 (N_8469,N_8081,N_7690);
or U8470 (N_8470,N_7818,N_7792);
nand U8471 (N_8471,N_7795,N_7741);
or U8472 (N_8472,N_7679,N_7558);
nand U8473 (N_8473,N_7542,N_7933);
xor U8474 (N_8474,N_7552,N_7810);
or U8475 (N_8475,N_7950,N_7987);
nand U8476 (N_8476,N_7663,N_7679);
nor U8477 (N_8477,N_7773,N_7837);
or U8478 (N_8478,N_7705,N_7935);
and U8479 (N_8479,N_8056,N_7563);
nand U8480 (N_8480,N_7910,N_7584);
and U8481 (N_8481,N_7532,N_7568);
or U8482 (N_8482,N_7974,N_8043);
nor U8483 (N_8483,N_7952,N_8020);
or U8484 (N_8484,N_7872,N_7935);
xor U8485 (N_8485,N_8066,N_8071);
and U8486 (N_8486,N_8032,N_8113);
and U8487 (N_8487,N_7997,N_8020);
nand U8488 (N_8488,N_7569,N_7630);
nand U8489 (N_8489,N_7571,N_7983);
nor U8490 (N_8490,N_7903,N_8060);
nand U8491 (N_8491,N_7902,N_7901);
xnor U8492 (N_8492,N_7746,N_7649);
nand U8493 (N_8493,N_7948,N_7838);
nor U8494 (N_8494,N_7705,N_8064);
nand U8495 (N_8495,N_7751,N_7904);
nand U8496 (N_8496,N_8082,N_7841);
nand U8497 (N_8497,N_7927,N_7938);
nor U8498 (N_8498,N_7836,N_8068);
and U8499 (N_8499,N_8022,N_8059);
or U8500 (N_8500,N_7501,N_7901);
or U8501 (N_8501,N_7538,N_7625);
and U8502 (N_8502,N_7848,N_7621);
xor U8503 (N_8503,N_7588,N_7707);
nand U8504 (N_8504,N_7654,N_7726);
or U8505 (N_8505,N_7530,N_7670);
and U8506 (N_8506,N_7941,N_7665);
and U8507 (N_8507,N_7692,N_7950);
nor U8508 (N_8508,N_7913,N_7666);
and U8509 (N_8509,N_7636,N_7917);
nor U8510 (N_8510,N_7828,N_7739);
nor U8511 (N_8511,N_7935,N_7794);
nor U8512 (N_8512,N_7553,N_8025);
nand U8513 (N_8513,N_7691,N_7609);
nand U8514 (N_8514,N_7747,N_7667);
nand U8515 (N_8515,N_7746,N_7718);
and U8516 (N_8516,N_8116,N_7583);
or U8517 (N_8517,N_8041,N_7895);
and U8518 (N_8518,N_7897,N_7564);
or U8519 (N_8519,N_7599,N_7831);
nor U8520 (N_8520,N_8020,N_7826);
and U8521 (N_8521,N_8038,N_7534);
nand U8522 (N_8522,N_7971,N_7743);
nand U8523 (N_8523,N_7944,N_7824);
nor U8524 (N_8524,N_7692,N_7670);
xnor U8525 (N_8525,N_7860,N_7889);
xor U8526 (N_8526,N_7959,N_7729);
or U8527 (N_8527,N_7974,N_7986);
xor U8528 (N_8528,N_7940,N_7521);
nor U8529 (N_8529,N_7660,N_7848);
xnor U8530 (N_8530,N_7763,N_8034);
nand U8531 (N_8531,N_7587,N_7929);
nor U8532 (N_8532,N_8096,N_8078);
xnor U8533 (N_8533,N_8015,N_7733);
and U8534 (N_8534,N_8048,N_7801);
and U8535 (N_8535,N_7719,N_7537);
and U8536 (N_8536,N_7866,N_7961);
xnor U8537 (N_8537,N_8095,N_8085);
or U8538 (N_8538,N_8001,N_8012);
nor U8539 (N_8539,N_7716,N_8076);
xnor U8540 (N_8540,N_7627,N_8000);
or U8541 (N_8541,N_7671,N_7980);
nand U8542 (N_8542,N_7821,N_8117);
nand U8543 (N_8543,N_7792,N_7692);
or U8544 (N_8544,N_7758,N_7512);
or U8545 (N_8545,N_7969,N_7781);
nand U8546 (N_8546,N_7961,N_7798);
or U8547 (N_8547,N_7631,N_7566);
xor U8548 (N_8548,N_7744,N_8027);
or U8549 (N_8549,N_7588,N_7580);
xor U8550 (N_8550,N_7674,N_8123);
and U8551 (N_8551,N_7568,N_8074);
nor U8552 (N_8552,N_7519,N_7767);
nand U8553 (N_8553,N_8095,N_7832);
xnor U8554 (N_8554,N_8098,N_8071);
nor U8555 (N_8555,N_7939,N_7934);
and U8556 (N_8556,N_7608,N_7708);
or U8557 (N_8557,N_7714,N_7742);
or U8558 (N_8558,N_7762,N_7893);
and U8559 (N_8559,N_7600,N_7976);
or U8560 (N_8560,N_7843,N_7742);
xor U8561 (N_8561,N_7976,N_7667);
nor U8562 (N_8562,N_7750,N_8064);
and U8563 (N_8563,N_8028,N_7519);
and U8564 (N_8564,N_7641,N_7850);
nor U8565 (N_8565,N_7896,N_7700);
and U8566 (N_8566,N_7793,N_7740);
or U8567 (N_8567,N_7577,N_7881);
xnor U8568 (N_8568,N_7618,N_7640);
nor U8569 (N_8569,N_7643,N_7724);
xnor U8570 (N_8570,N_8047,N_7718);
and U8571 (N_8571,N_7613,N_7524);
nor U8572 (N_8572,N_7769,N_7741);
or U8573 (N_8573,N_7666,N_7616);
xnor U8574 (N_8574,N_7808,N_7965);
nand U8575 (N_8575,N_7871,N_7504);
or U8576 (N_8576,N_7939,N_7970);
and U8577 (N_8577,N_7770,N_7989);
and U8578 (N_8578,N_7830,N_7709);
xnor U8579 (N_8579,N_7538,N_7629);
or U8580 (N_8580,N_7662,N_7550);
and U8581 (N_8581,N_7755,N_7942);
nor U8582 (N_8582,N_7914,N_7642);
xnor U8583 (N_8583,N_7746,N_7759);
or U8584 (N_8584,N_7563,N_7965);
or U8585 (N_8585,N_7676,N_8044);
nor U8586 (N_8586,N_7678,N_8112);
nor U8587 (N_8587,N_7547,N_8062);
and U8588 (N_8588,N_8095,N_7791);
nor U8589 (N_8589,N_7971,N_8024);
or U8590 (N_8590,N_7743,N_7591);
or U8591 (N_8591,N_7831,N_7510);
nand U8592 (N_8592,N_7570,N_7937);
and U8593 (N_8593,N_7806,N_7550);
xor U8594 (N_8594,N_7652,N_7699);
and U8595 (N_8595,N_8056,N_8071);
xnor U8596 (N_8596,N_7798,N_7785);
xor U8597 (N_8597,N_7505,N_7638);
nor U8598 (N_8598,N_8111,N_7884);
nand U8599 (N_8599,N_8012,N_8084);
and U8600 (N_8600,N_8066,N_7988);
nor U8601 (N_8601,N_7861,N_7675);
nand U8602 (N_8602,N_8000,N_8013);
xor U8603 (N_8603,N_7747,N_7742);
nand U8604 (N_8604,N_7550,N_7660);
and U8605 (N_8605,N_7714,N_7543);
nand U8606 (N_8606,N_7665,N_7742);
xnor U8607 (N_8607,N_8086,N_7811);
or U8608 (N_8608,N_7676,N_7997);
nand U8609 (N_8609,N_7833,N_7783);
nand U8610 (N_8610,N_8067,N_7825);
and U8611 (N_8611,N_7995,N_8059);
xnor U8612 (N_8612,N_7972,N_7512);
or U8613 (N_8613,N_7931,N_8117);
or U8614 (N_8614,N_7640,N_7623);
xor U8615 (N_8615,N_7939,N_8015);
xnor U8616 (N_8616,N_7762,N_8012);
and U8617 (N_8617,N_7652,N_8116);
xor U8618 (N_8618,N_7903,N_7562);
or U8619 (N_8619,N_7505,N_7550);
and U8620 (N_8620,N_7901,N_7506);
and U8621 (N_8621,N_7534,N_7883);
and U8622 (N_8622,N_7927,N_7683);
nor U8623 (N_8623,N_8065,N_7560);
and U8624 (N_8624,N_7521,N_8086);
nand U8625 (N_8625,N_7791,N_7945);
and U8626 (N_8626,N_7933,N_7950);
xor U8627 (N_8627,N_7882,N_8025);
xor U8628 (N_8628,N_7986,N_7980);
xnor U8629 (N_8629,N_7852,N_7647);
and U8630 (N_8630,N_7950,N_7929);
xnor U8631 (N_8631,N_7840,N_7597);
xor U8632 (N_8632,N_7975,N_7542);
and U8633 (N_8633,N_7645,N_7818);
xnor U8634 (N_8634,N_7719,N_7857);
nor U8635 (N_8635,N_7617,N_7672);
xor U8636 (N_8636,N_7922,N_7516);
xor U8637 (N_8637,N_7797,N_7905);
nor U8638 (N_8638,N_7730,N_8076);
and U8639 (N_8639,N_8123,N_7578);
or U8640 (N_8640,N_7983,N_8120);
nor U8641 (N_8641,N_7530,N_7718);
xnor U8642 (N_8642,N_7779,N_7961);
nor U8643 (N_8643,N_7599,N_7795);
nor U8644 (N_8644,N_7984,N_7682);
nor U8645 (N_8645,N_7500,N_8013);
or U8646 (N_8646,N_7505,N_8079);
nor U8647 (N_8647,N_7868,N_8037);
xnor U8648 (N_8648,N_7915,N_8105);
xnor U8649 (N_8649,N_7988,N_7834);
and U8650 (N_8650,N_7938,N_8046);
or U8651 (N_8651,N_7926,N_8103);
or U8652 (N_8652,N_7714,N_7967);
and U8653 (N_8653,N_7815,N_7937);
or U8654 (N_8654,N_7534,N_8063);
xor U8655 (N_8655,N_7908,N_7823);
or U8656 (N_8656,N_7691,N_7849);
or U8657 (N_8657,N_7662,N_7988);
nand U8658 (N_8658,N_8068,N_7983);
nand U8659 (N_8659,N_7614,N_8019);
and U8660 (N_8660,N_7761,N_7557);
nand U8661 (N_8661,N_7994,N_7741);
nor U8662 (N_8662,N_8029,N_7821);
nand U8663 (N_8663,N_7872,N_7993);
nand U8664 (N_8664,N_8094,N_8042);
nor U8665 (N_8665,N_7652,N_7703);
or U8666 (N_8666,N_7696,N_7603);
nand U8667 (N_8667,N_7687,N_7739);
or U8668 (N_8668,N_7713,N_7678);
nor U8669 (N_8669,N_7900,N_7672);
nand U8670 (N_8670,N_7676,N_7993);
xnor U8671 (N_8671,N_7741,N_7764);
nand U8672 (N_8672,N_7539,N_7910);
or U8673 (N_8673,N_7541,N_7936);
or U8674 (N_8674,N_7772,N_7874);
and U8675 (N_8675,N_8035,N_7710);
and U8676 (N_8676,N_7565,N_7869);
nand U8677 (N_8677,N_7580,N_8009);
nor U8678 (N_8678,N_7913,N_7804);
nor U8679 (N_8679,N_8074,N_7826);
and U8680 (N_8680,N_7814,N_7532);
or U8681 (N_8681,N_7952,N_7611);
and U8682 (N_8682,N_7886,N_7500);
xnor U8683 (N_8683,N_8012,N_7994);
nor U8684 (N_8684,N_7971,N_7796);
and U8685 (N_8685,N_8034,N_7761);
and U8686 (N_8686,N_7608,N_8037);
nor U8687 (N_8687,N_8006,N_7720);
xor U8688 (N_8688,N_7797,N_7801);
or U8689 (N_8689,N_7504,N_7859);
and U8690 (N_8690,N_8092,N_7878);
nand U8691 (N_8691,N_7786,N_7662);
xor U8692 (N_8692,N_7517,N_7811);
nor U8693 (N_8693,N_7834,N_7804);
nand U8694 (N_8694,N_7887,N_7962);
nand U8695 (N_8695,N_7574,N_7542);
nor U8696 (N_8696,N_8039,N_8057);
nor U8697 (N_8697,N_7884,N_7867);
and U8698 (N_8698,N_8027,N_7712);
and U8699 (N_8699,N_8099,N_8034);
or U8700 (N_8700,N_7902,N_7576);
xor U8701 (N_8701,N_7896,N_8078);
nand U8702 (N_8702,N_7689,N_7662);
nor U8703 (N_8703,N_7537,N_7701);
or U8704 (N_8704,N_7910,N_8084);
xnor U8705 (N_8705,N_7585,N_7624);
xor U8706 (N_8706,N_7895,N_7969);
nand U8707 (N_8707,N_7841,N_7745);
or U8708 (N_8708,N_7760,N_7510);
or U8709 (N_8709,N_7650,N_7649);
xor U8710 (N_8710,N_7936,N_7856);
nor U8711 (N_8711,N_7810,N_7916);
and U8712 (N_8712,N_7568,N_7866);
and U8713 (N_8713,N_7773,N_7665);
nand U8714 (N_8714,N_7671,N_8067);
and U8715 (N_8715,N_7945,N_7882);
nor U8716 (N_8716,N_7863,N_7505);
nand U8717 (N_8717,N_8108,N_7543);
and U8718 (N_8718,N_7834,N_7661);
and U8719 (N_8719,N_7861,N_7600);
nand U8720 (N_8720,N_8096,N_7821);
or U8721 (N_8721,N_7944,N_7908);
and U8722 (N_8722,N_8036,N_7744);
nor U8723 (N_8723,N_7628,N_8071);
nand U8724 (N_8724,N_7548,N_7637);
nor U8725 (N_8725,N_8003,N_7853);
or U8726 (N_8726,N_7540,N_7720);
xor U8727 (N_8727,N_7735,N_7864);
nand U8728 (N_8728,N_7977,N_7958);
xnor U8729 (N_8729,N_7656,N_7767);
and U8730 (N_8730,N_7589,N_7523);
or U8731 (N_8731,N_7940,N_7910);
nand U8732 (N_8732,N_7533,N_7881);
or U8733 (N_8733,N_7677,N_7544);
or U8734 (N_8734,N_7982,N_7678);
nor U8735 (N_8735,N_7591,N_7855);
xnor U8736 (N_8736,N_7732,N_7944);
or U8737 (N_8737,N_7907,N_7713);
or U8738 (N_8738,N_7682,N_7731);
and U8739 (N_8739,N_7887,N_7892);
nand U8740 (N_8740,N_7514,N_7630);
xnor U8741 (N_8741,N_7689,N_8003);
and U8742 (N_8742,N_8101,N_7980);
nand U8743 (N_8743,N_8054,N_7848);
and U8744 (N_8744,N_7751,N_7589);
nor U8745 (N_8745,N_8020,N_7569);
or U8746 (N_8746,N_7648,N_7745);
or U8747 (N_8747,N_7976,N_7944);
xor U8748 (N_8748,N_7569,N_8086);
nor U8749 (N_8749,N_7729,N_7528);
and U8750 (N_8750,N_8533,N_8666);
and U8751 (N_8751,N_8284,N_8517);
xnor U8752 (N_8752,N_8360,N_8403);
nor U8753 (N_8753,N_8322,N_8499);
nand U8754 (N_8754,N_8727,N_8735);
nand U8755 (N_8755,N_8694,N_8373);
and U8756 (N_8756,N_8189,N_8527);
nand U8757 (N_8757,N_8326,N_8623);
nand U8758 (N_8758,N_8270,N_8140);
and U8759 (N_8759,N_8594,N_8621);
nand U8760 (N_8760,N_8178,N_8530);
xor U8761 (N_8761,N_8170,N_8225);
xnor U8762 (N_8762,N_8131,N_8400);
or U8763 (N_8763,N_8325,N_8337);
nor U8764 (N_8764,N_8241,N_8726);
nand U8765 (N_8765,N_8229,N_8637);
nand U8766 (N_8766,N_8260,N_8399);
xor U8767 (N_8767,N_8192,N_8612);
and U8768 (N_8768,N_8142,N_8515);
and U8769 (N_8769,N_8504,N_8136);
or U8770 (N_8770,N_8458,N_8453);
nand U8771 (N_8771,N_8611,N_8181);
xor U8772 (N_8772,N_8314,N_8704);
xor U8773 (N_8773,N_8473,N_8245);
or U8774 (N_8774,N_8149,N_8375);
nor U8775 (N_8775,N_8304,N_8432);
and U8776 (N_8776,N_8626,N_8214);
xnor U8777 (N_8777,N_8223,N_8576);
or U8778 (N_8778,N_8289,N_8269);
or U8779 (N_8779,N_8205,N_8548);
or U8780 (N_8780,N_8424,N_8737);
nand U8781 (N_8781,N_8363,N_8426);
or U8782 (N_8782,N_8238,N_8460);
xnor U8783 (N_8783,N_8572,N_8457);
nand U8784 (N_8784,N_8575,N_8454);
xnor U8785 (N_8785,N_8605,N_8497);
and U8786 (N_8786,N_8438,N_8348);
and U8787 (N_8787,N_8372,N_8509);
or U8788 (N_8788,N_8210,N_8675);
nor U8789 (N_8789,N_8640,N_8321);
nor U8790 (N_8790,N_8423,N_8182);
xnor U8791 (N_8791,N_8428,N_8561);
nand U8792 (N_8792,N_8741,N_8294);
nand U8793 (N_8793,N_8166,N_8511);
nor U8794 (N_8794,N_8642,N_8307);
xnor U8795 (N_8795,N_8303,N_8630);
or U8796 (N_8796,N_8316,N_8243);
nor U8797 (N_8797,N_8491,N_8686);
or U8798 (N_8798,N_8343,N_8518);
nor U8799 (N_8799,N_8606,N_8707);
nor U8800 (N_8800,N_8146,N_8132);
nor U8801 (N_8801,N_8297,N_8451);
xor U8802 (N_8802,N_8401,N_8393);
nand U8803 (N_8803,N_8434,N_8180);
nand U8804 (N_8804,N_8455,N_8267);
and U8805 (N_8805,N_8128,N_8165);
nand U8806 (N_8806,N_8160,N_8582);
and U8807 (N_8807,N_8351,N_8660);
nand U8808 (N_8808,N_8620,N_8163);
xnor U8809 (N_8809,N_8639,N_8285);
nor U8810 (N_8810,N_8731,N_8577);
xnor U8811 (N_8811,N_8494,N_8204);
nand U8812 (N_8812,N_8602,N_8683);
xnor U8813 (N_8813,N_8668,N_8654);
and U8814 (N_8814,N_8155,N_8526);
or U8815 (N_8815,N_8328,N_8317);
nor U8816 (N_8816,N_8616,N_8130);
and U8817 (N_8817,N_8129,N_8462);
nor U8818 (N_8818,N_8498,N_8468);
or U8819 (N_8819,N_8471,N_8436);
or U8820 (N_8820,N_8638,N_8701);
xor U8821 (N_8821,N_8696,N_8265);
nor U8822 (N_8822,N_8540,N_8254);
nor U8823 (N_8823,N_8440,N_8280);
nor U8824 (N_8824,N_8185,N_8174);
or U8825 (N_8825,N_8421,N_8306);
or U8826 (N_8826,N_8550,N_8693);
and U8827 (N_8827,N_8720,N_8619);
xnor U8828 (N_8828,N_8302,N_8566);
xnor U8829 (N_8829,N_8747,N_8547);
xnor U8830 (N_8830,N_8456,N_8341);
nand U8831 (N_8831,N_8300,N_8587);
xnor U8832 (N_8832,N_8588,N_8217);
nor U8833 (N_8833,N_8557,N_8717);
or U8834 (N_8834,N_8299,N_8725);
nor U8835 (N_8835,N_8493,N_8629);
xor U8836 (N_8836,N_8201,N_8376);
xnor U8837 (N_8837,N_8586,N_8344);
xnor U8838 (N_8838,N_8569,N_8695);
nor U8839 (N_8839,N_8233,N_8161);
or U8840 (N_8840,N_8703,N_8571);
and U8841 (N_8841,N_8203,N_8239);
or U8842 (N_8842,N_8329,N_8653);
nand U8843 (N_8843,N_8641,N_8417);
nor U8844 (N_8844,N_8295,N_8216);
nor U8845 (N_8845,N_8480,N_8397);
xnor U8846 (N_8846,N_8259,N_8676);
and U8847 (N_8847,N_8362,N_8150);
xnor U8848 (N_8848,N_8614,N_8476);
nor U8849 (N_8849,N_8710,N_8742);
nor U8850 (N_8850,N_8601,N_8157);
xor U8851 (N_8851,N_8247,N_8315);
nor U8852 (N_8852,N_8382,N_8371);
nand U8853 (N_8853,N_8420,N_8353);
nor U8854 (N_8854,N_8173,N_8554);
nor U8855 (N_8855,N_8425,N_8221);
and U8856 (N_8856,N_8222,N_8176);
nand U8857 (N_8857,N_8251,N_8231);
nor U8858 (N_8858,N_8633,N_8711);
or U8859 (N_8859,N_8593,N_8127);
and U8860 (N_8860,N_8169,N_8396);
xor U8861 (N_8861,N_8481,N_8364);
nor U8862 (N_8862,N_8628,N_8740);
nand U8863 (N_8863,N_8368,N_8411);
nor U8864 (N_8864,N_8336,N_8689);
or U8865 (N_8865,N_8230,N_8383);
or U8866 (N_8866,N_8137,N_8565);
and U8867 (N_8867,N_8690,N_8592);
or U8868 (N_8868,N_8392,N_8532);
nand U8869 (N_8869,N_8244,N_8543);
nand U8870 (N_8870,N_8598,N_8470);
nand U8871 (N_8871,N_8749,N_8198);
xnor U8872 (N_8872,N_8282,N_8590);
nor U8873 (N_8873,N_8171,N_8207);
or U8874 (N_8874,N_8283,N_8391);
xnor U8875 (N_8875,N_8332,N_8679);
xnor U8876 (N_8876,N_8609,N_8542);
nor U8877 (N_8877,N_8447,N_8736);
xnor U8878 (N_8878,N_8320,N_8734);
xnor U8879 (N_8879,N_8708,N_8746);
and U8880 (N_8880,N_8183,N_8579);
and U8881 (N_8881,N_8319,N_8730);
nand U8882 (N_8882,N_8715,N_8313);
nor U8883 (N_8883,N_8719,N_8305);
and U8884 (N_8884,N_8537,N_8429);
and U8885 (N_8885,N_8656,N_8702);
nand U8886 (N_8886,N_8416,N_8404);
nor U8887 (N_8887,N_8333,N_8144);
xor U8888 (N_8888,N_8597,N_8272);
and U8889 (N_8889,N_8208,N_8482);
nand U8890 (N_8890,N_8648,N_8452);
xnor U8891 (N_8891,N_8188,N_8591);
or U8892 (N_8892,N_8624,N_8414);
or U8893 (N_8893,N_8549,N_8248);
xor U8894 (N_8894,N_8716,N_8669);
nand U8895 (N_8895,N_8257,N_8552);
xnor U8896 (N_8896,N_8342,N_8290);
and U8897 (N_8897,N_8264,N_8151);
xnor U8898 (N_8898,N_8534,N_8308);
xnor U8899 (N_8899,N_8387,N_8158);
or U8900 (N_8900,N_8418,N_8148);
or U8901 (N_8901,N_8356,N_8227);
xor U8902 (N_8902,N_8293,N_8525);
xnor U8903 (N_8903,N_8268,N_8627);
nor U8904 (N_8904,N_8379,N_8724);
nor U8905 (N_8905,N_8651,N_8266);
xnor U8906 (N_8906,N_8159,N_8522);
or U8907 (N_8907,N_8141,N_8406);
or U8908 (N_8908,N_8665,N_8256);
or U8909 (N_8909,N_8309,N_8433);
nor U8910 (N_8910,N_8202,N_8435);
or U8911 (N_8911,N_8240,N_8439);
and U8912 (N_8912,N_8437,N_8622);
or U8913 (N_8913,N_8279,N_8374);
and U8914 (N_8914,N_8562,N_8249);
or U8915 (N_8915,N_8486,N_8528);
xor U8916 (N_8916,N_8446,N_8512);
and U8917 (N_8917,N_8459,N_8712);
or U8918 (N_8918,N_8327,N_8347);
or U8919 (N_8919,N_8478,N_8196);
and U8920 (N_8920,N_8650,N_8263);
or U8921 (N_8921,N_8496,N_8408);
nor U8922 (N_8922,N_8224,N_8258);
nor U8923 (N_8923,N_8236,N_8212);
xor U8924 (N_8924,N_8466,N_8324);
or U8925 (N_8925,N_8632,N_8748);
or U8926 (N_8926,N_8663,N_8728);
or U8927 (N_8927,N_8595,N_8469);
nor U8928 (N_8928,N_8490,N_8539);
and U8929 (N_8929,N_8464,N_8145);
nor U8930 (N_8930,N_8402,N_8358);
nand U8931 (N_8931,N_8652,N_8262);
nand U8932 (N_8932,N_8154,N_8535);
and U8933 (N_8933,N_8500,N_8580);
nand U8934 (N_8934,N_8443,N_8366);
nor U8935 (N_8935,N_8168,N_8430);
nand U8936 (N_8936,N_8134,N_8226);
nand U8937 (N_8937,N_8555,N_8330);
or U8938 (N_8938,N_8508,N_8688);
nand U8939 (N_8939,N_8489,N_8187);
or U8940 (N_8940,N_8261,N_8487);
nor U8941 (N_8941,N_8677,N_8381);
nor U8942 (N_8942,N_8655,N_8377);
or U8943 (N_8943,N_8485,N_8475);
nor U8944 (N_8944,N_8386,N_8618);
nand U8945 (N_8945,N_8448,N_8413);
nand U8946 (N_8946,N_8514,N_8444);
and U8947 (N_8947,N_8199,N_8125);
xnor U8948 (N_8948,N_8743,N_8567);
or U8949 (N_8949,N_8681,N_8422);
xor U8950 (N_8950,N_8472,N_8732);
nor U8951 (N_8951,N_8474,N_8349);
nand U8952 (N_8952,N_8583,N_8296);
nand U8953 (N_8953,N_8220,N_8488);
xnor U8954 (N_8954,N_8560,N_8699);
nor U8955 (N_8955,N_8415,N_8722);
or U8956 (N_8956,N_8367,N_8389);
and U8957 (N_8957,N_8193,N_8311);
nand U8958 (N_8958,N_8186,N_8179);
or U8959 (N_8959,N_8335,N_8190);
or U8960 (N_8960,N_8278,N_8318);
or U8961 (N_8961,N_8301,N_8310);
and U8962 (N_8962,N_8698,N_8143);
xor U8963 (N_8963,N_8599,N_8610);
and U8964 (N_8964,N_8503,N_8551);
nor U8965 (N_8965,N_8733,N_8331);
nor U8966 (N_8966,N_8209,N_8345);
nand U8967 (N_8967,N_8723,N_8152);
or U8968 (N_8968,N_8250,N_8662);
and U8969 (N_8969,N_8684,N_8649);
nor U8970 (N_8970,N_8273,N_8570);
nor U8971 (N_8971,N_8369,N_8645);
xor U8972 (N_8972,N_8573,N_8242);
and U8973 (N_8973,N_8409,N_8553);
nand U8974 (N_8974,N_8147,N_8680);
xnor U8975 (N_8975,N_8584,N_8219);
nor U8976 (N_8976,N_8431,N_8359);
nand U8977 (N_8977,N_8461,N_8643);
or U8978 (N_8978,N_8339,N_8410);
nor U8979 (N_8979,N_8213,N_8276);
or U8980 (N_8980,N_8625,N_8275);
and U8981 (N_8981,N_8556,N_8352);
nor U8982 (N_8982,N_8390,N_8510);
nor U8983 (N_8983,N_8538,N_8636);
nand U8984 (N_8984,N_8589,N_8340);
and U8985 (N_8985,N_8412,N_8613);
nor U8986 (N_8986,N_8398,N_8234);
or U8987 (N_8987,N_8361,N_8745);
xor U8988 (N_8988,N_8175,N_8477);
xnor U8989 (N_8989,N_8380,N_8427);
xor U8990 (N_8990,N_8667,N_8277);
or U8991 (N_8991,N_8644,N_8346);
xor U8992 (N_8992,N_8661,N_8388);
and U8993 (N_8993,N_8647,N_8281);
and U8994 (N_8994,N_8228,N_8657);
nor U8995 (N_8995,N_8568,N_8607);
or U8996 (N_8996,N_8558,N_8384);
nor U8997 (N_8997,N_8139,N_8274);
nor U8998 (N_8998,N_8292,N_8354);
nand U8999 (N_8999,N_8338,N_8287);
xnor U9000 (N_9000,N_8523,N_8739);
or U9001 (N_9001,N_8670,N_8578);
nand U9002 (N_9002,N_8673,N_8718);
or U9003 (N_9003,N_8237,N_8394);
xnor U9004 (N_9004,N_8246,N_8298);
nand U9005 (N_9005,N_8585,N_8206);
nor U9006 (N_9006,N_8172,N_8646);
nor U9007 (N_9007,N_8365,N_8729);
nand U9008 (N_9008,N_8323,N_8546);
nor U9009 (N_9009,N_8215,N_8659);
xor U9010 (N_9010,N_8378,N_8167);
or U9011 (N_9011,N_8442,N_8467);
nand U9012 (N_9012,N_8484,N_8501);
xor U9013 (N_9013,N_8545,N_8685);
xnor U9014 (N_9014,N_8706,N_8581);
nor U9015 (N_9015,N_8232,N_8355);
nand U9016 (N_9016,N_8574,N_8463);
xnor U9017 (N_9017,N_8407,N_8744);
or U9018 (N_9018,N_8634,N_8253);
and U9019 (N_9019,N_8153,N_8138);
or U9020 (N_9020,N_8291,N_8615);
xnor U9021 (N_9021,N_8559,N_8483);
and U9022 (N_9022,N_8691,N_8700);
nor U9023 (N_9023,N_8495,N_8156);
xnor U9024 (N_9024,N_8513,N_8164);
or U9025 (N_9025,N_8692,N_8564);
xor U9026 (N_9026,N_8596,N_8544);
nor U9027 (N_9027,N_8520,N_8162);
or U9028 (N_9028,N_8419,N_8713);
or U9029 (N_9029,N_8521,N_8405);
nand U9030 (N_9030,N_8721,N_8536);
nor U9031 (N_9031,N_8255,N_8505);
or U9032 (N_9032,N_8631,N_8312);
and U9033 (N_9033,N_8271,N_8671);
or U9034 (N_9034,N_8714,N_8195);
and U9035 (N_9035,N_8709,N_8286);
xnor U9036 (N_9036,N_8672,N_8126);
xnor U9037 (N_9037,N_8502,N_8541);
or U9038 (N_9038,N_8697,N_8738);
nor U9039 (N_9039,N_8617,N_8370);
nand U9040 (N_9040,N_8445,N_8135);
xnor U9041 (N_9041,N_8529,N_8705);
nor U9042 (N_9042,N_8608,N_8177);
or U9043 (N_9043,N_8516,N_8674);
nand U9044 (N_9044,N_8519,N_8235);
or U9045 (N_9045,N_8600,N_8531);
or U9046 (N_9046,N_8450,N_8218);
and U9047 (N_9047,N_8252,N_8664);
nand U9048 (N_9048,N_8492,N_8211);
xnor U9049 (N_9049,N_8288,N_8385);
xor U9050 (N_9050,N_8191,N_8687);
nand U9051 (N_9051,N_8506,N_8604);
nand U9052 (N_9052,N_8658,N_8479);
xor U9053 (N_9053,N_8184,N_8563);
and U9054 (N_9054,N_8395,N_8133);
nor U9055 (N_9055,N_8507,N_8350);
and U9056 (N_9056,N_8194,N_8357);
nand U9057 (N_9057,N_8197,N_8682);
nand U9058 (N_9058,N_8449,N_8635);
nor U9059 (N_9059,N_8200,N_8441);
xor U9060 (N_9060,N_8465,N_8334);
and U9061 (N_9061,N_8603,N_8678);
and U9062 (N_9062,N_8524,N_8648);
nor U9063 (N_9063,N_8139,N_8136);
nand U9064 (N_9064,N_8455,N_8554);
xnor U9065 (N_9065,N_8620,N_8342);
or U9066 (N_9066,N_8385,N_8300);
nor U9067 (N_9067,N_8282,N_8293);
xnor U9068 (N_9068,N_8209,N_8182);
or U9069 (N_9069,N_8246,N_8368);
and U9070 (N_9070,N_8177,N_8288);
and U9071 (N_9071,N_8589,N_8467);
or U9072 (N_9072,N_8609,N_8423);
nand U9073 (N_9073,N_8374,N_8194);
or U9074 (N_9074,N_8331,N_8606);
and U9075 (N_9075,N_8672,N_8421);
xor U9076 (N_9076,N_8649,N_8403);
or U9077 (N_9077,N_8383,N_8653);
and U9078 (N_9078,N_8152,N_8186);
nand U9079 (N_9079,N_8578,N_8480);
nor U9080 (N_9080,N_8503,N_8674);
or U9081 (N_9081,N_8523,N_8148);
nor U9082 (N_9082,N_8462,N_8474);
nand U9083 (N_9083,N_8455,N_8289);
xnor U9084 (N_9084,N_8282,N_8678);
and U9085 (N_9085,N_8185,N_8262);
and U9086 (N_9086,N_8722,N_8304);
or U9087 (N_9087,N_8236,N_8482);
and U9088 (N_9088,N_8686,N_8238);
or U9089 (N_9089,N_8374,N_8597);
nor U9090 (N_9090,N_8454,N_8135);
xor U9091 (N_9091,N_8196,N_8163);
or U9092 (N_9092,N_8125,N_8637);
or U9093 (N_9093,N_8131,N_8575);
and U9094 (N_9094,N_8156,N_8535);
xnor U9095 (N_9095,N_8125,N_8342);
nor U9096 (N_9096,N_8221,N_8306);
nor U9097 (N_9097,N_8558,N_8523);
nor U9098 (N_9098,N_8150,N_8604);
nor U9099 (N_9099,N_8492,N_8231);
nor U9100 (N_9100,N_8727,N_8558);
and U9101 (N_9101,N_8316,N_8261);
xnor U9102 (N_9102,N_8216,N_8260);
xor U9103 (N_9103,N_8597,N_8740);
xnor U9104 (N_9104,N_8705,N_8154);
and U9105 (N_9105,N_8242,N_8274);
nand U9106 (N_9106,N_8346,N_8576);
or U9107 (N_9107,N_8163,N_8705);
nor U9108 (N_9108,N_8483,N_8186);
and U9109 (N_9109,N_8386,N_8490);
and U9110 (N_9110,N_8257,N_8247);
or U9111 (N_9111,N_8440,N_8578);
nand U9112 (N_9112,N_8359,N_8546);
or U9113 (N_9113,N_8646,N_8701);
xor U9114 (N_9114,N_8279,N_8250);
or U9115 (N_9115,N_8221,N_8453);
or U9116 (N_9116,N_8133,N_8365);
nand U9117 (N_9117,N_8587,N_8396);
nor U9118 (N_9118,N_8632,N_8518);
xor U9119 (N_9119,N_8668,N_8345);
or U9120 (N_9120,N_8461,N_8688);
xnor U9121 (N_9121,N_8414,N_8359);
nand U9122 (N_9122,N_8193,N_8212);
or U9123 (N_9123,N_8491,N_8619);
nand U9124 (N_9124,N_8601,N_8545);
nor U9125 (N_9125,N_8483,N_8430);
nor U9126 (N_9126,N_8735,N_8206);
and U9127 (N_9127,N_8732,N_8398);
nor U9128 (N_9128,N_8199,N_8647);
xor U9129 (N_9129,N_8185,N_8698);
xnor U9130 (N_9130,N_8188,N_8126);
nor U9131 (N_9131,N_8191,N_8732);
and U9132 (N_9132,N_8359,N_8399);
nand U9133 (N_9133,N_8424,N_8708);
and U9134 (N_9134,N_8329,N_8146);
and U9135 (N_9135,N_8245,N_8744);
or U9136 (N_9136,N_8195,N_8247);
nand U9137 (N_9137,N_8595,N_8313);
and U9138 (N_9138,N_8306,N_8679);
xor U9139 (N_9139,N_8703,N_8331);
and U9140 (N_9140,N_8363,N_8634);
nand U9141 (N_9141,N_8689,N_8412);
nand U9142 (N_9142,N_8161,N_8695);
xor U9143 (N_9143,N_8575,N_8700);
or U9144 (N_9144,N_8496,N_8220);
or U9145 (N_9145,N_8249,N_8257);
nand U9146 (N_9146,N_8295,N_8727);
nor U9147 (N_9147,N_8674,N_8206);
or U9148 (N_9148,N_8381,N_8447);
and U9149 (N_9149,N_8356,N_8337);
nor U9150 (N_9150,N_8684,N_8666);
and U9151 (N_9151,N_8154,N_8252);
xor U9152 (N_9152,N_8558,N_8564);
nor U9153 (N_9153,N_8171,N_8165);
or U9154 (N_9154,N_8456,N_8393);
and U9155 (N_9155,N_8449,N_8735);
nor U9156 (N_9156,N_8625,N_8279);
nor U9157 (N_9157,N_8737,N_8547);
nor U9158 (N_9158,N_8159,N_8350);
and U9159 (N_9159,N_8693,N_8451);
nand U9160 (N_9160,N_8647,N_8515);
nand U9161 (N_9161,N_8562,N_8510);
or U9162 (N_9162,N_8225,N_8546);
and U9163 (N_9163,N_8652,N_8177);
nand U9164 (N_9164,N_8269,N_8630);
xor U9165 (N_9165,N_8291,N_8319);
nor U9166 (N_9166,N_8738,N_8512);
nor U9167 (N_9167,N_8163,N_8296);
and U9168 (N_9168,N_8269,N_8723);
nand U9169 (N_9169,N_8131,N_8191);
or U9170 (N_9170,N_8462,N_8329);
or U9171 (N_9171,N_8221,N_8434);
nand U9172 (N_9172,N_8620,N_8502);
nand U9173 (N_9173,N_8710,N_8551);
nand U9174 (N_9174,N_8513,N_8672);
nor U9175 (N_9175,N_8126,N_8449);
nor U9176 (N_9176,N_8488,N_8530);
or U9177 (N_9177,N_8310,N_8187);
or U9178 (N_9178,N_8153,N_8401);
or U9179 (N_9179,N_8271,N_8207);
xnor U9180 (N_9180,N_8622,N_8653);
or U9181 (N_9181,N_8338,N_8147);
nand U9182 (N_9182,N_8696,N_8433);
nand U9183 (N_9183,N_8264,N_8715);
and U9184 (N_9184,N_8677,N_8609);
or U9185 (N_9185,N_8491,N_8180);
nor U9186 (N_9186,N_8247,N_8688);
nor U9187 (N_9187,N_8228,N_8738);
or U9188 (N_9188,N_8709,N_8257);
xnor U9189 (N_9189,N_8329,N_8529);
or U9190 (N_9190,N_8286,N_8492);
and U9191 (N_9191,N_8145,N_8381);
nor U9192 (N_9192,N_8141,N_8417);
nand U9193 (N_9193,N_8280,N_8592);
and U9194 (N_9194,N_8482,N_8263);
nand U9195 (N_9195,N_8420,N_8183);
or U9196 (N_9196,N_8568,N_8146);
and U9197 (N_9197,N_8454,N_8278);
nand U9198 (N_9198,N_8597,N_8196);
xor U9199 (N_9199,N_8302,N_8202);
and U9200 (N_9200,N_8387,N_8718);
or U9201 (N_9201,N_8238,N_8422);
or U9202 (N_9202,N_8387,N_8376);
or U9203 (N_9203,N_8503,N_8194);
nand U9204 (N_9204,N_8217,N_8415);
xor U9205 (N_9205,N_8181,N_8574);
xor U9206 (N_9206,N_8321,N_8371);
nor U9207 (N_9207,N_8362,N_8653);
xnor U9208 (N_9208,N_8574,N_8326);
xor U9209 (N_9209,N_8716,N_8210);
and U9210 (N_9210,N_8669,N_8595);
xnor U9211 (N_9211,N_8361,N_8404);
nand U9212 (N_9212,N_8331,N_8699);
nand U9213 (N_9213,N_8240,N_8345);
or U9214 (N_9214,N_8615,N_8483);
nor U9215 (N_9215,N_8592,N_8585);
or U9216 (N_9216,N_8468,N_8476);
and U9217 (N_9217,N_8550,N_8663);
nand U9218 (N_9218,N_8614,N_8513);
nand U9219 (N_9219,N_8200,N_8704);
xor U9220 (N_9220,N_8331,N_8527);
nor U9221 (N_9221,N_8684,N_8405);
and U9222 (N_9222,N_8151,N_8258);
nor U9223 (N_9223,N_8248,N_8260);
xor U9224 (N_9224,N_8492,N_8266);
nand U9225 (N_9225,N_8166,N_8636);
xor U9226 (N_9226,N_8334,N_8172);
nor U9227 (N_9227,N_8406,N_8601);
xor U9228 (N_9228,N_8198,N_8223);
xor U9229 (N_9229,N_8371,N_8323);
nor U9230 (N_9230,N_8254,N_8327);
nand U9231 (N_9231,N_8477,N_8683);
nand U9232 (N_9232,N_8265,N_8170);
nand U9233 (N_9233,N_8215,N_8447);
xor U9234 (N_9234,N_8534,N_8174);
nor U9235 (N_9235,N_8738,N_8624);
nand U9236 (N_9236,N_8166,N_8694);
xor U9237 (N_9237,N_8223,N_8305);
nand U9238 (N_9238,N_8689,N_8532);
nand U9239 (N_9239,N_8499,N_8412);
xor U9240 (N_9240,N_8355,N_8606);
and U9241 (N_9241,N_8427,N_8448);
nor U9242 (N_9242,N_8282,N_8205);
xor U9243 (N_9243,N_8583,N_8578);
xor U9244 (N_9244,N_8218,N_8129);
nand U9245 (N_9245,N_8188,N_8371);
or U9246 (N_9246,N_8633,N_8650);
nor U9247 (N_9247,N_8307,N_8415);
or U9248 (N_9248,N_8646,N_8237);
and U9249 (N_9249,N_8232,N_8230);
or U9250 (N_9250,N_8736,N_8139);
nor U9251 (N_9251,N_8682,N_8499);
nand U9252 (N_9252,N_8125,N_8308);
xnor U9253 (N_9253,N_8330,N_8308);
nor U9254 (N_9254,N_8593,N_8600);
and U9255 (N_9255,N_8559,N_8227);
xor U9256 (N_9256,N_8425,N_8656);
xor U9257 (N_9257,N_8475,N_8582);
xor U9258 (N_9258,N_8633,N_8543);
or U9259 (N_9259,N_8220,N_8745);
nor U9260 (N_9260,N_8318,N_8606);
xor U9261 (N_9261,N_8250,N_8374);
xor U9262 (N_9262,N_8146,N_8376);
nand U9263 (N_9263,N_8198,N_8288);
or U9264 (N_9264,N_8301,N_8213);
or U9265 (N_9265,N_8126,N_8231);
nor U9266 (N_9266,N_8462,N_8243);
or U9267 (N_9267,N_8386,N_8638);
or U9268 (N_9268,N_8421,N_8341);
and U9269 (N_9269,N_8474,N_8153);
and U9270 (N_9270,N_8162,N_8741);
and U9271 (N_9271,N_8267,N_8738);
nand U9272 (N_9272,N_8297,N_8189);
nand U9273 (N_9273,N_8624,N_8513);
nor U9274 (N_9274,N_8523,N_8506);
nor U9275 (N_9275,N_8242,N_8255);
xnor U9276 (N_9276,N_8424,N_8640);
nand U9277 (N_9277,N_8364,N_8387);
or U9278 (N_9278,N_8140,N_8654);
and U9279 (N_9279,N_8397,N_8462);
nor U9280 (N_9280,N_8304,N_8163);
or U9281 (N_9281,N_8676,N_8430);
nor U9282 (N_9282,N_8719,N_8369);
and U9283 (N_9283,N_8621,N_8488);
and U9284 (N_9284,N_8584,N_8341);
nand U9285 (N_9285,N_8158,N_8509);
xor U9286 (N_9286,N_8591,N_8326);
and U9287 (N_9287,N_8451,N_8243);
nand U9288 (N_9288,N_8375,N_8638);
and U9289 (N_9289,N_8181,N_8651);
nand U9290 (N_9290,N_8421,N_8169);
nor U9291 (N_9291,N_8423,N_8229);
xnor U9292 (N_9292,N_8170,N_8141);
nand U9293 (N_9293,N_8605,N_8662);
nor U9294 (N_9294,N_8161,N_8377);
nor U9295 (N_9295,N_8237,N_8614);
xnor U9296 (N_9296,N_8283,N_8137);
nand U9297 (N_9297,N_8562,N_8448);
nor U9298 (N_9298,N_8356,N_8474);
nand U9299 (N_9299,N_8238,N_8306);
nor U9300 (N_9300,N_8515,N_8518);
and U9301 (N_9301,N_8538,N_8458);
nor U9302 (N_9302,N_8487,N_8262);
nor U9303 (N_9303,N_8361,N_8356);
nand U9304 (N_9304,N_8455,N_8735);
or U9305 (N_9305,N_8659,N_8125);
or U9306 (N_9306,N_8336,N_8528);
or U9307 (N_9307,N_8463,N_8447);
xnor U9308 (N_9308,N_8283,N_8532);
and U9309 (N_9309,N_8274,N_8541);
nor U9310 (N_9310,N_8139,N_8233);
or U9311 (N_9311,N_8269,N_8558);
nor U9312 (N_9312,N_8182,N_8567);
xor U9313 (N_9313,N_8745,N_8306);
and U9314 (N_9314,N_8316,N_8306);
nor U9315 (N_9315,N_8423,N_8262);
and U9316 (N_9316,N_8710,N_8248);
nor U9317 (N_9317,N_8595,N_8279);
or U9318 (N_9318,N_8333,N_8326);
nand U9319 (N_9319,N_8237,N_8363);
and U9320 (N_9320,N_8304,N_8392);
xnor U9321 (N_9321,N_8238,N_8575);
nand U9322 (N_9322,N_8456,N_8605);
and U9323 (N_9323,N_8420,N_8220);
nand U9324 (N_9324,N_8527,N_8612);
or U9325 (N_9325,N_8446,N_8629);
xnor U9326 (N_9326,N_8245,N_8729);
nor U9327 (N_9327,N_8221,N_8672);
and U9328 (N_9328,N_8356,N_8192);
xnor U9329 (N_9329,N_8598,N_8674);
and U9330 (N_9330,N_8575,N_8341);
nand U9331 (N_9331,N_8445,N_8154);
nor U9332 (N_9332,N_8517,N_8158);
nor U9333 (N_9333,N_8735,N_8165);
xnor U9334 (N_9334,N_8316,N_8511);
nor U9335 (N_9335,N_8164,N_8595);
nor U9336 (N_9336,N_8363,N_8696);
nor U9337 (N_9337,N_8576,N_8548);
nor U9338 (N_9338,N_8239,N_8166);
or U9339 (N_9339,N_8286,N_8668);
or U9340 (N_9340,N_8670,N_8333);
and U9341 (N_9341,N_8657,N_8464);
nand U9342 (N_9342,N_8574,N_8170);
xor U9343 (N_9343,N_8413,N_8446);
xor U9344 (N_9344,N_8745,N_8421);
nand U9345 (N_9345,N_8410,N_8235);
nand U9346 (N_9346,N_8253,N_8651);
or U9347 (N_9347,N_8333,N_8287);
nor U9348 (N_9348,N_8355,N_8418);
and U9349 (N_9349,N_8424,N_8503);
and U9350 (N_9350,N_8129,N_8410);
xor U9351 (N_9351,N_8410,N_8672);
nand U9352 (N_9352,N_8600,N_8153);
xor U9353 (N_9353,N_8358,N_8619);
nor U9354 (N_9354,N_8674,N_8217);
xnor U9355 (N_9355,N_8669,N_8166);
nand U9356 (N_9356,N_8152,N_8493);
xnor U9357 (N_9357,N_8497,N_8636);
xor U9358 (N_9358,N_8451,N_8315);
nand U9359 (N_9359,N_8422,N_8640);
or U9360 (N_9360,N_8501,N_8558);
xnor U9361 (N_9361,N_8535,N_8273);
and U9362 (N_9362,N_8346,N_8684);
and U9363 (N_9363,N_8184,N_8325);
xnor U9364 (N_9364,N_8597,N_8246);
or U9365 (N_9365,N_8306,N_8148);
or U9366 (N_9366,N_8638,N_8717);
nand U9367 (N_9367,N_8432,N_8394);
xor U9368 (N_9368,N_8639,N_8215);
nor U9369 (N_9369,N_8616,N_8318);
and U9370 (N_9370,N_8271,N_8593);
xnor U9371 (N_9371,N_8426,N_8545);
nor U9372 (N_9372,N_8415,N_8237);
or U9373 (N_9373,N_8677,N_8519);
nor U9374 (N_9374,N_8529,N_8188);
or U9375 (N_9375,N_9073,N_9319);
xnor U9376 (N_9376,N_9272,N_9138);
or U9377 (N_9377,N_8949,N_9051);
nand U9378 (N_9378,N_8967,N_8866);
and U9379 (N_9379,N_9140,N_9150);
xnor U9380 (N_9380,N_9347,N_9168);
or U9381 (N_9381,N_9317,N_9214);
nor U9382 (N_9382,N_9079,N_9224);
nand U9383 (N_9383,N_8905,N_9042);
nand U9384 (N_9384,N_9131,N_8880);
nand U9385 (N_9385,N_8830,N_9287);
nand U9386 (N_9386,N_9100,N_9164);
nor U9387 (N_9387,N_9335,N_8878);
and U9388 (N_9388,N_8773,N_9193);
nand U9389 (N_9389,N_8785,N_8851);
xnor U9390 (N_9390,N_8844,N_9093);
or U9391 (N_9391,N_8887,N_9273);
or U9392 (N_9392,N_8817,N_8863);
nand U9393 (N_9393,N_8794,N_9284);
nand U9394 (N_9394,N_8852,N_9212);
xor U9395 (N_9395,N_8791,N_8959);
or U9396 (N_9396,N_9230,N_9312);
xnor U9397 (N_9397,N_9313,N_8806);
xnor U9398 (N_9398,N_9155,N_9291);
nand U9399 (N_9399,N_9298,N_8804);
xor U9400 (N_9400,N_9369,N_9267);
nand U9401 (N_9401,N_9173,N_8893);
or U9402 (N_9402,N_9070,N_9081);
nor U9403 (N_9403,N_9075,N_9277);
and U9404 (N_9404,N_8882,N_9204);
xnor U9405 (N_9405,N_9135,N_9196);
nor U9406 (N_9406,N_8774,N_9185);
and U9407 (N_9407,N_8853,N_9221);
xor U9408 (N_9408,N_9141,N_9182);
or U9409 (N_9409,N_8936,N_8793);
or U9410 (N_9410,N_8931,N_8819);
and U9411 (N_9411,N_9342,N_9310);
nor U9412 (N_9412,N_9304,N_9199);
or U9413 (N_9413,N_9016,N_9340);
xnor U9414 (N_9414,N_9231,N_8858);
nand U9415 (N_9415,N_9015,N_9159);
and U9416 (N_9416,N_9156,N_8833);
nor U9417 (N_9417,N_9315,N_9142);
and U9418 (N_9418,N_9103,N_9048);
or U9419 (N_9419,N_8836,N_9053);
nand U9420 (N_9420,N_8977,N_8862);
and U9421 (N_9421,N_9363,N_8846);
nand U9422 (N_9422,N_9184,N_9002);
nand U9423 (N_9423,N_9239,N_8764);
or U9424 (N_9424,N_9368,N_9106);
nand U9425 (N_9425,N_8891,N_9054);
or U9426 (N_9426,N_9288,N_8903);
or U9427 (N_9427,N_9228,N_8921);
and U9428 (N_9428,N_9191,N_9326);
nand U9429 (N_9429,N_9175,N_9060);
nor U9430 (N_9430,N_8937,N_9167);
and U9431 (N_9431,N_8890,N_8986);
nand U9432 (N_9432,N_9353,N_9086);
nor U9433 (N_9433,N_8834,N_8990);
xor U9434 (N_9434,N_9307,N_9332);
nand U9435 (N_9435,N_8790,N_9233);
or U9436 (N_9436,N_9139,N_9323);
or U9437 (N_9437,N_8816,N_8910);
nand U9438 (N_9438,N_8953,N_9321);
xor U9439 (N_9439,N_9157,N_8795);
nor U9440 (N_9440,N_9041,N_9349);
nand U9441 (N_9441,N_8814,N_8783);
nor U9442 (N_9442,N_9072,N_8975);
nand U9443 (N_9443,N_9311,N_9244);
nand U9444 (N_9444,N_9163,N_9009);
nor U9445 (N_9445,N_8984,N_9198);
nand U9446 (N_9446,N_8849,N_8762);
or U9447 (N_9447,N_9074,N_9035);
xnor U9448 (N_9448,N_9005,N_8820);
or U9449 (N_9449,N_8904,N_8818);
and U9450 (N_9450,N_8923,N_8756);
and U9451 (N_9451,N_9000,N_8796);
or U9452 (N_9452,N_9028,N_8831);
nand U9453 (N_9453,N_8964,N_9125);
xnor U9454 (N_9454,N_9356,N_8750);
xor U9455 (N_9455,N_9308,N_8874);
or U9456 (N_9456,N_8974,N_9271);
nor U9457 (N_9457,N_9264,N_8875);
nor U9458 (N_9458,N_8883,N_8767);
or U9459 (N_9459,N_8811,N_9099);
nor U9460 (N_9460,N_9047,N_8754);
nor U9461 (N_9461,N_9314,N_9145);
nor U9462 (N_9462,N_9056,N_8792);
xor U9463 (N_9463,N_9297,N_9202);
nor U9464 (N_9464,N_8763,N_9011);
xor U9465 (N_9465,N_9306,N_9300);
nand U9466 (N_9466,N_9110,N_8752);
and U9467 (N_9467,N_9189,N_9275);
nand U9468 (N_9468,N_8802,N_9205);
or U9469 (N_9469,N_9077,N_8934);
nand U9470 (N_9470,N_8938,N_9339);
nand U9471 (N_9471,N_9024,N_9136);
xor U9472 (N_9472,N_9213,N_9087);
nor U9473 (N_9473,N_9153,N_8789);
nand U9474 (N_9474,N_8917,N_9301);
and U9475 (N_9475,N_8998,N_8927);
nor U9476 (N_9476,N_9065,N_8787);
xor U9477 (N_9477,N_9248,N_9219);
or U9478 (N_9478,N_9200,N_9345);
xnor U9479 (N_9479,N_8856,N_9082);
nand U9480 (N_9480,N_9088,N_8869);
or U9481 (N_9481,N_8919,N_8876);
xor U9482 (N_9482,N_9098,N_9172);
xor U9483 (N_9483,N_9115,N_9021);
xnor U9484 (N_9484,N_9063,N_8902);
xor U9485 (N_9485,N_8886,N_8993);
xor U9486 (N_9486,N_8784,N_9260);
xor U9487 (N_9487,N_8825,N_8980);
and U9488 (N_9488,N_9147,N_9289);
xnor U9489 (N_9489,N_8994,N_8845);
nor U9490 (N_9490,N_9162,N_9188);
and U9491 (N_9491,N_8900,N_8924);
xor U9492 (N_9492,N_9045,N_9170);
xnor U9493 (N_9493,N_8872,N_8847);
nand U9494 (N_9494,N_8956,N_9226);
or U9495 (N_9495,N_8981,N_8935);
and U9496 (N_9496,N_8828,N_9201);
xor U9497 (N_9497,N_9338,N_8757);
and U9498 (N_9498,N_9371,N_9357);
nand U9499 (N_9499,N_9374,N_9303);
nand U9500 (N_9500,N_8838,N_8929);
xor U9501 (N_9501,N_8861,N_9364);
or U9502 (N_9502,N_8772,N_8803);
nor U9503 (N_9503,N_8835,N_8865);
nand U9504 (N_9504,N_8871,N_9361);
nand U9505 (N_9505,N_8827,N_9178);
nand U9506 (N_9506,N_8766,N_9302);
nand U9507 (N_9507,N_9322,N_8780);
nor U9508 (N_9508,N_9169,N_9092);
nand U9509 (N_9509,N_8822,N_8751);
xnor U9510 (N_9510,N_9194,N_8988);
and U9511 (N_9511,N_9254,N_9033);
xnor U9512 (N_9512,N_9324,N_9211);
nor U9513 (N_9513,N_8765,N_9362);
xnor U9514 (N_9514,N_9071,N_8832);
nand U9515 (N_9515,N_8896,N_9066);
nand U9516 (N_9516,N_8776,N_8992);
or U9517 (N_9517,N_8800,N_9117);
nand U9518 (N_9518,N_9285,N_9293);
nand U9519 (N_9519,N_8989,N_9179);
xnor U9520 (N_9520,N_8952,N_9278);
nand U9521 (N_9521,N_9001,N_8841);
nor U9522 (N_9522,N_8837,N_9069);
nand U9523 (N_9523,N_9111,N_9240);
nor U9524 (N_9524,N_8920,N_8962);
nor U9525 (N_9525,N_9032,N_9127);
nand U9526 (N_9526,N_8909,N_8840);
and U9527 (N_9527,N_9274,N_8928);
or U9528 (N_9528,N_8985,N_9327);
nor U9529 (N_9529,N_9107,N_8813);
xor U9530 (N_9530,N_9052,N_8755);
nand U9531 (N_9531,N_9197,N_9358);
nor U9532 (N_9532,N_8864,N_8848);
and U9533 (N_9533,N_9121,N_9031);
xnor U9534 (N_9534,N_9160,N_9243);
and U9535 (N_9535,N_9090,N_9216);
nor U9536 (N_9536,N_9108,N_8758);
nor U9537 (N_9537,N_9143,N_9355);
nand U9538 (N_9538,N_9190,N_8951);
and U9539 (N_9539,N_8771,N_8940);
nand U9540 (N_9540,N_9220,N_9206);
or U9541 (N_9541,N_8976,N_9083);
nor U9542 (N_9542,N_9006,N_9113);
xor U9543 (N_9543,N_8970,N_9116);
nor U9544 (N_9544,N_9286,N_9067);
xnor U9545 (N_9545,N_9252,N_9114);
xnor U9546 (N_9546,N_9146,N_8892);
and U9547 (N_9547,N_9084,N_8799);
nand U9548 (N_9548,N_9018,N_9064);
nor U9549 (N_9549,N_8769,N_9367);
or U9550 (N_9550,N_8788,N_9038);
nand U9551 (N_9551,N_9091,N_8973);
and U9552 (N_9552,N_9095,N_8798);
nand U9553 (N_9553,N_9257,N_8925);
or U9554 (N_9554,N_9266,N_9341);
or U9555 (N_9555,N_9010,N_8942);
xnor U9556 (N_9556,N_9078,N_9330);
xor U9557 (N_9557,N_9246,N_9129);
xnor U9558 (N_9558,N_8944,N_9229);
xor U9559 (N_9559,N_9186,N_9105);
and U9560 (N_9560,N_8808,N_9180);
nand U9561 (N_9561,N_8963,N_8760);
or U9562 (N_9562,N_9046,N_9023);
or U9563 (N_9563,N_9373,N_8885);
nor U9564 (N_9564,N_9109,N_8997);
and U9565 (N_9565,N_8888,N_9027);
and U9566 (N_9566,N_9334,N_9112);
and U9567 (N_9567,N_8979,N_8908);
nor U9568 (N_9568,N_8812,N_9352);
and U9569 (N_9569,N_8809,N_9176);
and U9570 (N_9570,N_8932,N_9158);
xor U9571 (N_9571,N_9265,N_9259);
xnor U9572 (N_9572,N_8913,N_8759);
and U9573 (N_9573,N_8971,N_9346);
nand U9574 (N_9574,N_9370,N_8950);
and U9575 (N_9575,N_9250,N_9296);
xor U9576 (N_9576,N_8842,N_9183);
nand U9577 (N_9577,N_9034,N_9025);
nor U9578 (N_9578,N_9089,N_8941);
nand U9579 (N_9579,N_9133,N_9208);
nor U9580 (N_9580,N_8968,N_8912);
and U9581 (N_9581,N_9037,N_9059);
nor U9582 (N_9582,N_9101,N_9165);
nand U9583 (N_9583,N_8982,N_9359);
or U9584 (N_9584,N_9057,N_8895);
nand U9585 (N_9585,N_9350,N_9122);
nor U9586 (N_9586,N_8915,N_9030);
xnor U9587 (N_9587,N_9149,N_9119);
and U9588 (N_9588,N_9007,N_9043);
nand U9589 (N_9589,N_9049,N_8824);
xor U9590 (N_9590,N_9294,N_9062);
nand U9591 (N_9591,N_9004,N_8933);
xnor U9592 (N_9592,N_9130,N_8983);
xor U9593 (N_9593,N_9268,N_8995);
and U9594 (N_9594,N_9360,N_8914);
or U9595 (N_9595,N_9068,N_9343);
and U9596 (N_9596,N_9245,N_9282);
or U9597 (N_9597,N_8854,N_9058);
nand U9598 (N_9598,N_9192,N_8778);
nand U9599 (N_9599,N_8839,N_8801);
nor U9600 (N_9600,N_9123,N_8881);
nand U9601 (N_9601,N_8901,N_8957);
and U9602 (N_9602,N_8960,N_9209);
nor U9603 (N_9603,N_8829,N_9217);
and U9604 (N_9604,N_9012,N_9242);
or U9605 (N_9605,N_9351,N_9094);
and U9606 (N_9606,N_8961,N_9085);
nor U9607 (N_9607,N_9124,N_9325);
and U9608 (N_9608,N_8906,N_9174);
xor U9609 (N_9609,N_9336,N_8922);
and U9610 (N_9610,N_9225,N_8899);
nand U9611 (N_9611,N_9040,N_9365);
nand U9612 (N_9612,N_8916,N_9097);
xnor U9613 (N_9613,N_9237,N_9218);
or U9614 (N_9614,N_8969,N_8860);
or U9615 (N_9615,N_9281,N_8991);
and U9616 (N_9616,N_9014,N_8907);
nand U9617 (N_9617,N_8873,N_8850);
and U9618 (N_9618,N_8753,N_9137);
nor U9619 (N_9619,N_9029,N_9171);
or U9620 (N_9620,N_9247,N_8946);
nand U9621 (N_9621,N_8879,N_9102);
nor U9622 (N_9622,N_9305,N_9235);
nand U9623 (N_9623,N_9234,N_9372);
and U9624 (N_9624,N_9207,N_9316);
xor U9625 (N_9625,N_9050,N_9195);
and U9626 (N_9626,N_9061,N_8898);
xnor U9627 (N_9627,N_8897,N_9256);
nand U9628 (N_9628,N_9299,N_9263);
nor U9629 (N_9629,N_8855,N_8884);
and U9630 (N_9630,N_8889,N_9166);
nor U9631 (N_9631,N_8786,N_9203);
xnor U9632 (N_9632,N_9227,N_9348);
nor U9633 (N_9633,N_9161,N_8807);
nor U9634 (N_9634,N_9026,N_9290);
xnor U9635 (N_9635,N_8877,N_9295);
nand U9636 (N_9636,N_8954,N_9238);
and U9637 (N_9637,N_9019,N_9013);
nor U9638 (N_9638,N_9276,N_9181);
nor U9639 (N_9639,N_9255,N_9261);
or U9640 (N_9640,N_9253,N_9279);
nand U9641 (N_9641,N_9236,N_9223);
nor U9642 (N_9642,N_8857,N_8987);
nand U9643 (N_9643,N_8821,N_8965);
nand U9644 (N_9644,N_9320,N_8972);
nor U9645 (N_9645,N_8868,N_8805);
and U9646 (N_9646,N_9118,N_8761);
nand U9647 (N_9647,N_9134,N_9022);
nor U9648 (N_9648,N_8978,N_9333);
xor U9649 (N_9649,N_8826,N_9262);
and U9650 (N_9650,N_9144,N_8797);
or U9651 (N_9651,N_8943,N_9003);
and U9652 (N_9652,N_8966,N_8823);
and U9653 (N_9653,N_9337,N_9309);
or U9654 (N_9654,N_9020,N_8999);
nor U9655 (N_9655,N_9039,N_9222);
xnor U9656 (N_9656,N_8939,N_9258);
nand U9657 (N_9657,N_9044,N_9154);
and U9658 (N_9658,N_8867,N_9076);
or U9659 (N_9659,N_9152,N_8870);
nor U9660 (N_9660,N_9126,N_8777);
and U9661 (N_9661,N_9232,N_9148);
xnor U9662 (N_9662,N_9151,N_9366);
xnor U9663 (N_9663,N_8930,N_8770);
and U9664 (N_9664,N_9187,N_8768);
nor U9665 (N_9665,N_8782,N_9120);
nor U9666 (N_9666,N_9017,N_9055);
nor U9667 (N_9667,N_9132,N_8911);
nand U9668 (N_9668,N_9104,N_9241);
and U9669 (N_9669,N_8859,N_9177);
nand U9670 (N_9670,N_9249,N_8894);
nor U9671 (N_9671,N_9331,N_8958);
and U9672 (N_9672,N_9292,N_9128);
xnor U9673 (N_9673,N_8775,N_9328);
or U9674 (N_9674,N_9318,N_8918);
nand U9675 (N_9675,N_9096,N_8779);
xor U9676 (N_9676,N_9269,N_8926);
xor U9677 (N_9677,N_9283,N_9036);
xor U9678 (N_9678,N_9354,N_9251);
nand U9679 (N_9679,N_8948,N_9080);
xor U9680 (N_9680,N_8843,N_8945);
and U9681 (N_9681,N_9215,N_8810);
nor U9682 (N_9682,N_8781,N_9210);
xor U9683 (N_9683,N_9344,N_9008);
and U9684 (N_9684,N_8815,N_8955);
xnor U9685 (N_9685,N_9280,N_8947);
and U9686 (N_9686,N_8996,N_9270);
nor U9687 (N_9687,N_9329,N_9101);
xor U9688 (N_9688,N_8878,N_8892);
nor U9689 (N_9689,N_9236,N_9185);
or U9690 (N_9690,N_8815,N_9181);
and U9691 (N_9691,N_9207,N_9029);
or U9692 (N_9692,N_8938,N_9136);
and U9693 (N_9693,N_8997,N_9127);
and U9694 (N_9694,N_9288,N_9336);
or U9695 (N_9695,N_8972,N_9277);
nor U9696 (N_9696,N_9226,N_9111);
and U9697 (N_9697,N_9087,N_8859);
nand U9698 (N_9698,N_9286,N_8883);
xnor U9699 (N_9699,N_9086,N_9294);
or U9700 (N_9700,N_8958,N_9155);
xnor U9701 (N_9701,N_9152,N_8886);
xor U9702 (N_9702,N_9338,N_8922);
nand U9703 (N_9703,N_8877,N_8757);
nor U9704 (N_9704,N_9121,N_9082);
or U9705 (N_9705,N_8996,N_8855);
xor U9706 (N_9706,N_9227,N_8787);
nor U9707 (N_9707,N_9111,N_9035);
nand U9708 (N_9708,N_9091,N_8873);
nand U9709 (N_9709,N_9245,N_9242);
xnor U9710 (N_9710,N_9053,N_9371);
nor U9711 (N_9711,N_9214,N_9019);
nand U9712 (N_9712,N_9048,N_8969);
xor U9713 (N_9713,N_9141,N_9018);
nor U9714 (N_9714,N_8976,N_9030);
xor U9715 (N_9715,N_8992,N_9167);
xnor U9716 (N_9716,N_9372,N_8976);
xnor U9717 (N_9717,N_9030,N_8993);
nor U9718 (N_9718,N_8761,N_8866);
nor U9719 (N_9719,N_9061,N_9078);
and U9720 (N_9720,N_8878,N_9177);
and U9721 (N_9721,N_8992,N_9373);
nand U9722 (N_9722,N_9202,N_9047);
nand U9723 (N_9723,N_8785,N_8944);
or U9724 (N_9724,N_8936,N_8922);
or U9725 (N_9725,N_9223,N_9161);
nand U9726 (N_9726,N_8997,N_9073);
and U9727 (N_9727,N_9207,N_9290);
nand U9728 (N_9728,N_9189,N_8823);
and U9729 (N_9729,N_9282,N_9084);
and U9730 (N_9730,N_9235,N_8973);
nand U9731 (N_9731,N_9250,N_9135);
xor U9732 (N_9732,N_8888,N_8863);
and U9733 (N_9733,N_8775,N_9138);
xor U9734 (N_9734,N_8872,N_8911);
nand U9735 (N_9735,N_8983,N_9211);
or U9736 (N_9736,N_8871,N_9371);
and U9737 (N_9737,N_8825,N_8918);
or U9738 (N_9738,N_8982,N_8813);
or U9739 (N_9739,N_9297,N_9268);
nor U9740 (N_9740,N_9268,N_8859);
and U9741 (N_9741,N_9270,N_9220);
nand U9742 (N_9742,N_9230,N_8950);
nor U9743 (N_9743,N_9154,N_8891);
nor U9744 (N_9744,N_9334,N_8949);
or U9745 (N_9745,N_9083,N_9135);
nand U9746 (N_9746,N_9158,N_9112);
nand U9747 (N_9747,N_8841,N_9191);
and U9748 (N_9748,N_8977,N_9349);
and U9749 (N_9749,N_9259,N_9241);
nand U9750 (N_9750,N_9325,N_8872);
xor U9751 (N_9751,N_9217,N_9241);
xor U9752 (N_9752,N_9225,N_9068);
and U9753 (N_9753,N_9372,N_9133);
or U9754 (N_9754,N_9307,N_9349);
xnor U9755 (N_9755,N_8825,N_9297);
nor U9756 (N_9756,N_8947,N_9279);
and U9757 (N_9757,N_8924,N_9319);
nor U9758 (N_9758,N_9300,N_9155);
and U9759 (N_9759,N_8894,N_9033);
nor U9760 (N_9760,N_8845,N_9030);
xnor U9761 (N_9761,N_9111,N_9215);
and U9762 (N_9762,N_9223,N_9309);
nor U9763 (N_9763,N_9302,N_8932);
nor U9764 (N_9764,N_8762,N_8898);
nand U9765 (N_9765,N_8826,N_9201);
nand U9766 (N_9766,N_9297,N_9172);
and U9767 (N_9767,N_8886,N_9124);
or U9768 (N_9768,N_8918,N_9178);
nor U9769 (N_9769,N_8809,N_9356);
and U9770 (N_9770,N_9081,N_9285);
nand U9771 (N_9771,N_9020,N_9124);
and U9772 (N_9772,N_8962,N_9010);
nor U9773 (N_9773,N_8861,N_9208);
and U9774 (N_9774,N_9168,N_9133);
nand U9775 (N_9775,N_8906,N_9199);
nor U9776 (N_9776,N_9131,N_8836);
nor U9777 (N_9777,N_8861,N_9227);
xor U9778 (N_9778,N_9299,N_8786);
and U9779 (N_9779,N_8875,N_9234);
and U9780 (N_9780,N_9176,N_8911);
nor U9781 (N_9781,N_9032,N_8754);
nand U9782 (N_9782,N_8909,N_8978);
nor U9783 (N_9783,N_8854,N_8999);
or U9784 (N_9784,N_9226,N_9355);
xnor U9785 (N_9785,N_9080,N_9171);
nor U9786 (N_9786,N_9013,N_9364);
or U9787 (N_9787,N_9322,N_8943);
or U9788 (N_9788,N_8834,N_8924);
nor U9789 (N_9789,N_8889,N_9331);
nor U9790 (N_9790,N_8954,N_8933);
or U9791 (N_9791,N_9114,N_9087);
or U9792 (N_9792,N_9354,N_8880);
and U9793 (N_9793,N_8999,N_8792);
or U9794 (N_9794,N_9350,N_9256);
nor U9795 (N_9795,N_8873,N_9368);
xnor U9796 (N_9796,N_9329,N_9016);
or U9797 (N_9797,N_9296,N_9161);
and U9798 (N_9798,N_9179,N_8850);
and U9799 (N_9799,N_8757,N_9215);
xnor U9800 (N_9800,N_9264,N_9221);
xor U9801 (N_9801,N_9245,N_9097);
xor U9802 (N_9802,N_9044,N_8918);
or U9803 (N_9803,N_9267,N_9104);
nand U9804 (N_9804,N_9056,N_9050);
nand U9805 (N_9805,N_9129,N_9145);
and U9806 (N_9806,N_8870,N_9352);
or U9807 (N_9807,N_8765,N_9066);
xnor U9808 (N_9808,N_9027,N_9326);
nor U9809 (N_9809,N_9090,N_9366);
nand U9810 (N_9810,N_9203,N_8852);
xor U9811 (N_9811,N_9333,N_9195);
nor U9812 (N_9812,N_9099,N_9096);
xnor U9813 (N_9813,N_9122,N_8859);
nand U9814 (N_9814,N_9157,N_9159);
and U9815 (N_9815,N_9287,N_8847);
nor U9816 (N_9816,N_9352,N_8756);
and U9817 (N_9817,N_9078,N_8759);
xnor U9818 (N_9818,N_9145,N_9293);
or U9819 (N_9819,N_9215,N_9145);
xnor U9820 (N_9820,N_9030,N_8814);
nand U9821 (N_9821,N_8753,N_8912);
and U9822 (N_9822,N_9045,N_8809);
or U9823 (N_9823,N_8907,N_9105);
nand U9824 (N_9824,N_9032,N_8903);
nand U9825 (N_9825,N_9038,N_9097);
nor U9826 (N_9826,N_9204,N_9218);
or U9827 (N_9827,N_8892,N_9248);
nand U9828 (N_9828,N_8849,N_8909);
and U9829 (N_9829,N_8842,N_8897);
nor U9830 (N_9830,N_9244,N_9044);
and U9831 (N_9831,N_9021,N_8895);
nand U9832 (N_9832,N_9335,N_8847);
and U9833 (N_9833,N_9342,N_9347);
xor U9834 (N_9834,N_9288,N_9071);
nor U9835 (N_9835,N_9112,N_9109);
nand U9836 (N_9836,N_9220,N_9338);
nor U9837 (N_9837,N_9209,N_8937);
xnor U9838 (N_9838,N_8763,N_8958);
and U9839 (N_9839,N_8948,N_8982);
nor U9840 (N_9840,N_8825,N_9090);
xor U9841 (N_9841,N_9011,N_9267);
xnor U9842 (N_9842,N_9112,N_9201);
nand U9843 (N_9843,N_8757,N_8945);
nor U9844 (N_9844,N_9109,N_8908);
and U9845 (N_9845,N_8951,N_9290);
and U9846 (N_9846,N_9113,N_8908);
xor U9847 (N_9847,N_8898,N_9297);
nand U9848 (N_9848,N_8822,N_8962);
or U9849 (N_9849,N_9273,N_9143);
nand U9850 (N_9850,N_8903,N_8971);
xnor U9851 (N_9851,N_8969,N_9287);
and U9852 (N_9852,N_8844,N_9083);
and U9853 (N_9853,N_9224,N_9168);
or U9854 (N_9854,N_8791,N_8906);
or U9855 (N_9855,N_8940,N_8912);
or U9856 (N_9856,N_8887,N_9326);
and U9857 (N_9857,N_9211,N_9009);
xnor U9858 (N_9858,N_8899,N_9273);
nand U9859 (N_9859,N_8773,N_8925);
nor U9860 (N_9860,N_9031,N_8770);
and U9861 (N_9861,N_8851,N_9029);
and U9862 (N_9862,N_9147,N_9326);
or U9863 (N_9863,N_8821,N_8943);
nand U9864 (N_9864,N_9111,N_8948);
nor U9865 (N_9865,N_8750,N_8945);
or U9866 (N_9866,N_9257,N_8787);
xnor U9867 (N_9867,N_9231,N_8969);
and U9868 (N_9868,N_8825,N_9298);
nand U9869 (N_9869,N_8861,N_9024);
nand U9870 (N_9870,N_9132,N_9301);
nand U9871 (N_9871,N_9347,N_9179);
or U9872 (N_9872,N_9354,N_9350);
nor U9873 (N_9873,N_9196,N_9117);
or U9874 (N_9874,N_9235,N_8981);
nor U9875 (N_9875,N_9258,N_9326);
or U9876 (N_9876,N_9059,N_9305);
nor U9877 (N_9877,N_8971,N_9010);
nor U9878 (N_9878,N_9074,N_9197);
nand U9879 (N_9879,N_9185,N_9359);
or U9880 (N_9880,N_8960,N_8826);
or U9881 (N_9881,N_9175,N_9124);
xor U9882 (N_9882,N_8872,N_8894);
nor U9883 (N_9883,N_9119,N_9009);
and U9884 (N_9884,N_9086,N_8954);
nand U9885 (N_9885,N_9108,N_9068);
xor U9886 (N_9886,N_8778,N_8814);
nor U9887 (N_9887,N_9073,N_8946);
and U9888 (N_9888,N_9219,N_8856);
nand U9889 (N_9889,N_8876,N_9151);
or U9890 (N_9890,N_8987,N_9269);
nor U9891 (N_9891,N_8974,N_8958);
nor U9892 (N_9892,N_9075,N_9216);
nand U9893 (N_9893,N_8791,N_9038);
and U9894 (N_9894,N_9062,N_9035);
xor U9895 (N_9895,N_9324,N_8761);
or U9896 (N_9896,N_9122,N_8958);
and U9897 (N_9897,N_9163,N_8948);
nor U9898 (N_9898,N_9136,N_9281);
xnor U9899 (N_9899,N_8976,N_8926);
or U9900 (N_9900,N_8794,N_9160);
nor U9901 (N_9901,N_9009,N_9270);
and U9902 (N_9902,N_9196,N_9063);
nand U9903 (N_9903,N_8970,N_8829);
xor U9904 (N_9904,N_8885,N_9039);
or U9905 (N_9905,N_9145,N_8793);
nor U9906 (N_9906,N_9191,N_8943);
or U9907 (N_9907,N_8920,N_9020);
xor U9908 (N_9908,N_9019,N_8942);
and U9909 (N_9909,N_8966,N_9209);
or U9910 (N_9910,N_8933,N_9124);
nand U9911 (N_9911,N_9037,N_9303);
xor U9912 (N_9912,N_8960,N_9002);
nor U9913 (N_9913,N_8908,N_9039);
nand U9914 (N_9914,N_9330,N_9152);
xor U9915 (N_9915,N_8805,N_9227);
nor U9916 (N_9916,N_8761,N_9156);
nand U9917 (N_9917,N_8852,N_9254);
xnor U9918 (N_9918,N_8756,N_8985);
nor U9919 (N_9919,N_9064,N_9057);
and U9920 (N_9920,N_9135,N_9125);
and U9921 (N_9921,N_8896,N_9134);
and U9922 (N_9922,N_8828,N_9108);
and U9923 (N_9923,N_9017,N_9206);
or U9924 (N_9924,N_9114,N_9158);
xor U9925 (N_9925,N_9017,N_9300);
xnor U9926 (N_9926,N_8900,N_8993);
nand U9927 (N_9927,N_9132,N_8810);
nor U9928 (N_9928,N_9050,N_8976);
or U9929 (N_9929,N_9267,N_8977);
nor U9930 (N_9930,N_9169,N_9062);
nand U9931 (N_9931,N_8949,N_8964);
or U9932 (N_9932,N_8848,N_8868);
nand U9933 (N_9933,N_9291,N_9237);
nand U9934 (N_9934,N_9322,N_8872);
nor U9935 (N_9935,N_8851,N_9065);
xor U9936 (N_9936,N_9109,N_9290);
and U9937 (N_9937,N_8930,N_9246);
or U9938 (N_9938,N_8950,N_9101);
or U9939 (N_9939,N_9049,N_8814);
or U9940 (N_9940,N_8836,N_9057);
or U9941 (N_9941,N_8767,N_8933);
nor U9942 (N_9942,N_9301,N_9357);
or U9943 (N_9943,N_8904,N_9138);
or U9944 (N_9944,N_9080,N_8819);
or U9945 (N_9945,N_9335,N_9117);
and U9946 (N_9946,N_8922,N_8820);
xnor U9947 (N_9947,N_9010,N_9140);
nand U9948 (N_9948,N_9356,N_9336);
and U9949 (N_9949,N_9169,N_9053);
or U9950 (N_9950,N_8840,N_9004);
or U9951 (N_9951,N_8932,N_8883);
and U9952 (N_9952,N_8784,N_9251);
or U9953 (N_9953,N_9310,N_9272);
nor U9954 (N_9954,N_9116,N_9224);
nor U9955 (N_9955,N_8929,N_9185);
nor U9956 (N_9956,N_8785,N_8961);
and U9957 (N_9957,N_8942,N_9023);
or U9958 (N_9958,N_9280,N_9087);
and U9959 (N_9959,N_8841,N_9091);
nor U9960 (N_9960,N_9020,N_9303);
xor U9961 (N_9961,N_8808,N_9183);
and U9962 (N_9962,N_8883,N_9216);
nand U9963 (N_9963,N_9041,N_9302);
xnor U9964 (N_9964,N_9068,N_9203);
and U9965 (N_9965,N_8963,N_9118);
nand U9966 (N_9966,N_9240,N_9003);
nor U9967 (N_9967,N_9182,N_8808);
nor U9968 (N_9968,N_8893,N_8913);
nor U9969 (N_9969,N_8908,N_8913);
xor U9970 (N_9970,N_9346,N_8759);
nor U9971 (N_9971,N_9145,N_9200);
or U9972 (N_9972,N_9028,N_9022);
xnor U9973 (N_9973,N_9072,N_9012);
and U9974 (N_9974,N_9340,N_9019);
xnor U9975 (N_9975,N_9208,N_9121);
and U9976 (N_9976,N_9328,N_8930);
xor U9977 (N_9977,N_8808,N_8782);
nor U9978 (N_9978,N_9205,N_9122);
xor U9979 (N_9979,N_9334,N_8858);
or U9980 (N_9980,N_9138,N_8794);
nor U9981 (N_9981,N_8841,N_9273);
or U9982 (N_9982,N_8889,N_8815);
and U9983 (N_9983,N_8820,N_9034);
and U9984 (N_9984,N_8947,N_9136);
xor U9985 (N_9985,N_8793,N_8878);
nand U9986 (N_9986,N_9235,N_8833);
or U9987 (N_9987,N_9073,N_8851);
and U9988 (N_9988,N_9114,N_8847);
and U9989 (N_9989,N_8887,N_8952);
nor U9990 (N_9990,N_9347,N_8907);
and U9991 (N_9991,N_8825,N_9091);
nor U9992 (N_9992,N_9266,N_9313);
nand U9993 (N_9993,N_9327,N_8800);
or U9994 (N_9994,N_8790,N_9277);
nand U9995 (N_9995,N_9208,N_8875);
and U9996 (N_9996,N_8757,N_9206);
xor U9997 (N_9997,N_9011,N_9348);
xnor U9998 (N_9998,N_9200,N_9339);
or U9999 (N_9999,N_9341,N_8979);
xor U10000 (N_10000,N_9833,N_9499);
or U10001 (N_10001,N_9970,N_9486);
nand U10002 (N_10002,N_9607,N_9450);
nand U10003 (N_10003,N_9581,N_9571);
nand U10004 (N_10004,N_9604,N_9826);
nand U10005 (N_10005,N_9477,N_9395);
xnor U10006 (N_10006,N_9967,N_9564);
and U10007 (N_10007,N_9965,N_9904);
nand U10008 (N_10008,N_9543,N_9753);
xnor U10009 (N_10009,N_9678,N_9404);
or U10010 (N_10010,N_9540,N_9768);
nand U10011 (N_10011,N_9628,N_9759);
nor U10012 (N_10012,N_9595,N_9929);
xor U10013 (N_10013,N_9875,N_9443);
nor U10014 (N_10014,N_9563,N_9415);
nand U10015 (N_10015,N_9862,N_9626);
nand U10016 (N_10016,N_9890,N_9547);
nand U10017 (N_10017,N_9987,N_9925);
nand U10018 (N_10018,N_9984,N_9602);
and U10019 (N_10019,N_9774,N_9732);
or U10020 (N_10020,N_9746,N_9534);
xnor U10021 (N_10021,N_9501,N_9658);
nor U10022 (N_10022,N_9898,N_9961);
xor U10023 (N_10023,N_9691,N_9418);
xor U10024 (N_10024,N_9428,N_9813);
nor U10025 (N_10025,N_9420,N_9682);
or U10026 (N_10026,N_9570,N_9684);
nor U10027 (N_10027,N_9951,N_9893);
nand U10028 (N_10028,N_9829,N_9432);
nor U10029 (N_10029,N_9757,N_9671);
nand U10030 (N_10030,N_9505,N_9489);
or U10031 (N_10031,N_9593,N_9895);
or U10032 (N_10032,N_9897,N_9990);
and U10033 (N_10033,N_9692,N_9778);
or U10034 (N_10034,N_9963,N_9407);
nor U10035 (N_10035,N_9905,N_9846);
nand U10036 (N_10036,N_9789,N_9780);
or U10037 (N_10037,N_9527,N_9726);
or U10038 (N_10038,N_9818,N_9456);
and U10039 (N_10039,N_9383,N_9594);
nor U10040 (N_10040,N_9988,N_9663);
nor U10041 (N_10041,N_9931,N_9569);
nor U10042 (N_10042,N_9971,N_9978);
or U10043 (N_10043,N_9464,N_9969);
or U10044 (N_10044,N_9831,N_9666);
nand U10045 (N_10045,N_9613,N_9400);
nand U10046 (N_10046,N_9561,N_9766);
nand U10047 (N_10047,N_9730,N_9565);
nor U10048 (N_10048,N_9463,N_9975);
nand U10049 (N_10049,N_9665,N_9655);
or U10050 (N_10050,N_9956,N_9530);
nand U10051 (N_10051,N_9474,N_9412);
and U10052 (N_10052,N_9492,N_9388);
and U10053 (N_10053,N_9508,N_9851);
or U10054 (N_10054,N_9745,N_9725);
and U10055 (N_10055,N_9762,N_9586);
nor U10056 (N_10056,N_9488,N_9957);
nor U10057 (N_10057,N_9502,N_9484);
nand U10058 (N_10058,N_9651,N_9389);
and U10059 (N_10059,N_9493,N_9381);
xor U10060 (N_10060,N_9913,N_9834);
nor U10061 (N_10061,N_9847,N_9782);
and U10062 (N_10062,N_9504,N_9932);
or U10063 (N_10063,N_9906,N_9601);
xnor U10064 (N_10064,N_9771,N_9703);
or U10065 (N_10065,N_9473,N_9427);
or U10066 (N_10066,N_9619,N_9770);
nand U10067 (N_10067,N_9668,N_9852);
xnor U10068 (N_10068,N_9809,N_9659);
nand U10069 (N_10069,N_9868,N_9618);
and U10070 (N_10070,N_9399,N_9724);
and U10071 (N_10071,N_9680,N_9924);
nor U10072 (N_10072,N_9424,N_9883);
nand U10073 (N_10073,N_9825,N_9958);
nor U10074 (N_10074,N_9927,N_9878);
or U10075 (N_10075,N_9838,N_9796);
nand U10076 (N_10076,N_9792,N_9396);
and U10077 (N_10077,N_9624,N_9806);
nor U10078 (N_10078,N_9576,N_9741);
and U10079 (N_10079,N_9882,N_9797);
nand U10080 (N_10080,N_9532,N_9814);
and U10081 (N_10081,N_9944,N_9977);
nand U10082 (N_10082,N_9920,N_9572);
and U10083 (N_10083,N_9791,N_9495);
nand U10084 (N_10084,N_9860,N_9476);
or U10085 (N_10085,N_9526,N_9794);
nor U10086 (N_10086,N_9661,N_9907);
xor U10087 (N_10087,N_9636,N_9445);
or U10088 (N_10088,N_9781,N_9981);
nand U10089 (N_10089,N_9616,N_9674);
nor U10090 (N_10090,N_9715,N_9550);
nor U10091 (N_10091,N_9717,N_9462);
and U10092 (N_10092,N_9598,N_9630);
nor U10093 (N_10093,N_9644,N_9740);
or U10094 (N_10094,N_9700,N_9475);
nand U10095 (N_10095,N_9437,N_9603);
nor U10096 (N_10096,N_9764,N_9631);
and U10097 (N_10097,N_9448,N_9800);
xnor U10098 (N_10098,N_9687,N_9386);
xnor U10099 (N_10099,N_9917,N_9683);
or U10100 (N_10100,N_9681,N_9954);
nand U10101 (N_10101,N_9888,N_9402);
and U10102 (N_10102,N_9544,N_9596);
and U10103 (N_10103,N_9719,N_9634);
and U10104 (N_10104,N_9694,N_9514);
or U10105 (N_10105,N_9449,N_9701);
nor U10106 (N_10106,N_9799,N_9994);
and U10107 (N_10107,N_9812,N_9537);
nor U10108 (N_10108,N_9894,N_9858);
or U10109 (N_10109,N_9410,N_9490);
xor U10110 (N_10110,N_9458,N_9417);
nand U10111 (N_10111,N_9664,N_9747);
nand U10112 (N_10112,N_9620,N_9454);
xnor U10113 (N_10113,N_9453,N_9699);
and U10114 (N_10114,N_9803,N_9704);
nand U10115 (N_10115,N_9845,N_9459);
and U10116 (N_10116,N_9784,N_9641);
nor U10117 (N_10117,N_9881,N_9714);
and U10118 (N_10118,N_9853,N_9436);
nand U10119 (N_10119,N_9506,N_9720);
nor U10120 (N_10120,N_9431,N_9478);
nor U10121 (N_10121,N_9708,N_9827);
xor U10122 (N_10122,N_9850,N_9621);
and U10123 (N_10123,N_9529,N_9891);
nor U10124 (N_10124,N_9541,N_9949);
nand U10125 (N_10125,N_9483,N_9980);
nand U10126 (N_10126,N_9640,N_9941);
or U10127 (N_10127,N_9836,N_9467);
nor U10128 (N_10128,N_9642,N_9440);
or U10129 (N_10129,N_9710,N_9997);
or U10130 (N_10130,N_9662,N_9556);
or U10131 (N_10131,N_9919,N_9837);
xor U10132 (N_10132,N_9752,N_9592);
or U10133 (N_10133,N_9999,N_9549);
xor U10134 (N_10134,N_9643,N_9646);
nand U10135 (N_10135,N_9817,N_9554);
and U10136 (N_10136,N_9401,N_9713);
or U10137 (N_10137,N_9657,N_9828);
xnor U10138 (N_10138,N_9783,N_9496);
nand U10139 (N_10139,N_9393,N_9545);
or U10140 (N_10140,N_9568,N_9785);
nor U10141 (N_10141,N_9937,N_9413);
nand U10142 (N_10142,N_9955,N_9712);
nand U10143 (N_10143,N_9938,N_9736);
nor U10144 (N_10144,N_9964,N_9871);
or U10145 (N_10145,N_9911,N_9481);
nand U10146 (N_10146,N_9434,N_9669);
nor U10147 (N_10147,N_9385,N_9989);
and U10148 (N_10148,N_9790,N_9756);
or U10149 (N_10149,N_9578,N_9697);
nor U10150 (N_10150,N_9709,N_9686);
nand U10151 (N_10151,N_9832,N_9900);
or U10152 (N_10152,N_9525,N_9579);
nor U10153 (N_10153,N_9482,N_9805);
xnor U10154 (N_10154,N_9749,N_9648);
nor U10155 (N_10155,N_9435,N_9652);
and U10156 (N_10156,N_9899,N_9728);
nor U10157 (N_10157,N_9562,N_9441);
xor U10158 (N_10158,N_9901,N_9439);
or U10159 (N_10159,N_9382,N_9754);
nand U10160 (N_10160,N_9972,N_9808);
or U10161 (N_10161,N_9469,N_9559);
nor U10162 (N_10162,N_9982,N_9419);
nor U10163 (N_10163,N_9429,N_9487);
and U10164 (N_10164,N_9468,N_9580);
xnor U10165 (N_10165,N_9926,N_9660);
nor U10166 (N_10166,N_9876,N_9597);
nand U10167 (N_10167,N_9654,N_9952);
xnor U10168 (N_10168,N_9821,N_9460);
or U10169 (N_10169,N_9688,N_9497);
nor U10170 (N_10170,N_9696,N_9776);
xor U10171 (N_10171,N_9535,N_9892);
nand U10172 (N_10172,N_9903,N_9423);
and U10173 (N_10173,N_9575,N_9908);
xor U10174 (N_10174,N_9479,N_9896);
xor U10175 (N_10175,N_9558,N_9416);
nor U10176 (N_10176,N_9810,N_9695);
and U10177 (N_10177,N_9509,N_9998);
and U10178 (N_10178,N_9380,N_9617);
xor U10179 (N_10179,N_9553,N_9748);
nor U10180 (N_10180,N_9976,N_9819);
nor U10181 (N_10181,N_9614,N_9974);
or U10182 (N_10182,N_9743,N_9472);
nand U10183 (N_10183,N_9447,N_9555);
or U10184 (N_10184,N_9645,N_9706);
or U10185 (N_10185,N_9933,N_9889);
nor U10186 (N_10186,N_9995,N_9992);
and U10187 (N_10187,N_9446,N_9722);
or U10188 (N_10188,N_9649,N_9676);
or U10189 (N_10189,N_9887,N_9507);
or U10190 (N_10190,N_9795,N_9962);
nand U10191 (N_10191,N_9914,N_9408);
nand U10192 (N_10192,N_9633,N_9874);
or U10193 (N_10193,N_9414,N_9873);
or U10194 (N_10194,N_9635,N_9584);
and U10195 (N_10195,N_9653,N_9779);
and U10196 (N_10196,N_9455,N_9582);
and U10197 (N_10197,N_9859,N_9566);
nor U10198 (N_10198,N_9379,N_9466);
and U10199 (N_10199,N_9375,N_9667);
nor U10200 (N_10200,N_9968,N_9909);
nor U10201 (N_10201,N_9915,N_9787);
nand U10202 (N_10202,N_9921,N_9936);
and U10203 (N_10203,N_9923,N_9793);
and U10204 (N_10204,N_9539,N_9711);
nand U10205 (N_10205,N_9823,N_9461);
or U10206 (N_10206,N_9639,N_9433);
nand U10207 (N_10207,N_9716,N_9879);
nor U10208 (N_10208,N_9376,N_9928);
nor U10209 (N_10209,N_9848,N_9991);
nand U10210 (N_10210,N_9811,N_9672);
xor U10211 (N_10211,N_9524,N_9528);
nor U10212 (N_10212,N_9629,N_9442);
and U10213 (N_10213,N_9996,N_9841);
xnor U10214 (N_10214,N_9538,N_9609);
or U10215 (N_10215,N_9993,N_9758);
nor U10216 (N_10216,N_9727,N_9480);
xor U10217 (N_10217,N_9839,N_9922);
nor U10218 (N_10218,N_9422,N_9930);
nand U10219 (N_10219,N_9542,N_9511);
xor U10220 (N_10220,N_9391,N_9677);
xnor U10221 (N_10221,N_9403,N_9767);
and U10222 (N_10222,N_9465,N_9503);
xor U10223 (N_10223,N_9548,N_9605);
nor U10224 (N_10224,N_9421,N_9470);
xnor U10225 (N_10225,N_9775,N_9471);
and U10226 (N_10226,N_9457,N_9405);
nand U10227 (N_10227,N_9761,N_9769);
nand U10228 (N_10228,N_9869,N_9590);
nand U10229 (N_10229,N_9986,N_9679);
nor U10230 (N_10230,N_9397,N_9411);
nand U10231 (N_10231,N_9721,N_9786);
nand U10232 (N_10232,N_9521,N_9392);
nor U10233 (N_10233,N_9409,N_9863);
nand U10234 (N_10234,N_9765,N_9650);
and U10235 (N_10235,N_9877,N_9567);
nor U10236 (N_10236,N_9546,N_9498);
or U10237 (N_10237,N_9606,N_9406);
or U10238 (N_10238,N_9512,N_9430);
and U10239 (N_10239,N_9425,N_9656);
nor U10240 (N_10240,N_9522,N_9934);
or U10241 (N_10241,N_9760,N_9788);
and U10242 (N_10242,N_9763,N_9918);
and U10243 (N_10243,N_9378,N_9485);
and U10244 (N_10244,N_9985,N_9739);
or U10245 (N_10245,N_9491,N_9815);
xor U10246 (N_10246,N_9557,N_9623);
nand U10247 (N_10247,N_9856,N_9777);
and U10248 (N_10248,N_9438,N_9885);
and U10249 (N_10249,N_9844,N_9599);
nand U10250 (N_10250,N_9520,N_9637);
and U10251 (N_10251,N_9690,N_9872);
xnor U10252 (N_10252,N_9772,N_9854);
xnor U10253 (N_10253,N_9750,N_9588);
or U10254 (N_10254,N_9519,N_9560);
and U10255 (N_10255,N_9517,N_9510);
xnor U10256 (N_10256,N_9959,N_9902);
xor U10257 (N_10257,N_9583,N_9723);
nand U10258 (N_10258,N_9835,N_9533);
and U10259 (N_10259,N_9622,N_9600);
and U10260 (N_10260,N_9820,N_9611);
or U10261 (N_10261,N_9531,N_9735);
nand U10262 (N_10262,N_9377,N_9802);
nand U10263 (N_10263,N_9855,N_9685);
xnor U10264 (N_10264,N_9864,N_9625);
nor U10265 (N_10265,N_9966,N_9807);
and U10266 (N_10266,N_9830,N_9494);
nand U10267 (N_10267,N_9946,N_9816);
nand U10268 (N_10268,N_9587,N_9870);
or U10269 (N_10269,N_9387,N_9612);
nand U10270 (N_10270,N_9647,N_9591);
or U10271 (N_10271,N_9733,N_9729);
xor U10272 (N_10272,N_9861,N_9577);
nor U10273 (N_10273,N_9773,N_9515);
xor U10274 (N_10274,N_9513,N_9950);
nand U10275 (N_10275,N_9500,N_9451);
xor U10276 (N_10276,N_9737,N_9536);
or U10277 (N_10277,N_9673,N_9983);
nand U10278 (N_10278,N_9865,N_9880);
or U10279 (N_10279,N_9574,N_9444);
nand U10280 (N_10280,N_9675,N_9973);
or U10281 (N_10281,N_9585,N_9670);
and U10282 (N_10282,N_9705,N_9693);
nand U10283 (N_10283,N_9940,N_9638);
nor U10284 (N_10284,N_9551,N_9948);
or U10285 (N_10285,N_9804,N_9615);
or U10286 (N_10286,N_9801,N_9943);
nor U10287 (N_10287,N_9912,N_9518);
xor U10288 (N_10288,N_9798,N_9866);
xnor U10289 (N_10289,N_9942,N_9718);
nand U10290 (N_10290,N_9384,N_9573);
and U10291 (N_10291,N_9632,N_9751);
and U10292 (N_10292,N_9945,N_9610);
nand U10293 (N_10293,N_9744,N_9390);
or U10294 (N_10294,N_9824,N_9822);
nand U10295 (N_10295,N_9867,N_9755);
or U10296 (N_10296,N_9939,N_9608);
nor U10297 (N_10297,N_9426,N_9589);
nor U10298 (N_10298,N_9516,N_9935);
nand U10299 (N_10299,N_9849,N_9857);
nand U10300 (N_10300,N_9916,N_9960);
or U10301 (N_10301,N_9886,N_9707);
nor U10302 (N_10302,N_9947,N_9523);
nor U10303 (N_10303,N_9627,N_9398);
nor U10304 (N_10304,N_9884,N_9843);
nand U10305 (N_10305,N_9731,N_9742);
nor U10306 (N_10306,N_9840,N_9910);
nand U10307 (N_10307,N_9394,N_9452);
and U10308 (N_10308,N_9979,N_9689);
or U10309 (N_10309,N_9953,N_9702);
nor U10310 (N_10310,N_9738,N_9552);
nor U10311 (N_10311,N_9698,N_9734);
xor U10312 (N_10312,N_9842,N_9521);
nand U10313 (N_10313,N_9595,N_9979);
xnor U10314 (N_10314,N_9928,N_9397);
xnor U10315 (N_10315,N_9547,N_9987);
nand U10316 (N_10316,N_9504,N_9458);
nor U10317 (N_10317,N_9840,N_9950);
or U10318 (N_10318,N_9897,N_9940);
and U10319 (N_10319,N_9962,N_9878);
nand U10320 (N_10320,N_9426,N_9692);
nand U10321 (N_10321,N_9482,N_9712);
xnor U10322 (N_10322,N_9453,N_9652);
xor U10323 (N_10323,N_9762,N_9452);
or U10324 (N_10324,N_9989,N_9927);
or U10325 (N_10325,N_9871,N_9480);
and U10326 (N_10326,N_9965,N_9822);
nor U10327 (N_10327,N_9527,N_9667);
nand U10328 (N_10328,N_9890,N_9576);
nand U10329 (N_10329,N_9656,N_9561);
and U10330 (N_10330,N_9988,N_9667);
or U10331 (N_10331,N_9441,N_9493);
and U10332 (N_10332,N_9810,N_9417);
or U10333 (N_10333,N_9600,N_9859);
xnor U10334 (N_10334,N_9478,N_9799);
nor U10335 (N_10335,N_9928,N_9578);
nor U10336 (N_10336,N_9877,N_9753);
nor U10337 (N_10337,N_9947,N_9737);
xor U10338 (N_10338,N_9523,N_9626);
nand U10339 (N_10339,N_9379,N_9977);
and U10340 (N_10340,N_9732,N_9961);
and U10341 (N_10341,N_9494,N_9540);
and U10342 (N_10342,N_9694,N_9695);
or U10343 (N_10343,N_9788,N_9385);
nor U10344 (N_10344,N_9841,N_9705);
and U10345 (N_10345,N_9950,N_9967);
nor U10346 (N_10346,N_9866,N_9822);
nor U10347 (N_10347,N_9724,N_9677);
xnor U10348 (N_10348,N_9398,N_9758);
or U10349 (N_10349,N_9895,N_9477);
nand U10350 (N_10350,N_9631,N_9469);
nand U10351 (N_10351,N_9796,N_9378);
xnor U10352 (N_10352,N_9714,N_9414);
and U10353 (N_10353,N_9601,N_9947);
and U10354 (N_10354,N_9594,N_9859);
nor U10355 (N_10355,N_9524,N_9943);
or U10356 (N_10356,N_9483,N_9393);
and U10357 (N_10357,N_9388,N_9675);
and U10358 (N_10358,N_9937,N_9644);
nor U10359 (N_10359,N_9992,N_9613);
xnor U10360 (N_10360,N_9681,N_9853);
nor U10361 (N_10361,N_9484,N_9438);
nor U10362 (N_10362,N_9926,N_9679);
xnor U10363 (N_10363,N_9503,N_9655);
xor U10364 (N_10364,N_9497,N_9397);
xor U10365 (N_10365,N_9842,N_9387);
nand U10366 (N_10366,N_9579,N_9691);
xor U10367 (N_10367,N_9466,N_9561);
and U10368 (N_10368,N_9611,N_9975);
and U10369 (N_10369,N_9504,N_9653);
or U10370 (N_10370,N_9694,N_9604);
nor U10371 (N_10371,N_9743,N_9403);
nand U10372 (N_10372,N_9648,N_9642);
or U10373 (N_10373,N_9470,N_9966);
xor U10374 (N_10374,N_9398,N_9837);
or U10375 (N_10375,N_9477,N_9481);
or U10376 (N_10376,N_9739,N_9693);
nor U10377 (N_10377,N_9666,N_9500);
xnor U10378 (N_10378,N_9779,N_9455);
or U10379 (N_10379,N_9512,N_9858);
nand U10380 (N_10380,N_9938,N_9871);
nand U10381 (N_10381,N_9836,N_9760);
nand U10382 (N_10382,N_9433,N_9507);
xor U10383 (N_10383,N_9840,N_9421);
and U10384 (N_10384,N_9796,N_9444);
or U10385 (N_10385,N_9405,N_9910);
and U10386 (N_10386,N_9874,N_9980);
and U10387 (N_10387,N_9990,N_9400);
xnor U10388 (N_10388,N_9749,N_9576);
and U10389 (N_10389,N_9823,N_9536);
nor U10390 (N_10390,N_9789,N_9617);
nand U10391 (N_10391,N_9885,N_9835);
xor U10392 (N_10392,N_9895,N_9891);
and U10393 (N_10393,N_9380,N_9787);
and U10394 (N_10394,N_9686,N_9598);
xnor U10395 (N_10395,N_9957,N_9609);
nand U10396 (N_10396,N_9694,N_9497);
xnor U10397 (N_10397,N_9927,N_9676);
or U10398 (N_10398,N_9648,N_9524);
nand U10399 (N_10399,N_9906,N_9658);
or U10400 (N_10400,N_9856,N_9700);
nor U10401 (N_10401,N_9613,N_9523);
and U10402 (N_10402,N_9912,N_9591);
or U10403 (N_10403,N_9926,N_9642);
nor U10404 (N_10404,N_9568,N_9551);
and U10405 (N_10405,N_9849,N_9789);
xnor U10406 (N_10406,N_9388,N_9599);
and U10407 (N_10407,N_9717,N_9451);
or U10408 (N_10408,N_9996,N_9505);
and U10409 (N_10409,N_9775,N_9473);
and U10410 (N_10410,N_9481,N_9955);
nor U10411 (N_10411,N_9635,N_9863);
and U10412 (N_10412,N_9511,N_9683);
and U10413 (N_10413,N_9535,N_9981);
nor U10414 (N_10414,N_9519,N_9434);
or U10415 (N_10415,N_9799,N_9516);
nand U10416 (N_10416,N_9882,N_9820);
or U10417 (N_10417,N_9712,N_9491);
and U10418 (N_10418,N_9805,N_9816);
nand U10419 (N_10419,N_9981,N_9652);
and U10420 (N_10420,N_9648,N_9402);
nor U10421 (N_10421,N_9433,N_9831);
nor U10422 (N_10422,N_9629,N_9518);
and U10423 (N_10423,N_9982,N_9847);
or U10424 (N_10424,N_9385,N_9474);
or U10425 (N_10425,N_9928,N_9799);
xnor U10426 (N_10426,N_9690,N_9480);
and U10427 (N_10427,N_9832,N_9750);
nor U10428 (N_10428,N_9735,N_9576);
nor U10429 (N_10429,N_9871,N_9743);
or U10430 (N_10430,N_9626,N_9528);
nor U10431 (N_10431,N_9510,N_9456);
or U10432 (N_10432,N_9991,N_9548);
or U10433 (N_10433,N_9725,N_9715);
and U10434 (N_10434,N_9881,N_9473);
nand U10435 (N_10435,N_9479,N_9857);
nand U10436 (N_10436,N_9720,N_9408);
or U10437 (N_10437,N_9759,N_9417);
nor U10438 (N_10438,N_9626,N_9462);
or U10439 (N_10439,N_9762,N_9612);
and U10440 (N_10440,N_9687,N_9776);
or U10441 (N_10441,N_9421,N_9931);
or U10442 (N_10442,N_9963,N_9980);
and U10443 (N_10443,N_9905,N_9454);
nand U10444 (N_10444,N_9949,N_9849);
nand U10445 (N_10445,N_9753,N_9794);
and U10446 (N_10446,N_9991,N_9441);
xnor U10447 (N_10447,N_9739,N_9650);
xnor U10448 (N_10448,N_9411,N_9534);
xnor U10449 (N_10449,N_9453,N_9752);
xor U10450 (N_10450,N_9422,N_9927);
nor U10451 (N_10451,N_9621,N_9487);
xnor U10452 (N_10452,N_9392,N_9670);
or U10453 (N_10453,N_9910,N_9861);
xor U10454 (N_10454,N_9400,N_9583);
xnor U10455 (N_10455,N_9613,N_9568);
or U10456 (N_10456,N_9425,N_9488);
xnor U10457 (N_10457,N_9771,N_9770);
and U10458 (N_10458,N_9877,N_9818);
or U10459 (N_10459,N_9877,N_9792);
nand U10460 (N_10460,N_9671,N_9916);
or U10461 (N_10461,N_9392,N_9746);
xor U10462 (N_10462,N_9903,N_9863);
xnor U10463 (N_10463,N_9795,N_9839);
and U10464 (N_10464,N_9931,N_9714);
and U10465 (N_10465,N_9462,N_9902);
xor U10466 (N_10466,N_9447,N_9931);
nor U10467 (N_10467,N_9497,N_9437);
and U10468 (N_10468,N_9389,N_9429);
and U10469 (N_10469,N_9808,N_9863);
nor U10470 (N_10470,N_9386,N_9458);
and U10471 (N_10471,N_9738,N_9416);
nor U10472 (N_10472,N_9503,N_9697);
and U10473 (N_10473,N_9506,N_9664);
xnor U10474 (N_10474,N_9824,N_9682);
nand U10475 (N_10475,N_9472,N_9547);
nand U10476 (N_10476,N_9726,N_9667);
nor U10477 (N_10477,N_9719,N_9539);
nor U10478 (N_10478,N_9918,N_9903);
xor U10479 (N_10479,N_9996,N_9506);
and U10480 (N_10480,N_9801,N_9987);
xor U10481 (N_10481,N_9591,N_9405);
and U10482 (N_10482,N_9871,N_9758);
nand U10483 (N_10483,N_9539,N_9485);
or U10484 (N_10484,N_9398,N_9545);
xor U10485 (N_10485,N_9759,N_9825);
nor U10486 (N_10486,N_9671,N_9434);
or U10487 (N_10487,N_9392,N_9609);
nor U10488 (N_10488,N_9385,N_9538);
nor U10489 (N_10489,N_9920,N_9928);
xnor U10490 (N_10490,N_9956,N_9463);
nor U10491 (N_10491,N_9588,N_9419);
and U10492 (N_10492,N_9823,N_9546);
nand U10493 (N_10493,N_9720,N_9561);
xnor U10494 (N_10494,N_9823,N_9449);
or U10495 (N_10495,N_9838,N_9485);
nand U10496 (N_10496,N_9838,N_9594);
or U10497 (N_10497,N_9671,N_9894);
and U10498 (N_10498,N_9449,N_9868);
nand U10499 (N_10499,N_9815,N_9690);
or U10500 (N_10500,N_9709,N_9646);
and U10501 (N_10501,N_9567,N_9951);
or U10502 (N_10502,N_9958,N_9882);
nor U10503 (N_10503,N_9645,N_9541);
xnor U10504 (N_10504,N_9826,N_9859);
nand U10505 (N_10505,N_9461,N_9900);
xor U10506 (N_10506,N_9714,N_9547);
nor U10507 (N_10507,N_9760,N_9620);
nor U10508 (N_10508,N_9548,N_9877);
or U10509 (N_10509,N_9438,N_9417);
nand U10510 (N_10510,N_9746,N_9601);
and U10511 (N_10511,N_9688,N_9979);
or U10512 (N_10512,N_9493,N_9455);
xnor U10513 (N_10513,N_9547,N_9833);
and U10514 (N_10514,N_9879,N_9965);
nor U10515 (N_10515,N_9911,N_9654);
or U10516 (N_10516,N_9953,N_9630);
nand U10517 (N_10517,N_9490,N_9476);
nand U10518 (N_10518,N_9617,N_9929);
or U10519 (N_10519,N_9862,N_9802);
or U10520 (N_10520,N_9619,N_9846);
xnor U10521 (N_10521,N_9644,N_9710);
nor U10522 (N_10522,N_9405,N_9713);
nor U10523 (N_10523,N_9485,N_9849);
nand U10524 (N_10524,N_9905,N_9894);
nand U10525 (N_10525,N_9385,N_9825);
or U10526 (N_10526,N_9380,N_9857);
and U10527 (N_10527,N_9611,N_9731);
xnor U10528 (N_10528,N_9583,N_9962);
xnor U10529 (N_10529,N_9834,N_9549);
or U10530 (N_10530,N_9506,N_9829);
nand U10531 (N_10531,N_9768,N_9844);
and U10532 (N_10532,N_9856,N_9512);
or U10533 (N_10533,N_9912,N_9724);
nand U10534 (N_10534,N_9414,N_9582);
and U10535 (N_10535,N_9987,N_9973);
nand U10536 (N_10536,N_9813,N_9465);
or U10537 (N_10537,N_9630,N_9376);
nand U10538 (N_10538,N_9867,N_9694);
nand U10539 (N_10539,N_9872,N_9998);
xnor U10540 (N_10540,N_9680,N_9687);
nand U10541 (N_10541,N_9718,N_9564);
and U10542 (N_10542,N_9759,N_9410);
or U10543 (N_10543,N_9739,N_9957);
nand U10544 (N_10544,N_9437,N_9402);
nand U10545 (N_10545,N_9945,N_9792);
and U10546 (N_10546,N_9619,N_9808);
nor U10547 (N_10547,N_9689,N_9882);
and U10548 (N_10548,N_9720,N_9826);
xor U10549 (N_10549,N_9469,N_9820);
and U10550 (N_10550,N_9389,N_9465);
or U10551 (N_10551,N_9808,N_9763);
or U10552 (N_10552,N_9920,N_9556);
and U10553 (N_10553,N_9842,N_9817);
and U10554 (N_10554,N_9808,N_9470);
xnor U10555 (N_10555,N_9616,N_9682);
nand U10556 (N_10556,N_9728,N_9923);
nand U10557 (N_10557,N_9805,N_9977);
nor U10558 (N_10558,N_9393,N_9757);
or U10559 (N_10559,N_9873,N_9613);
and U10560 (N_10560,N_9908,N_9624);
and U10561 (N_10561,N_9924,N_9704);
xnor U10562 (N_10562,N_9678,N_9727);
nand U10563 (N_10563,N_9946,N_9712);
nand U10564 (N_10564,N_9628,N_9622);
nor U10565 (N_10565,N_9857,N_9591);
nor U10566 (N_10566,N_9472,N_9463);
or U10567 (N_10567,N_9567,N_9494);
xnor U10568 (N_10568,N_9662,N_9978);
or U10569 (N_10569,N_9457,N_9869);
or U10570 (N_10570,N_9382,N_9971);
nand U10571 (N_10571,N_9405,N_9550);
or U10572 (N_10572,N_9930,N_9650);
nor U10573 (N_10573,N_9389,N_9704);
nor U10574 (N_10574,N_9571,N_9646);
nor U10575 (N_10575,N_9554,N_9957);
xnor U10576 (N_10576,N_9828,N_9857);
nand U10577 (N_10577,N_9483,N_9707);
nand U10578 (N_10578,N_9786,N_9619);
nand U10579 (N_10579,N_9513,N_9841);
and U10580 (N_10580,N_9616,N_9854);
or U10581 (N_10581,N_9577,N_9515);
xnor U10582 (N_10582,N_9602,N_9776);
nor U10583 (N_10583,N_9493,N_9426);
nor U10584 (N_10584,N_9759,N_9758);
nor U10585 (N_10585,N_9716,N_9883);
nand U10586 (N_10586,N_9550,N_9523);
nor U10587 (N_10587,N_9970,N_9902);
or U10588 (N_10588,N_9426,N_9393);
xnor U10589 (N_10589,N_9694,N_9984);
nor U10590 (N_10590,N_9940,N_9545);
nor U10591 (N_10591,N_9783,N_9520);
xor U10592 (N_10592,N_9751,N_9799);
nand U10593 (N_10593,N_9624,N_9586);
nor U10594 (N_10594,N_9675,N_9745);
and U10595 (N_10595,N_9621,N_9983);
xnor U10596 (N_10596,N_9506,N_9432);
nor U10597 (N_10597,N_9858,N_9897);
xnor U10598 (N_10598,N_9454,N_9996);
xor U10599 (N_10599,N_9607,N_9993);
nor U10600 (N_10600,N_9517,N_9740);
nor U10601 (N_10601,N_9434,N_9565);
and U10602 (N_10602,N_9560,N_9989);
and U10603 (N_10603,N_9986,N_9902);
and U10604 (N_10604,N_9384,N_9563);
or U10605 (N_10605,N_9960,N_9554);
and U10606 (N_10606,N_9871,N_9892);
or U10607 (N_10607,N_9671,N_9971);
nor U10608 (N_10608,N_9765,N_9885);
or U10609 (N_10609,N_9629,N_9440);
nor U10610 (N_10610,N_9441,N_9766);
nand U10611 (N_10611,N_9477,N_9713);
nand U10612 (N_10612,N_9725,N_9716);
or U10613 (N_10613,N_9814,N_9816);
and U10614 (N_10614,N_9420,N_9473);
xor U10615 (N_10615,N_9756,N_9814);
or U10616 (N_10616,N_9395,N_9419);
nand U10617 (N_10617,N_9438,N_9447);
nor U10618 (N_10618,N_9931,N_9892);
or U10619 (N_10619,N_9793,N_9386);
and U10620 (N_10620,N_9600,N_9375);
nand U10621 (N_10621,N_9889,N_9567);
and U10622 (N_10622,N_9384,N_9969);
or U10623 (N_10623,N_9492,N_9394);
or U10624 (N_10624,N_9556,N_9517);
and U10625 (N_10625,N_10164,N_10222);
nand U10626 (N_10626,N_10409,N_10534);
or U10627 (N_10627,N_10444,N_10615);
and U10628 (N_10628,N_10330,N_10600);
xnor U10629 (N_10629,N_10249,N_10064);
or U10630 (N_10630,N_10225,N_10036);
or U10631 (N_10631,N_10583,N_10536);
nand U10632 (N_10632,N_10071,N_10176);
and U10633 (N_10633,N_10174,N_10067);
or U10634 (N_10634,N_10013,N_10492);
nand U10635 (N_10635,N_10120,N_10396);
or U10636 (N_10636,N_10541,N_10196);
or U10637 (N_10637,N_10571,N_10488);
nor U10638 (N_10638,N_10066,N_10579);
or U10639 (N_10639,N_10292,N_10574);
xor U10640 (N_10640,N_10234,N_10267);
nand U10641 (N_10641,N_10148,N_10135);
or U10642 (N_10642,N_10158,N_10080);
xor U10643 (N_10643,N_10549,N_10086);
or U10644 (N_10644,N_10075,N_10026);
and U10645 (N_10645,N_10326,N_10424);
nor U10646 (N_10646,N_10531,N_10042);
or U10647 (N_10647,N_10498,N_10096);
nor U10648 (N_10648,N_10505,N_10493);
nand U10649 (N_10649,N_10281,N_10261);
nand U10650 (N_10650,N_10320,N_10394);
nand U10651 (N_10651,N_10468,N_10475);
xor U10652 (N_10652,N_10608,N_10489);
nand U10653 (N_10653,N_10291,N_10322);
xor U10654 (N_10654,N_10464,N_10461);
or U10655 (N_10655,N_10348,N_10278);
and U10656 (N_10656,N_10374,N_10573);
or U10657 (N_10657,N_10430,N_10546);
or U10658 (N_10658,N_10392,N_10597);
and U10659 (N_10659,N_10051,N_10177);
and U10660 (N_10660,N_10443,N_10325);
nand U10661 (N_10661,N_10271,N_10366);
and U10662 (N_10662,N_10074,N_10447);
nand U10663 (N_10663,N_10437,N_10308);
or U10664 (N_10664,N_10577,N_10385);
xnor U10665 (N_10665,N_10124,N_10091);
nor U10666 (N_10666,N_10083,N_10060);
nand U10667 (N_10667,N_10545,N_10016);
or U10668 (N_10668,N_10250,N_10204);
nor U10669 (N_10669,N_10300,N_10045);
nor U10670 (N_10670,N_10119,N_10537);
and U10671 (N_10671,N_10128,N_10034);
or U10672 (N_10672,N_10215,N_10359);
xor U10673 (N_10673,N_10479,N_10340);
or U10674 (N_10674,N_10205,N_10237);
xnor U10675 (N_10675,N_10193,N_10252);
or U10676 (N_10676,N_10092,N_10155);
or U10677 (N_10677,N_10570,N_10024);
xor U10678 (N_10678,N_10483,N_10514);
or U10679 (N_10679,N_10232,N_10547);
xnor U10680 (N_10680,N_10001,N_10548);
nor U10681 (N_10681,N_10018,N_10550);
nor U10682 (N_10682,N_10360,N_10065);
and U10683 (N_10683,N_10185,N_10414);
nor U10684 (N_10684,N_10527,N_10460);
nand U10685 (N_10685,N_10353,N_10207);
nor U10686 (N_10686,N_10298,N_10614);
xnor U10687 (N_10687,N_10616,N_10401);
or U10688 (N_10688,N_10059,N_10596);
xor U10689 (N_10689,N_10297,N_10442);
xnor U10690 (N_10690,N_10568,N_10469);
nand U10691 (N_10691,N_10180,N_10594);
nand U10692 (N_10692,N_10603,N_10429);
and U10693 (N_10693,N_10313,N_10287);
nand U10694 (N_10694,N_10613,N_10317);
xor U10695 (N_10695,N_10288,N_10258);
xnor U10696 (N_10696,N_10318,N_10482);
or U10697 (N_10697,N_10395,N_10111);
xnor U10698 (N_10698,N_10099,N_10110);
or U10699 (N_10699,N_10123,N_10587);
and U10700 (N_10700,N_10147,N_10463);
and U10701 (N_10701,N_10428,N_10166);
xnor U10702 (N_10702,N_10139,N_10520);
and U10703 (N_10703,N_10262,N_10380);
xnor U10704 (N_10704,N_10049,N_10303);
xor U10705 (N_10705,N_10585,N_10364);
and U10706 (N_10706,N_10019,N_10542);
nor U10707 (N_10707,N_10555,N_10199);
or U10708 (N_10708,N_10529,N_10617);
and U10709 (N_10709,N_10077,N_10312);
nand U10710 (N_10710,N_10612,N_10211);
nor U10711 (N_10711,N_10253,N_10324);
nor U10712 (N_10712,N_10143,N_10150);
nor U10713 (N_10713,N_10333,N_10566);
xnor U10714 (N_10714,N_10512,N_10445);
xor U10715 (N_10715,N_10532,N_10623);
nor U10716 (N_10716,N_10336,N_10495);
nand U10717 (N_10717,N_10456,N_10501);
nand U10718 (N_10718,N_10126,N_10112);
or U10719 (N_10719,N_10089,N_10040);
nor U10720 (N_10720,N_10522,N_10131);
nand U10721 (N_10721,N_10478,N_10342);
nand U10722 (N_10722,N_10470,N_10053);
nand U10723 (N_10723,N_10393,N_10524);
and U10724 (N_10724,N_10104,N_10384);
nand U10725 (N_10725,N_10552,N_10163);
xor U10726 (N_10726,N_10179,N_10423);
xor U10727 (N_10727,N_10419,N_10358);
or U10728 (N_10728,N_10029,N_10233);
nor U10729 (N_10729,N_10219,N_10014);
nand U10730 (N_10730,N_10153,N_10408);
or U10731 (N_10731,N_10149,N_10012);
nor U10732 (N_10732,N_10102,N_10416);
nor U10733 (N_10733,N_10356,N_10343);
nor U10734 (N_10734,N_10210,N_10285);
or U10735 (N_10735,N_10457,N_10523);
or U10736 (N_10736,N_10004,N_10236);
nand U10737 (N_10737,N_10455,N_10076);
xor U10738 (N_10738,N_10321,N_10008);
and U10739 (N_10739,N_10011,N_10589);
nor U10740 (N_10740,N_10183,N_10269);
nor U10741 (N_10741,N_10251,N_10095);
nand U10742 (N_10742,N_10412,N_10432);
or U10743 (N_10743,N_10376,N_10454);
and U10744 (N_10744,N_10165,N_10159);
xnor U10745 (N_10745,N_10068,N_10404);
xor U10746 (N_10746,N_10553,N_10473);
and U10747 (N_10747,N_10097,N_10031);
and U10748 (N_10748,N_10256,N_10239);
or U10749 (N_10749,N_10050,N_10306);
nor U10750 (N_10750,N_10030,N_10338);
nand U10751 (N_10751,N_10494,N_10178);
or U10752 (N_10752,N_10441,N_10244);
nor U10753 (N_10753,N_10301,N_10103);
nor U10754 (N_10754,N_10508,N_10000);
nor U10755 (N_10755,N_10094,N_10586);
xor U10756 (N_10756,N_10341,N_10216);
and U10757 (N_10757,N_10304,N_10369);
or U10758 (N_10758,N_10069,N_10381);
nand U10759 (N_10759,N_10611,N_10604);
nand U10760 (N_10760,N_10388,N_10551);
and U10761 (N_10761,N_10472,N_10184);
or U10762 (N_10762,N_10602,N_10487);
xor U10763 (N_10763,N_10310,N_10363);
nand U10764 (N_10764,N_10228,N_10367);
nor U10765 (N_10765,N_10593,N_10476);
nand U10766 (N_10766,N_10323,N_10302);
or U10767 (N_10767,N_10161,N_10521);
nor U10768 (N_10768,N_10515,N_10117);
xor U10769 (N_10769,N_10023,N_10564);
and U10770 (N_10770,N_10160,N_10209);
nor U10771 (N_10771,N_10349,N_10020);
nand U10772 (N_10772,N_10450,N_10328);
nor U10773 (N_10773,N_10466,N_10339);
and U10774 (N_10774,N_10506,N_10263);
nand U10775 (N_10775,N_10499,N_10538);
nand U10776 (N_10776,N_10197,N_10544);
nor U10777 (N_10777,N_10195,N_10079);
nand U10778 (N_10778,N_10191,N_10061);
and U10779 (N_10779,N_10332,N_10130);
nand U10780 (N_10780,N_10418,N_10295);
or U10781 (N_10781,N_10151,N_10556);
or U10782 (N_10782,N_10025,N_10425);
or U10783 (N_10783,N_10471,N_10224);
xor U10784 (N_10784,N_10055,N_10557);
or U10785 (N_10785,N_10462,N_10115);
nand U10786 (N_10786,N_10560,N_10052);
and U10787 (N_10787,N_10398,N_10279);
or U10788 (N_10788,N_10081,N_10144);
nand U10789 (N_10789,N_10214,N_10563);
or U10790 (N_10790,N_10280,N_10235);
and U10791 (N_10791,N_10022,N_10543);
xor U10792 (N_10792,N_10352,N_10006);
xor U10793 (N_10793,N_10203,N_10386);
nor U10794 (N_10794,N_10426,N_10569);
or U10795 (N_10795,N_10427,N_10605);
nand U10796 (N_10796,N_10518,N_10109);
or U10797 (N_10797,N_10175,N_10435);
and U10798 (N_10798,N_10403,N_10245);
xor U10799 (N_10799,N_10167,N_10129);
and U10800 (N_10800,N_10516,N_10098);
xnor U10801 (N_10801,N_10491,N_10397);
nor U10802 (N_10802,N_10265,N_10351);
or U10803 (N_10803,N_10005,N_10345);
xor U10804 (N_10804,N_10503,N_10584);
and U10805 (N_10805,N_10504,N_10255);
and U10806 (N_10806,N_10226,N_10609);
xor U10807 (N_10807,N_10477,N_10361);
and U10808 (N_10808,N_10347,N_10156);
and U10809 (N_10809,N_10186,N_10433);
and U10810 (N_10810,N_10519,N_10284);
or U10811 (N_10811,N_10474,N_10282);
and U10812 (N_10812,N_10459,N_10411);
xor U10813 (N_10813,N_10192,N_10598);
or U10814 (N_10814,N_10276,N_10277);
nor U10815 (N_10815,N_10422,N_10171);
xnor U10816 (N_10816,N_10283,N_10290);
or U10817 (N_10817,N_10554,N_10062);
and U10818 (N_10818,N_10043,N_10315);
and U10819 (N_10819,N_10314,N_10619);
xor U10820 (N_10820,N_10572,N_10621);
and U10821 (N_10821,N_10558,N_10057);
or U10822 (N_10822,N_10188,N_10595);
or U10823 (N_10823,N_10122,N_10389);
nor U10824 (N_10824,N_10327,N_10046);
nand U10825 (N_10825,N_10223,N_10116);
nor U10826 (N_10826,N_10382,N_10420);
xnor U10827 (N_10827,N_10449,N_10257);
or U10828 (N_10828,N_10041,N_10017);
xor U10829 (N_10829,N_10421,N_10350);
nand U10830 (N_10830,N_10507,N_10480);
and U10831 (N_10831,N_10434,N_10208);
nor U10832 (N_10832,N_10132,N_10481);
nor U10833 (N_10833,N_10243,N_10073);
nor U10834 (N_10834,N_10375,N_10142);
nand U10835 (N_10835,N_10458,N_10200);
or U10836 (N_10836,N_10490,N_10502);
nor U10837 (N_10837,N_10198,N_10329);
and U10838 (N_10838,N_10113,N_10357);
and U10839 (N_10839,N_10599,N_10294);
nor U10840 (N_10840,N_10344,N_10168);
and U10841 (N_10841,N_10513,N_10436);
nand U10842 (N_10842,N_10540,N_10446);
nand U10843 (N_10843,N_10453,N_10582);
nor U10844 (N_10844,N_10248,N_10334);
nor U10845 (N_10845,N_10189,N_10610);
nor U10846 (N_10846,N_10133,N_10108);
nor U10847 (N_10847,N_10264,N_10181);
or U10848 (N_10848,N_10335,N_10173);
or U10849 (N_10849,N_10268,N_10134);
and U10850 (N_10850,N_10009,N_10511);
or U10851 (N_10851,N_10090,N_10027);
and U10852 (N_10852,N_10274,N_10624);
nand U10853 (N_10853,N_10035,N_10368);
nand U10854 (N_10854,N_10247,N_10601);
or U10855 (N_10855,N_10202,N_10525);
nand U10856 (N_10856,N_10390,N_10377);
or U10857 (N_10857,N_10530,N_10141);
or U10858 (N_10858,N_10561,N_10154);
and U10859 (N_10859,N_10606,N_10137);
xnor U10860 (N_10860,N_10362,N_10145);
nor U10861 (N_10861,N_10170,N_10127);
xor U10862 (N_10862,N_10319,N_10213);
and U10863 (N_10863,N_10093,N_10015);
and U10864 (N_10864,N_10565,N_10270);
and U10865 (N_10865,N_10162,N_10227);
xnor U10866 (N_10866,N_10497,N_10106);
or U10867 (N_10867,N_10048,N_10286);
xor U10868 (N_10868,N_10365,N_10010);
nor U10869 (N_10869,N_10088,N_10407);
nor U10870 (N_10870,N_10033,N_10372);
and U10871 (N_10871,N_10438,N_10187);
xor U10872 (N_10872,N_10331,N_10509);
nor U10873 (N_10873,N_10138,N_10405);
and U10874 (N_10874,N_10379,N_10229);
nand U10875 (N_10875,N_10212,N_10622);
nand U10876 (N_10876,N_10273,N_10201);
nand U10877 (N_10877,N_10576,N_10539);
xnor U10878 (N_10878,N_10528,N_10221);
and U10879 (N_10879,N_10305,N_10535);
and U10880 (N_10880,N_10039,N_10021);
or U10881 (N_10881,N_10242,N_10559);
nand U10882 (N_10882,N_10580,N_10087);
nand U10883 (N_10883,N_10496,N_10581);
nand U10884 (N_10884,N_10410,N_10114);
or U10885 (N_10885,N_10440,N_10002);
and U10886 (N_10886,N_10220,N_10070);
and U10887 (N_10887,N_10607,N_10452);
and U10888 (N_10888,N_10620,N_10378);
and U10889 (N_10889,N_10590,N_10371);
nor U10890 (N_10890,N_10417,N_10575);
xnor U10891 (N_10891,N_10406,N_10231);
nor U10892 (N_10892,N_10084,N_10309);
and U10893 (N_10893,N_10217,N_10299);
xnor U10894 (N_10894,N_10238,N_10240);
or U10895 (N_10895,N_10439,N_10346);
xor U10896 (N_10896,N_10260,N_10485);
xnor U10897 (N_10897,N_10063,N_10078);
and U10898 (N_10898,N_10275,N_10467);
or U10899 (N_10899,N_10038,N_10044);
nand U10900 (N_10900,N_10028,N_10451);
or U10901 (N_10901,N_10391,N_10272);
xnor U10902 (N_10902,N_10157,N_10056);
or U10903 (N_10903,N_10105,N_10289);
xor U10904 (N_10904,N_10591,N_10431);
or U10905 (N_10905,N_10413,N_10293);
xor U10906 (N_10906,N_10003,N_10383);
nor U10907 (N_10907,N_10121,N_10307);
or U10908 (N_10908,N_10387,N_10533);
nand U10909 (N_10909,N_10246,N_10500);
nand U10910 (N_10910,N_10190,N_10588);
nand U10911 (N_10911,N_10136,N_10047);
or U10912 (N_10912,N_10402,N_10567);
nand U10913 (N_10913,N_10007,N_10241);
nand U10914 (N_10914,N_10316,N_10072);
xnor U10915 (N_10915,N_10296,N_10218);
or U10916 (N_10916,N_10259,N_10169);
nand U10917 (N_10917,N_10517,N_10254);
or U10918 (N_10918,N_10118,N_10152);
or U10919 (N_10919,N_10592,N_10037);
xnor U10920 (N_10920,N_10182,N_10526);
nand U10921 (N_10921,N_10415,N_10194);
xnor U10922 (N_10922,N_10146,N_10354);
and U10923 (N_10923,N_10578,N_10370);
xnor U10924 (N_10924,N_10101,N_10100);
nor U10925 (N_10925,N_10400,N_10486);
and U10926 (N_10926,N_10562,N_10484);
nor U10927 (N_10927,N_10510,N_10085);
and U10928 (N_10928,N_10140,N_10230);
and U10929 (N_10929,N_10058,N_10082);
nand U10930 (N_10930,N_10618,N_10355);
nand U10931 (N_10931,N_10399,N_10125);
xnor U10932 (N_10932,N_10311,N_10448);
and U10933 (N_10933,N_10337,N_10107);
xor U10934 (N_10934,N_10032,N_10054);
or U10935 (N_10935,N_10266,N_10172);
or U10936 (N_10936,N_10206,N_10373);
or U10937 (N_10937,N_10465,N_10226);
xor U10938 (N_10938,N_10382,N_10388);
nor U10939 (N_10939,N_10043,N_10221);
nand U10940 (N_10940,N_10511,N_10237);
and U10941 (N_10941,N_10482,N_10071);
nand U10942 (N_10942,N_10130,N_10335);
or U10943 (N_10943,N_10466,N_10485);
nor U10944 (N_10944,N_10122,N_10195);
nand U10945 (N_10945,N_10615,N_10386);
and U10946 (N_10946,N_10018,N_10160);
xor U10947 (N_10947,N_10035,N_10456);
and U10948 (N_10948,N_10336,N_10083);
nand U10949 (N_10949,N_10324,N_10018);
xor U10950 (N_10950,N_10484,N_10104);
nand U10951 (N_10951,N_10024,N_10539);
xor U10952 (N_10952,N_10069,N_10039);
or U10953 (N_10953,N_10331,N_10365);
xnor U10954 (N_10954,N_10321,N_10177);
and U10955 (N_10955,N_10135,N_10356);
xnor U10956 (N_10956,N_10428,N_10226);
nand U10957 (N_10957,N_10194,N_10134);
nand U10958 (N_10958,N_10411,N_10009);
nand U10959 (N_10959,N_10028,N_10173);
nor U10960 (N_10960,N_10188,N_10439);
or U10961 (N_10961,N_10148,N_10005);
nand U10962 (N_10962,N_10261,N_10118);
and U10963 (N_10963,N_10171,N_10187);
and U10964 (N_10964,N_10613,N_10577);
xor U10965 (N_10965,N_10589,N_10009);
xnor U10966 (N_10966,N_10541,N_10274);
xor U10967 (N_10967,N_10522,N_10181);
and U10968 (N_10968,N_10247,N_10005);
and U10969 (N_10969,N_10499,N_10386);
nand U10970 (N_10970,N_10569,N_10281);
xnor U10971 (N_10971,N_10170,N_10184);
xor U10972 (N_10972,N_10391,N_10091);
and U10973 (N_10973,N_10311,N_10532);
xor U10974 (N_10974,N_10471,N_10569);
and U10975 (N_10975,N_10617,N_10089);
or U10976 (N_10976,N_10061,N_10319);
nor U10977 (N_10977,N_10209,N_10149);
xor U10978 (N_10978,N_10224,N_10221);
nand U10979 (N_10979,N_10343,N_10009);
xor U10980 (N_10980,N_10442,N_10061);
xor U10981 (N_10981,N_10033,N_10253);
nor U10982 (N_10982,N_10562,N_10476);
and U10983 (N_10983,N_10260,N_10553);
nor U10984 (N_10984,N_10539,N_10607);
or U10985 (N_10985,N_10477,N_10169);
nand U10986 (N_10986,N_10575,N_10005);
and U10987 (N_10987,N_10161,N_10379);
nor U10988 (N_10988,N_10002,N_10075);
and U10989 (N_10989,N_10201,N_10001);
or U10990 (N_10990,N_10249,N_10301);
nand U10991 (N_10991,N_10326,N_10206);
xnor U10992 (N_10992,N_10493,N_10187);
nor U10993 (N_10993,N_10005,N_10400);
xor U10994 (N_10994,N_10405,N_10105);
xnor U10995 (N_10995,N_10427,N_10020);
and U10996 (N_10996,N_10466,N_10125);
and U10997 (N_10997,N_10255,N_10605);
nand U10998 (N_10998,N_10262,N_10124);
and U10999 (N_10999,N_10055,N_10553);
nand U11000 (N_11000,N_10207,N_10246);
and U11001 (N_11001,N_10168,N_10074);
nor U11002 (N_11002,N_10554,N_10607);
or U11003 (N_11003,N_10527,N_10423);
xor U11004 (N_11004,N_10002,N_10435);
or U11005 (N_11005,N_10600,N_10405);
and U11006 (N_11006,N_10523,N_10082);
nand U11007 (N_11007,N_10185,N_10602);
and U11008 (N_11008,N_10171,N_10177);
and U11009 (N_11009,N_10273,N_10023);
nand U11010 (N_11010,N_10414,N_10197);
nor U11011 (N_11011,N_10473,N_10534);
nand U11012 (N_11012,N_10084,N_10012);
nor U11013 (N_11013,N_10399,N_10523);
or U11014 (N_11014,N_10235,N_10041);
nor U11015 (N_11015,N_10287,N_10190);
nand U11016 (N_11016,N_10512,N_10543);
nor U11017 (N_11017,N_10265,N_10224);
xnor U11018 (N_11018,N_10442,N_10409);
xnor U11019 (N_11019,N_10548,N_10063);
or U11020 (N_11020,N_10410,N_10330);
or U11021 (N_11021,N_10526,N_10232);
or U11022 (N_11022,N_10038,N_10068);
and U11023 (N_11023,N_10581,N_10147);
xnor U11024 (N_11024,N_10088,N_10056);
or U11025 (N_11025,N_10275,N_10321);
or U11026 (N_11026,N_10157,N_10212);
xor U11027 (N_11027,N_10160,N_10318);
or U11028 (N_11028,N_10230,N_10203);
or U11029 (N_11029,N_10057,N_10305);
and U11030 (N_11030,N_10300,N_10284);
and U11031 (N_11031,N_10186,N_10479);
nor U11032 (N_11032,N_10601,N_10518);
nand U11033 (N_11033,N_10255,N_10004);
xnor U11034 (N_11034,N_10040,N_10395);
xnor U11035 (N_11035,N_10581,N_10260);
nand U11036 (N_11036,N_10200,N_10561);
nand U11037 (N_11037,N_10139,N_10100);
nand U11038 (N_11038,N_10458,N_10584);
xor U11039 (N_11039,N_10609,N_10400);
nand U11040 (N_11040,N_10301,N_10404);
xor U11041 (N_11041,N_10169,N_10262);
xor U11042 (N_11042,N_10251,N_10135);
nand U11043 (N_11043,N_10556,N_10538);
or U11044 (N_11044,N_10140,N_10129);
xnor U11045 (N_11045,N_10539,N_10416);
nand U11046 (N_11046,N_10591,N_10036);
or U11047 (N_11047,N_10433,N_10351);
xnor U11048 (N_11048,N_10314,N_10342);
and U11049 (N_11049,N_10067,N_10298);
or U11050 (N_11050,N_10482,N_10294);
nor U11051 (N_11051,N_10272,N_10069);
nor U11052 (N_11052,N_10437,N_10099);
xor U11053 (N_11053,N_10210,N_10313);
nand U11054 (N_11054,N_10501,N_10098);
xnor U11055 (N_11055,N_10557,N_10309);
nor U11056 (N_11056,N_10217,N_10022);
or U11057 (N_11057,N_10371,N_10403);
or U11058 (N_11058,N_10284,N_10196);
or U11059 (N_11059,N_10355,N_10034);
xor U11060 (N_11060,N_10157,N_10613);
xnor U11061 (N_11061,N_10498,N_10094);
and U11062 (N_11062,N_10614,N_10173);
xor U11063 (N_11063,N_10539,N_10166);
nor U11064 (N_11064,N_10344,N_10411);
xor U11065 (N_11065,N_10575,N_10227);
nor U11066 (N_11066,N_10198,N_10324);
nor U11067 (N_11067,N_10482,N_10237);
xnor U11068 (N_11068,N_10410,N_10438);
or U11069 (N_11069,N_10262,N_10333);
nor U11070 (N_11070,N_10010,N_10228);
or U11071 (N_11071,N_10260,N_10295);
nor U11072 (N_11072,N_10303,N_10510);
or U11073 (N_11073,N_10419,N_10294);
xnor U11074 (N_11074,N_10616,N_10128);
nor U11075 (N_11075,N_10148,N_10596);
or U11076 (N_11076,N_10590,N_10338);
and U11077 (N_11077,N_10040,N_10126);
nand U11078 (N_11078,N_10547,N_10427);
nor U11079 (N_11079,N_10502,N_10501);
xnor U11080 (N_11080,N_10204,N_10426);
and U11081 (N_11081,N_10183,N_10531);
and U11082 (N_11082,N_10289,N_10235);
xnor U11083 (N_11083,N_10145,N_10055);
nor U11084 (N_11084,N_10477,N_10371);
or U11085 (N_11085,N_10465,N_10477);
nor U11086 (N_11086,N_10439,N_10605);
and U11087 (N_11087,N_10023,N_10160);
nand U11088 (N_11088,N_10137,N_10140);
nor U11089 (N_11089,N_10086,N_10368);
xor U11090 (N_11090,N_10319,N_10350);
xnor U11091 (N_11091,N_10607,N_10566);
nand U11092 (N_11092,N_10061,N_10175);
nand U11093 (N_11093,N_10238,N_10183);
or U11094 (N_11094,N_10373,N_10550);
nor U11095 (N_11095,N_10085,N_10445);
xor U11096 (N_11096,N_10347,N_10120);
nand U11097 (N_11097,N_10134,N_10360);
xor U11098 (N_11098,N_10328,N_10449);
nand U11099 (N_11099,N_10052,N_10133);
or U11100 (N_11100,N_10419,N_10620);
and U11101 (N_11101,N_10012,N_10248);
nand U11102 (N_11102,N_10303,N_10469);
xor U11103 (N_11103,N_10624,N_10450);
xnor U11104 (N_11104,N_10252,N_10600);
nand U11105 (N_11105,N_10362,N_10514);
and U11106 (N_11106,N_10551,N_10155);
and U11107 (N_11107,N_10353,N_10260);
nand U11108 (N_11108,N_10482,N_10039);
nand U11109 (N_11109,N_10580,N_10183);
and U11110 (N_11110,N_10064,N_10613);
nor U11111 (N_11111,N_10415,N_10120);
nor U11112 (N_11112,N_10521,N_10581);
xnor U11113 (N_11113,N_10348,N_10074);
nor U11114 (N_11114,N_10238,N_10236);
or U11115 (N_11115,N_10304,N_10343);
nand U11116 (N_11116,N_10570,N_10133);
or U11117 (N_11117,N_10337,N_10474);
or U11118 (N_11118,N_10118,N_10566);
or U11119 (N_11119,N_10317,N_10146);
or U11120 (N_11120,N_10464,N_10216);
nand U11121 (N_11121,N_10172,N_10478);
and U11122 (N_11122,N_10506,N_10294);
nand U11123 (N_11123,N_10521,N_10623);
or U11124 (N_11124,N_10232,N_10176);
nor U11125 (N_11125,N_10261,N_10121);
xor U11126 (N_11126,N_10341,N_10470);
nor U11127 (N_11127,N_10083,N_10561);
and U11128 (N_11128,N_10420,N_10012);
nand U11129 (N_11129,N_10239,N_10012);
xnor U11130 (N_11130,N_10219,N_10207);
nor U11131 (N_11131,N_10409,N_10472);
nor U11132 (N_11132,N_10506,N_10553);
nor U11133 (N_11133,N_10620,N_10339);
nand U11134 (N_11134,N_10369,N_10195);
or U11135 (N_11135,N_10255,N_10092);
nor U11136 (N_11136,N_10183,N_10328);
nand U11137 (N_11137,N_10210,N_10572);
and U11138 (N_11138,N_10279,N_10210);
or U11139 (N_11139,N_10319,N_10432);
xnor U11140 (N_11140,N_10204,N_10180);
nor U11141 (N_11141,N_10569,N_10615);
nand U11142 (N_11142,N_10353,N_10176);
xnor U11143 (N_11143,N_10164,N_10161);
and U11144 (N_11144,N_10542,N_10456);
xor U11145 (N_11145,N_10047,N_10072);
nand U11146 (N_11146,N_10552,N_10321);
xnor U11147 (N_11147,N_10449,N_10249);
nor U11148 (N_11148,N_10012,N_10167);
nand U11149 (N_11149,N_10167,N_10615);
or U11150 (N_11150,N_10399,N_10174);
xnor U11151 (N_11151,N_10418,N_10369);
nor U11152 (N_11152,N_10204,N_10388);
or U11153 (N_11153,N_10506,N_10239);
xor U11154 (N_11154,N_10590,N_10103);
or U11155 (N_11155,N_10267,N_10013);
nor U11156 (N_11156,N_10335,N_10552);
and U11157 (N_11157,N_10216,N_10329);
nor U11158 (N_11158,N_10489,N_10464);
or U11159 (N_11159,N_10053,N_10317);
nand U11160 (N_11160,N_10136,N_10092);
nor U11161 (N_11161,N_10198,N_10474);
and U11162 (N_11162,N_10427,N_10385);
nor U11163 (N_11163,N_10492,N_10340);
xnor U11164 (N_11164,N_10443,N_10065);
xnor U11165 (N_11165,N_10364,N_10414);
and U11166 (N_11166,N_10350,N_10422);
and U11167 (N_11167,N_10267,N_10132);
nor U11168 (N_11168,N_10473,N_10288);
xor U11169 (N_11169,N_10484,N_10309);
xor U11170 (N_11170,N_10037,N_10421);
or U11171 (N_11171,N_10208,N_10178);
and U11172 (N_11172,N_10517,N_10142);
and U11173 (N_11173,N_10598,N_10266);
xnor U11174 (N_11174,N_10442,N_10331);
nand U11175 (N_11175,N_10486,N_10251);
xor U11176 (N_11176,N_10434,N_10312);
xor U11177 (N_11177,N_10187,N_10620);
or U11178 (N_11178,N_10076,N_10025);
xnor U11179 (N_11179,N_10268,N_10609);
or U11180 (N_11180,N_10063,N_10222);
nand U11181 (N_11181,N_10318,N_10520);
nor U11182 (N_11182,N_10573,N_10574);
or U11183 (N_11183,N_10187,N_10615);
nand U11184 (N_11184,N_10265,N_10092);
nand U11185 (N_11185,N_10008,N_10390);
and U11186 (N_11186,N_10558,N_10139);
or U11187 (N_11187,N_10163,N_10166);
and U11188 (N_11188,N_10239,N_10176);
and U11189 (N_11189,N_10398,N_10145);
nand U11190 (N_11190,N_10208,N_10277);
nor U11191 (N_11191,N_10228,N_10544);
nor U11192 (N_11192,N_10010,N_10257);
nor U11193 (N_11193,N_10428,N_10048);
and U11194 (N_11194,N_10220,N_10118);
xor U11195 (N_11195,N_10006,N_10065);
xnor U11196 (N_11196,N_10395,N_10350);
and U11197 (N_11197,N_10542,N_10274);
nand U11198 (N_11198,N_10585,N_10037);
or U11199 (N_11199,N_10034,N_10200);
nand U11200 (N_11200,N_10101,N_10515);
or U11201 (N_11201,N_10334,N_10547);
xor U11202 (N_11202,N_10481,N_10153);
or U11203 (N_11203,N_10426,N_10507);
or U11204 (N_11204,N_10193,N_10395);
or U11205 (N_11205,N_10133,N_10576);
or U11206 (N_11206,N_10139,N_10000);
and U11207 (N_11207,N_10302,N_10607);
and U11208 (N_11208,N_10152,N_10068);
xnor U11209 (N_11209,N_10131,N_10470);
and U11210 (N_11210,N_10363,N_10419);
or U11211 (N_11211,N_10313,N_10178);
or U11212 (N_11212,N_10463,N_10454);
and U11213 (N_11213,N_10073,N_10487);
or U11214 (N_11214,N_10177,N_10011);
and U11215 (N_11215,N_10190,N_10342);
nand U11216 (N_11216,N_10165,N_10535);
or U11217 (N_11217,N_10174,N_10048);
nor U11218 (N_11218,N_10335,N_10249);
nand U11219 (N_11219,N_10036,N_10493);
xor U11220 (N_11220,N_10044,N_10164);
nand U11221 (N_11221,N_10238,N_10477);
or U11222 (N_11222,N_10136,N_10572);
or U11223 (N_11223,N_10137,N_10193);
or U11224 (N_11224,N_10596,N_10223);
xor U11225 (N_11225,N_10569,N_10380);
nor U11226 (N_11226,N_10348,N_10099);
or U11227 (N_11227,N_10304,N_10540);
xor U11228 (N_11228,N_10049,N_10468);
or U11229 (N_11229,N_10351,N_10017);
xor U11230 (N_11230,N_10124,N_10602);
nor U11231 (N_11231,N_10246,N_10040);
and U11232 (N_11232,N_10116,N_10090);
or U11233 (N_11233,N_10255,N_10190);
or U11234 (N_11234,N_10167,N_10565);
nor U11235 (N_11235,N_10347,N_10234);
and U11236 (N_11236,N_10384,N_10563);
nor U11237 (N_11237,N_10088,N_10521);
and U11238 (N_11238,N_10040,N_10196);
nor U11239 (N_11239,N_10333,N_10359);
nand U11240 (N_11240,N_10055,N_10085);
nand U11241 (N_11241,N_10005,N_10169);
nand U11242 (N_11242,N_10298,N_10578);
or U11243 (N_11243,N_10003,N_10263);
xor U11244 (N_11244,N_10597,N_10229);
nand U11245 (N_11245,N_10394,N_10383);
and U11246 (N_11246,N_10087,N_10181);
or U11247 (N_11247,N_10396,N_10162);
and U11248 (N_11248,N_10297,N_10049);
xnor U11249 (N_11249,N_10159,N_10579);
or U11250 (N_11250,N_11237,N_10970);
nor U11251 (N_11251,N_10932,N_11200);
or U11252 (N_11252,N_11225,N_10662);
nor U11253 (N_11253,N_10660,N_10656);
xor U11254 (N_11254,N_10736,N_11047);
or U11255 (N_11255,N_11178,N_11034);
nor U11256 (N_11256,N_10680,N_11060);
or U11257 (N_11257,N_10746,N_11196);
and U11258 (N_11258,N_10698,N_10849);
nor U11259 (N_11259,N_10887,N_10985);
or U11260 (N_11260,N_10813,N_11040);
and U11261 (N_11261,N_10979,N_10818);
xnor U11262 (N_11262,N_10768,N_10635);
nand U11263 (N_11263,N_10878,N_10799);
or U11264 (N_11264,N_10930,N_10800);
nor U11265 (N_11265,N_10784,N_10923);
or U11266 (N_11266,N_10865,N_10657);
and U11267 (N_11267,N_11003,N_11062);
xnor U11268 (N_11268,N_11142,N_11104);
nand U11269 (N_11269,N_10793,N_10689);
nand U11270 (N_11270,N_11024,N_11232);
and U11271 (N_11271,N_10670,N_10926);
nor U11272 (N_11272,N_10872,N_11145);
and U11273 (N_11273,N_10762,N_11091);
nand U11274 (N_11274,N_10980,N_11005);
nor U11275 (N_11275,N_11241,N_11072);
nand U11276 (N_11276,N_11075,N_10888);
nor U11277 (N_11277,N_11103,N_10847);
and U11278 (N_11278,N_11243,N_10783);
or U11279 (N_11279,N_10911,N_10904);
or U11280 (N_11280,N_10673,N_10733);
nand U11281 (N_11281,N_11012,N_11121);
or U11282 (N_11282,N_10919,N_10642);
and U11283 (N_11283,N_10961,N_10627);
and U11284 (N_11284,N_10927,N_10871);
nand U11285 (N_11285,N_10896,N_10755);
nand U11286 (N_11286,N_11132,N_11038);
or U11287 (N_11287,N_11147,N_10890);
and U11288 (N_11288,N_10972,N_11112);
nand U11289 (N_11289,N_10902,N_10722);
nand U11290 (N_11290,N_10839,N_10907);
and U11291 (N_11291,N_10988,N_10664);
xnor U11292 (N_11292,N_11079,N_10837);
nor U11293 (N_11293,N_11146,N_10761);
or U11294 (N_11294,N_10922,N_11156);
xor U11295 (N_11295,N_10681,N_10801);
nor U11296 (N_11296,N_10967,N_11052);
or U11297 (N_11297,N_11213,N_10672);
nor U11298 (N_11298,N_10986,N_10987);
or U11299 (N_11299,N_11209,N_10853);
and U11300 (N_11300,N_11080,N_11114);
and U11301 (N_11301,N_10645,N_10936);
xor U11302 (N_11302,N_10869,N_11195);
xnor U11303 (N_11303,N_10994,N_11119);
nor U11304 (N_11304,N_11013,N_11063);
and U11305 (N_11305,N_10991,N_10727);
nand U11306 (N_11306,N_10631,N_10637);
xnor U11307 (N_11307,N_10639,N_11223);
and U11308 (N_11308,N_11204,N_11070);
xor U11309 (N_11309,N_10968,N_11214);
nor U11310 (N_11310,N_10906,N_10905);
nand U11311 (N_11311,N_11236,N_10992);
nor U11312 (N_11312,N_10862,N_10823);
xor U11313 (N_11313,N_10777,N_10993);
nand U11314 (N_11314,N_10965,N_10696);
xnor U11315 (N_11315,N_11211,N_10735);
nor U11316 (N_11316,N_10854,N_10759);
nor U11317 (N_11317,N_10725,N_10648);
or U11318 (N_11318,N_10921,N_10719);
xnor U11319 (N_11319,N_11217,N_10834);
or U11320 (N_11320,N_10866,N_10705);
and U11321 (N_11321,N_11144,N_10644);
xor U11322 (N_11322,N_10816,N_11078);
nor U11323 (N_11323,N_10663,N_11248);
xnor U11324 (N_11324,N_11022,N_10952);
or U11325 (N_11325,N_11152,N_11051);
xnor U11326 (N_11326,N_10821,N_10721);
and U11327 (N_11327,N_10828,N_10729);
xnor U11328 (N_11328,N_10815,N_10638);
and U11329 (N_11329,N_11056,N_10717);
xor U11330 (N_11330,N_10899,N_10751);
and U11331 (N_11331,N_11073,N_11122);
or U11332 (N_11332,N_11138,N_10875);
nor U11333 (N_11333,N_11007,N_10962);
nand U11334 (N_11334,N_11045,N_10773);
xor U11335 (N_11335,N_10646,N_11172);
or U11336 (N_11336,N_10937,N_10728);
xnor U11337 (N_11337,N_10702,N_10626);
nand U11338 (N_11338,N_11126,N_11127);
or U11339 (N_11339,N_10889,N_10687);
xor U11340 (N_11340,N_10797,N_10860);
or U11341 (N_11341,N_11203,N_11210);
nand U11342 (N_11342,N_10963,N_10830);
or U11343 (N_11343,N_10658,N_10882);
xor U11344 (N_11344,N_10842,N_11099);
or U11345 (N_11345,N_11109,N_10769);
nor U11346 (N_11346,N_11090,N_10858);
or U11347 (N_11347,N_10706,N_11238);
xnor U11348 (N_11348,N_10838,N_11016);
xor U11349 (N_11349,N_10951,N_11035);
xnor U11350 (N_11350,N_11100,N_10977);
and U11351 (N_11351,N_10855,N_11027);
and U11352 (N_11352,N_10812,N_10683);
nor U11353 (N_11353,N_11066,N_10678);
xor U11354 (N_11354,N_10647,N_10792);
and U11355 (N_11355,N_10750,N_10807);
nor U11356 (N_11356,N_11183,N_11086);
xor U11357 (N_11357,N_11131,N_10959);
xor U11358 (N_11358,N_10629,N_11023);
xnor U11359 (N_11359,N_11006,N_10774);
xor U11360 (N_11360,N_11031,N_10739);
xor U11361 (N_11361,N_10822,N_11092);
and U11362 (N_11362,N_11094,N_10841);
nor U11363 (N_11363,N_11067,N_10669);
or U11364 (N_11364,N_10894,N_10666);
or U11365 (N_11365,N_10796,N_11048);
xor U11366 (N_11366,N_10643,N_10641);
nand U11367 (N_11367,N_11186,N_11185);
nor U11368 (N_11368,N_10873,N_11245);
and U11369 (N_11369,N_10715,N_11088);
nor U11370 (N_11370,N_10982,N_10667);
or U11371 (N_11371,N_10892,N_11054);
and U11372 (N_11372,N_11097,N_10798);
nor U11373 (N_11373,N_11188,N_11149);
or U11374 (N_11374,N_10741,N_10795);
or U11375 (N_11375,N_11219,N_11148);
xnor U11376 (N_11376,N_10928,N_10956);
nor U11377 (N_11377,N_11076,N_10883);
or U11378 (N_11378,N_11116,N_10835);
or U11379 (N_11379,N_10820,N_11227);
and U11380 (N_11380,N_10943,N_10753);
and U11381 (N_11381,N_10805,N_10953);
or U11382 (N_11382,N_11115,N_10668);
xnor U11383 (N_11383,N_11244,N_11162);
or U11384 (N_11384,N_11030,N_11019);
nor U11385 (N_11385,N_11230,N_10730);
nor U11386 (N_11386,N_10942,N_11120);
nand U11387 (N_11387,N_11102,N_11032);
xnor U11388 (N_11388,N_11137,N_10900);
or U11389 (N_11389,N_10918,N_11201);
nand U11390 (N_11390,N_10895,N_10964);
nand U11391 (N_11391,N_10778,N_10747);
and U11392 (N_11392,N_10946,N_11096);
and U11393 (N_11393,N_10861,N_10945);
nor U11394 (N_11394,N_10659,N_11176);
nand U11395 (N_11395,N_10754,N_10694);
nor U11396 (N_11396,N_10917,N_11157);
and U11397 (N_11397,N_11057,N_11105);
nand U11398 (N_11398,N_11033,N_10787);
nor U11399 (N_11399,N_11123,N_10874);
nor U11400 (N_11400,N_10654,N_10857);
nor U11401 (N_11401,N_10675,N_10740);
nand U11402 (N_11402,N_10949,N_10877);
nor U11403 (N_11403,N_10884,N_10756);
nor U11404 (N_11404,N_11050,N_10910);
nand U11405 (N_11405,N_11240,N_10863);
or U11406 (N_11406,N_10832,N_11010);
nand U11407 (N_11407,N_11160,N_10650);
nor U11408 (N_11408,N_11163,N_10786);
nand U11409 (N_11409,N_10674,N_10825);
or U11410 (N_11410,N_11184,N_10710);
or U11411 (N_11411,N_10652,N_10737);
and U11412 (N_11412,N_11018,N_11068);
nor U11413 (N_11413,N_10726,N_11216);
xnor U11414 (N_11414,N_11134,N_10939);
nor U11415 (N_11415,N_10709,N_11058);
nand U11416 (N_11416,N_10802,N_11009);
or U11417 (N_11417,N_10731,N_11205);
or U11418 (N_11418,N_10628,N_11193);
nor U11419 (N_11419,N_11174,N_10843);
and U11420 (N_11420,N_11191,N_10886);
xor U11421 (N_11421,N_10976,N_11029);
and U11422 (N_11422,N_10819,N_10814);
nor U11423 (N_11423,N_10732,N_11233);
xnor U11424 (N_11424,N_11222,N_11011);
xor U11425 (N_11425,N_11190,N_10749);
and U11426 (N_11426,N_10685,N_10898);
xor U11427 (N_11427,N_11041,N_10772);
or U11428 (N_11428,N_11008,N_10782);
and U11429 (N_11429,N_11089,N_10879);
and U11430 (N_11430,N_10776,N_10996);
nor U11431 (N_11431,N_11061,N_11218);
nand U11432 (N_11432,N_10984,N_10636);
or U11433 (N_11433,N_11036,N_11049);
nand U11434 (N_11434,N_10914,N_10840);
nand U11435 (N_11435,N_10780,N_10633);
and U11436 (N_11436,N_10651,N_10995);
nand U11437 (N_11437,N_11177,N_11231);
nand U11438 (N_11438,N_10859,N_11081);
or U11439 (N_11439,N_10938,N_10954);
or U11440 (N_11440,N_10950,N_10817);
and U11441 (N_11441,N_10974,N_10891);
or U11442 (N_11442,N_10711,N_10738);
nand U11443 (N_11443,N_11180,N_10897);
nor U11444 (N_11444,N_10708,N_11095);
xnor U11445 (N_11445,N_10844,N_10810);
xor U11446 (N_11446,N_11140,N_10720);
and U11447 (N_11447,N_10682,N_11065);
nand U11448 (N_11448,N_11000,N_10809);
xnor U11449 (N_11449,N_10999,N_10966);
nor U11450 (N_11450,N_10723,N_10661);
xnor U11451 (N_11451,N_10909,N_11242);
and U11452 (N_11452,N_10925,N_11069);
or U11453 (N_11453,N_11197,N_10941);
and U11454 (N_11454,N_11130,N_11004);
and U11455 (N_11455,N_11110,N_11084);
nand U11456 (N_11456,N_11085,N_11226);
xor U11457 (N_11457,N_10791,N_10748);
xor U11458 (N_11458,N_11077,N_11207);
or U11459 (N_11459,N_11124,N_10912);
or U11460 (N_11460,N_11020,N_10692);
nor U11461 (N_11461,N_10690,N_11199);
and U11462 (N_11462,N_11133,N_11150);
and U11463 (N_11463,N_10948,N_10864);
xnor U11464 (N_11464,N_10718,N_10929);
and U11465 (N_11465,N_10688,N_10893);
xor U11466 (N_11466,N_10625,N_10653);
nand U11467 (N_11467,N_10908,N_10655);
nand U11468 (N_11468,N_10881,N_10649);
and U11469 (N_11469,N_11247,N_11039);
or U11470 (N_11470,N_11161,N_10960);
and U11471 (N_11471,N_10707,N_11015);
xor U11472 (N_11472,N_10920,N_11171);
nand U11473 (N_11473,N_11229,N_10744);
or U11474 (N_11474,N_11064,N_10699);
and U11475 (N_11475,N_11082,N_10679);
nand U11476 (N_11476,N_10700,N_11037);
or U11477 (N_11477,N_11141,N_11143);
nand U11478 (N_11478,N_10763,N_10713);
and U11479 (N_11479,N_11192,N_10885);
xor U11480 (N_11480,N_11206,N_10671);
nor U11481 (N_11481,N_10806,N_10634);
or U11482 (N_11482,N_11055,N_10931);
nand U11483 (N_11483,N_10788,N_11044);
or U11484 (N_11484,N_11098,N_10981);
xor U11485 (N_11485,N_10836,N_10846);
nor U11486 (N_11486,N_10940,N_11167);
or U11487 (N_11487,N_11175,N_10803);
nand U11488 (N_11488,N_11046,N_11128);
xor U11489 (N_11489,N_11169,N_11151);
nand U11490 (N_11490,N_11111,N_10901);
nand U11491 (N_11491,N_10990,N_10947);
and U11492 (N_11492,N_11166,N_10851);
nor U11493 (N_11493,N_10676,N_11083);
nand U11494 (N_11494,N_10848,N_11106);
and U11495 (N_11495,N_11117,N_11059);
or U11496 (N_11496,N_10831,N_11042);
and U11497 (N_11497,N_10880,N_11028);
xor U11498 (N_11498,N_11014,N_10826);
nor U11499 (N_11499,N_10934,N_11165);
nand U11500 (N_11500,N_10716,N_10785);
and U11501 (N_11501,N_11074,N_11187);
nor U11502 (N_11502,N_11139,N_11136);
nand U11503 (N_11503,N_11235,N_11212);
or U11504 (N_11504,N_10824,N_11021);
or U11505 (N_11505,N_10829,N_11221);
nor U11506 (N_11506,N_10789,N_11170);
or U11507 (N_11507,N_10876,N_10975);
xnor U11508 (N_11508,N_11164,N_10916);
nand U11509 (N_11509,N_10760,N_10758);
nor U11510 (N_11510,N_10852,N_10804);
nand U11511 (N_11511,N_10998,N_11208);
nand U11512 (N_11512,N_11001,N_10845);
xor U11513 (N_11513,N_10765,N_10969);
and U11514 (N_11514,N_11179,N_11125);
xor U11515 (N_11515,N_11093,N_10989);
or U11516 (N_11516,N_11025,N_11154);
nor U11517 (N_11517,N_10734,N_10933);
or U11518 (N_11518,N_10915,N_11168);
nor U11519 (N_11519,N_10640,N_11108);
nand U11520 (N_11520,N_10973,N_11198);
xnor U11521 (N_11521,N_11239,N_10766);
nor U11522 (N_11522,N_11173,N_10971);
and U11523 (N_11523,N_11129,N_10697);
xnor U11524 (N_11524,N_10752,N_10868);
and U11525 (N_11525,N_10850,N_10903);
xor U11526 (N_11526,N_10983,N_11053);
xor U11527 (N_11527,N_11194,N_10935);
and U11528 (N_11528,N_11159,N_10745);
nor U11529 (N_11529,N_10957,N_10827);
nand U11530 (N_11530,N_10704,N_10714);
or U11531 (N_11531,N_10997,N_11153);
nand U11532 (N_11532,N_10684,N_10924);
xnor U11533 (N_11533,N_10913,N_11026);
nand U11534 (N_11534,N_10779,N_10794);
xor U11535 (N_11535,N_10712,N_10958);
or U11536 (N_11536,N_10944,N_10743);
nand U11537 (N_11537,N_10703,N_10693);
xor U11538 (N_11538,N_10781,N_11155);
xor U11539 (N_11539,N_11118,N_11220);
nor U11540 (N_11540,N_11158,N_10856);
or U11541 (N_11541,N_11181,N_11215);
nor U11542 (N_11542,N_11224,N_10771);
xor U11543 (N_11543,N_10665,N_10691);
xnor U11544 (N_11544,N_10686,N_11087);
nand U11545 (N_11545,N_10790,N_11071);
xnor U11546 (N_11546,N_11234,N_11101);
nor U11547 (N_11547,N_10701,N_10632);
xnor U11548 (N_11548,N_10867,N_10742);
and U11549 (N_11549,N_11202,N_10764);
xor U11550 (N_11550,N_11228,N_11249);
nand U11551 (N_11551,N_10775,N_11017);
nand U11552 (N_11552,N_10808,N_11182);
nor U11553 (N_11553,N_10833,N_10724);
nor U11554 (N_11554,N_10770,N_10757);
xor U11555 (N_11555,N_10767,N_11043);
nand U11556 (N_11556,N_10695,N_10811);
nand U11557 (N_11557,N_10870,N_11246);
nor U11558 (N_11558,N_11113,N_11002);
or U11559 (N_11559,N_10630,N_11189);
nor U11560 (N_11560,N_10955,N_11135);
nor U11561 (N_11561,N_10677,N_11107);
xnor U11562 (N_11562,N_10978,N_11134);
nor U11563 (N_11563,N_10729,N_10676);
xnor U11564 (N_11564,N_11082,N_10896);
and U11565 (N_11565,N_10874,N_10861);
nor U11566 (N_11566,N_11216,N_10815);
nand U11567 (N_11567,N_10780,N_10734);
or U11568 (N_11568,N_11131,N_11249);
nor U11569 (N_11569,N_10758,N_10855);
and U11570 (N_11570,N_11156,N_10976);
nor U11571 (N_11571,N_11100,N_10642);
and U11572 (N_11572,N_11060,N_10848);
nand U11573 (N_11573,N_10869,N_10934);
nor U11574 (N_11574,N_11176,N_11039);
and U11575 (N_11575,N_10649,N_10841);
or U11576 (N_11576,N_10793,N_10937);
and U11577 (N_11577,N_10784,N_10637);
xor U11578 (N_11578,N_10695,N_10839);
nor U11579 (N_11579,N_11050,N_11193);
nand U11580 (N_11580,N_11091,N_11010);
nand U11581 (N_11581,N_10973,N_10809);
nand U11582 (N_11582,N_10629,N_11156);
nor U11583 (N_11583,N_10658,N_10849);
nand U11584 (N_11584,N_10901,N_10645);
xnor U11585 (N_11585,N_10937,N_10752);
and U11586 (N_11586,N_11225,N_10974);
nand U11587 (N_11587,N_10810,N_11162);
nand U11588 (N_11588,N_10841,N_10635);
or U11589 (N_11589,N_10973,N_10968);
nand U11590 (N_11590,N_10736,N_10670);
nand U11591 (N_11591,N_11187,N_10952);
and U11592 (N_11592,N_11216,N_11244);
and U11593 (N_11593,N_10990,N_10979);
xnor U11594 (N_11594,N_11034,N_10949);
or U11595 (N_11595,N_11176,N_10700);
nor U11596 (N_11596,N_11249,N_11152);
nand U11597 (N_11597,N_10630,N_11135);
nor U11598 (N_11598,N_10790,N_10791);
and U11599 (N_11599,N_10745,N_10869);
and U11600 (N_11600,N_11096,N_10866);
nor U11601 (N_11601,N_10737,N_10936);
or U11602 (N_11602,N_10713,N_10870);
and U11603 (N_11603,N_11053,N_11154);
xor U11604 (N_11604,N_11099,N_11110);
or U11605 (N_11605,N_10782,N_10925);
nor U11606 (N_11606,N_10830,N_11223);
and U11607 (N_11607,N_10839,N_10775);
xor U11608 (N_11608,N_10731,N_10935);
or U11609 (N_11609,N_11142,N_10644);
xnor U11610 (N_11610,N_10631,N_10817);
or U11611 (N_11611,N_11151,N_10760);
nor U11612 (N_11612,N_11226,N_10993);
or U11613 (N_11613,N_11106,N_10757);
or U11614 (N_11614,N_10797,N_10658);
or U11615 (N_11615,N_11182,N_10976);
nand U11616 (N_11616,N_11078,N_10928);
and U11617 (N_11617,N_10992,N_10810);
nand U11618 (N_11618,N_10679,N_10898);
nand U11619 (N_11619,N_10988,N_10982);
and U11620 (N_11620,N_10728,N_10961);
nand U11621 (N_11621,N_10868,N_11036);
and U11622 (N_11622,N_11056,N_10990);
nand U11623 (N_11623,N_11010,N_10716);
nand U11624 (N_11624,N_10721,N_10997);
nor U11625 (N_11625,N_11183,N_11231);
nor U11626 (N_11626,N_11221,N_10786);
nand U11627 (N_11627,N_11179,N_11048);
xor U11628 (N_11628,N_10898,N_11202);
nand U11629 (N_11629,N_11089,N_11104);
xor U11630 (N_11630,N_11211,N_11042);
nand U11631 (N_11631,N_11170,N_10950);
nand U11632 (N_11632,N_10807,N_11135);
xor U11633 (N_11633,N_10805,N_10718);
nor U11634 (N_11634,N_11119,N_10976);
nand U11635 (N_11635,N_10698,N_10903);
and U11636 (N_11636,N_10666,N_10917);
or U11637 (N_11637,N_11050,N_11072);
nand U11638 (N_11638,N_11234,N_10920);
nor U11639 (N_11639,N_11054,N_11032);
xnor U11640 (N_11640,N_10766,N_11206);
or U11641 (N_11641,N_11141,N_10815);
nand U11642 (N_11642,N_10948,N_10808);
xnor U11643 (N_11643,N_10784,N_10898);
and U11644 (N_11644,N_11214,N_11099);
or U11645 (N_11645,N_11201,N_10638);
nand U11646 (N_11646,N_10676,N_10967);
and U11647 (N_11647,N_10887,N_10797);
nand U11648 (N_11648,N_11194,N_10835);
xnor U11649 (N_11649,N_10819,N_10809);
xor U11650 (N_11650,N_10747,N_10944);
nand U11651 (N_11651,N_11094,N_10716);
xnor U11652 (N_11652,N_10771,N_10987);
and U11653 (N_11653,N_11210,N_10960);
and U11654 (N_11654,N_10897,N_10721);
nand U11655 (N_11655,N_11143,N_10755);
nand U11656 (N_11656,N_10956,N_11140);
and U11657 (N_11657,N_11106,N_11082);
nor U11658 (N_11658,N_11163,N_10647);
nand U11659 (N_11659,N_10912,N_10923);
or U11660 (N_11660,N_11027,N_11028);
or U11661 (N_11661,N_11036,N_10873);
and U11662 (N_11662,N_10779,N_10781);
or U11663 (N_11663,N_10723,N_10837);
or U11664 (N_11664,N_10830,N_10827);
xor U11665 (N_11665,N_10797,N_10790);
xnor U11666 (N_11666,N_11066,N_10764);
nand U11667 (N_11667,N_11144,N_10728);
and U11668 (N_11668,N_10737,N_10759);
or U11669 (N_11669,N_10871,N_10649);
or U11670 (N_11670,N_10871,N_10891);
or U11671 (N_11671,N_10698,N_10828);
nor U11672 (N_11672,N_10906,N_10776);
or U11673 (N_11673,N_11048,N_10744);
or U11674 (N_11674,N_11216,N_10705);
or U11675 (N_11675,N_11017,N_11141);
nand U11676 (N_11676,N_11024,N_10966);
nor U11677 (N_11677,N_10986,N_10868);
xnor U11678 (N_11678,N_10712,N_11162);
and U11679 (N_11679,N_10784,N_11082);
xnor U11680 (N_11680,N_10719,N_10875);
or U11681 (N_11681,N_10910,N_11216);
nand U11682 (N_11682,N_11233,N_10927);
or U11683 (N_11683,N_10786,N_10947);
nand U11684 (N_11684,N_10981,N_10784);
nor U11685 (N_11685,N_10725,N_10865);
nand U11686 (N_11686,N_11213,N_11166);
or U11687 (N_11687,N_11237,N_11078);
nor U11688 (N_11688,N_10803,N_11238);
and U11689 (N_11689,N_10886,N_10743);
xnor U11690 (N_11690,N_10665,N_10848);
nand U11691 (N_11691,N_11109,N_11039);
xnor U11692 (N_11692,N_10945,N_10974);
and U11693 (N_11693,N_10986,N_10940);
and U11694 (N_11694,N_10771,N_11171);
xor U11695 (N_11695,N_11165,N_10952);
nand U11696 (N_11696,N_10794,N_10639);
and U11697 (N_11697,N_10753,N_10991);
nand U11698 (N_11698,N_10995,N_10850);
xor U11699 (N_11699,N_11070,N_10760);
nor U11700 (N_11700,N_11178,N_10862);
or U11701 (N_11701,N_10762,N_11051);
nand U11702 (N_11702,N_10860,N_11190);
or U11703 (N_11703,N_11201,N_10866);
nor U11704 (N_11704,N_10700,N_10994);
or U11705 (N_11705,N_10827,N_11195);
or U11706 (N_11706,N_10926,N_10635);
or U11707 (N_11707,N_11102,N_10841);
nor U11708 (N_11708,N_11240,N_11102);
and U11709 (N_11709,N_10990,N_10931);
xnor U11710 (N_11710,N_11196,N_10647);
or U11711 (N_11711,N_10723,N_10708);
xor U11712 (N_11712,N_10770,N_11182);
nor U11713 (N_11713,N_10873,N_10909);
and U11714 (N_11714,N_11212,N_11083);
and U11715 (N_11715,N_10765,N_11037);
and U11716 (N_11716,N_10782,N_10911);
and U11717 (N_11717,N_11159,N_10746);
and U11718 (N_11718,N_11005,N_10811);
or U11719 (N_11719,N_10758,N_10780);
or U11720 (N_11720,N_11160,N_11200);
nand U11721 (N_11721,N_10984,N_10690);
nand U11722 (N_11722,N_11177,N_11067);
xor U11723 (N_11723,N_11004,N_11088);
and U11724 (N_11724,N_10996,N_10730);
nor U11725 (N_11725,N_10670,N_10795);
nor U11726 (N_11726,N_10899,N_11017);
nor U11727 (N_11727,N_11080,N_11082);
nand U11728 (N_11728,N_10683,N_11102);
nand U11729 (N_11729,N_10633,N_10736);
nor U11730 (N_11730,N_11017,N_10953);
nand U11731 (N_11731,N_11157,N_10791);
nand U11732 (N_11732,N_11181,N_10997);
nor U11733 (N_11733,N_10936,N_10872);
nand U11734 (N_11734,N_10690,N_10920);
and U11735 (N_11735,N_10866,N_11018);
or U11736 (N_11736,N_11194,N_10678);
xnor U11737 (N_11737,N_10776,N_11194);
or U11738 (N_11738,N_11025,N_11116);
or U11739 (N_11739,N_10864,N_11165);
or U11740 (N_11740,N_10940,N_10841);
nand U11741 (N_11741,N_11235,N_11105);
and U11742 (N_11742,N_10820,N_10779);
nand U11743 (N_11743,N_10733,N_11243);
nor U11744 (N_11744,N_11015,N_11089);
nand U11745 (N_11745,N_10703,N_11043);
nand U11746 (N_11746,N_11022,N_10678);
xnor U11747 (N_11747,N_10858,N_10820);
nor U11748 (N_11748,N_10919,N_10741);
xor U11749 (N_11749,N_11079,N_11015);
nor U11750 (N_11750,N_11146,N_10801);
nand U11751 (N_11751,N_11170,N_10697);
nand U11752 (N_11752,N_10910,N_10680);
nand U11753 (N_11753,N_11041,N_10764);
or U11754 (N_11754,N_11043,N_10932);
xnor U11755 (N_11755,N_10718,N_10722);
xor U11756 (N_11756,N_10739,N_10792);
or U11757 (N_11757,N_11106,N_11113);
or U11758 (N_11758,N_10719,N_11133);
nor U11759 (N_11759,N_10876,N_11023);
or U11760 (N_11760,N_10701,N_11246);
or U11761 (N_11761,N_10890,N_10639);
or U11762 (N_11762,N_11155,N_11212);
xnor U11763 (N_11763,N_11193,N_10977);
and U11764 (N_11764,N_10805,N_10822);
nor U11765 (N_11765,N_11080,N_11211);
and U11766 (N_11766,N_11167,N_10842);
and U11767 (N_11767,N_10972,N_10638);
nor U11768 (N_11768,N_10903,N_10834);
xor U11769 (N_11769,N_10808,N_10981);
nand U11770 (N_11770,N_11153,N_11139);
nor U11771 (N_11771,N_11134,N_10771);
nand U11772 (N_11772,N_11025,N_10787);
nor U11773 (N_11773,N_11055,N_11143);
xnor U11774 (N_11774,N_10648,N_11127);
or U11775 (N_11775,N_11022,N_11171);
and U11776 (N_11776,N_11018,N_10925);
xor U11777 (N_11777,N_11090,N_11186);
and U11778 (N_11778,N_11100,N_11206);
or U11779 (N_11779,N_11042,N_10892);
nand U11780 (N_11780,N_10891,N_11042);
and U11781 (N_11781,N_10645,N_11197);
xor U11782 (N_11782,N_10928,N_11134);
or U11783 (N_11783,N_10692,N_11076);
and U11784 (N_11784,N_10813,N_10868);
xnor U11785 (N_11785,N_10789,N_11020);
or U11786 (N_11786,N_10799,N_11053);
or U11787 (N_11787,N_11034,N_11226);
or U11788 (N_11788,N_10773,N_10888);
or U11789 (N_11789,N_10792,N_10913);
nand U11790 (N_11790,N_11174,N_10795);
nand U11791 (N_11791,N_11040,N_11003);
nand U11792 (N_11792,N_10955,N_10672);
or U11793 (N_11793,N_10997,N_10831);
and U11794 (N_11794,N_10751,N_10664);
or U11795 (N_11795,N_10691,N_10956);
and U11796 (N_11796,N_11030,N_10818);
nand U11797 (N_11797,N_10880,N_10716);
xnor U11798 (N_11798,N_10979,N_10951);
and U11799 (N_11799,N_10976,N_11057);
and U11800 (N_11800,N_11204,N_10782);
xnor U11801 (N_11801,N_11057,N_10809);
nand U11802 (N_11802,N_10786,N_11145);
nor U11803 (N_11803,N_10915,N_11027);
or U11804 (N_11804,N_11147,N_11162);
or U11805 (N_11805,N_11133,N_11171);
and U11806 (N_11806,N_10687,N_11059);
or U11807 (N_11807,N_10978,N_10625);
nand U11808 (N_11808,N_10646,N_11209);
xnor U11809 (N_11809,N_10848,N_10997);
xnor U11810 (N_11810,N_11015,N_10909);
xor U11811 (N_11811,N_10991,N_10700);
nand U11812 (N_11812,N_10845,N_11109);
or U11813 (N_11813,N_11227,N_10764);
and U11814 (N_11814,N_11197,N_11193);
or U11815 (N_11815,N_11247,N_10887);
xor U11816 (N_11816,N_10936,N_10712);
nor U11817 (N_11817,N_11081,N_10870);
and U11818 (N_11818,N_10669,N_11075);
nor U11819 (N_11819,N_11053,N_10914);
xnor U11820 (N_11820,N_10888,N_10690);
nor U11821 (N_11821,N_10812,N_11163);
nand U11822 (N_11822,N_11218,N_10890);
xnor U11823 (N_11823,N_10823,N_11135);
xnor U11824 (N_11824,N_10810,N_11003);
nand U11825 (N_11825,N_10927,N_10883);
xnor U11826 (N_11826,N_11008,N_10649);
xor U11827 (N_11827,N_11050,N_11042);
or U11828 (N_11828,N_10916,N_11096);
xor U11829 (N_11829,N_11030,N_10648);
or U11830 (N_11830,N_10630,N_11169);
nand U11831 (N_11831,N_11194,N_10833);
nand U11832 (N_11832,N_11149,N_10660);
and U11833 (N_11833,N_10870,N_11019);
nand U11834 (N_11834,N_10801,N_10831);
nand U11835 (N_11835,N_11049,N_10787);
xor U11836 (N_11836,N_11103,N_10915);
and U11837 (N_11837,N_11016,N_10778);
xnor U11838 (N_11838,N_11057,N_10749);
xor U11839 (N_11839,N_10904,N_11135);
nand U11840 (N_11840,N_10914,N_10779);
nor U11841 (N_11841,N_10810,N_11099);
or U11842 (N_11842,N_11188,N_10887);
and U11843 (N_11843,N_11197,N_10958);
nor U11844 (N_11844,N_11213,N_11101);
or U11845 (N_11845,N_10838,N_11141);
nor U11846 (N_11846,N_10649,N_10795);
xnor U11847 (N_11847,N_10851,N_10871);
nor U11848 (N_11848,N_10998,N_10987);
nand U11849 (N_11849,N_11161,N_10642);
or U11850 (N_11850,N_10872,N_10738);
or U11851 (N_11851,N_11004,N_11143);
nor U11852 (N_11852,N_10959,N_10648);
nand U11853 (N_11853,N_10932,N_11231);
xnor U11854 (N_11854,N_10923,N_10643);
nor U11855 (N_11855,N_10684,N_11151);
xor U11856 (N_11856,N_10718,N_10809);
xor U11857 (N_11857,N_10671,N_10937);
nor U11858 (N_11858,N_10664,N_10733);
and U11859 (N_11859,N_11217,N_10917);
nand U11860 (N_11860,N_10870,N_11075);
nor U11861 (N_11861,N_10899,N_10851);
or U11862 (N_11862,N_10812,N_10647);
nor U11863 (N_11863,N_11158,N_10962);
nor U11864 (N_11864,N_10957,N_11159);
and U11865 (N_11865,N_11238,N_11103);
or U11866 (N_11866,N_11233,N_10886);
nand U11867 (N_11867,N_10718,N_11206);
nor U11868 (N_11868,N_11037,N_10969);
nand U11869 (N_11869,N_10829,N_10934);
and U11870 (N_11870,N_10796,N_11009);
nor U11871 (N_11871,N_10941,N_10975);
xor U11872 (N_11872,N_10811,N_11056);
nor U11873 (N_11873,N_10714,N_11102);
nor U11874 (N_11874,N_11111,N_11203);
nand U11875 (N_11875,N_11817,N_11427);
or U11876 (N_11876,N_11772,N_11323);
nand U11877 (N_11877,N_11691,N_11429);
and U11878 (N_11878,N_11497,N_11456);
xnor U11879 (N_11879,N_11699,N_11484);
xor U11880 (N_11880,N_11807,N_11819);
and U11881 (N_11881,N_11339,N_11540);
or U11882 (N_11882,N_11758,N_11658);
nor U11883 (N_11883,N_11558,N_11336);
and U11884 (N_11884,N_11356,N_11349);
or U11885 (N_11885,N_11255,N_11655);
nor U11886 (N_11886,N_11347,N_11635);
xnor U11887 (N_11887,N_11622,N_11768);
nor U11888 (N_11888,N_11637,N_11867);
nand U11889 (N_11889,N_11866,N_11763);
xnor U11890 (N_11890,N_11673,N_11783);
nand U11891 (N_11891,N_11472,N_11495);
xor U11892 (N_11892,N_11443,N_11494);
or U11893 (N_11893,N_11551,N_11390);
or U11894 (N_11894,N_11613,N_11611);
and U11895 (N_11895,N_11771,N_11756);
nor U11896 (N_11896,N_11409,N_11646);
or U11897 (N_11897,N_11471,N_11759);
xor U11898 (N_11898,N_11440,N_11853);
and U11899 (N_11899,N_11786,N_11822);
nand U11900 (N_11900,N_11376,N_11684);
or U11901 (N_11901,N_11873,N_11703);
xor U11902 (N_11902,N_11568,N_11617);
or U11903 (N_11903,N_11451,N_11803);
or U11904 (N_11904,N_11659,N_11348);
or U11905 (N_11905,N_11424,N_11357);
nand U11906 (N_11906,N_11683,N_11340);
nor U11907 (N_11907,N_11672,N_11770);
nand U11908 (N_11908,N_11396,N_11530);
or U11909 (N_11909,N_11282,N_11315);
xnor U11910 (N_11910,N_11739,N_11687);
xnor U11911 (N_11911,N_11270,N_11671);
or U11912 (N_11912,N_11562,N_11620);
nand U11913 (N_11913,N_11810,N_11350);
xnor U11914 (N_11914,N_11793,N_11678);
or U11915 (N_11915,N_11736,N_11656);
and U11916 (N_11916,N_11734,N_11490);
and U11917 (N_11917,N_11438,N_11836);
and U11918 (N_11918,N_11820,N_11652);
or U11919 (N_11919,N_11859,N_11346);
nand U11920 (N_11920,N_11441,N_11846);
and U11921 (N_11921,N_11277,N_11697);
xor U11922 (N_11922,N_11838,N_11757);
xor U11923 (N_11923,N_11461,N_11405);
nor U11924 (N_11924,N_11774,N_11358);
nand U11925 (N_11925,N_11462,N_11640);
and U11926 (N_11926,N_11344,N_11552);
and U11927 (N_11927,N_11466,N_11401);
nor U11928 (N_11928,N_11851,N_11491);
and U11929 (N_11929,N_11636,N_11468);
xor U11930 (N_11930,N_11342,N_11860);
or U11931 (N_11931,N_11273,N_11510);
and U11932 (N_11932,N_11400,N_11581);
nor U11933 (N_11933,N_11605,N_11665);
nand U11934 (N_11934,N_11855,N_11333);
and U11935 (N_11935,N_11477,N_11526);
or U11936 (N_11936,N_11292,N_11385);
nor U11937 (N_11937,N_11492,N_11863);
and U11938 (N_11938,N_11577,N_11566);
nand U11939 (N_11939,N_11589,N_11585);
and U11940 (N_11940,N_11704,N_11445);
nand U11941 (N_11941,N_11775,N_11812);
or U11942 (N_11942,N_11378,N_11413);
nor U11943 (N_11943,N_11728,N_11579);
nand U11944 (N_11944,N_11741,N_11573);
or U11945 (N_11945,N_11353,N_11564);
or U11946 (N_11946,N_11834,N_11571);
and U11947 (N_11947,N_11723,N_11548);
and U11948 (N_11948,N_11436,N_11785);
xnor U11949 (N_11949,N_11604,N_11523);
xor U11950 (N_11950,N_11519,N_11354);
nand U11951 (N_11951,N_11864,N_11307);
nor U11952 (N_11952,N_11508,N_11708);
xnor U11953 (N_11953,N_11433,N_11667);
and U11954 (N_11954,N_11743,N_11865);
xnor U11955 (N_11955,N_11261,N_11686);
and U11956 (N_11956,N_11476,N_11749);
or U11957 (N_11957,N_11457,N_11489);
nor U11958 (N_11958,N_11818,N_11676);
xor U11959 (N_11959,N_11352,N_11750);
nor U11960 (N_11960,N_11787,N_11259);
xor U11961 (N_11961,N_11474,N_11572);
nand U11962 (N_11962,N_11709,N_11381);
or U11963 (N_11963,N_11502,N_11721);
xnor U11964 (N_11964,N_11693,N_11710);
nor U11965 (N_11965,N_11782,N_11610);
or U11966 (N_11966,N_11393,N_11389);
or U11967 (N_11967,N_11872,N_11811);
and U11968 (N_11968,N_11360,N_11318);
nand U11969 (N_11969,N_11284,N_11871);
and U11970 (N_11970,N_11647,N_11574);
xnor U11971 (N_11971,N_11501,N_11844);
or U11972 (N_11972,N_11722,N_11805);
and U11973 (N_11973,N_11290,N_11712);
nor U11974 (N_11974,N_11375,N_11618);
nand U11975 (N_11975,N_11773,N_11583);
or U11976 (N_11976,N_11415,N_11266);
nand U11977 (N_11977,N_11685,N_11293);
or U11978 (N_11978,N_11857,N_11275);
nor U11979 (N_11979,N_11764,N_11383);
nand U11980 (N_11980,N_11535,N_11412);
nand U11981 (N_11981,N_11660,N_11328);
xor U11982 (N_11982,N_11330,N_11578);
or U11983 (N_11983,N_11711,N_11299);
nor U11984 (N_11984,N_11285,N_11602);
or U11985 (N_11985,N_11372,N_11274);
and U11986 (N_11986,N_11780,N_11794);
or U11987 (N_11987,N_11406,N_11762);
or U11988 (N_11988,N_11725,N_11629);
or U11989 (N_11989,N_11254,N_11802);
nor U11990 (N_11990,N_11576,N_11317);
and U11991 (N_11991,N_11777,N_11545);
and U11992 (N_11992,N_11554,N_11781);
nand U11993 (N_11993,N_11487,N_11479);
xor U11994 (N_11994,N_11439,N_11262);
and U11995 (N_11995,N_11541,N_11707);
nor U11996 (N_11996,N_11475,N_11688);
and U11997 (N_11997,N_11861,N_11595);
nand U11998 (N_11998,N_11796,N_11531);
nor U11999 (N_11999,N_11386,N_11366);
or U12000 (N_12000,N_11669,N_11345);
and U12001 (N_12001,N_11628,N_11563);
xnor U12002 (N_12002,N_11464,N_11705);
xnor U12003 (N_12003,N_11550,N_11294);
nand U12004 (N_12004,N_11421,N_11446);
nand U12005 (N_12005,N_11341,N_11465);
nor U12006 (N_12006,N_11437,N_11649);
nand U12007 (N_12007,N_11623,N_11542);
and U12008 (N_12008,N_11694,N_11615);
xnor U12009 (N_12009,N_11403,N_11305);
nand U12010 (N_12010,N_11792,N_11858);
nor U12011 (N_12011,N_11674,N_11856);
xor U12012 (N_12012,N_11634,N_11624);
nor U12013 (N_12013,N_11766,N_11744);
and U12014 (N_12014,N_11263,N_11753);
or U12015 (N_12015,N_11594,N_11483);
nand U12016 (N_12016,N_11874,N_11411);
nor U12017 (N_12017,N_11513,N_11829);
or U12018 (N_12018,N_11279,N_11361);
nand U12019 (N_12019,N_11544,N_11575);
or U12020 (N_12020,N_11458,N_11848);
and U12021 (N_12021,N_11524,N_11603);
nor U12022 (N_12022,N_11256,N_11698);
xnor U12023 (N_12023,N_11364,N_11518);
nand U12024 (N_12024,N_11561,N_11500);
nand U12025 (N_12025,N_11833,N_11387);
or U12026 (N_12026,N_11504,N_11382);
nor U12027 (N_12027,N_11823,N_11809);
or U12028 (N_12028,N_11496,N_11632);
and U12029 (N_12029,N_11546,N_11444);
nand U12030 (N_12030,N_11742,N_11379);
or U12031 (N_12031,N_11486,N_11313);
nor U12032 (N_12032,N_11425,N_11837);
nand U12033 (N_12033,N_11337,N_11702);
nand U12034 (N_12034,N_11407,N_11303);
xor U12035 (N_12035,N_11334,N_11418);
nand U12036 (N_12036,N_11601,N_11512);
and U12037 (N_12037,N_11559,N_11816);
xnor U12038 (N_12038,N_11539,N_11616);
nor U12039 (N_12039,N_11469,N_11265);
or U12040 (N_12040,N_11402,N_11419);
or U12041 (N_12041,N_11748,N_11268);
and U12042 (N_12042,N_11591,N_11729);
nand U12043 (N_12043,N_11830,N_11827);
nor U12044 (N_12044,N_11410,N_11459);
and U12045 (N_12045,N_11482,N_11804);
and U12046 (N_12046,N_11434,N_11831);
nor U12047 (N_12047,N_11297,N_11302);
and U12048 (N_12048,N_11845,N_11841);
nand U12049 (N_12049,N_11362,N_11529);
and U12050 (N_12050,N_11304,N_11499);
nand U12051 (N_12051,N_11662,N_11450);
xnor U12052 (N_12052,N_11276,N_11760);
xor U12053 (N_12053,N_11593,N_11731);
nor U12054 (N_12054,N_11257,N_11849);
or U12055 (N_12055,N_11677,N_11543);
nor U12056 (N_12056,N_11633,N_11310);
or U12057 (N_12057,N_11556,N_11296);
xnor U12058 (N_12058,N_11808,N_11291);
xnor U12059 (N_12059,N_11253,N_11498);
and U12060 (N_12060,N_11625,N_11847);
xnor U12061 (N_12061,N_11680,N_11306);
nor U12062 (N_12062,N_11626,N_11517);
nand U12063 (N_12063,N_11870,N_11631);
nor U12064 (N_12064,N_11286,N_11735);
and U12065 (N_12065,N_11740,N_11448);
and U12066 (N_12066,N_11319,N_11692);
nor U12067 (N_12067,N_11600,N_11399);
xnor U12068 (N_12068,N_11596,N_11325);
and U12069 (N_12069,N_11797,N_11534);
nand U12070 (N_12070,N_11314,N_11798);
or U12071 (N_12071,N_11716,N_11832);
xor U12072 (N_12072,N_11283,N_11321);
nor U12073 (N_12073,N_11547,N_11668);
and U12074 (N_12074,N_11643,N_11806);
nand U12075 (N_12075,N_11582,N_11642);
nand U12076 (N_12076,N_11839,N_11675);
or U12077 (N_12077,N_11592,N_11638);
nor U12078 (N_12078,N_11663,N_11449);
nand U12079 (N_12079,N_11460,N_11384);
and U12080 (N_12080,N_11507,N_11869);
nor U12081 (N_12081,N_11453,N_11470);
and U12082 (N_12082,N_11567,N_11506);
nor U12083 (N_12083,N_11281,N_11821);
and U12084 (N_12084,N_11532,N_11367);
xnor U12085 (N_12085,N_11799,N_11473);
xnor U12086 (N_12086,N_11258,N_11769);
nor U12087 (N_12087,N_11509,N_11351);
or U12088 (N_12088,N_11516,N_11627);
and U12089 (N_12089,N_11478,N_11287);
xor U12090 (N_12090,N_11395,N_11398);
and U12091 (N_12091,N_11761,N_11250);
nor U12092 (N_12092,N_11428,N_11430);
xnor U12093 (N_12093,N_11363,N_11298);
nor U12094 (N_12094,N_11590,N_11755);
and U12095 (N_12095,N_11732,N_11850);
nand U12096 (N_12096,N_11511,N_11752);
or U12097 (N_12097,N_11852,N_11784);
xor U12098 (N_12098,N_11380,N_11788);
nor U12099 (N_12099,N_11653,N_11713);
nor U12100 (N_12100,N_11730,N_11840);
xor U12101 (N_12101,N_11278,N_11326);
xnor U12102 (N_12102,N_11790,N_11666);
or U12103 (N_12103,N_11414,N_11815);
xor U12104 (N_12104,N_11480,N_11733);
and U12105 (N_12105,N_11377,N_11488);
xnor U12106 (N_12106,N_11431,N_11522);
nand U12107 (N_12107,N_11289,N_11271);
xnor U12108 (N_12108,N_11335,N_11426);
or U12109 (N_12109,N_11701,N_11828);
xor U12110 (N_12110,N_11588,N_11689);
or U12111 (N_12111,N_11447,N_11813);
nor U12112 (N_12112,N_11404,N_11417);
xor U12113 (N_12113,N_11370,N_11654);
or U12114 (N_12114,N_11300,N_11826);
nand U12115 (N_12115,N_11862,N_11714);
and U12116 (N_12116,N_11650,N_11842);
nor U12117 (N_12117,N_11316,N_11570);
xnor U12118 (N_12118,N_11536,N_11681);
and U12119 (N_12119,N_11408,N_11778);
or U12120 (N_12120,N_11814,N_11641);
nor U12121 (N_12121,N_11538,N_11776);
or U12122 (N_12122,N_11715,N_11442);
or U12123 (N_12123,N_11267,N_11565);
xnor U12124 (N_12124,N_11555,N_11288);
xnor U12125 (N_12125,N_11269,N_11422);
xnor U12126 (N_12126,N_11868,N_11651);
and U12127 (N_12127,N_11416,N_11331);
nor U12128 (N_12128,N_11737,N_11843);
and U12129 (N_12129,N_11598,N_11607);
nand U12130 (N_12130,N_11301,N_11724);
nor U12131 (N_12131,N_11392,N_11824);
nor U12132 (N_12132,N_11560,N_11308);
nor U12133 (N_12133,N_11369,N_11423);
and U12134 (N_12134,N_11619,N_11854);
or U12135 (N_12135,N_11648,N_11309);
and U12136 (N_12136,N_11493,N_11549);
nand U12137 (N_12137,N_11679,N_11251);
or U12138 (N_12138,N_11612,N_11719);
or U12139 (N_12139,N_11690,N_11630);
and U12140 (N_12140,N_11779,N_11746);
xor U12141 (N_12141,N_11608,N_11454);
xor U12142 (N_12142,N_11553,N_11738);
xor U12143 (N_12143,N_11745,N_11609);
nor U12144 (N_12144,N_11700,N_11432);
xnor U12145 (N_12145,N_11343,N_11801);
nor U12146 (N_12146,N_11260,N_11751);
or U12147 (N_12147,N_11365,N_11295);
nand U12148 (N_12148,N_11528,N_11329);
xor U12149 (N_12149,N_11320,N_11569);
nor U12150 (N_12150,N_11706,N_11597);
nand U12151 (N_12151,N_11645,N_11557);
nor U12152 (N_12152,N_11332,N_11505);
nor U12153 (N_12153,N_11825,N_11515);
nand U12154 (N_12154,N_11599,N_11614);
nor U12155 (N_12155,N_11388,N_11606);
or U12156 (N_12156,N_11312,N_11391);
nor U12157 (N_12157,N_11727,N_11720);
or U12158 (N_12158,N_11311,N_11795);
xor U12159 (N_12159,N_11252,N_11503);
nand U12160 (N_12160,N_11359,N_11420);
xnor U12161 (N_12161,N_11695,N_11435);
or U12162 (N_12162,N_11767,N_11835);
nor U12163 (N_12163,N_11264,N_11520);
or U12164 (N_12164,N_11327,N_11657);
nor U12165 (N_12165,N_11485,N_11586);
nand U12166 (N_12166,N_11718,N_11324);
nor U12167 (N_12167,N_11726,N_11747);
xor U12168 (N_12168,N_11355,N_11467);
and U12169 (N_12169,N_11521,N_11717);
nand U12170 (N_12170,N_11639,N_11664);
and U12171 (N_12171,N_11765,N_11644);
or U12172 (N_12172,N_11525,N_11527);
and U12173 (N_12173,N_11791,N_11800);
or U12174 (N_12174,N_11481,N_11587);
nor U12175 (N_12175,N_11452,N_11537);
xnor U12176 (N_12176,N_11754,N_11533);
and U12177 (N_12177,N_11580,N_11373);
nand U12178 (N_12178,N_11455,N_11789);
nand U12179 (N_12179,N_11338,N_11661);
or U12180 (N_12180,N_11394,N_11514);
and U12181 (N_12181,N_11584,N_11670);
xnor U12182 (N_12182,N_11621,N_11696);
nor U12183 (N_12183,N_11397,N_11463);
and U12184 (N_12184,N_11322,N_11371);
nand U12185 (N_12185,N_11682,N_11280);
and U12186 (N_12186,N_11374,N_11272);
xor U12187 (N_12187,N_11368,N_11588);
nor U12188 (N_12188,N_11870,N_11421);
or U12189 (N_12189,N_11712,N_11801);
or U12190 (N_12190,N_11747,N_11614);
nor U12191 (N_12191,N_11350,N_11544);
and U12192 (N_12192,N_11420,N_11623);
or U12193 (N_12193,N_11317,N_11437);
nor U12194 (N_12194,N_11814,N_11705);
nand U12195 (N_12195,N_11587,N_11301);
or U12196 (N_12196,N_11317,N_11256);
xor U12197 (N_12197,N_11819,N_11725);
and U12198 (N_12198,N_11646,N_11496);
xor U12199 (N_12199,N_11652,N_11673);
nand U12200 (N_12200,N_11268,N_11397);
nor U12201 (N_12201,N_11285,N_11495);
xnor U12202 (N_12202,N_11730,N_11478);
nand U12203 (N_12203,N_11424,N_11684);
nand U12204 (N_12204,N_11709,N_11673);
or U12205 (N_12205,N_11854,N_11843);
xor U12206 (N_12206,N_11284,N_11394);
nand U12207 (N_12207,N_11746,N_11553);
xor U12208 (N_12208,N_11667,N_11284);
or U12209 (N_12209,N_11444,N_11423);
xor U12210 (N_12210,N_11865,N_11606);
nand U12211 (N_12211,N_11814,N_11868);
or U12212 (N_12212,N_11263,N_11422);
or U12213 (N_12213,N_11569,N_11757);
xnor U12214 (N_12214,N_11398,N_11708);
nand U12215 (N_12215,N_11664,N_11327);
nand U12216 (N_12216,N_11810,N_11490);
nand U12217 (N_12217,N_11422,N_11725);
and U12218 (N_12218,N_11617,N_11326);
or U12219 (N_12219,N_11381,N_11404);
or U12220 (N_12220,N_11331,N_11843);
nand U12221 (N_12221,N_11338,N_11480);
and U12222 (N_12222,N_11707,N_11417);
nor U12223 (N_12223,N_11366,N_11673);
or U12224 (N_12224,N_11803,N_11794);
and U12225 (N_12225,N_11563,N_11433);
or U12226 (N_12226,N_11526,N_11832);
nor U12227 (N_12227,N_11434,N_11709);
and U12228 (N_12228,N_11532,N_11783);
nand U12229 (N_12229,N_11381,N_11478);
and U12230 (N_12230,N_11711,N_11770);
nor U12231 (N_12231,N_11332,N_11785);
or U12232 (N_12232,N_11650,N_11588);
nor U12233 (N_12233,N_11457,N_11809);
nor U12234 (N_12234,N_11816,N_11429);
nor U12235 (N_12235,N_11546,N_11463);
and U12236 (N_12236,N_11637,N_11582);
nor U12237 (N_12237,N_11300,N_11287);
and U12238 (N_12238,N_11767,N_11691);
nor U12239 (N_12239,N_11747,N_11399);
and U12240 (N_12240,N_11568,N_11640);
nor U12241 (N_12241,N_11260,N_11324);
nand U12242 (N_12242,N_11413,N_11471);
xnor U12243 (N_12243,N_11433,N_11369);
and U12244 (N_12244,N_11318,N_11527);
nor U12245 (N_12245,N_11725,N_11827);
xor U12246 (N_12246,N_11824,N_11298);
and U12247 (N_12247,N_11734,N_11569);
nor U12248 (N_12248,N_11402,N_11523);
nor U12249 (N_12249,N_11448,N_11610);
nand U12250 (N_12250,N_11558,N_11724);
xor U12251 (N_12251,N_11677,N_11712);
xnor U12252 (N_12252,N_11857,N_11657);
xor U12253 (N_12253,N_11334,N_11652);
and U12254 (N_12254,N_11632,N_11413);
nand U12255 (N_12255,N_11275,N_11782);
xor U12256 (N_12256,N_11755,N_11738);
nand U12257 (N_12257,N_11556,N_11761);
and U12258 (N_12258,N_11787,N_11554);
nor U12259 (N_12259,N_11649,N_11594);
nor U12260 (N_12260,N_11798,N_11386);
and U12261 (N_12261,N_11640,N_11629);
nor U12262 (N_12262,N_11832,N_11742);
nand U12263 (N_12263,N_11517,N_11814);
and U12264 (N_12264,N_11835,N_11322);
nand U12265 (N_12265,N_11852,N_11773);
or U12266 (N_12266,N_11481,N_11357);
or U12267 (N_12267,N_11357,N_11263);
and U12268 (N_12268,N_11541,N_11711);
nor U12269 (N_12269,N_11397,N_11295);
or U12270 (N_12270,N_11379,N_11773);
or U12271 (N_12271,N_11335,N_11266);
nor U12272 (N_12272,N_11658,N_11744);
nand U12273 (N_12273,N_11663,N_11262);
or U12274 (N_12274,N_11611,N_11767);
or U12275 (N_12275,N_11334,N_11686);
and U12276 (N_12276,N_11283,N_11733);
nand U12277 (N_12277,N_11493,N_11629);
xnor U12278 (N_12278,N_11822,N_11403);
nand U12279 (N_12279,N_11673,N_11432);
or U12280 (N_12280,N_11724,N_11503);
and U12281 (N_12281,N_11743,N_11695);
or U12282 (N_12282,N_11604,N_11732);
xnor U12283 (N_12283,N_11800,N_11298);
xnor U12284 (N_12284,N_11462,N_11632);
or U12285 (N_12285,N_11509,N_11404);
nor U12286 (N_12286,N_11675,N_11607);
nor U12287 (N_12287,N_11803,N_11582);
nand U12288 (N_12288,N_11611,N_11352);
nor U12289 (N_12289,N_11556,N_11860);
nor U12290 (N_12290,N_11492,N_11342);
nand U12291 (N_12291,N_11751,N_11691);
nor U12292 (N_12292,N_11871,N_11597);
nand U12293 (N_12293,N_11721,N_11366);
or U12294 (N_12294,N_11400,N_11792);
nor U12295 (N_12295,N_11861,N_11524);
and U12296 (N_12296,N_11513,N_11576);
xnor U12297 (N_12297,N_11494,N_11290);
nand U12298 (N_12298,N_11418,N_11347);
and U12299 (N_12299,N_11379,N_11524);
and U12300 (N_12300,N_11874,N_11408);
or U12301 (N_12301,N_11332,N_11689);
nand U12302 (N_12302,N_11517,N_11360);
xnor U12303 (N_12303,N_11842,N_11825);
nor U12304 (N_12304,N_11568,N_11506);
nor U12305 (N_12305,N_11841,N_11664);
and U12306 (N_12306,N_11388,N_11519);
nand U12307 (N_12307,N_11586,N_11531);
nand U12308 (N_12308,N_11470,N_11742);
nor U12309 (N_12309,N_11364,N_11817);
nand U12310 (N_12310,N_11515,N_11460);
nor U12311 (N_12311,N_11448,N_11253);
or U12312 (N_12312,N_11414,N_11676);
nand U12313 (N_12313,N_11338,N_11576);
and U12314 (N_12314,N_11847,N_11352);
and U12315 (N_12315,N_11318,N_11839);
xor U12316 (N_12316,N_11537,N_11611);
nor U12317 (N_12317,N_11778,N_11728);
and U12318 (N_12318,N_11609,N_11552);
and U12319 (N_12319,N_11561,N_11729);
xor U12320 (N_12320,N_11258,N_11650);
and U12321 (N_12321,N_11414,N_11538);
and U12322 (N_12322,N_11308,N_11556);
nor U12323 (N_12323,N_11255,N_11695);
nand U12324 (N_12324,N_11347,N_11330);
and U12325 (N_12325,N_11521,N_11655);
and U12326 (N_12326,N_11757,N_11873);
and U12327 (N_12327,N_11359,N_11303);
and U12328 (N_12328,N_11442,N_11750);
nor U12329 (N_12329,N_11457,N_11334);
xor U12330 (N_12330,N_11741,N_11321);
nand U12331 (N_12331,N_11262,N_11831);
and U12332 (N_12332,N_11874,N_11748);
or U12333 (N_12333,N_11545,N_11410);
and U12334 (N_12334,N_11304,N_11368);
or U12335 (N_12335,N_11686,N_11840);
or U12336 (N_12336,N_11718,N_11386);
xnor U12337 (N_12337,N_11448,N_11715);
nor U12338 (N_12338,N_11429,N_11253);
or U12339 (N_12339,N_11747,N_11548);
and U12340 (N_12340,N_11639,N_11460);
or U12341 (N_12341,N_11676,N_11614);
and U12342 (N_12342,N_11362,N_11850);
nor U12343 (N_12343,N_11585,N_11617);
or U12344 (N_12344,N_11741,N_11700);
xor U12345 (N_12345,N_11274,N_11365);
nand U12346 (N_12346,N_11695,N_11331);
or U12347 (N_12347,N_11269,N_11520);
xnor U12348 (N_12348,N_11384,N_11730);
nor U12349 (N_12349,N_11709,N_11602);
or U12350 (N_12350,N_11744,N_11256);
nand U12351 (N_12351,N_11718,N_11860);
nor U12352 (N_12352,N_11819,N_11597);
or U12353 (N_12353,N_11608,N_11714);
nand U12354 (N_12354,N_11845,N_11717);
or U12355 (N_12355,N_11847,N_11517);
nand U12356 (N_12356,N_11678,N_11477);
or U12357 (N_12357,N_11385,N_11427);
xor U12358 (N_12358,N_11852,N_11494);
or U12359 (N_12359,N_11798,N_11769);
or U12360 (N_12360,N_11357,N_11717);
or U12361 (N_12361,N_11844,N_11705);
nand U12362 (N_12362,N_11673,N_11583);
and U12363 (N_12363,N_11366,N_11492);
nand U12364 (N_12364,N_11811,N_11406);
or U12365 (N_12365,N_11838,N_11543);
and U12366 (N_12366,N_11525,N_11575);
xnor U12367 (N_12367,N_11811,N_11487);
or U12368 (N_12368,N_11495,N_11580);
or U12369 (N_12369,N_11408,N_11707);
nor U12370 (N_12370,N_11745,N_11382);
or U12371 (N_12371,N_11847,N_11519);
xnor U12372 (N_12372,N_11395,N_11598);
nor U12373 (N_12373,N_11675,N_11832);
or U12374 (N_12374,N_11748,N_11326);
xnor U12375 (N_12375,N_11555,N_11473);
nand U12376 (N_12376,N_11721,N_11479);
xor U12377 (N_12377,N_11848,N_11645);
or U12378 (N_12378,N_11453,N_11389);
xor U12379 (N_12379,N_11531,N_11264);
nand U12380 (N_12380,N_11841,N_11268);
nand U12381 (N_12381,N_11625,N_11453);
and U12382 (N_12382,N_11868,N_11808);
and U12383 (N_12383,N_11708,N_11689);
or U12384 (N_12384,N_11545,N_11414);
and U12385 (N_12385,N_11289,N_11404);
nor U12386 (N_12386,N_11631,N_11607);
nor U12387 (N_12387,N_11308,N_11797);
xor U12388 (N_12388,N_11613,N_11621);
nor U12389 (N_12389,N_11709,N_11809);
nand U12390 (N_12390,N_11544,N_11412);
nand U12391 (N_12391,N_11502,N_11717);
xnor U12392 (N_12392,N_11499,N_11671);
nand U12393 (N_12393,N_11505,N_11522);
nor U12394 (N_12394,N_11805,N_11695);
xnor U12395 (N_12395,N_11588,N_11299);
and U12396 (N_12396,N_11602,N_11418);
nand U12397 (N_12397,N_11447,N_11848);
or U12398 (N_12398,N_11500,N_11839);
nand U12399 (N_12399,N_11802,N_11599);
or U12400 (N_12400,N_11326,N_11284);
nor U12401 (N_12401,N_11471,N_11552);
nor U12402 (N_12402,N_11686,N_11700);
nor U12403 (N_12403,N_11699,N_11383);
and U12404 (N_12404,N_11775,N_11296);
xor U12405 (N_12405,N_11775,N_11791);
nand U12406 (N_12406,N_11866,N_11301);
xnor U12407 (N_12407,N_11662,N_11424);
nor U12408 (N_12408,N_11417,N_11693);
xor U12409 (N_12409,N_11839,N_11374);
xor U12410 (N_12410,N_11691,N_11709);
xnor U12411 (N_12411,N_11433,N_11740);
xnor U12412 (N_12412,N_11393,N_11859);
nand U12413 (N_12413,N_11485,N_11593);
xor U12414 (N_12414,N_11378,N_11503);
and U12415 (N_12415,N_11802,N_11682);
nor U12416 (N_12416,N_11435,N_11696);
xor U12417 (N_12417,N_11336,N_11835);
and U12418 (N_12418,N_11623,N_11630);
xor U12419 (N_12419,N_11441,N_11311);
or U12420 (N_12420,N_11470,N_11258);
nor U12421 (N_12421,N_11272,N_11522);
nand U12422 (N_12422,N_11565,N_11413);
nand U12423 (N_12423,N_11489,N_11829);
nand U12424 (N_12424,N_11582,N_11306);
nor U12425 (N_12425,N_11303,N_11512);
or U12426 (N_12426,N_11768,N_11776);
nor U12427 (N_12427,N_11750,N_11849);
and U12428 (N_12428,N_11253,N_11421);
nand U12429 (N_12429,N_11273,N_11514);
nor U12430 (N_12430,N_11289,N_11629);
and U12431 (N_12431,N_11856,N_11738);
xnor U12432 (N_12432,N_11848,N_11342);
or U12433 (N_12433,N_11848,N_11751);
and U12434 (N_12434,N_11856,N_11847);
nor U12435 (N_12435,N_11337,N_11395);
and U12436 (N_12436,N_11699,N_11453);
or U12437 (N_12437,N_11318,N_11253);
xnor U12438 (N_12438,N_11271,N_11864);
nor U12439 (N_12439,N_11464,N_11323);
nor U12440 (N_12440,N_11643,N_11803);
or U12441 (N_12441,N_11291,N_11801);
nand U12442 (N_12442,N_11308,N_11369);
xnor U12443 (N_12443,N_11558,N_11874);
and U12444 (N_12444,N_11653,N_11561);
and U12445 (N_12445,N_11835,N_11811);
xnor U12446 (N_12446,N_11728,N_11646);
nand U12447 (N_12447,N_11331,N_11357);
nand U12448 (N_12448,N_11365,N_11342);
and U12449 (N_12449,N_11724,N_11389);
and U12450 (N_12450,N_11527,N_11302);
xnor U12451 (N_12451,N_11843,N_11730);
xor U12452 (N_12452,N_11393,N_11429);
or U12453 (N_12453,N_11365,N_11390);
nand U12454 (N_12454,N_11469,N_11718);
nor U12455 (N_12455,N_11515,N_11569);
or U12456 (N_12456,N_11470,N_11590);
and U12457 (N_12457,N_11278,N_11451);
or U12458 (N_12458,N_11846,N_11640);
or U12459 (N_12459,N_11491,N_11813);
nor U12460 (N_12460,N_11832,N_11788);
nand U12461 (N_12461,N_11479,N_11419);
or U12462 (N_12462,N_11381,N_11669);
nand U12463 (N_12463,N_11405,N_11507);
or U12464 (N_12464,N_11834,N_11551);
or U12465 (N_12465,N_11462,N_11368);
and U12466 (N_12466,N_11682,N_11413);
nand U12467 (N_12467,N_11291,N_11732);
nand U12468 (N_12468,N_11399,N_11675);
nor U12469 (N_12469,N_11667,N_11514);
xor U12470 (N_12470,N_11872,N_11673);
nand U12471 (N_12471,N_11323,N_11475);
xnor U12472 (N_12472,N_11604,N_11677);
and U12473 (N_12473,N_11394,N_11663);
nor U12474 (N_12474,N_11558,N_11395);
or U12475 (N_12475,N_11386,N_11321);
nor U12476 (N_12476,N_11529,N_11479);
or U12477 (N_12477,N_11355,N_11775);
or U12478 (N_12478,N_11815,N_11833);
nand U12479 (N_12479,N_11436,N_11565);
nand U12480 (N_12480,N_11391,N_11500);
and U12481 (N_12481,N_11352,N_11335);
nor U12482 (N_12482,N_11349,N_11673);
or U12483 (N_12483,N_11805,N_11675);
and U12484 (N_12484,N_11659,N_11629);
or U12485 (N_12485,N_11652,N_11776);
nor U12486 (N_12486,N_11818,N_11850);
nor U12487 (N_12487,N_11574,N_11275);
and U12488 (N_12488,N_11708,N_11612);
nand U12489 (N_12489,N_11708,N_11562);
xor U12490 (N_12490,N_11302,N_11781);
and U12491 (N_12491,N_11393,N_11802);
xor U12492 (N_12492,N_11460,N_11733);
nor U12493 (N_12493,N_11669,N_11257);
and U12494 (N_12494,N_11389,N_11792);
and U12495 (N_12495,N_11828,N_11625);
or U12496 (N_12496,N_11539,N_11818);
nor U12497 (N_12497,N_11332,N_11790);
and U12498 (N_12498,N_11757,N_11575);
nand U12499 (N_12499,N_11768,N_11501);
and U12500 (N_12500,N_11948,N_12170);
or U12501 (N_12501,N_12154,N_12251);
or U12502 (N_12502,N_12125,N_11938);
xnor U12503 (N_12503,N_11943,N_12305);
nor U12504 (N_12504,N_12107,N_12211);
nor U12505 (N_12505,N_12065,N_12172);
nand U12506 (N_12506,N_11889,N_11959);
nand U12507 (N_12507,N_12481,N_12057);
and U12508 (N_12508,N_11932,N_12127);
nor U12509 (N_12509,N_12344,N_12167);
and U12510 (N_12510,N_11883,N_12488);
and U12511 (N_12511,N_12383,N_12165);
xor U12512 (N_12512,N_12108,N_11970);
and U12513 (N_12513,N_12077,N_11980);
nand U12514 (N_12514,N_11913,N_12494);
and U12515 (N_12515,N_12327,N_12298);
or U12516 (N_12516,N_11891,N_12166);
nor U12517 (N_12517,N_12053,N_12087);
xnor U12518 (N_12518,N_11965,N_12338);
or U12519 (N_12519,N_11890,N_12006);
xor U12520 (N_12520,N_11964,N_12121);
nand U12521 (N_12521,N_12234,N_12236);
nor U12522 (N_12522,N_12004,N_12394);
xor U12523 (N_12523,N_12267,N_12348);
xnor U12524 (N_12524,N_11976,N_12059);
xnor U12525 (N_12525,N_12384,N_12212);
or U12526 (N_12526,N_12005,N_12188);
nor U12527 (N_12527,N_12213,N_12418);
nor U12528 (N_12528,N_11956,N_11928);
xnor U12529 (N_12529,N_12099,N_11933);
and U12530 (N_12530,N_12264,N_12209);
nor U12531 (N_12531,N_12388,N_12037);
nor U12532 (N_12532,N_12490,N_12200);
or U12533 (N_12533,N_12438,N_12149);
and U12534 (N_12534,N_12069,N_12473);
nand U12535 (N_12535,N_11963,N_11885);
nand U12536 (N_12536,N_12233,N_12133);
nor U12537 (N_12537,N_12277,N_12462);
xor U12538 (N_12538,N_12095,N_12412);
nor U12539 (N_12539,N_12335,N_12416);
and U12540 (N_12540,N_12495,N_12193);
xor U12541 (N_12541,N_12238,N_12269);
nor U12542 (N_12542,N_12480,N_11896);
nor U12543 (N_12543,N_12284,N_12300);
and U12544 (N_12544,N_12157,N_12011);
and U12545 (N_12545,N_11934,N_12080);
nor U12546 (N_12546,N_12458,N_11916);
xor U12547 (N_12547,N_12406,N_12390);
nor U12548 (N_12548,N_12337,N_12359);
and U12549 (N_12549,N_12422,N_11990);
nand U12550 (N_12550,N_11882,N_12449);
or U12551 (N_12551,N_11892,N_12202);
nor U12552 (N_12552,N_12393,N_12180);
nor U12553 (N_12553,N_12022,N_11901);
or U12554 (N_12554,N_11881,N_12361);
or U12555 (N_12555,N_12281,N_12242);
nor U12556 (N_12556,N_12181,N_12185);
xnor U12557 (N_12557,N_12253,N_12472);
nand U12558 (N_12558,N_12447,N_12258);
and U12559 (N_12559,N_12444,N_12278);
or U12560 (N_12560,N_12227,N_11972);
xnor U12561 (N_12561,N_12243,N_12102);
nor U12562 (N_12562,N_12340,N_12270);
nand U12563 (N_12563,N_11936,N_12461);
nor U12564 (N_12564,N_12023,N_12455);
xnor U12565 (N_12565,N_12312,N_12222);
nand U12566 (N_12566,N_12179,N_12194);
or U12567 (N_12567,N_12308,N_11981);
or U12568 (N_12568,N_12366,N_12064);
and U12569 (N_12569,N_12235,N_11971);
nor U12570 (N_12570,N_12483,N_12082);
nand U12571 (N_12571,N_12097,N_12345);
and U12572 (N_12572,N_12214,N_12413);
or U12573 (N_12573,N_12441,N_12228);
nor U12574 (N_12574,N_12294,N_12025);
nor U12575 (N_12575,N_11947,N_12096);
or U12576 (N_12576,N_12199,N_12035);
xnor U12577 (N_12577,N_12311,N_12192);
nand U12578 (N_12578,N_12079,N_12475);
and U12579 (N_12579,N_11921,N_12171);
and U12580 (N_12580,N_11878,N_12105);
or U12581 (N_12581,N_12248,N_12293);
nor U12582 (N_12582,N_12104,N_12431);
and U12583 (N_12583,N_11908,N_12452);
and U12584 (N_12584,N_12319,N_12245);
xnor U12585 (N_12585,N_12147,N_12026);
and U12586 (N_12586,N_12349,N_12400);
nor U12587 (N_12587,N_12119,N_12411);
nor U12588 (N_12588,N_12460,N_12223);
or U12589 (N_12589,N_12442,N_12259);
or U12590 (N_12590,N_12457,N_12008);
nand U12591 (N_12591,N_12292,N_12356);
nor U12592 (N_12592,N_11995,N_12168);
xnor U12593 (N_12593,N_11950,N_12144);
or U12594 (N_12594,N_12191,N_11988);
or U12595 (N_12595,N_12479,N_12268);
nand U12596 (N_12596,N_12027,N_12407);
and U12597 (N_12597,N_11898,N_12249);
nor U12598 (N_12598,N_12395,N_11912);
and U12599 (N_12599,N_12226,N_12201);
and U12600 (N_12600,N_12210,N_12252);
or U12601 (N_12601,N_12204,N_12419);
or U12602 (N_12602,N_12331,N_12369);
xnor U12603 (N_12603,N_12357,N_12063);
nand U12604 (N_12604,N_12208,N_11909);
and U12605 (N_12605,N_12015,N_11904);
nor U12606 (N_12606,N_12332,N_11922);
and U12607 (N_12607,N_12471,N_12030);
nand U12608 (N_12608,N_12049,N_12244);
xnor U12609 (N_12609,N_12113,N_12048);
and U12610 (N_12610,N_12336,N_12169);
xnor U12611 (N_12611,N_11924,N_11925);
nor U12612 (N_12612,N_12138,N_12066);
or U12613 (N_12613,N_12318,N_12274);
nand U12614 (N_12614,N_12368,N_12387);
nand U12615 (N_12615,N_12177,N_12134);
nand U12616 (N_12616,N_12362,N_12158);
and U12617 (N_12617,N_12085,N_12060);
or U12618 (N_12618,N_12040,N_12489);
and U12619 (N_12619,N_12010,N_12364);
nor U12620 (N_12620,N_11888,N_11911);
or U12621 (N_12621,N_12056,N_12143);
and U12622 (N_12622,N_12146,N_12456);
or U12623 (N_12623,N_12405,N_12067);
nand U12624 (N_12624,N_12100,N_12290);
nor U12625 (N_12625,N_12353,N_12478);
xor U12626 (N_12626,N_12189,N_12091);
or U12627 (N_12627,N_12289,N_11975);
nor U12628 (N_12628,N_12280,N_12246);
or U12629 (N_12629,N_11879,N_12306);
nand U12630 (N_12630,N_12225,N_12002);
and U12631 (N_12631,N_12469,N_11905);
xnor U12632 (N_12632,N_12196,N_12164);
and U12633 (N_12633,N_12162,N_12072);
and U12634 (N_12634,N_12482,N_12279);
or U12635 (N_12635,N_12429,N_11914);
nor U12636 (N_12636,N_12250,N_12358);
xnor U12637 (N_12637,N_12145,N_12001);
xnor U12638 (N_12638,N_12135,N_12093);
and U12639 (N_12639,N_12173,N_11931);
and U12640 (N_12640,N_11877,N_12302);
xnor U12641 (N_12641,N_12052,N_12451);
or U12642 (N_12642,N_12117,N_12351);
nand U12643 (N_12643,N_12382,N_12313);
xnor U12644 (N_12644,N_12486,N_12379);
xor U12645 (N_12645,N_12326,N_12101);
or U12646 (N_12646,N_11876,N_12114);
and U12647 (N_12647,N_11953,N_12291);
xor U12648 (N_12648,N_12012,N_12432);
or U12649 (N_12649,N_12041,N_12074);
or U12650 (N_12650,N_12425,N_11967);
or U12651 (N_12651,N_12402,N_12355);
or U12652 (N_12652,N_12375,N_12070);
xnor U12653 (N_12653,N_11983,N_12151);
and U12654 (N_12654,N_12215,N_12054);
xor U12655 (N_12655,N_11942,N_12083);
or U12656 (N_12656,N_12078,N_12203);
or U12657 (N_12657,N_12218,N_12286);
nor U12658 (N_12658,N_12029,N_12389);
nor U12659 (N_12659,N_12304,N_12414);
nor U12660 (N_12660,N_12019,N_12403);
nor U12661 (N_12661,N_12423,N_12299);
or U12662 (N_12662,N_12000,N_12071);
nor U12663 (N_12663,N_12352,N_11902);
nor U12664 (N_12664,N_12437,N_12485);
or U12665 (N_12665,N_11917,N_12288);
nand U12666 (N_12666,N_12496,N_12325);
nor U12667 (N_12667,N_12273,N_12229);
or U12668 (N_12668,N_12266,N_12230);
nor U12669 (N_12669,N_12016,N_12263);
and U12670 (N_12670,N_12370,N_12322);
nand U12671 (N_12671,N_11999,N_12276);
or U12672 (N_12672,N_12476,N_12090);
and U12673 (N_12673,N_11895,N_11974);
nand U12674 (N_12674,N_12068,N_12257);
nor U12675 (N_12675,N_12062,N_11982);
nor U12676 (N_12676,N_12498,N_11915);
or U12677 (N_12677,N_12392,N_12161);
xor U12678 (N_12678,N_12426,N_12130);
or U12679 (N_12679,N_12073,N_12217);
and U12680 (N_12680,N_12148,N_11984);
and U12681 (N_12681,N_12014,N_12081);
nor U12682 (N_12682,N_11962,N_12155);
xnor U12683 (N_12683,N_11961,N_11944);
nor U12684 (N_12684,N_12373,N_12465);
nand U12685 (N_12685,N_11919,N_12031);
or U12686 (N_12686,N_12381,N_12347);
and U12687 (N_12687,N_12317,N_12434);
xor U12688 (N_12688,N_11958,N_12424);
and U12689 (N_12689,N_12047,N_12131);
xnor U12690 (N_12690,N_12391,N_12420);
and U12691 (N_12691,N_12315,N_11875);
nor U12692 (N_12692,N_12109,N_12198);
nand U12693 (N_12693,N_12129,N_12285);
and U12694 (N_12694,N_12474,N_12184);
or U12695 (N_12695,N_11969,N_12183);
nand U12696 (N_12696,N_12409,N_12241);
or U12697 (N_12697,N_12443,N_11968);
xnor U12698 (N_12698,N_12466,N_11960);
nand U12699 (N_12699,N_11899,N_12058);
nor U12700 (N_12700,N_11997,N_12163);
or U12701 (N_12701,N_11989,N_11987);
nand U12702 (N_12702,N_11957,N_12282);
xor U12703 (N_12703,N_12231,N_12240);
xor U12704 (N_12704,N_12174,N_12399);
or U12705 (N_12705,N_12024,N_11923);
and U12706 (N_12706,N_12003,N_12275);
xor U12707 (N_12707,N_12430,N_11941);
xnor U12708 (N_12708,N_12120,N_12497);
nand U12709 (N_12709,N_11897,N_11979);
xor U12710 (N_12710,N_12197,N_12116);
xor U12711 (N_12711,N_12132,N_12178);
xnor U12712 (N_12712,N_11954,N_12372);
xnor U12713 (N_12713,N_12086,N_12247);
nand U12714 (N_12714,N_12321,N_12459);
xor U12715 (N_12715,N_12287,N_12360);
nor U12716 (N_12716,N_11951,N_11966);
or U12717 (N_12717,N_12112,N_11952);
xor U12718 (N_12718,N_12484,N_12219);
or U12719 (N_12719,N_12160,N_12470);
nand U12720 (N_12720,N_12050,N_12187);
and U12721 (N_12721,N_12126,N_12297);
or U12722 (N_12722,N_12009,N_12115);
nor U12723 (N_12723,N_12295,N_12141);
nor U12724 (N_12724,N_12255,N_11927);
nor U12725 (N_12725,N_12254,N_12468);
nor U12726 (N_12726,N_11992,N_12310);
xor U12727 (N_12727,N_12377,N_12224);
nor U12728 (N_12728,N_12123,N_12477);
and U12729 (N_12729,N_12028,N_11996);
or U12730 (N_12730,N_11910,N_12262);
xor U12731 (N_12731,N_12415,N_12256);
nand U12732 (N_12732,N_12453,N_11945);
or U12733 (N_12733,N_12440,N_12427);
nand U12734 (N_12734,N_12467,N_12320);
nor U12735 (N_12735,N_12324,N_11993);
nand U12736 (N_12736,N_12385,N_12445);
nand U12737 (N_12737,N_12195,N_12491);
and U12738 (N_12738,N_12398,N_11900);
or U12739 (N_12739,N_12499,N_11929);
xnor U12740 (N_12740,N_12448,N_12111);
nand U12741 (N_12741,N_12307,N_11887);
and U12742 (N_12742,N_11935,N_12020);
and U12743 (N_12743,N_11906,N_12103);
and U12744 (N_12744,N_12261,N_12487);
xnor U12745 (N_12745,N_12367,N_12371);
nand U12746 (N_12746,N_11918,N_11886);
nor U12747 (N_12747,N_12216,N_12186);
nor U12748 (N_12748,N_12021,N_12118);
and U12749 (N_12749,N_12110,N_12376);
or U12750 (N_12750,N_12239,N_11893);
nor U12751 (N_12751,N_12314,N_12493);
and U12752 (N_12752,N_12386,N_12436);
and U12753 (N_12753,N_12150,N_12220);
and U12754 (N_12754,N_12350,N_12396);
or U12755 (N_12755,N_12032,N_12334);
xnor U12756 (N_12756,N_12044,N_11940);
or U12757 (N_12757,N_11930,N_12205);
xnor U12758 (N_12758,N_12088,N_12036);
or U12759 (N_12759,N_11955,N_12207);
nand U12760 (N_12760,N_12076,N_11920);
and U12761 (N_12761,N_12341,N_11949);
xor U12762 (N_12762,N_12045,N_12124);
and U12763 (N_12763,N_12378,N_12221);
nor U12764 (N_12764,N_12128,N_12136);
nand U12765 (N_12765,N_12043,N_12175);
or U12766 (N_12766,N_12046,N_11991);
nand U12767 (N_12767,N_12137,N_12232);
xor U12768 (N_12768,N_12404,N_12042);
or U12769 (N_12769,N_12039,N_11994);
or U12770 (N_12770,N_12374,N_12343);
and U12771 (N_12771,N_11880,N_12152);
nand U12772 (N_12772,N_12346,N_12446);
nor U12773 (N_12773,N_12408,N_12007);
xnor U12774 (N_12774,N_12092,N_12309);
and U12775 (N_12775,N_12272,N_11939);
xor U12776 (N_12776,N_11946,N_12098);
nand U12777 (N_12777,N_12463,N_12034);
or U12778 (N_12778,N_12339,N_12354);
and U12779 (N_12779,N_11884,N_12061);
or U12780 (N_12780,N_12139,N_12089);
or U12781 (N_12781,N_12142,N_12365);
nor U12782 (N_12782,N_12421,N_12435);
or U12783 (N_12783,N_12303,N_12323);
xor U12784 (N_12784,N_11973,N_12018);
nand U12785 (N_12785,N_12159,N_11907);
nand U12786 (N_12786,N_12492,N_12055);
and U12787 (N_12787,N_12401,N_12140);
and U12788 (N_12788,N_12450,N_12329);
nand U12789 (N_12789,N_12265,N_12316);
and U12790 (N_12790,N_12237,N_12417);
xor U12791 (N_12791,N_11986,N_12106);
xnor U12792 (N_12792,N_12296,N_12033);
and U12793 (N_12793,N_12363,N_11985);
or U12794 (N_12794,N_12342,N_12176);
xor U12795 (N_12795,N_12301,N_11977);
and U12796 (N_12796,N_12464,N_12428);
nand U12797 (N_12797,N_12439,N_12260);
and U12798 (N_12798,N_12380,N_12156);
and U12799 (N_12799,N_11937,N_12094);
xnor U12800 (N_12800,N_12206,N_12283);
and U12801 (N_12801,N_12153,N_12017);
xor U12802 (N_12802,N_11978,N_12333);
nand U12803 (N_12803,N_12038,N_12075);
or U12804 (N_12804,N_12182,N_12271);
nand U12805 (N_12805,N_11926,N_12051);
or U12806 (N_12806,N_12410,N_11894);
nand U12807 (N_12807,N_12433,N_12013);
nand U12808 (N_12808,N_12122,N_12397);
or U12809 (N_12809,N_12190,N_12454);
nand U12810 (N_12810,N_12328,N_12084);
xnor U12811 (N_12811,N_11998,N_11903);
nand U12812 (N_12812,N_12330,N_12391);
xnor U12813 (N_12813,N_12419,N_12343);
and U12814 (N_12814,N_12426,N_12321);
or U12815 (N_12815,N_12355,N_12177);
xnor U12816 (N_12816,N_12341,N_12120);
nand U12817 (N_12817,N_12109,N_12443);
and U12818 (N_12818,N_11895,N_11968);
and U12819 (N_12819,N_12350,N_12299);
xor U12820 (N_12820,N_11922,N_11904);
and U12821 (N_12821,N_12207,N_11960);
or U12822 (N_12822,N_12392,N_12039);
or U12823 (N_12823,N_11883,N_11985);
nand U12824 (N_12824,N_12082,N_12065);
or U12825 (N_12825,N_12211,N_11877);
and U12826 (N_12826,N_11929,N_12010);
or U12827 (N_12827,N_12221,N_12471);
nand U12828 (N_12828,N_12257,N_11909);
nand U12829 (N_12829,N_12466,N_12497);
nor U12830 (N_12830,N_11991,N_12159);
and U12831 (N_12831,N_12219,N_12399);
or U12832 (N_12832,N_12006,N_11958);
or U12833 (N_12833,N_12089,N_12359);
nor U12834 (N_12834,N_12407,N_11927);
or U12835 (N_12835,N_12226,N_12463);
xnor U12836 (N_12836,N_12447,N_12489);
nor U12837 (N_12837,N_12202,N_12013);
xor U12838 (N_12838,N_12085,N_12182);
nand U12839 (N_12839,N_12240,N_12480);
nor U12840 (N_12840,N_12194,N_12386);
nor U12841 (N_12841,N_12451,N_11994);
or U12842 (N_12842,N_12494,N_12361);
nor U12843 (N_12843,N_11953,N_12212);
or U12844 (N_12844,N_12053,N_12028);
nand U12845 (N_12845,N_12205,N_12097);
and U12846 (N_12846,N_11942,N_11955);
and U12847 (N_12847,N_12192,N_11963);
nand U12848 (N_12848,N_12491,N_12107);
nor U12849 (N_12849,N_12053,N_12255);
or U12850 (N_12850,N_12347,N_12252);
nor U12851 (N_12851,N_12285,N_12082);
nand U12852 (N_12852,N_12044,N_12401);
nor U12853 (N_12853,N_12089,N_12043);
and U12854 (N_12854,N_12318,N_12457);
nand U12855 (N_12855,N_12292,N_12317);
xnor U12856 (N_12856,N_12001,N_12265);
nand U12857 (N_12857,N_12409,N_12363);
nand U12858 (N_12858,N_12100,N_12350);
xor U12859 (N_12859,N_12266,N_12348);
or U12860 (N_12860,N_12375,N_12168);
nor U12861 (N_12861,N_12002,N_11883);
and U12862 (N_12862,N_12409,N_12038);
nor U12863 (N_12863,N_12390,N_12387);
nor U12864 (N_12864,N_11944,N_12154);
nand U12865 (N_12865,N_12415,N_11942);
nor U12866 (N_12866,N_11878,N_12122);
or U12867 (N_12867,N_12308,N_12376);
nand U12868 (N_12868,N_12253,N_12373);
xor U12869 (N_12869,N_11947,N_11920);
xnor U12870 (N_12870,N_12484,N_11927);
or U12871 (N_12871,N_12110,N_12067);
xor U12872 (N_12872,N_11974,N_12259);
and U12873 (N_12873,N_12074,N_12403);
and U12874 (N_12874,N_12302,N_11876);
xnor U12875 (N_12875,N_12420,N_11993);
xnor U12876 (N_12876,N_11884,N_11952);
nand U12877 (N_12877,N_12148,N_12276);
xnor U12878 (N_12878,N_12334,N_12393);
or U12879 (N_12879,N_12195,N_12016);
and U12880 (N_12880,N_12371,N_12079);
xnor U12881 (N_12881,N_12214,N_12403);
nor U12882 (N_12882,N_12358,N_11915);
nand U12883 (N_12883,N_12202,N_12010);
xor U12884 (N_12884,N_12308,N_12244);
nand U12885 (N_12885,N_12154,N_12458);
and U12886 (N_12886,N_12248,N_11941);
or U12887 (N_12887,N_12079,N_12106);
nand U12888 (N_12888,N_12093,N_12358);
nand U12889 (N_12889,N_12462,N_11980);
nand U12890 (N_12890,N_12101,N_12393);
and U12891 (N_12891,N_12032,N_12255);
nand U12892 (N_12892,N_12257,N_12394);
nor U12893 (N_12893,N_11957,N_11911);
xnor U12894 (N_12894,N_12226,N_11910);
or U12895 (N_12895,N_11910,N_12198);
xnor U12896 (N_12896,N_12487,N_12191);
nand U12897 (N_12897,N_12425,N_12131);
xor U12898 (N_12898,N_12250,N_12329);
nand U12899 (N_12899,N_11923,N_12182);
nor U12900 (N_12900,N_12416,N_12007);
nand U12901 (N_12901,N_11962,N_11972);
xor U12902 (N_12902,N_12090,N_12250);
and U12903 (N_12903,N_12498,N_12315);
or U12904 (N_12904,N_12265,N_12465);
xnor U12905 (N_12905,N_11926,N_12417);
nor U12906 (N_12906,N_12235,N_12340);
nor U12907 (N_12907,N_12191,N_12478);
xnor U12908 (N_12908,N_12337,N_12159);
xnor U12909 (N_12909,N_12360,N_12446);
or U12910 (N_12910,N_12124,N_12041);
or U12911 (N_12911,N_12271,N_11935);
nor U12912 (N_12912,N_12489,N_11939);
nor U12913 (N_12913,N_12210,N_11966);
xnor U12914 (N_12914,N_11941,N_11912);
xnor U12915 (N_12915,N_12404,N_12433);
or U12916 (N_12916,N_12153,N_12395);
and U12917 (N_12917,N_12488,N_11988);
nor U12918 (N_12918,N_12379,N_11886);
and U12919 (N_12919,N_12224,N_12302);
nor U12920 (N_12920,N_11943,N_11897);
or U12921 (N_12921,N_12331,N_12140);
nor U12922 (N_12922,N_12059,N_12117);
and U12923 (N_12923,N_11970,N_12439);
nand U12924 (N_12924,N_11939,N_12229);
nand U12925 (N_12925,N_12249,N_12343);
nand U12926 (N_12926,N_12045,N_12386);
nor U12927 (N_12927,N_11923,N_12361);
nand U12928 (N_12928,N_12235,N_12106);
or U12929 (N_12929,N_11891,N_12216);
nand U12930 (N_12930,N_12065,N_11927);
nand U12931 (N_12931,N_11894,N_12015);
or U12932 (N_12932,N_12418,N_12443);
xnor U12933 (N_12933,N_12449,N_11888);
xor U12934 (N_12934,N_12243,N_12362);
nand U12935 (N_12935,N_12418,N_12080);
nor U12936 (N_12936,N_12105,N_12004);
and U12937 (N_12937,N_12268,N_12054);
and U12938 (N_12938,N_12321,N_12072);
nand U12939 (N_12939,N_12134,N_12371);
nand U12940 (N_12940,N_11975,N_12324);
or U12941 (N_12941,N_12321,N_12469);
xnor U12942 (N_12942,N_11951,N_12032);
and U12943 (N_12943,N_12476,N_12303);
or U12944 (N_12944,N_11926,N_12319);
and U12945 (N_12945,N_12277,N_12106);
and U12946 (N_12946,N_12276,N_12174);
nor U12947 (N_12947,N_12220,N_12167);
and U12948 (N_12948,N_11911,N_12031);
nor U12949 (N_12949,N_12232,N_12456);
or U12950 (N_12950,N_12124,N_12139);
nor U12951 (N_12951,N_12031,N_12398);
nor U12952 (N_12952,N_11926,N_12457);
xnor U12953 (N_12953,N_12481,N_12407);
nor U12954 (N_12954,N_12438,N_12235);
and U12955 (N_12955,N_12272,N_12050);
nor U12956 (N_12956,N_12092,N_12479);
nand U12957 (N_12957,N_12253,N_12099);
xor U12958 (N_12958,N_12481,N_12187);
and U12959 (N_12959,N_12091,N_12424);
and U12960 (N_12960,N_12115,N_12114);
nand U12961 (N_12961,N_11894,N_12448);
nor U12962 (N_12962,N_11910,N_12164);
and U12963 (N_12963,N_12158,N_11895);
xnor U12964 (N_12964,N_12263,N_12014);
and U12965 (N_12965,N_11887,N_11982);
nand U12966 (N_12966,N_12303,N_12209);
nor U12967 (N_12967,N_12295,N_12078);
xor U12968 (N_12968,N_12217,N_12486);
or U12969 (N_12969,N_12153,N_12032);
nand U12970 (N_12970,N_12407,N_12241);
nor U12971 (N_12971,N_12443,N_11919);
and U12972 (N_12972,N_12200,N_12069);
xor U12973 (N_12973,N_12361,N_12488);
nor U12974 (N_12974,N_11898,N_12421);
xor U12975 (N_12975,N_12142,N_11894);
nand U12976 (N_12976,N_12474,N_12057);
nor U12977 (N_12977,N_12291,N_12144);
xor U12978 (N_12978,N_12017,N_12089);
and U12979 (N_12979,N_12190,N_12077);
xor U12980 (N_12980,N_12093,N_12482);
nor U12981 (N_12981,N_11924,N_12061);
nand U12982 (N_12982,N_12493,N_12040);
and U12983 (N_12983,N_12032,N_12189);
or U12984 (N_12984,N_12084,N_12053);
or U12985 (N_12985,N_12259,N_12211);
and U12986 (N_12986,N_12469,N_11886);
nor U12987 (N_12987,N_11926,N_11914);
or U12988 (N_12988,N_12074,N_12199);
nand U12989 (N_12989,N_12383,N_12289);
xnor U12990 (N_12990,N_12346,N_11976);
nor U12991 (N_12991,N_12001,N_12096);
nor U12992 (N_12992,N_12250,N_12179);
or U12993 (N_12993,N_12462,N_12014);
and U12994 (N_12994,N_12295,N_11886);
and U12995 (N_12995,N_12480,N_12317);
or U12996 (N_12996,N_11930,N_12200);
xor U12997 (N_12997,N_12451,N_11976);
nor U12998 (N_12998,N_11989,N_12475);
nor U12999 (N_12999,N_12407,N_12339);
nor U13000 (N_13000,N_12258,N_12022);
xnor U13001 (N_13001,N_12243,N_12440);
xor U13002 (N_13002,N_12469,N_12056);
nand U13003 (N_13003,N_11892,N_12347);
and U13004 (N_13004,N_12196,N_12015);
or U13005 (N_13005,N_12177,N_12268);
xor U13006 (N_13006,N_11962,N_12368);
nor U13007 (N_13007,N_12250,N_12010);
nand U13008 (N_13008,N_12436,N_12115);
nor U13009 (N_13009,N_12283,N_12392);
or U13010 (N_13010,N_12478,N_12415);
and U13011 (N_13011,N_12133,N_12385);
or U13012 (N_13012,N_12180,N_12025);
xor U13013 (N_13013,N_11976,N_12403);
nor U13014 (N_13014,N_12452,N_12258);
xor U13015 (N_13015,N_12015,N_12155);
nand U13016 (N_13016,N_12386,N_12301);
nand U13017 (N_13017,N_12495,N_12475);
xnor U13018 (N_13018,N_12353,N_12318);
or U13019 (N_13019,N_12208,N_11875);
xor U13020 (N_13020,N_12075,N_12216);
and U13021 (N_13021,N_12329,N_12365);
and U13022 (N_13022,N_12007,N_11944);
xnor U13023 (N_13023,N_12353,N_12076);
nor U13024 (N_13024,N_12335,N_12460);
and U13025 (N_13025,N_11907,N_12436);
nand U13026 (N_13026,N_12262,N_12356);
nor U13027 (N_13027,N_12467,N_12160);
or U13028 (N_13028,N_11997,N_12283);
nand U13029 (N_13029,N_11900,N_12019);
xor U13030 (N_13030,N_11932,N_12425);
nand U13031 (N_13031,N_12436,N_12159);
nor U13032 (N_13032,N_12387,N_11934);
xor U13033 (N_13033,N_12238,N_12237);
nand U13034 (N_13034,N_12440,N_11971);
and U13035 (N_13035,N_11928,N_12462);
xor U13036 (N_13036,N_12084,N_12301);
nor U13037 (N_13037,N_12285,N_12343);
nor U13038 (N_13038,N_12155,N_11932);
nor U13039 (N_13039,N_12276,N_12240);
nor U13040 (N_13040,N_12022,N_12035);
nor U13041 (N_13041,N_12063,N_12482);
or U13042 (N_13042,N_12364,N_12325);
nor U13043 (N_13043,N_12467,N_12495);
nor U13044 (N_13044,N_11922,N_12043);
and U13045 (N_13045,N_12201,N_12389);
and U13046 (N_13046,N_12292,N_11922);
or U13047 (N_13047,N_12187,N_12208);
nor U13048 (N_13048,N_12155,N_12121);
or U13049 (N_13049,N_12210,N_12298);
xnor U13050 (N_13050,N_12244,N_12395);
nor U13051 (N_13051,N_12138,N_11912);
nand U13052 (N_13052,N_12478,N_12278);
nand U13053 (N_13053,N_12436,N_12183);
nor U13054 (N_13054,N_11998,N_12158);
or U13055 (N_13055,N_11916,N_12034);
nand U13056 (N_13056,N_12451,N_12351);
nand U13057 (N_13057,N_12146,N_12402);
nand U13058 (N_13058,N_12304,N_12303);
or U13059 (N_13059,N_11938,N_12398);
xnor U13060 (N_13060,N_12391,N_12476);
nand U13061 (N_13061,N_12386,N_12407);
nand U13062 (N_13062,N_11891,N_12388);
nand U13063 (N_13063,N_11949,N_11964);
xor U13064 (N_13064,N_12017,N_12199);
nand U13065 (N_13065,N_11882,N_12313);
nand U13066 (N_13066,N_12120,N_12086);
nor U13067 (N_13067,N_12039,N_12275);
nor U13068 (N_13068,N_12259,N_12348);
and U13069 (N_13069,N_12045,N_11903);
nor U13070 (N_13070,N_12194,N_11878);
xor U13071 (N_13071,N_12073,N_12235);
xnor U13072 (N_13072,N_12195,N_12103);
and U13073 (N_13073,N_11959,N_12281);
nor U13074 (N_13074,N_12396,N_11921);
or U13075 (N_13075,N_12360,N_11924);
nor U13076 (N_13076,N_12441,N_12020);
or U13077 (N_13077,N_12485,N_12087);
or U13078 (N_13078,N_12255,N_12007);
xor U13079 (N_13079,N_12226,N_12294);
or U13080 (N_13080,N_12491,N_12197);
nor U13081 (N_13081,N_11938,N_12325);
nor U13082 (N_13082,N_12330,N_12437);
and U13083 (N_13083,N_12189,N_12047);
nand U13084 (N_13084,N_12414,N_12388);
nand U13085 (N_13085,N_12211,N_12149);
xor U13086 (N_13086,N_12033,N_12088);
nand U13087 (N_13087,N_12229,N_12346);
or U13088 (N_13088,N_11960,N_12383);
nand U13089 (N_13089,N_12368,N_12028);
nand U13090 (N_13090,N_11913,N_12455);
nand U13091 (N_13091,N_11894,N_12041);
nand U13092 (N_13092,N_12224,N_12316);
nor U13093 (N_13093,N_12298,N_11905);
nor U13094 (N_13094,N_11963,N_12479);
or U13095 (N_13095,N_11957,N_12054);
and U13096 (N_13096,N_12370,N_12004);
nand U13097 (N_13097,N_12353,N_12396);
or U13098 (N_13098,N_12224,N_12156);
and U13099 (N_13099,N_11894,N_12323);
xor U13100 (N_13100,N_12374,N_12443);
xnor U13101 (N_13101,N_12476,N_12081);
xor U13102 (N_13102,N_12404,N_12266);
xor U13103 (N_13103,N_12378,N_12428);
xnor U13104 (N_13104,N_11956,N_11980);
nor U13105 (N_13105,N_11970,N_11952);
and U13106 (N_13106,N_11901,N_11983);
xnor U13107 (N_13107,N_12116,N_12278);
nand U13108 (N_13108,N_12141,N_12350);
nand U13109 (N_13109,N_11890,N_12043);
xor U13110 (N_13110,N_12300,N_12024);
or U13111 (N_13111,N_12020,N_11876);
nand U13112 (N_13112,N_12448,N_11933);
xnor U13113 (N_13113,N_12119,N_12442);
xnor U13114 (N_13114,N_12003,N_12086);
or U13115 (N_13115,N_12184,N_12017);
xnor U13116 (N_13116,N_12244,N_12372);
nand U13117 (N_13117,N_12454,N_12302);
or U13118 (N_13118,N_12163,N_12326);
nor U13119 (N_13119,N_11893,N_12044);
or U13120 (N_13120,N_12284,N_12242);
and U13121 (N_13121,N_12486,N_12265);
or U13122 (N_13122,N_12287,N_12007);
nand U13123 (N_13123,N_11918,N_12300);
or U13124 (N_13124,N_11978,N_12374);
xnor U13125 (N_13125,N_12654,N_13042);
or U13126 (N_13126,N_13010,N_12607);
nand U13127 (N_13127,N_12627,N_12759);
and U13128 (N_13128,N_12534,N_12705);
nand U13129 (N_13129,N_12750,N_12777);
and U13130 (N_13130,N_12771,N_12787);
or U13131 (N_13131,N_12743,N_12990);
nand U13132 (N_13132,N_12576,N_12852);
nor U13133 (N_13133,N_13002,N_12675);
and U13134 (N_13134,N_12506,N_13078);
and U13135 (N_13135,N_12543,N_12657);
and U13136 (N_13136,N_12755,N_12826);
nand U13137 (N_13137,N_13004,N_12805);
nor U13138 (N_13138,N_12742,N_12925);
and U13139 (N_13139,N_13061,N_12979);
nand U13140 (N_13140,N_12850,N_12948);
and U13141 (N_13141,N_12545,N_12954);
xor U13142 (N_13142,N_12996,N_12728);
xor U13143 (N_13143,N_13031,N_13067);
xnor U13144 (N_13144,N_12942,N_12868);
nor U13145 (N_13145,N_12569,N_12514);
and U13146 (N_13146,N_12516,N_12571);
xor U13147 (N_13147,N_12653,N_12773);
and U13148 (N_13148,N_12770,N_12873);
nor U13149 (N_13149,N_12790,N_12574);
or U13150 (N_13150,N_13100,N_12587);
and U13151 (N_13151,N_12918,N_12929);
and U13152 (N_13152,N_12685,N_12949);
nand U13153 (N_13153,N_13083,N_12781);
nand U13154 (N_13154,N_12508,N_12647);
nor U13155 (N_13155,N_12941,N_12798);
nor U13156 (N_13156,N_13107,N_12839);
and U13157 (N_13157,N_13124,N_12994);
nand U13158 (N_13158,N_12749,N_12557);
nand U13159 (N_13159,N_13085,N_13000);
xnor U13160 (N_13160,N_12503,N_13068);
or U13161 (N_13161,N_13087,N_13081);
xnor U13162 (N_13162,N_12811,N_12993);
and U13163 (N_13163,N_13027,N_12582);
or U13164 (N_13164,N_12519,N_12875);
nor U13165 (N_13165,N_12695,N_13065);
nor U13166 (N_13166,N_12637,N_12776);
or U13167 (N_13167,N_12639,N_12783);
and U13168 (N_13168,N_12565,N_12830);
or U13169 (N_13169,N_12838,N_12870);
nor U13170 (N_13170,N_12718,N_12761);
xnor U13171 (N_13171,N_12558,N_12601);
and U13172 (N_13172,N_13096,N_13095);
and U13173 (N_13173,N_12577,N_12735);
xor U13174 (N_13174,N_12959,N_12936);
and U13175 (N_13175,N_12600,N_12694);
or U13176 (N_13176,N_12589,N_12943);
or U13177 (N_13177,N_12917,N_12691);
and U13178 (N_13178,N_12524,N_12840);
and U13179 (N_13179,N_12765,N_13059);
nor U13180 (N_13180,N_12902,N_12832);
nand U13181 (N_13181,N_12843,N_12779);
nor U13182 (N_13182,N_13074,N_12853);
nor U13183 (N_13183,N_12976,N_12937);
and U13184 (N_13184,N_12624,N_12640);
nor U13185 (N_13185,N_12592,N_12769);
or U13186 (N_13186,N_12611,N_12971);
and U13187 (N_13187,N_13036,N_12594);
or U13188 (N_13188,N_12899,N_12872);
or U13189 (N_13189,N_12904,N_12740);
xnor U13190 (N_13190,N_13051,N_12803);
or U13191 (N_13191,N_12836,N_12615);
or U13192 (N_13192,N_13043,N_12860);
nor U13193 (N_13193,N_12752,N_13120);
nand U13194 (N_13194,N_12513,N_12580);
or U13195 (N_13195,N_12597,N_12766);
nor U13196 (N_13196,N_12876,N_12586);
and U13197 (N_13197,N_13073,N_13116);
and U13198 (N_13198,N_12567,N_12633);
xnor U13199 (N_13199,N_12612,N_12505);
nor U13200 (N_13200,N_13017,N_12704);
nand U13201 (N_13201,N_12537,N_12609);
nor U13202 (N_13202,N_12914,N_12856);
xnor U13203 (N_13203,N_12699,N_12896);
xnor U13204 (N_13204,N_12898,N_13021);
nand U13205 (N_13205,N_12989,N_12882);
xnor U13206 (N_13206,N_12634,N_13114);
or U13207 (N_13207,N_12613,N_12813);
nor U13208 (N_13208,N_12707,N_12712);
nand U13209 (N_13209,N_12523,N_12730);
or U13210 (N_13210,N_12906,N_12664);
xnor U13211 (N_13211,N_12665,N_12668);
or U13212 (N_13212,N_12884,N_12900);
nand U13213 (N_13213,N_12683,N_13121);
nor U13214 (N_13214,N_12784,N_12982);
nand U13215 (N_13215,N_12760,N_12926);
nand U13216 (N_13216,N_12854,N_12525);
nor U13217 (N_13217,N_12945,N_12541);
xnor U13218 (N_13218,N_12535,N_12867);
xor U13219 (N_13219,N_12628,N_12751);
xor U13220 (N_13220,N_13039,N_12590);
or U13221 (N_13221,N_12824,N_12630);
nor U13222 (N_13222,N_13093,N_12967);
nor U13223 (N_13223,N_12602,N_12720);
xnor U13224 (N_13224,N_13052,N_12794);
xor U13225 (N_13225,N_13032,N_12999);
and U13226 (N_13226,N_12593,N_12905);
nor U13227 (N_13227,N_12969,N_12828);
xor U13228 (N_13228,N_12673,N_13006);
xor U13229 (N_13229,N_12754,N_13025);
nand U13230 (N_13230,N_13101,N_12814);
and U13231 (N_13231,N_12762,N_12666);
nor U13232 (N_13232,N_12578,N_12809);
or U13233 (N_13233,N_12672,N_12964);
xor U13234 (N_13234,N_13047,N_12539);
and U13235 (N_13235,N_12901,N_12572);
or U13236 (N_13236,N_12745,N_12913);
or U13237 (N_13237,N_12864,N_12570);
or U13238 (N_13238,N_12625,N_12866);
and U13239 (N_13239,N_12512,N_12804);
or U13240 (N_13240,N_12818,N_12642);
xnor U13241 (N_13241,N_13038,N_13044);
and U13242 (N_13242,N_12502,N_12616);
or U13243 (N_13243,N_13098,N_13086);
or U13244 (N_13244,N_12983,N_12738);
nand U13245 (N_13245,N_12603,N_12975);
nor U13246 (N_13246,N_13020,N_12529);
nor U13247 (N_13247,N_12518,N_12833);
nand U13248 (N_13248,N_13123,N_12658);
and U13249 (N_13249,N_12885,N_12903);
and U13250 (N_13250,N_12509,N_12511);
and U13251 (N_13251,N_12845,N_13056);
and U13252 (N_13252,N_13001,N_12617);
or U13253 (N_13253,N_12897,N_12656);
or U13254 (N_13254,N_13041,N_13058);
nand U13255 (N_13255,N_12895,N_12931);
nand U13256 (N_13256,N_12693,N_13069);
xnor U13257 (N_13257,N_12702,N_12561);
nor U13258 (N_13258,N_12563,N_12659);
or U13259 (N_13259,N_12552,N_12566);
or U13260 (N_13260,N_12528,N_13024);
or U13261 (N_13261,N_12802,N_12973);
and U13262 (N_13262,N_12504,N_12823);
and U13263 (N_13263,N_12962,N_12927);
xor U13264 (N_13264,N_12646,N_12662);
nand U13265 (N_13265,N_12741,N_12579);
or U13266 (N_13266,N_12692,N_12938);
nor U13267 (N_13267,N_13048,N_13111);
and U13268 (N_13268,N_12965,N_12972);
nand U13269 (N_13269,N_12756,N_12871);
and U13270 (N_13270,N_12584,N_12661);
xnor U13271 (N_13271,N_12689,N_12889);
nand U13272 (N_13272,N_12588,N_12928);
nand U13273 (N_13273,N_12799,N_13018);
nand U13274 (N_13274,N_13094,N_12961);
xnor U13275 (N_13275,N_12677,N_12977);
nand U13276 (N_13276,N_12690,N_12688);
and U13277 (N_13277,N_12785,N_12703);
or U13278 (N_13278,N_12869,N_12786);
or U13279 (N_13279,N_12599,N_12955);
xnor U13280 (N_13280,N_12556,N_12985);
and U13281 (N_13281,N_12651,N_12890);
nor U13282 (N_13282,N_12851,N_12550);
or U13283 (N_13283,N_12546,N_12669);
and U13284 (N_13284,N_12924,N_12939);
nand U13285 (N_13285,N_12713,N_12758);
nand U13286 (N_13286,N_12629,N_13060);
and U13287 (N_13287,N_12731,N_12923);
and U13288 (N_13288,N_12829,N_12841);
and U13289 (N_13289,N_12831,N_12547);
and U13290 (N_13290,N_13102,N_13072);
xnor U13291 (N_13291,N_12536,N_12636);
nand U13292 (N_13292,N_12951,N_12892);
nor U13293 (N_13293,N_12700,N_12966);
or U13294 (N_13294,N_12595,N_13029);
xor U13295 (N_13295,N_13092,N_12746);
and U13296 (N_13296,N_12734,N_13105);
xnor U13297 (N_13297,N_13099,N_13091);
and U13298 (N_13298,N_12626,N_12963);
and U13299 (N_13299,N_13108,N_13033);
nor U13300 (N_13300,N_13028,N_12655);
and U13301 (N_13301,N_12709,N_12729);
nor U13302 (N_13302,N_12825,N_12801);
nor U13303 (N_13303,N_12527,N_12606);
nor U13304 (N_13304,N_12988,N_13050);
nand U13305 (N_13305,N_13035,N_12846);
xor U13306 (N_13306,N_12957,N_12844);
xnor U13307 (N_13307,N_12810,N_13084);
nor U13308 (N_13308,N_12671,N_12544);
or U13309 (N_13309,N_12522,N_13109);
or U13310 (N_13310,N_12879,N_12849);
or U13311 (N_13311,N_12553,N_12820);
nand U13312 (N_13312,N_13112,N_12681);
nor U13313 (N_13313,N_12568,N_13070);
xor U13314 (N_13314,N_12797,N_13103);
xnor U13315 (N_13315,N_12862,N_12632);
xnor U13316 (N_13316,N_13122,N_12583);
or U13317 (N_13317,N_12863,N_12932);
nor U13318 (N_13318,N_12916,N_13012);
nand U13319 (N_13319,N_12521,N_12542);
nand U13320 (N_13320,N_13030,N_12748);
nor U13321 (N_13321,N_12861,N_13057);
nor U13322 (N_13322,N_12591,N_12791);
xnor U13323 (N_13323,N_12944,N_13113);
and U13324 (N_13324,N_12698,N_12974);
and U13325 (N_13325,N_12635,N_12778);
nand U13326 (N_13326,N_12995,N_13045);
nor U13327 (N_13327,N_12554,N_12819);
and U13328 (N_13328,N_12711,N_12922);
nand U13329 (N_13329,N_13079,N_13104);
nor U13330 (N_13330,N_12510,N_12827);
nor U13331 (N_13331,N_12947,N_12621);
and U13332 (N_13332,N_12956,N_12724);
nand U13333 (N_13333,N_13046,N_12559);
nor U13334 (N_13334,N_12598,N_13075);
or U13335 (N_13335,N_12822,N_12644);
nand U13336 (N_13336,N_12912,N_12910);
and U13337 (N_13337,N_12878,N_13117);
or U13338 (N_13338,N_12920,N_12953);
and U13339 (N_13339,N_12782,N_12533);
nand U13340 (N_13340,N_12678,N_12835);
nor U13341 (N_13341,N_12650,N_12806);
or U13342 (N_13342,N_12911,N_13023);
or U13343 (N_13343,N_12847,N_12857);
and U13344 (N_13344,N_12865,N_13082);
nand U13345 (N_13345,N_12997,N_12701);
xor U13346 (N_13346,N_12881,N_12520);
nor U13347 (N_13347,N_12952,N_12915);
or U13348 (N_13348,N_12909,N_12517);
nand U13349 (N_13349,N_13119,N_13040);
nor U13350 (N_13350,N_12680,N_13016);
and U13351 (N_13351,N_13049,N_12793);
xor U13352 (N_13352,N_12788,N_12620);
nor U13353 (N_13353,N_12501,N_12987);
or U13354 (N_13354,N_12774,N_12679);
nand U13355 (N_13355,N_12645,N_12684);
xor U13356 (N_13356,N_12796,N_12618);
nand U13357 (N_13357,N_12807,N_12721);
nand U13358 (N_13358,N_12723,N_12815);
and U13359 (N_13359,N_12652,N_13077);
or U13360 (N_13360,N_12744,N_12562);
nor U13361 (N_13361,N_12682,N_13011);
xnor U13362 (N_13362,N_12880,N_12772);
or U13363 (N_13363,N_12667,N_13106);
nor U13364 (N_13364,N_12812,N_12526);
and U13365 (N_13365,N_12581,N_12716);
and U13366 (N_13366,N_13064,N_12883);
xor U13367 (N_13367,N_12792,N_12888);
nor U13368 (N_13368,N_12935,N_13003);
or U13369 (N_13369,N_12708,N_13089);
or U13370 (N_13370,N_12780,N_12834);
xor U13371 (N_13371,N_12732,N_12855);
nor U13372 (N_13372,N_13110,N_12631);
nand U13373 (N_13373,N_13009,N_12757);
and U13374 (N_13374,N_12960,N_12560);
xnor U13375 (N_13375,N_12767,N_12687);
or U13376 (N_13376,N_12604,N_13053);
and U13377 (N_13377,N_13054,N_12837);
nand U13378 (N_13378,N_12737,N_12725);
or U13379 (N_13379,N_12727,N_13022);
xor U13380 (N_13380,N_13076,N_12649);
or U13381 (N_13381,N_12808,N_12891);
nand U13382 (N_13382,N_12940,N_12821);
or U13383 (N_13383,N_12697,N_12933);
nor U13384 (N_13384,N_13014,N_12763);
nand U13385 (N_13385,N_12585,N_12764);
xor U13386 (N_13386,N_12573,N_12970);
nor U13387 (N_13387,N_12548,N_13097);
or U13388 (N_13388,N_13088,N_12893);
xnor U13389 (N_13389,N_13034,N_12921);
nand U13390 (N_13390,N_12946,N_12877);
or U13391 (N_13391,N_13007,N_12719);
nand U13392 (N_13392,N_12596,N_13063);
xor U13393 (N_13393,N_13015,N_12842);
or U13394 (N_13394,N_12722,N_12978);
nand U13395 (N_13395,N_12874,N_12747);
and U13396 (N_13396,N_12575,N_13037);
nand U13397 (N_13397,N_12980,N_12641);
xnor U13398 (N_13398,N_12991,N_12610);
nor U13399 (N_13399,N_12789,N_12998);
or U13400 (N_13400,N_12551,N_12908);
or U13401 (N_13401,N_12858,N_12660);
nand U13402 (N_13402,N_12564,N_13090);
xor U13403 (N_13403,N_12753,N_12958);
nand U13404 (N_13404,N_13080,N_12739);
nand U13405 (N_13405,N_12984,N_12530);
nor U13406 (N_13406,N_12859,N_12726);
nand U13407 (N_13407,N_12816,N_12608);
or U13408 (N_13408,N_13013,N_12919);
xnor U13409 (N_13409,N_12614,N_13066);
or U13410 (N_13410,N_12696,N_12515);
nand U13411 (N_13411,N_12733,N_12894);
or U13412 (N_13412,N_12538,N_12605);
and U13413 (N_13413,N_12531,N_12670);
and U13414 (N_13414,N_12714,N_12992);
and U13415 (N_13415,N_12706,N_12887);
nor U13416 (N_13416,N_12950,N_13008);
or U13417 (N_13417,N_12817,N_12930);
nor U13418 (N_13418,N_12768,N_12549);
nand U13419 (N_13419,N_12500,N_12507);
or U13420 (N_13420,N_12986,N_12619);
or U13421 (N_13421,N_12800,N_12968);
or U13422 (N_13422,N_12622,N_12686);
or U13423 (N_13423,N_13118,N_13005);
xnor U13424 (N_13424,N_13055,N_13062);
and U13425 (N_13425,N_13115,N_12848);
and U13426 (N_13426,N_12648,N_12907);
or U13427 (N_13427,N_12663,N_12643);
and U13428 (N_13428,N_12532,N_12555);
or U13429 (N_13429,N_13019,N_12715);
or U13430 (N_13430,N_12717,N_12676);
or U13431 (N_13431,N_12795,N_12736);
nor U13432 (N_13432,N_12623,N_12934);
nor U13433 (N_13433,N_12775,N_12886);
xnor U13434 (N_13434,N_12674,N_12638);
xor U13435 (N_13435,N_13026,N_12710);
and U13436 (N_13436,N_12981,N_13071);
or U13437 (N_13437,N_12540,N_12849);
xnor U13438 (N_13438,N_12543,N_13095);
and U13439 (N_13439,N_12501,N_12635);
or U13440 (N_13440,N_12917,N_13040);
or U13441 (N_13441,N_12729,N_12849);
nand U13442 (N_13442,N_12688,N_13121);
and U13443 (N_13443,N_12945,N_12549);
nand U13444 (N_13444,N_12818,N_13105);
nor U13445 (N_13445,N_12567,N_12710);
nor U13446 (N_13446,N_12799,N_12961);
and U13447 (N_13447,N_13097,N_12885);
xnor U13448 (N_13448,N_12847,N_12885);
xnor U13449 (N_13449,N_13054,N_12513);
xnor U13450 (N_13450,N_12772,N_12825);
nor U13451 (N_13451,N_12983,N_12876);
xnor U13452 (N_13452,N_12603,N_12922);
nor U13453 (N_13453,N_12917,N_12631);
or U13454 (N_13454,N_12799,N_12516);
and U13455 (N_13455,N_12857,N_12723);
nor U13456 (N_13456,N_12852,N_12745);
or U13457 (N_13457,N_13035,N_12778);
or U13458 (N_13458,N_12529,N_13035);
nand U13459 (N_13459,N_13091,N_13052);
and U13460 (N_13460,N_12740,N_13041);
nor U13461 (N_13461,N_12538,N_12694);
nor U13462 (N_13462,N_12935,N_12893);
or U13463 (N_13463,N_13117,N_12994);
xnor U13464 (N_13464,N_13039,N_12980);
and U13465 (N_13465,N_12717,N_13045);
nor U13466 (N_13466,N_12541,N_12881);
nor U13467 (N_13467,N_12716,N_13046);
nand U13468 (N_13468,N_12625,N_12565);
or U13469 (N_13469,N_12936,N_12968);
nand U13470 (N_13470,N_12951,N_12829);
and U13471 (N_13471,N_12678,N_12988);
xnor U13472 (N_13472,N_12976,N_13089);
and U13473 (N_13473,N_12809,N_12550);
xor U13474 (N_13474,N_13003,N_12951);
or U13475 (N_13475,N_12690,N_12518);
xor U13476 (N_13476,N_12553,N_12940);
nand U13477 (N_13477,N_12961,N_12526);
and U13478 (N_13478,N_13017,N_12702);
and U13479 (N_13479,N_12683,N_12658);
and U13480 (N_13480,N_12998,N_12923);
nor U13481 (N_13481,N_12954,N_12914);
nand U13482 (N_13482,N_12618,N_12828);
xor U13483 (N_13483,N_13084,N_12756);
or U13484 (N_13484,N_13115,N_12664);
or U13485 (N_13485,N_12949,N_12771);
or U13486 (N_13486,N_12872,N_13058);
and U13487 (N_13487,N_12647,N_12628);
xnor U13488 (N_13488,N_12501,N_12917);
xnor U13489 (N_13489,N_12559,N_13063);
nand U13490 (N_13490,N_13061,N_13031);
nor U13491 (N_13491,N_12987,N_12537);
nand U13492 (N_13492,N_12542,N_13103);
xor U13493 (N_13493,N_12902,N_12759);
and U13494 (N_13494,N_12573,N_12601);
xor U13495 (N_13495,N_12594,N_12710);
nor U13496 (N_13496,N_12553,N_12548);
xnor U13497 (N_13497,N_12531,N_12754);
or U13498 (N_13498,N_12976,N_13109);
or U13499 (N_13499,N_13028,N_12927);
nand U13500 (N_13500,N_12620,N_13064);
xor U13501 (N_13501,N_13063,N_12796);
or U13502 (N_13502,N_12923,N_13045);
or U13503 (N_13503,N_12658,N_12538);
or U13504 (N_13504,N_12560,N_13102);
nand U13505 (N_13505,N_12529,N_12934);
nand U13506 (N_13506,N_12862,N_12796);
or U13507 (N_13507,N_12706,N_12755);
or U13508 (N_13508,N_12565,N_12980);
or U13509 (N_13509,N_13045,N_13059);
nor U13510 (N_13510,N_12666,N_13113);
or U13511 (N_13511,N_12616,N_12713);
nand U13512 (N_13512,N_12854,N_12699);
or U13513 (N_13513,N_13053,N_12605);
xnor U13514 (N_13514,N_12726,N_12933);
xor U13515 (N_13515,N_12872,N_13027);
nand U13516 (N_13516,N_12904,N_12620);
nand U13517 (N_13517,N_13050,N_12555);
nand U13518 (N_13518,N_12698,N_12863);
or U13519 (N_13519,N_13091,N_13020);
xnor U13520 (N_13520,N_12854,N_12712);
and U13521 (N_13521,N_12685,N_12867);
nand U13522 (N_13522,N_12517,N_12866);
xnor U13523 (N_13523,N_12673,N_13068);
or U13524 (N_13524,N_13058,N_12854);
nand U13525 (N_13525,N_12762,N_12936);
xor U13526 (N_13526,N_12870,N_12726);
or U13527 (N_13527,N_12568,N_12680);
nand U13528 (N_13528,N_13108,N_12618);
nand U13529 (N_13529,N_12814,N_12507);
xor U13530 (N_13530,N_12760,N_12546);
xor U13531 (N_13531,N_12615,N_12997);
nand U13532 (N_13532,N_12847,N_13084);
or U13533 (N_13533,N_12674,N_12592);
or U13534 (N_13534,N_12863,N_13037);
and U13535 (N_13535,N_12614,N_12815);
or U13536 (N_13536,N_13091,N_12528);
xor U13537 (N_13537,N_12704,N_13035);
nand U13538 (N_13538,N_12737,N_12639);
nand U13539 (N_13539,N_12548,N_12515);
nor U13540 (N_13540,N_12826,N_12943);
and U13541 (N_13541,N_13090,N_12867);
nor U13542 (N_13542,N_12622,N_12811);
xnor U13543 (N_13543,N_13015,N_12973);
or U13544 (N_13544,N_12993,N_12519);
or U13545 (N_13545,N_12667,N_13080);
nand U13546 (N_13546,N_12793,N_12504);
xnor U13547 (N_13547,N_12525,N_13068);
xnor U13548 (N_13548,N_12990,N_12700);
and U13549 (N_13549,N_12893,N_12547);
and U13550 (N_13550,N_12859,N_12509);
or U13551 (N_13551,N_12862,N_12783);
xnor U13552 (N_13552,N_12655,N_13005);
nor U13553 (N_13553,N_12508,N_12701);
and U13554 (N_13554,N_13056,N_13111);
and U13555 (N_13555,N_12587,N_12701);
nor U13556 (N_13556,N_12836,N_12621);
nor U13557 (N_13557,N_12844,N_12850);
nand U13558 (N_13558,N_13122,N_13058);
nor U13559 (N_13559,N_12794,N_12715);
or U13560 (N_13560,N_12708,N_12547);
nor U13561 (N_13561,N_12654,N_12722);
nand U13562 (N_13562,N_12737,N_12795);
nand U13563 (N_13563,N_12640,N_13097);
xor U13564 (N_13564,N_12926,N_12850);
nand U13565 (N_13565,N_12868,N_13114);
nor U13566 (N_13566,N_13076,N_12784);
or U13567 (N_13567,N_13060,N_12690);
xnor U13568 (N_13568,N_12671,N_12969);
nor U13569 (N_13569,N_12860,N_12841);
nand U13570 (N_13570,N_12997,N_12845);
or U13571 (N_13571,N_12590,N_12784);
or U13572 (N_13572,N_12795,N_12938);
nor U13573 (N_13573,N_12524,N_12694);
xor U13574 (N_13574,N_12770,N_12815);
or U13575 (N_13575,N_12997,N_12856);
nor U13576 (N_13576,N_12595,N_12826);
nand U13577 (N_13577,N_12729,N_13027);
and U13578 (N_13578,N_12672,N_12666);
xnor U13579 (N_13579,N_12715,N_12942);
nor U13580 (N_13580,N_12804,N_12653);
or U13581 (N_13581,N_12959,N_12882);
nand U13582 (N_13582,N_12639,N_12644);
xnor U13583 (N_13583,N_12658,N_12558);
xnor U13584 (N_13584,N_12508,N_12648);
nor U13585 (N_13585,N_13058,N_13026);
or U13586 (N_13586,N_12737,N_12713);
and U13587 (N_13587,N_12637,N_12729);
nor U13588 (N_13588,N_12795,N_12886);
nand U13589 (N_13589,N_12739,N_12833);
xnor U13590 (N_13590,N_12704,N_12835);
nor U13591 (N_13591,N_12999,N_13055);
nand U13592 (N_13592,N_12959,N_12892);
nor U13593 (N_13593,N_13083,N_12762);
and U13594 (N_13594,N_12796,N_12636);
xnor U13595 (N_13595,N_12717,N_12664);
xnor U13596 (N_13596,N_12711,N_12739);
and U13597 (N_13597,N_12835,N_12690);
or U13598 (N_13598,N_12936,N_12845);
nand U13599 (N_13599,N_12755,N_12998);
nand U13600 (N_13600,N_12951,N_12883);
nor U13601 (N_13601,N_12738,N_13110);
nand U13602 (N_13602,N_12851,N_12797);
or U13603 (N_13603,N_13017,N_12871);
or U13604 (N_13604,N_13025,N_13060);
or U13605 (N_13605,N_12958,N_12923);
and U13606 (N_13606,N_12906,N_12970);
and U13607 (N_13607,N_13025,N_12790);
and U13608 (N_13608,N_12988,N_12849);
or U13609 (N_13609,N_13064,N_12779);
xor U13610 (N_13610,N_12985,N_12908);
and U13611 (N_13611,N_13067,N_12506);
nor U13612 (N_13612,N_12579,N_12707);
and U13613 (N_13613,N_12925,N_13105);
and U13614 (N_13614,N_12615,N_12650);
and U13615 (N_13615,N_12662,N_12650);
and U13616 (N_13616,N_12607,N_12660);
or U13617 (N_13617,N_12867,N_12597);
nor U13618 (N_13618,N_12961,N_12767);
or U13619 (N_13619,N_12706,N_12962);
and U13620 (N_13620,N_12908,N_12859);
nor U13621 (N_13621,N_12535,N_12654);
xor U13622 (N_13622,N_12865,N_12610);
and U13623 (N_13623,N_12805,N_13064);
nor U13624 (N_13624,N_12840,N_12650);
xor U13625 (N_13625,N_12707,N_12876);
or U13626 (N_13626,N_13043,N_12591);
nor U13627 (N_13627,N_12645,N_12718);
nand U13628 (N_13628,N_13092,N_12711);
nand U13629 (N_13629,N_13013,N_12530);
or U13630 (N_13630,N_12604,N_12548);
or U13631 (N_13631,N_12778,N_12633);
xnor U13632 (N_13632,N_12746,N_12625);
xor U13633 (N_13633,N_12927,N_12712);
and U13634 (N_13634,N_12733,N_13083);
or U13635 (N_13635,N_12537,N_12662);
nand U13636 (N_13636,N_12946,N_12699);
nand U13637 (N_13637,N_13056,N_13076);
or U13638 (N_13638,N_12804,N_12974);
and U13639 (N_13639,N_13047,N_12577);
or U13640 (N_13640,N_12555,N_12593);
and U13641 (N_13641,N_12833,N_12906);
nand U13642 (N_13642,N_12562,N_12664);
or U13643 (N_13643,N_12815,N_12735);
nand U13644 (N_13644,N_12757,N_13015);
and U13645 (N_13645,N_12570,N_12693);
nor U13646 (N_13646,N_12958,N_12957);
or U13647 (N_13647,N_13021,N_12752);
or U13648 (N_13648,N_12929,N_12805);
and U13649 (N_13649,N_12710,N_12997);
and U13650 (N_13650,N_12832,N_13045);
and U13651 (N_13651,N_12811,N_12772);
nor U13652 (N_13652,N_12897,N_12503);
and U13653 (N_13653,N_12582,N_12765);
or U13654 (N_13654,N_12831,N_13115);
and U13655 (N_13655,N_12680,N_12821);
nor U13656 (N_13656,N_12961,N_12873);
nand U13657 (N_13657,N_12553,N_13001);
nand U13658 (N_13658,N_12549,N_12673);
nand U13659 (N_13659,N_12735,N_12779);
xnor U13660 (N_13660,N_12540,N_12652);
xor U13661 (N_13661,N_13033,N_12958);
xor U13662 (N_13662,N_13119,N_12586);
xnor U13663 (N_13663,N_12980,N_12796);
or U13664 (N_13664,N_12534,N_12864);
nand U13665 (N_13665,N_12576,N_12715);
nor U13666 (N_13666,N_12687,N_12515);
nor U13667 (N_13667,N_12945,N_12924);
nand U13668 (N_13668,N_12662,N_12626);
nor U13669 (N_13669,N_13068,N_12852);
and U13670 (N_13670,N_12773,N_12604);
xor U13671 (N_13671,N_12709,N_12734);
xnor U13672 (N_13672,N_13054,N_12656);
or U13673 (N_13673,N_12981,N_13047);
nand U13674 (N_13674,N_12961,N_13000);
or U13675 (N_13675,N_12569,N_13100);
or U13676 (N_13676,N_12995,N_12827);
nor U13677 (N_13677,N_12669,N_13073);
nand U13678 (N_13678,N_13027,N_12556);
or U13679 (N_13679,N_12983,N_12847);
nor U13680 (N_13680,N_13019,N_12865);
and U13681 (N_13681,N_12825,N_12708);
nand U13682 (N_13682,N_12970,N_12623);
or U13683 (N_13683,N_12924,N_12510);
nand U13684 (N_13684,N_13029,N_12612);
or U13685 (N_13685,N_12998,N_12653);
nand U13686 (N_13686,N_12758,N_12730);
nand U13687 (N_13687,N_13014,N_12748);
nor U13688 (N_13688,N_12641,N_12824);
and U13689 (N_13689,N_13068,N_13050);
nor U13690 (N_13690,N_12662,N_12671);
or U13691 (N_13691,N_12717,N_12653);
and U13692 (N_13692,N_12669,N_13094);
xor U13693 (N_13693,N_12699,N_12933);
or U13694 (N_13694,N_12925,N_12660);
nand U13695 (N_13695,N_12961,N_12561);
and U13696 (N_13696,N_12729,N_13111);
nor U13697 (N_13697,N_12668,N_12938);
xnor U13698 (N_13698,N_12756,N_12839);
or U13699 (N_13699,N_12870,N_12904);
nand U13700 (N_13700,N_12598,N_13080);
nor U13701 (N_13701,N_12932,N_12598);
or U13702 (N_13702,N_12709,N_13026);
nor U13703 (N_13703,N_12517,N_12857);
xnor U13704 (N_13704,N_12546,N_12983);
or U13705 (N_13705,N_12688,N_12536);
and U13706 (N_13706,N_12884,N_12815);
or U13707 (N_13707,N_12774,N_12917);
and U13708 (N_13708,N_12505,N_12788);
xor U13709 (N_13709,N_12640,N_12806);
and U13710 (N_13710,N_12784,N_12628);
xnor U13711 (N_13711,N_12669,N_13050);
and U13712 (N_13712,N_12959,N_12728);
nor U13713 (N_13713,N_12740,N_12578);
xnor U13714 (N_13714,N_12646,N_12626);
or U13715 (N_13715,N_13033,N_12572);
or U13716 (N_13716,N_13121,N_12829);
xnor U13717 (N_13717,N_12577,N_13024);
nand U13718 (N_13718,N_12995,N_13078);
or U13719 (N_13719,N_12899,N_12668);
and U13720 (N_13720,N_12523,N_12662);
nor U13721 (N_13721,N_13104,N_13011);
xnor U13722 (N_13722,N_12758,N_13067);
nand U13723 (N_13723,N_13056,N_12943);
nor U13724 (N_13724,N_12702,N_12797);
nand U13725 (N_13725,N_12614,N_13045);
xor U13726 (N_13726,N_13076,N_13060);
or U13727 (N_13727,N_12864,N_12780);
nand U13728 (N_13728,N_12987,N_12624);
nor U13729 (N_13729,N_12728,N_12660);
and U13730 (N_13730,N_12824,N_13049);
nor U13731 (N_13731,N_13080,N_12753);
nand U13732 (N_13732,N_12920,N_12826);
xor U13733 (N_13733,N_12592,N_13073);
and U13734 (N_13734,N_12893,N_12504);
or U13735 (N_13735,N_13003,N_12590);
nor U13736 (N_13736,N_12732,N_12692);
xnor U13737 (N_13737,N_12934,N_13058);
nand U13738 (N_13738,N_13055,N_13048);
nand U13739 (N_13739,N_12593,N_12930);
xnor U13740 (N_13740,N_12988,N_12842);
xnor U13741 (N_13741,N_12836,N_12833);
nor U13742 (N_13742,N_13091,N_12555);
xor U13743 (N_13743,N_12719,N_12976);
and U13744 (N_13744,N_12840,N_12726);
nand U13745 (N_13745,N_12556,N_13008);
and U13746 (N_13746,N_13016,N_13044);
and U13747 (N_13747,N_12756,N_12592);
and U13748 (N_13748,N_12672,N_12597);
nor U13749 (N_13749,N_12940,N_12935);
nor U13750 (N_13750,N_13325,N_13657);
or U13751 (N_13751,N_13350,N_13142);
xor U13752 (N_13752,N_13282,N_13633);
nand U13753 (N_13753,N_13223,N_13339);
or U13754 (N_13754,N_13500,N_13332);
nand U13755 (N_13755,N_13689,N_13433);
nor U13756 (N_13756,N_13712,N_13519);
nor U13757 (N_13757,N_13412,N_13192);
and U13758 (N_13758,N_13386,N_13366);
nand U13759 (N_13759,N_13479,N_13193);
nand U13760 (N_13760,N_13649,N_13640);
and U13761 (N_13761,N_13336,N_13306);
nand U13762 (N_13762,N_13362,N_13221);
nor U13763 (N_13763,N_13523,N_13129);
and U13764 (N_13764,N_13602,N_13165);
nand U13765 (N_13765,N_13213,N_13662);
xnor U13766 (N_13766,N_13367,N_13423);
xnor U13767 (N_13767,N_13608,N_13283);
nor U13768 (N_13768,N_13319,N_13243);
nor U13769 (N_13769,N_13540,N_13456);
nor U13770 (N_13770,N_13302,N_13260);
xnor U13771 (N_13771,N_13395,N_13530);
nand U13772 (N_13772,N_13704,N_13733);
nand U13773 (N_13773,N_13745,N_13295);
nor U13774 (N_13774,N_13399,N_13130);
nand U13775 (N_13775,N_13700,N_13131);
and U13776 (N_13776,N_13125,N_13132);
or U13777 (N_13777,N_13368,N_13443);
and U13778 (N_13778,N_13450,N_13714);
xnor U13779 (N_13779,N_13344,N_13385);
or U13780 (N_13780,N_13206,N_13564);
or U13781 (N_13781,N_13191,N_13588);
or U13782 (N_13782,N_13343,N_13749);
and U13783 (N_13783,N_13369,N_13577);
nor U13784 (N_13784,N_13422,N_13321);
xor U13785 (N_13785,N_13454,N_13446);
and U13786 (N_13786,N_13219,N_13693);
nor U13787 (N_13787,N_13436,N_13234);
nand U13788 (N_13788,N_13708,N_13641);
xnor U13789 (N_13789,N_13465,N_13155);
nand U13790 (N_13790,N_13555,N_13383);
nand U13791 (N_13791,N_13562,N_13727);
and U13792 (N_13792,N_13384,N_13146);
nor U13793 (N_13793,N_13374,N_13291);
nor U13794 (N_13794,N_13275,N_13718);
nor U13795 (N_13795,N_13480,N_13140);
or U13796 (N_13796,N_13136,N_13476);
nand U13797 (N_13797,N_13288,N_13609);
xor U13798 (N_13798,N_13630,N_13611);
nor U13799 (N_13799,N_13468,N_13341);
nor U13800 (N_13800,N_13655,N_13496);
nand U13801 (N_13801,N_13631,N_13667);
xnor U13802 (N_13802,N_13392,N_13563);
nand U13803 (N_13803,N_13499,N_13545);
xnor U13804 (N_13804,N_13444,N_13683);
nand U13805 (N_13805,N_13181,N_13618);
or U13806 (N_13806,N_13403,N_13228);
and U13807 (N_13807,N_13590,N_13520);
nand U13808 (N_13808,N_13415,N_13370);
and U13809 (N_13809,N_13244,N_13143);
xor U13810 (N_13810,N_13691,N_13642);
xor U13811 (N_13811,N_13679,N_13535);
xor U13812 (N_13812,N_13313,N_13317);
nand U13813 (N_13813,N_13429,N_13424);
nand U13814 (N_13814,N_13717,N_13330);
nand U13815 (N_13815,N_13196,N_13303);
or U13816 (N_13816,N_13498,N_13265);
xnor U13817 (N_13817,N_13510,N_13276);
xnor U13818 (N_13818,N_13159,N_13445);
nor U13819 (N_13819,N_13485,N_13627);
nand U13820 (N_13820,N_13232,N_13477);
nand U13821 (N_13821,N_13501,N_13204);
xor U13822 (N_13822,N_13154,N_13141);
or U13823 (N_13823,N_13730,N_13380);
and U13824 (N_13824,N_13307,N_13267);
nand U13825 (N_13825,N_13684,N_13709);
and U13826 (N_13826,N_13552,N_13144);
and U13827 (N_13827,N_13646,N_13194);
nor U13828 (N_13828,N_13372,N_13175);
nand U13829 (N_13829,N_13692,N_13453);
nor U13830 (N_13830,N_13725,N_13539);
xnor U13831 (N_13831,N_13638,N_13410);
or U13832 (N_13832,N_13647,N_13721);
and U13833 (N_13833,N_13728,N_13742);
nor U13834 (N_13834,N_13599,N_13208);
or U13835 (N_13835,N_13157,N_13526);
or U13836 (N_13836,N_13387,N_13170);
nor U13837 (N_13837,N_13461,N_13508);
and U13838 (N_13838,N_13224,N_13541);
and U13839 (N_13839,N_13470,N_13162);
nand U13840 (N_13840,N_13391,N_13357);
nand U13841 (N_13841,N_13506,N_13656);
nand U13842 (N_13842,N_13360,N_13671);
nor U13843 (N_13843,N_13713,N_13351);
nand U13844 (N_13844,N_13460,N_13305);
and U13845 (N_13845,N_13285,N_13637);
and U13846 (N_13846,N_13490,N_13229);
and U13847 (N_13847,N_13658,N_13212);
or U13848 (N_13848,N_13556,N_13166);
or U13849 (N_13849,N_13582,N_13706);
or U13850 (N_13850,N_13239,N_13571);
and U13851 (N_13851,N_13626,N_13148);
xor U13852 (N_13852,N_13334,N_13682);
xnor U13853 (N_13853,N_13492,N_13598);
nand U13854 (N_13854,N_13186,N_13137);
xnor U13855 (N_13855,N_13172,N_13398);
or U13856 (N_13856,N_13363,N_13371);
or U13857 (N_13857,N_13281,N_13469);
xor U13858 (N_13858,N_13699,N_13597);
and U13859 (N_13859,N_13549,N_13722);
or U13860 (N_13860,N_13411,N_13676);
xnor U13861 (N_13861,N_13743,N_13441);
or U13862 (N_13862,N_13680,N_13438);
nand U13863 (N_13863,N_13352,N_13396);
or U13864 (N_13864,N_13472,N_13624);
nor U13865 (N_13865,N_13365,N_13377);
xnor U13866 (N_13866,N_13720,N_13327);
and U13867 (N_13867,N_13557,N_13278);
nor U13868 (N_13868,N_13458,N_13426);
nand U13869 (N_13869,N_13437,N_13734);
and U13870 (N_13870,N_13747,N_13553);
and U13871 (N_13871,N_13511,N_13304);
nor U13872 (N_13872,N_13430,N_13575);
nor U13873 (N_13873,N_13202,N_13687);
or U13874 (N_13874,N_13629,N_13688);
and U13875 (N_13875,N_13723,N_13364);
nor U13876 (N_13876,N_13634,N_13616);
xor U13877 (N_13877,N_13405,N_13199);
nand U13878 (N_13878,N_13533,N_13561);
or U13879 (N_13879,N_13613,N_13551);
and U13880 (N_13880,N_13462,N_13390);
nand U13881 (N_13881,N_13653,N_13297);
xnor U13882 (N_13882,N_13376,N_13231);
xor U13883 (N_13883,N_13690,N_13241);
xnor U13884 (N_13884,N_13279,N_13173);
xor U13885 (N_13885,N_13284,N_13299);
or U13886 (N_13886,N_13126,N_13233);
nand U13887 (N_13887,N_13169,N_13505);
or U13888 (N_13888,N_13448,N_13719);
nor U13889 (N_13889,N_13558,N_13705);
xor U13890 (N_13890,N_13489,N_13628);
nand U13891 (N_13891,N_13413,N_13340);
and U13892 (N_13892,N_13335,N_13466);
nand U13893 (N_13893,N_13666,N_13277);
nor U13894 (N_13894,N_13495,N_13271);
xor U13895 (N_13895,N_13353,N_13548);
and U13896 (N_13896,N_13428,N_13158);
xnor U13897 (N_13897,N_13715,N_13435);
and U13898 (N_13898,N_13417,N_13731);
nor U13899 (N_13899,N_13197,N_13610);
and U13900 (N_13900,N_13205,N_13513);
or U13901 (N_13901,N_13612,N_13550);
or U13902 (N_13902,N_13314,N_13529);
nor U13903 (N_13903,N_13261,N_13230);
or U13904 (N_13904,N_13685,N_13574);
and U13905 (N_13905,N_13534,N_13289);
or U13906 (N_13906,N_13536,N_13152);
and U13907 (N_13907,N_13486,N_13257);
nor U13908 (N_13908,N_13207,N_13249);
and U13909 (N_13909,N_13587,N_13250);
nor U13910 (N_13910,N_13493,N_13678);
nor U13911 (N_13911,N_13748,N_13133);
or U13912 (N_13912,N_13525,N_13711);
and U13913 (N_13913,N_13147,N_13237);
nand U13914 (N_13914,N_13179,N_13674);
xor U13915 (N_13915,N_13246,N_13654);
nand U13916 (N_13916,N_13672,N_13245);
or U13917 (N_13917,N_13503,N_13635);
nand U13918 (N_13918,N_13128,N_13559);
and U13919 (N_13919,N_13361,N_13311);
nor U13920 (N_13920,N_13702,N_13315);
nor U13921 (N_13921,N_13606,N_13607);
xnor U13922 (N_13922,N_13620,N_13168);
and U13923 (N_13923,N_13509,N_13251);
xor U13924 (N_13924,N_13560,N_13664);
or U13925 (N_13925,N_13355,N_13404);
or U13926 (N_13926,N_13670,N_13138);
xnor U13927 (N_13927,N_13238,N_13595);
nand U13928 (N_13928,N_13594,N_13639);
and U13929 (N_13929,N_13473,N_13153);
or U13930 (N_13930,N_13650,N_13252);
or U13931 (N_13931,N_13333,N_13346);
nor U13932 (N_13932,N_13164,N_13729);
nand U13933 (N_13933,N_13222,N_13308);
nand U13934 (N_13934,N_13409,N_13215);
xor U13935 (N_13935,N_13686,N_13592);
or U13936 (N_13936,N_13292,N_13488);
nand U13937 (N_13937,N_13264,N_13174);
or U13938 (N_13938,N_13544,N_13464);
or U13939 (N_13939,N_13320,N_13494);
nor U13940 (N_13940,N_13201,N_13565);
and U13941 (N_13941,N_13586,N_13452);
nand U13942 (N_13942,N_13518,N_13402);
and U13943 (N_13943,N_13431,N_13216);
nor U13944 (N_13944,N_13178,N_13139);
and U13945 (N_13945,N_13347,N_13167);
nand U13946 (N_13946,N_13570,N_13603);
nand U13947 (N_13947,N_13467,N_13440);
nor U13948 (N_13948,N_13732,N_13736);
and U13949 (N_13949,N_13487,N_13268);
nand U13950 (N_13950,N_13584,N_13724);
nor U13951 (N_13951,N_13515,N_13567);
nand U13952 (N_13952,N_13324,N_13401);
nor U13953 (N_13953,N_13601,N_13695);
or U13954 (N_13954,N_13632,N_13585);
xnor U13955 (N_13955,N_13521,N_13580);
nor U13956 (N_13956,N_13359,N_13614);
nand U13957 (N_13957,N_13439,N_13378);
or U13958 (N_13958,N_13310,N_13400);
nand U13959 (N_13959,N_13531,N_13568);
nand U13960 (N_13960,N_13375,N_13696);
or U13961 (N_13961,N_13547,N_13478);
nor U13962 (N_13962,N_13681,N_13449);
or U13963 (N_13963,N_13741,N_13593);
nor U13964 (N_13964,N_13522,N_13406);
nand U13965 (N_13965,N_13190,N_13572);
and U13966 (N_13966,N_13726,N_13419);
and U13967 (N_13967,N_13738,N_13211);
xnor U13968 (N_13968,N_13484,N_13604);
or U13969 (N_13969,N_13290,N_13701);
or U13970 (N_13970,N_13242,N_13471);
and U13971 (N_13971,N_13644,N_13171);
nor U13972 (N_13972,N_13255,N_13524);
nor U13973 (N_13973,N_13455,N_13459);
xor U13974 (N_13974,N_13161,N_13482);
or U13975 (N_13975,N_13474,N_13150);
or U13976 (N_13976,N_13176,N_13183);
and U13977 (N_13977,N_13636,N_13262);
and U13978 (N_13978,N_13625,N_13342);
nand U13979 (N_13979,N_13698,N_13189);
nor U13980 (N_13980,N_13716,N_13326);
and U13981 (N_13981,N_13293,N_13348);
and U13982 (N_13982,N_13151,N_13660);
and U13983 (N_13983,N_13349,N_13483);
nor U13984 (N_13984,N_13739,N_13566);
nand U13985 (N_13985,N_13316,N_13596);
and U13986 (N_13986,N_13270,N_13414);
xnor U13987 (N_13987,N_13675,N_13187);
xor U13988 (N_13988,N_13744,N_13298);
nor U13989 (N_13989,N_13188,N_13434);
xnor U13990 (N_13990,N_13235,N_13694);
xnor U13991 (N_13991,N_13578,N_13589);
xor U13992 (N_13992,N_13502,N_13247);
xor U13993 (N_13993,N_13673,N_13287);
xnor U13994 (N_13994,N_13418,N_13280);
nand U13995 (N_13995,N_13200,N_13328);
xnor U13996 (N_13996,N_13301,N_13354);
or U13997 (N_13997,N_13256,N_13516);
nand U13998 (N_13998,N_13648,N_13240);
xnor U13999 (N_13999,N_13156,N_13740);
nor U14000 (N_14000,N_13546,N_13149);
xnor U14001 (N_14001,N_13703,N_13248);
xor U14002 (N_14002,N_13543,N_13210);
nand U14003 (N_14003,N_13504,N_13209);
xor U14004 (N_14004,N_13203,N_13331);
xnor U14005 (N_14005,N_13397,N_13569);
or U14006 (N_14006,N_13184,N_13218);
and U14007 (N_14007,N_13420,N_13579);
or U14008 (N_14008,N_13661,N_13318);
nand U14009 (N_14009,N_13442,N_13226);
nor U14010 (N_14010,N_13615,N_13266);
nand U14011 (N_14011,N_13145,N_13195);
xor U14012 (N_14012,N_13274,N_13312);
and U14013 (N_14013,N_13329,N_13425);
or U14014 (N_14014,N_13322,N_13447);
nor U14015 (N_14015,N_13177,N_13517);
nor U14016 (N_14016,N_13225,N_13622);
nand U14017 (N_14017,N_13617,N_13259);
or U14018 (N_14018,N_13457,N_13746);
nor U14019 (N_14019,N_13677,N_13227);
or U14020 (N_14020,N_13651,N_13481);
xor U14021 (N_14021,N_13220,N_13358);
nor U14022 (N_14022,N_13619,N_13697);
or U14023 (N_14023,N_13451,N_13269);
xor U14024 (N_14024,N_13323,N_13645);
or U14025 (N_14025,N_13393,N_13379);
nor U14026 (N_14026,N_13253,N_13337);
or U14027 (N_14027,N_13356,N_13659);
and U14028 (N_14028,N_13198,N_13160);
and U14029 (N_14029,N_13135,N_13180);
nor U14030 (N_14030,N_13382,N_13254);
xor U14031 (N_14031,N_13263,N_13463);
nand U14032 (N_14032,N_13514,N_13127);
or U14033 (N_14033,N_13527,N_13737);
nor U14034 (N_14034,N_13163,N_13345);
nand U14035 (N_14035,N_13432,N_13309);
and U14036 (N_14036,N_13296,N_13600);
and U14037 (N_14037,N_13576,N_13214);
xor U14038 (N_14038,N_13388,N_13581);
or U14039 (N_14039,N_13338,N_13652);
nand U14040 (N_14040,N_13497,N_13663);
xnor U14041 (N_14041,N_13573,N_13134);
and U14042 (N_14042,N_13668,N_13710);
nand U14043 (N_14043,N_13665,N_13507);
xor U14044 (N_14044,N_13537,N_13300);
xor U14045 (N_14045,N_13408,N_13421);
nor U14046 (N_14046,N_13528,N_13591);
or U14047 (N_14047,N_13273,N_13381);
and U14048 (N_14048,N_13394,N_13707);
xnor U14049 (N_14049,N_13554,N_13605);
and U14050 (N_14050,N_13491,N_13669);
nor U14051 (N_14051,N_13258,N_13538);
nor U14052 (N_14052,N_13427,N_13583);
nor U14053 (N_14053,N_13643,N_13185);
nor U14054 (N_14054,N_13532,N_13294);
xor U14055 (N_14055,N_13542,N_13512);
nand U14056 (N_14056,N_13735,N_13621);
nor U14057 (N_14057,N_13623,N_13272);
or U14058 (N_14058,N_13389,N_13236);
and U14059 (N_14059,N_13217,N_13475);
nor U14060 (N_14060,N_13182,N_13286);
xor U14061 (N_14061,N_13373,N_13407);
or U14062 (N_14062,N_13416,N_13402);
xor U14063 (N_14063,N_13742,N_13593);
or U14064 (N_14064,N_13454,N_13310);
nor U14065 (N_14065,N_13404,N_13250);
nor U14066 (N_14066,N_13579,N_13636);
nor U14067 (N_14067,N_13485,N_13425);
and U14068 (N_14068,N_13173,N_13205);
nand U14069 (N_14069,N_13624,N_13332);
or U14070 (N_14070,N_13653,N_13339);
xor U14071 (N_14071,N_13224,N_13732);
or U14072 (N_14072,N_13438,N_13222);
and U14073 (N_14073,N_13144,N_13669);
and U14074 (N_14074,N_13636,N_13742);
and U14075 (N_14075,N_13209,N_13435);
nor U14076 (N_14076,N_13544,N_13273);
and U14077 (N_14077,N_13303,N_13203);
or U14078 (N_14078,N_13540,N_13550);
xnor U14079 (N_14079,N_13299,N_13640);
or U14080 (N_14080,N_13502,N_13345);
xor U14081 (N_14081,N_13508,N_13293);
xor U14082 (N_14082,N_13553,N_13263);
nand U14083 (N_14083,N_13588,N_13147);
or U14084 (N_14084,N_13431,N_13649);
nor U14085 (N_14085,N_13129,N_13547);
nor U14086 (N_14086,N_13565,N_13748);
or U14087 (N_14087,N_13416,N_13617);
nor U14088 (N_14088,N_13288,N_13160);
and U14089 (N_14089,N_13681,N_13400);
xnor U14090 (N_14090,N_13280,N_13726);
nor U14091 (N_14091,N_13476,N_13310);
nor U14092 (N_14092,N_13456,N_13306);
xor U14093 (N_14093,N_13422,N_13630);
nor U14094 (N_14094,N_13355,N_13326);
nor U14095 (N_14095,N_13188,N_13141);
and U14096 (N_14096,N_13312,N_13401);
xnor U14097 (N_14097,N_13250,N_13247);
or U14098 (N_14098,N_13389,N_13748);
nor U14099 (N_14099,N_13577,N_13663);
nor U14100 (N_14100,N_13446,N_13290);
nor U14101 (N_14101,N_13747,N_13597);
or U14102 (N_14102,N_13429,N_13546);
nand U14103 (N_14103,N_13356,N_13308);
or U14104 (N_14104,N_13154,N_13631);
and U14105 (N_14105,N_13388,N_13342);
nor U14106 (N_14106,N_13497,N_13560);
and U14107 (N_14107,N_13420,N_13246);
and U14108 (N_14108,N_13448,N_13371);
xnor U14109 (N_14109,N_13725,N_13728);
nand U14110 (N_14110,N_13377,N_13384);
xnor U14111 (N_14111,N_13294,N_13507);
nand U14112 (N_14112,N_13626,N_13546);
xor U14113 (N_14113,N_13172,N_13354);
and U14114 (N_14114,N_13744,N_13521);
xnor U14115 (N_14115,N_13683,N_13452);
xor U14116 (N_14116,N_13746,N_13462);
and U14117 (N_14117,N_13602,N_13512);
and U14118 (N_14118,N_13466,N_13150);
xor U14119 (N_14119,N_13445,N_13689);
and U14120 (N_14120,N_13607,N_13521);
nor U14121 (N_14121,N_13138,N_13486);
nand U14122 (N_14122,N_13485,N_13668);
or U14123 (N_14123,N_13553,N_13480);
nor U14124 (N_14124,N_13523,N_13229);
xnor U14125 (N_14125,N_13322,N_13278);
or U14126 (N_14126,N_13403,N_13374);
xor U14127 (N_14127,N_13339,N_13427);
nor U14128 (N_14128,N_13184,N_13506);
xor U14129 (N_14129,N_13167,N_13434);
nor U14130 (N_14130,N_13418,N_13567);
and U14131 (N_14131,N_13231,N_13313);
or U14132 (N_14132,N_13638,N_13374);
nor U14133 (N_14133,N_13281,N_13196);
nand U14134 (N_14134,N_13579,N_13543);
nor U14135 (N_14135,N_13327,N_13331);
xor U14136 (N_14136,N_13703,N_13370);
xnor U14137 (N_14137,N_13322,N_13312);
and U14138 (N_14138,N_13228,N_13222);
nand U14139 (N_14139,N_13375,N_13526);
or U14140 (N_14140,N_13426,N_13252);
nand U14141 (N_14141,N_13635,N_13202);
xnor U14142 (N_14142,N_13283,N_13261);
nor U14143 (N_14143,N_13190,N_13630);
or U14144 (N_14144,N_13225,N_13545);
nand U14145 (N_14145,N_13128,N_13176);
nor U14146 (N_14146,N_13541,N_13289);
xnor U14147 (N_14147,N_13550,N_13392);
xnor U14148 (N_14148,N_13582,N_13217);
xnor U14149 (N_14149,N_13159,N_13187);
nand U14150 (N_14150,N_13445,N_13645);
or U14151 (N_14151,N_13615,N_13258);
nor U14152 (N_14152,N_13485,N_13536);
nor U14153 (N_14153,N_13692,N_13386);
or U14154 (N_14154,N_13475,N_13599);
nand U14155 (N_14155,N_13552,N_13355);
xnor U14156 (N_14156,N_13297,N_13358);
and U14157 (N_14157,N_13639,N_13279);
and U14158 (N_14158,N_13647,N_13275);
nor U14159 (N_14159,N_13643,N_13638);
or U14160 (N_14160,N_13678,N_13148);
xor U14161 (N_14161,N_13515,N_13399);
and U14162 (N_14162,N_13288,N_13211);
xnor U14163 (N_14163,N_13223,N_13477);
nand U14164 (N_14164,N_13267,N_13343);
and U14165 (N_14165,N_13569,N_13460);
or U14166 (N_14166,N_13657,N_13146);
nor U14167 (N_14167,N_13387,N_13178);
and U14168 (N_14168,N_13356,N_13653);
xnor U14169 (N_14169,N_13624,N_13165);
xnor U14170 (N_14170,N_13478,N_13319);
and U14171 (N_14171,N_13236,N_13409);
and U14172 (N_14172,N_13559,N_13276);
and U14173 (N_14173,N_13481,N_13655);
and U14174 (N_14174,N_13426,N_13219);
nand U14175 (N_14175,N_13370,N_13236);
nor U14176 (N_14176,N_13605,N_13188);
and U14177 (N_14177,N_13386,N_13499);
nor U14178 (N_14178,N_13693,N_13199);
xor U14179 (N_14179,N_13488,N_13251);
xnor U14180 (N_14180,N_13248,N_13554);
nand U14181 (N_14181,N_13283,N_13271);
and U14182 (N_14182,N_13260,N_13534);
and U14183 (N_14183,N_13516,N_13640);
and U14184 (N_14184,N_13305,N_13274);
and U14185 (N_14185,N_13540,N_13204);
xor U14186 (N_14186,N_13195,N_13528);
nor U14187 (N_14187,N_13688,N_13503);
and U14188 (N_14188,N_13601,N_13336);
xor U14189 (N_14189,N_13638,N_13637);
xnor U14190 (N_14190,N_13237,N_13424);
nor U14191 (N_14191,N_13469,N_13248);
nand U14192 (N_14192,N_13442,N_13730);
nand U14193 (N_14193,N_13581,N_13589);
nand U14194 (N_14194,N_13248,N_13145);
or U14195 (N_14195,N_13638,N_13214);
and U14196 (N_14196,N_13709,N_13149);
or U14197 (N_14197,N_13228,N_13199);
or U14198 (N_14198,N_13569,N_13635);
or U14199 (N_14199,N_13175,N_13564);
and U14200 (N_14200,N_13385,N_13200);
nor U14201 (N_14201,N_13399,N_13365);
xor U14202 (N_14202,N_13637,N_13651);
xor U14203 (N_14203,N_13725,N_13300);
nand U14204 (N_14204,N_13652,N_13630);
nand U14205 (N_14205,N_13562,N_13427);
or U14206 (N_14206,N_13640,N_13727);
or U14207 (N_14207,N_13544,N_13250);
and U14208 (N_14208,N_13554,N_13256);
xnor U14209 (N_14209,N_13262,N_13257);
nand U14210 (N_14210,N_13542,N_13299);
or U14211 (N_14211,N_13585,N_13614);
or U14212 (N_14212,N_13257,N_13134);
and U14213 (N_14213,N_13281,N_13629);
xnor U14214 (N_14214,N_13521,N_13413);
nor U14215 (N_14215,N_13612,N_13425);
nor U14216 (N_14216,N_13552,N_13187);
or U14217 (N_14217,N_13302,N_13543);
xnor U14218 (N_14218,N_13714,N_13426);
or U14219 (N_14219,N_13259,N_13693);
nand U14220 (N_14220,N_13466,N_13426);
or U14221 (N_14221,N_13679,N_13469);
or U14222 (N_14222,N_13410,N_13688);
or U14223 (N_14223,N_13138,N_13325);
nor U14224 (N_14224,N_13173,N_13253);
and U14225 (N_14225,N_13626,N_13686);
nand U14226 (N_14226,N_13184,N_13294);
xnor U14227 (N_14227,N_13635,N_13309);
nor U14228 (N_14228,N_13658,N_13669);
nor U14229 (N_14229,N_13310,N_13198);
xnor U14230 (N_14230,N_13428,N_13454);
nand U14231 (N_14231,N_13415,N_13537);
and U14232 (N_14232,N_13664,N_13696);
nand U14233 (N_14233,N_13447,N_13705);
and U14234 (N_14234,N_13665,N_13131);
and U14235 (N_14235,N_13279,N_13634);
and U14236 (N_14236,N_13349,N_13719);
and U14237 (N_14237,N_13402,N_13207);
and U14238 (N_14238,N_13390,N_13459);
xnor U14239 (N_14239,N_13370,N_13388);
or U14240 (N_14240,N_13681,N_13240);
nor U14241 (N_14241,N_13431,N_13505);
nand U14242 (N_14242,N_13698,N_13731);
nand U14243 (N_14243,N_13268,N_13663);
and U14244 (N_14244,N_13125,N_13274);
and U14245 (N_14245,N_13457,N_13526);
or U14246 (N_14246,N_13181,N_13460);
or U14247 (N_14247,N_13438,N_13449);
nor U14248 (N_14248,N_13507,N_13572);
xnor U14249 (N_14249,N_13398,N_13746);
nor U14250 (N_14250,N_13316,N_13126);
or U14251 (N_14251,N_13316,N_13239);
nor U14252 (N_14252,N_13493,N_13727);
xor U14253 (N_14253,N_13661,N_13511);
nor U14254 (N_14254,N_13396,N_13491);
xor U14255 (N_14255,N_13676,N_13311);
xnor U14256 (N_14256,N_13618,N_13158);
nand U14257 (N_14257,N_13745,N_13189);
nand U14258 (N_14258,N_13321,N_13507);
xor U14259 (N_14259,N_13383,N_13741);
xnor U14260 (N_14260,N_13348,N_13568);
or U14261 (N_14261,N_13588,N_13638);
nor U14262 (N_14262,N_13291,N_13488);
nor U14263 (N_14263,N_13310,N_13487);
or U14264 (N_14264,N_13729,N_13423);
xnor U14265 (N_14265,N_13166,N_13502);
nor U14266 (N_14266,N_13373,N_13240);
nor U14267 (N_14267,N_13657,N_13288);
nor U14268 (N_14268,N_13306,N_13258);
nor U14269 (N_14269,N_13239,N_13395);
and U14270 (N_14270,N_13442,N_13737);
and U14271 (N_14271,N_13527,N_13634);
nand U14272 (N_14272,N_13637,N_13476);
xor U14273 (N_14273,N_13140,N_13335);
xor U14274 (N_14274,N_13560,N_13584);
and U14275 (N_14275,N_13680,N_13433);
or U14276 (N_14276,N_13402,N_13266);
and U14277 (N_14277,N_13555,N_13215);
and U14278 (N_14278,N_13478,N_13212);
xor U14279 (N_14279,N_13156,N_13464);
nand U14280 (N_14280,N_13671,N_13677);
nand U14281 (N_14281,N_13626,N_13159);
nand U14282 (N_14282,N_13708,N_13471);
xor U14283 (N_14283,N_13254,N_13385);
xor U14284 (N_14284,N_13333,N_13357);
nand U14285 (N_14285,N_13233,N_13634);
or U14286 (N_14286,N_13184,N_13175);
nand U14287 (N_14287,N_13337,N_13561);
nand U14288 (N_14288,N_13436,N_13225);
or U14289 (N_14289,N_13730,N_13487);
nor U14290 (N_14290,N_13623,N_13139);
nor U14291 (N_14291,N_13246,N_13370);
or U14292 (N_14292,N_13555,N_13331);
and U14293 (N_14293,N_13440,N_13666);
nand U14294 (N_14294,N_13269,N_13714);
or U14295 (N_14295,N_13484,N_13450);
nor U14296 (N_14296,N_13467,N_13498);
and U14297 (N_14297,N_13327,N_13328);
nand U14298 (N_14298,N_13552,N_13659);
xor U14299 (N_14299,N_13662,N_13193);
nand U14300 (N_14300,N_13664,N_13648);
or U14301 (N_14301,N_13232,N_13401);
xor U14302 (N_14302,N_13611,N_13326);
nor U14303 (N_14303,N_13439,N_13624);
and U14304 (N_14304,N_13511,N_13204);
and U14305 (N_14305,N_13474,N_13277);
nand U14306 (N_14306,N_13543,N_13611);
xor U14307 (N_14307,N_13619,N_13689);
and U14308 (N_14308,N_13352,N_13695);
and U14309 (N_14309,N_13508,N_13231);
or U14310 (N_14310,N_13138,N_13131);
and U14311 (N_14311,N_13724,N_13494);
or U14312 (N_14312,N_13258,N_13442);
nor U14313 (N_14313,N_13738,N_13237);
or U14314 (N_14314,N_13478,N_13150);
and U14315 (N_14315,N_13228,N_13593);
nand U14316 (N_14316,N_13165,N_13607);
nand U14317 (N_14317,N_13318,N_13539);
xnor U14318 (N_14318,N_13272,N_13180);
xor U14319 (N_14319,N_13294,N_13432);
and U14320 (N_14320,N_13646,N_13685);
and U14321 (N_14321,N_13597,N_13445);
nand U14322 (N_14322,N_13272,N_13389);
xnor U14323 (N_14323,N_13683,N_13238);
and U14324 (N_14324,N_13173,N_13501);
nor U14325 (N_14325,N_13374,N_13652);
or U14326 (N_14326,N_13525,N_13476);
nor U14327 (N_14327,N_13332,N_13482);
nor U14328 (N_14328,N_13499,N_13366);
xnor U14329 (N_14329,N_13491,N_13661);
nor U14330 (N_14330,N_13339,N_13476);
and U14331 (N_14331,N_13561,N_13502);
nor U14332 (N_14332,N_13453,N_13693);
nor U14333 (N_14333,N_13449,N_13250);
nor U14334 (N_14334,N_13480,N_13381);
nor U14335 (N_14335,N_13589,N_13604);
xnor U14336 (N_14336,N_13431,N_13656);
and U14337 (N_14337,N_13330,N_13333);
or U14338 (N_14338,N_13299,N_13209);
xor U14339 (N_14339,N_13632,N_13128);
xor U14340 (N_14340,N_13440,N_13276);
or U14341 (N_14341,N_13185,N_13679);
or U14342 (N_14342,N_13404,N_13397);
nor U14343 (N_14343,N_13396,N_13327);
nand U14344 (N_14344,N_13377,N_13467);
nor U14345 (N_14345,N_13720,N_13376);
nand U14346 (N_14346,N_13694,N_13740);
and U14347 (N_14347,N_13572,N_13147);
xor U14348 (N_14348,N_13586,N_13681);
nand U14349 (N_14349,N_13265,N_13564);
nand U14350 (N_14350,N_13206,N_13547);
nor U14351 (N_14351,N_13191,N_13127);
xnor U14352 (N_14352,N_13261,N_13394);
or U14353 (N_14353,N_13658,N_13589);
nor U14354 (N_14354,N_13351,N_13317);
xor U14355 (N_14355,N_13431,N_13205);
or U14356 (N_14356,N_13388,N_13730);
xor U14357 (N_14357,N_13524,N_13238);
and U14358 (N_14358,N_13324,N_13208);
nand U14359 (N_14359,N_13225,N_13446);
nand U14360 (N_14360,N_13194,N_13640);
xor U14361 (N_14361,N_13269,N_13488);
nand U14362 (N_14362,N_13733,N_13681);
xnor U14363 (N_14363,N_13200,N_13609);
xor U14364 (N_14364,N_13629,N_13676);
and U14365 (N_14365,N_13424,N_13377);
or U14366 (N_14366,N_13278,N_13466);
or U14367 (N_14367,N_13422,N_13367);
xor U14368 (N_14368,N_13365,N_13191);
or U14369 (N_14369,N_13302,N_13349);
nand U14370 (N_14370,N_13670,N_13148);
nand U14371 (N_14371,N_13198,N_13469);
xor U14372 (N_14372,N_13581,N_13579);
and U14373 (N_14373,N_13238,N_13652);
nor U14374 (N_14374,N_13706,N_13389);
nor U14375 (N_14375,N_14070,N_14218);
xnor U14376 (N_14376,N_14098,N_13876);
xor U14377 (N_14377,N_14261,N_13814);
nand U14378 (N_14378,N_14367,N_14049);
or U14379 (N_14379,N_14300,N_14271);
or U14380 (N_14380,N_14132,N_13922);
or U14381 (N_14381,N_14291,N_14019);
and U14382 (N_14382,N_14133,N_14059);
nand U14383 (N_14383,N_13819,N_14328);
nand U14384 (N_14384,N_13896,N_14112);
and U14385 (N_14385,N_13797,N_13979);
nor U14386 (N_14386,N_14015,N_14018);
nand U14387 (N_14387,N_13902,N_14129);
or U14388 (N_14388,N_13769,N_14124);
xnor U14389 (N_14389,N_13994,N_13998);
xor U14390 (N_14390,N_14348,N_14313);
nand U14391 (N_14391,N_13976,N_14101);
or U14392 (N_14392,N_13755,N_13838);
nand U14393 (N_14393,N_14258,N_13907);
or U14394 (N_14394,N_13832,N_14270);
nor U14395 (N_14395,N_14297,N_14268);
nor U14396 (N_14396,N_13798,N_14180);
xnor U14397 (N_14397,N_13912,N_13826);
xor U14398 (N_14398,N_14182,N_14312);
nand U14399 (N_14399,N_13843,N_13770);
nand U14400 (N_14400,N_14050,N_14311);
nor U14401 (N_14401,N_13951,N_14203);
and U14402 (N_14402,N_13947,N_14318);
or U14403 (N_14403,N_13981,N_14316);
or U14404 (N_14404,N_14024,N_14248);
nor U14405 (N_14405,N_13844,N_14212);
xor U14406 (N_14406,N_14274,N_14037);
nand U14407 (N_14407,N_13815,N_14083);
xor U14408 (N_14408,N_14041,N_13888);
xor U14409 (N_14409,N_14062,N_13925);
xnor U14410 (N_14410,N_14090,N_13799);
nand U14411 (N_14411,N_13975,N_14119);
or U14412 (N_14412,N_14205,N_13884);
or U14413 (N_14413,N_14331,N_13861);
nor U14414 (N_14414,N_14255,N_14321);
and U14415 (N_14415,N_14094,N_13965);
nand U14416 (N_14416,N_14165,N_14307);
xnor U14417 (N_14417,N_14071,N_13862);
nor U14418 (N_14418,N_13791,N_14040);
and U14419 (N_14419,N_13850,N_13767);
nor U14420 (N_14420,N_13878,N_14078);
nand U14421 (N_14421,N_14104,N_14232);
xor U14422 (N_14422,N_14371,N_13978);
xnor U14423 (N_14423,N_14108,N_14156);
nand U14424 (N_14424,N_14202,N_13885);
and U14425 (N_14425,N_13822,N_13802);
nand U14426 (N_14426,N_14245,N_14235);
or U14427 (N_14427,N_14336,N_13758);
or U14428 (N_14428,N_14320,N_14206);
and U14429 (N_14429,N_14079,N_14177);
and U14430 (N_14430,N_14053,N_13857);
nor U14431 (N_14431,N_13833,N_14365);
nand U14432 (N_14432,N_14069,N_14178);
nor U14433 (N_14433,N_14077,N_14369);
and U14434 (N_14434,N_13946,N_13751);
and U14435 (N_14435,N_13794,N_14135);
nor U14436 (N_14436,N_13910,N_13768);
and U14437 (N_14437,N_13916,N_14020);
xor U14438 (N_14438,N_14342,N_14089);
and U14439 (N_14439,N_13904,N_14179);
nand U14440 (N_14440,N_14052,N_13996);
nor U14441 (N_14441,N_14087,N_13971);
and U14442 (N_14442,N_14225,N_14175);
nand U14443 (N_14443,N_13764,N_13892);
and U14444 (N_14444,N_13901,N_14047);
xnor U14445 (N_14445,N_13988,N_13874);
and U14446 (N_14446,N_13972,N_14334);
and U14447 (N_14447,N_13897,N_14257);
or U14448 (N_14448,N_14027,N_14106);
nor U14449 (N_14449,N_13911,N_13795);
xor U14450 (N_14450,N_14344,N_14296);
and U14451 (N_14451,N_13913,N_14359);
xor U14452 (N_14452,N_13997,N_13865);
and U14453 (N_14453,N_14193,N_14264);
xor U14454 (N_14454,N_14262,N_14332);
nand U14455 (N_14455,N_14249,N_14215);
nand U14456 (N_14456,N_14084,N_14373);
and U14457 (N_14457,N_14231,N_13957);
nand U14458 (N_14458,N_14242,N_13944);
nand U14459 (N_14459,N_14322,N_13811);
xnor U14460 (N_14460,N_14091,N_13835);
nand U14461 (N_14461,N_14067,N_14029);
and U14462 (N_14462,N_13959,N_14191);
and U14463 (N_14463,N_13984,N_13955);
xor U14464 (N_14464,N_14109,N_14176);
nand U14465 (N_14465,N_13923,N_13869);
xnor U14466 (N_14466,N_14014,N_13895);
xor U14467 (N_14467,N_13806,N_13827);
nand U14468 (N_14468,N_13929,N_14207);
nor U14469 (N_14469,N_13800,N_14240);
nand U14470 (N_14470,N_13858,N_14081);
nor U14471 (N_14471,N_14286,N_13841);
and U14472 (N_14472,N_13881,N_14173);
xor U14473 (N_14473,N_14181,N_14276);
and U14474 (N_14474,N_13870,N_14374);
nor U14475 (N_14475,N_14317,N_13785);
nand U14476 (N_14476,N_14337,N_13950);
nand U14477 (N_14477,N_14073,N_13966);
nand U14478 (N_14478,N_13898,N_13777);
nand U14479 (N_14479,N_13790,N_14120);
or U14480 (N_14480,N_14326,N_14309);
xor U14481 (N_14481,N_13808,N_13813);
nor U14482 (N_14482,N_14057,N_14241);
nand U14483 (N_14483,N_13852,N_14126);
or U14484 (N_14484,N_14278,N_14222);
or U14485 (N_14485,N_14021,N_14004);
nor U14486 (N_14486,N_13879,N_13940);
xor U14487 (N_14487,N_14330,N_13756);
or U14488 (N_14488,N_13831,N_14056);
or U14489 (N_14489,N_14158,N_14054);
and U14490 (N_14490,N_14030,N_13872);
or U14491 (N_14491,N_13866,N_13812);
and U14492 (N_14492,N_13757,N_13967);
nor U14493 (N_14493,N_14153,N_13823);
nor U14494 (N_14494,N_14017,N_14190);
or U14495 (N_14495,N_13809,N_13918);
or U14496 (N_14496,N_13779,N_14008);
nand U14497 (N_14497,N_14033,N_13945);
and U14498 (N_14498,N_14325,N_13842);
xor U14499 (N_14499,N_14290,N_13886);
and U14500 (N_14500,N_13942,N_14256);
nor U14501 (N_14501,N_14155,N_14259);
xor U14502 (N_14502,N_14095,N_14238);
nand U14503 (N_14503,N_14226,N_14055);
nand U14504 (N_14504,N_13864,N_14234);
and U14505 (N_14505,N_13938,N_13949);
nor U14506 (N_14506,N_13825,N_14251);
nand U14507 (N_14507,N_14269,N_14304);
nor U14508 (N_14508,N_14145,N_14099);
nor U14509 (N_14509,N_13840,N_14282);
xor U14510 (N_14510,N_13848,N_14142);
nand U14511 (N_14511,N_14186,N_14368);
and U14512 (N_14512,N_13860,N_13933);
and U14513 (N_14513,N_14005,N_13820);
nand U14514 (N_14514,N_13789,N_13854);
and U14515 (N_14515,N_14210,N_13889);
and U14516 (N_14516,N_13915,N_14370);
nand U14517 (N_14517,N_14157,N_14093);
nor U14518 (N_14518,N_14034,N_14149);
nand U14519 (N_14519,N_14340,N_13863);
nand U14520 (N_14520,N_13932,N_13778);
nand U14521 (N_14521,N_13867,N_14366);
and U14522 (N_14522,N_14338,N_14134);
or U14523 (N_14523,N_14220,N_14166);
or U14524 (N_14524,N_13919,N_14272);
or U14525 (N_14525,N_14045,N_14195);
nand U14526 (N_14526,N_14148,N_14111);
or U14527 (N_14527,N_13908,N_14250);
or U14528 (N_14528,N_14329,N_13900);
and U14529 (N_14529,N_14323,N_13807);
nor U14530 (N_14530,N_14364,N_14150);
nand U14531 (N_14531,N_13982,N_14183);
or U14532 (N_14532,N_13927,N_13928);
or U14533 (N_14533,N_14011,N_14038);
nand U14534 (N_14534,N_13759,N_13829);
nand U14535 (N_14535,N_14013,N_13763);
nor U14536 (N_14536,N_13987,N_14154);
and U14537 (N_14537,N_13917,N_14009);
and U14538 (N_14538,N_13761,N_14168);
nor U14539 (N_14539,N_13969,N_14061);
and U14540 (N_14540,N_14032,N_14324);
nand U14541 (N_14541,N_14299,N_14185);
or U14542 (N_14542,N_13845,N_14287);
or U14543 (N_14543,N_14302,N_13871);
and U14544 (N_14544,N_13891,N_13782);
or U14545 (N_14545,N_14341,N_14136);
and U14546 (N_14546,N_14113,N_14333);
nand U14547 (N_14547,N_14284,N_13973);
nand U14548 (N_14548,N_13937,N_14080);
and U14549 (N_14549,N_14114,N_14260);
xnor U14550 (N_14550,N_13853,N_14354);
xnor U14551 (N_14551,N_14065,N_14006);
nor U14552 (N_14552,N_14201,N_14327);
xnor U14553 (N_14553,N_14343,N_14265);
nor U14554 (N_14554,N_13754,N_14243);
xnor U14555 (N_14555,N_13766,N_13752);
and U14556 (N_14556,N_14066,N_13905);
or U14557 (N_14557,N_13855,N_14167);
xor U14558 (N_14558,N_14164,N_14163);
or U14559 (N_14559,N_14319,N_14228);
nor U14560 (N_14560,N_14127,N_14116);
nor U14561 (N_14561,N_13941,N_14360);
nor U14562 (N_14562,N_14012,N_13921);
and U14563 (N_14563,N_13953,N_14229);
xor U14564 (N_14564,N_13849,N_14289);
or U14565 (N_14565,N_14003,N_13803);
xor U14566 (N_14566,N_14292,N_14310);
nor U14567 (N_14567,N_13804,N_13788);
nand U14568 (N_14568,N_13989,N_13793);
xnor U14569 (N_14569,N_14253,N_14362);
or U14570 (N_14570,N_14097,N_14169);
or U14571 (N_14571,N_13780,N_13903);
and U14572 (N_14572,N_14345,N_14144);
and U14573 (N_14573,N_14188,N_14211);
nand U14574 (N_14574,N_13883,N_13762);
nor U14575 (N_14575,N_13890,N_14121);
nand U14576 (N_14576,N_13771,N_14075);
or U14577 (N_14577,N_14192,N_13784);
nor U14578 (N_14578,N_14146,N_14170);
and U14579 (N_14579,N_14039,N_14131);
xor U14580 (N_14580,N_13880,N_14224);
or U14581 (N_14581,N_14267,N_14352);
nor U14582 (N_14582,N_14102,N_14246);
and U14583 (N_14583,N_14074,N_14244);
or U14584 (N_14584,N_14349,N_14277);
or U14585 (N_14585,N_14221,N_14068);
nor U14586 (N_14586,N_13774,N_14092);
nand U14587 (N_14587,N_14285,N_14028);
or U14588 (N_14588,N_13924,N_13805);
or U14589 (N_14589,N_13961,N_14187);
nor U14590 (N_14590,N_14025,N_13801);
nand U14591 (N_14591,N_14130,N_14266);
or U14592 (N_14592,N_14350,N_14043);
and U14593 (N_14593,N_13836,N_13796);
nor U14594 (N_14594,N_14288,N_13992);
nand U14595 (N_14595,N_13772,N_13824);
nor U14596 (N_14596,N_14358,N_14036);
xnor U14597 (N_14597,N_14044,N_13851);
nand U14598 (N_14598,N_13760,N_13810);
or U14599 (N_14599,N_13783,N_13958);
xor U14600 (N_14600,N_14230,N_14273);
nand U14601 (N_14601,N_14247,N_13765);
and U14602 (N_14602,N_13977,N_13830);
nor U14603 (N_14603,N_13964,N_14058);
nor U14604 (N_14604,N_13963,N_14162);
nor U14605 (N_14605,N_14236,N_14347);
and U14606 (N_14606,N_14306,N_14356);
nor U14607 (N_14607,N_14016,N_14189);
nor U14608 (N_14608,N_14060,N_14363);
nand U14609 (N_14609,N_14122,N_14216);
xor U14610 (N_14610,N_14022,N_14063);
xor U14611 (N_14611,N_14196,N_13974);
and U14612 (N_14612,N_13909,N_14239);
xnor U14613 (N_14613,N_14096,N_13991);
or U14614 (N_14614,N_14147,N_13873);
nand U14615 (N_14615,N_13882,N_14076);
nor U14616 (N_14616,N_14308,N_14140);
xor U14617 (N_14617,N_13906,N_14048);
xnor U14618 (N_14618,N_14141,N_14031);
and U14619 (N_14619,N_13930,N_14283);
xnor U14620 (N_14620,N_13834,N_14293);
nand U14621 (N_14621,N_14233,N_13821);
xor U14622 (N_14622,N_13773,N_14357);
nand U14623 (N_14623,N_14125,N_14082);
nor U14624 (N_14624,N_14252,N_14000);
nor U14625 (N_14625,N_14294,N_13936);
nor U14626 (N_14626,N_14263,N_14115);
nor U14627 (N_14627,N_13934,N_14128);
or U14628 (N_14628,N_13948,N_13750);
nor U14629 (N_14629,N_13931,N_13775);
nand U14630 (N_14630,N_14281,N_14198);
or U14631 (N_14631,N_14010,N_14118);
nand U14632 (N_14632,N_14305,N_13970);
nand U14633 (N_14633,N_14171,N_14105);
xor U14634 (N_14634,N_13786,N_13893);
xor U14635 (N_14635,N_13914,N_14139);
nor U14636 (N_14636,N_14361,N_13776);
nor U14637 (N_14637,N_14100,N_13939);
nand U14638 (N_14638,N_14023,N_14197);
xor U14639 (N_14639,N_14103,N_13995);
nor U14640 (N_14640,N_13956,N_14174);
nor U14641 (N_14641,N_13943,N_14117);
xnor U14642 (N_14642,N_14301,N_14279);
xor U14643 (N_14643,N_13792,N_13868);
nand U14644 (N_14644,N_14208,N_13920);
nand U14645 (N_14645,N_13935,N_14143);
or U14646 (N_14646,N_14209,N_13875);
nor U14647 (N_14647,N_13816,N_13968);
nand U14648 (N_14648,N_14372,N_14351);
xnor U14649 (N_14649,N_14007,N_13990);
or U14650 (N_14650,N_13817,N_13846);
xor U14651 (N_14651,N_14064,N_14217);
xor U14652 (N_14652,N_14295,N_14072);
nand U14653 (N_14653,N_14219,N_13887);
xor U14654 (N_14654,N_13962,N_14172);
and U14655 (N_14655,N_14137,N_13985);
nor U14656 (N_14656,N_14086,N_14314);
nor U14657 (N_14657,N_14152,N_13952);
nand U14658 (N_14658,N_14275,N_14339);
nand U14659 (N_14659,N_14051,N_13999);
and U14660 (N_14660,N_13986,N_13818);
xor U14661 (N_14661,N_14298,N_13787);
nor U14662 (N_14662,N_14194,N_14160);
and U14663 (N_14663,N_14088,N_14001);
and U14664 (N_14664,N_14200,N_13753);
and U14665 (N_14665,N_14085,N_13983);
nor U14666 (N_14666,N_13839,N_13993);
nor U14667 (N_14667,N_14254,N_14213);
nor U14668 (N_14668,N_14107,N_14280);
xnor U14669 (N_14669,N_13781,N_14046);
and U14670 (N_14670,N_13828,N_14042);
or U14671 (N_14671,N_14227,N_13954);
xor U14672 (N_14672,N_14159,N_13859);
nand U14673 (N_14673,N_13894,N_14151);
nand U14674 (N_14674,N_13856,N_14315);
and U14675 (N_14675,N_14161,N_14204);
xor U14676 (N_14676,N_14335,N_14199);
and U14677 (N_14677,N_13899,N_14138);
nand U14678 (N_14678,N_13980,N_14353);
xnor U14679 (N_14679,N_14110,N_14002);
nor U14680 (N_14680,N_14184,N_14026);
and U14681 (N_14681,N_13877,N_13837);
nor U14682 (N_14682,N_14303,N_14223);
or U14683 (N_14683,N_14346,N_14237);
nor U14684 (N_14684,N_14355,N_14035);
nand U14685 (N_14685,N_14123,N_13960);
nand U14686 (N_14686,N_13847,N_14214);
nand U14687 (N_14687,N_13926,N_14174);
nand U14688 (N_14688,N_13924,N_14181);
nor U14689 (N_14689,N_13946,N_14248);
xor U14690 (N_14690,N_13753,N_14312);
or U14691 (N_14691,N_13851,N_13859);
and U14692 (N_14692,N_14332,N_13985);
and U14693 (N_14693,N_13928,N_14005);
and U14694 (N_14694,N_13850,N_14284);
nand U14695 (N_14695,N_13898,N_14022);
nand U14696 (N_14696,N_13996,N_14300);
xnor U14697 (N_14697,N_14285,N_14083);
xor U14698 (N_14698,N_14166,N_13769);
and U14699 (N_14699,N_13844,N_14138);
nand U14700 (N_14700,N_14341,N_14225);
nor U14701 (N_14701,N_13846,N_14081);
nand U14702 (N_14702,N_14060,N_13955);
xor U14703 (N_14703,N_13763,N_14021);
xnor U14704 (N_14704,N_14347,N_13807);
and U14705 (N_14705,N_14160,N_13832);
nor U14706 (N_14706,N_13793,N_13834);
and U14707 (N_14707,N_14250,N_14199);
and U14708 (N_14708,N_13762,N_14162);
nor U14709 (N_14709,N_13851,N_14215);
nor U14710 (N_14710,N_14050,N_13782);
nor U14711 (N_14711,N_13761,N_13868);
and U14712 (N_14712,N_14163,N_13878);
or U14713 (N_14713,N_13899,N_14282);
nand U14714 (N_14714,N_14068,N_14004);
or U14715 (N_14715,N_14366,N_13826);
and U14716 (N_14716,N_14216,N_14324);
xor U14717 (N_14717,N_13856,N_13787);
and U14718 (N_14718,N_14357,N_13922);
xor U14719 (N_14719,N_13953,N_14073);
nand U14720 (N_14720,N_14298,N_14248);
nor U14721 (N_14721,N_14244,N_13962);
and U14722 (N_14722,N_13876,N_14142);
nand U14723 (N_14723,N_14352,N_13885);
nor U14724 (N_14724,N_14054,N_14097);
or U14725 (N_14725,N_13875,N_14148);
or U14726 (N_14726,N_13932,N_13948);
or U14727 (N_14727,N_13965,N_14061);
or U14728 (N_14728,N_13828,N_14067);
and U14729 (N_14729,N_14193,N_13858);
and U14730 (N_14730,N_14267,N_13964);
xor U14731 (N_14731,N_13803,N_14372);
and U14732 (N_14732,N_13832,N_14317);
nor U14733 (N_14733,N_14034,N_13836);
xnor U14734 (N_14734,N_13859,N_13960);
nor U14735 (N_14735,N_14180,N_14072);
nand U14736 (N_14736,N_14237,N_14103);
xnor U14737 (N_14737,N_14327,N_14158);
nand U14738 (N_14738,N_13834,N_14286);
nand U14739 (N_14739,N_14259,N_13851);
or U14740 (N_14740,N_14337,N_14364);
and U14741 (N_14741,N_14168,N_14303);
nor U14742 (N_14742,N_14069,N_14201);
xnor U14743 (N_14743,N_14194,N_14307);
and U14744 (N_14744,N_14079,N_14020);
xor U14745 (N_14745,N_14363,N_14318);
or U14746 (N_14746,N_14104,N_13881);
and U14747 (N_14747,N_13873,N_14341);
or U14748 (N_14748,N_14363,N_14186);
and U14749 (N_14749,N_14360,N_13770);
or U14750 (N_14750,N_14261,N_14279);
nor U14751 (N_14751,N_14322,N_13867);
or U14752 (N_14752,N_14275,N_14017);
or U14753 (N_14753,N_14153,N_14223);
xor U14754 (N_14754,N_14242,N_14337);
and U14755 (N_14755,N_14036,N_14066);
nand U14756 (N_14756,N_13783,N_14329);
or U14757 (N_14757,N_14235,N_13874);
nand U14758 (N_14758,N_14199,N_13946);
and U14759 (N_14759,N_13870,N_14365);
nand U14760 (N_14760,N_14307,N_14002);
and U14761 (N_14761,N_13868,N_14178);
xor U14762 (N_14762,N_14131,N_14213);
xnor U14763 (N_14763,N_14198,N_13763);
or U14764 (N_14764,N_13994,N_14187);
and U14765 (N_14765,N_14113,N_14215);
or U14766 (N_14766,N_14305,N_14286);
nor U14767 (N_14767,N_14078,N_14270);
or U14768 (N_14768,N_14135,N_14040);
xnor U14769 (N_14769,N_14042,N_14170);
and U14770 (N_14770,N_14246,N_13929);
and U14771 (N_14771,N_13820,N_14361);
xor U14772 (N_14772,N_14287,N_13902);
nand U14773 (N_14773,N_14086,N_13815);
and U14774 (N_14774,N_14069,N_14145);
and U14775 (N_14775,N_14231,N_14317);
xnor U14776 (N_14776,N_14348,N_13804);
and U14777 (N_14777,N_13872,N_14212);
or U14778 (N_14778,N_13802,N_13859);
or U14779 (N_14779,N_13822,N_14268);
nand U14780 (N_14780,N_14248,N_13862);
or U14781 (N_14781,N_14039,N_13889);
nor U14782 (N_14782,N_14277,N_14170);
xnor U14783 (N_14783,N_14201,N_13889);
xnor U14784 (N_14784,N_14036,N_13836);
xnor U14785 (N_14785,N_13860,N_14179);
and U14786 (N_14786,N_13854,N_14180);
and U14787 (N_14787,N_14015,N_13905);
and U14788 (N_14788,N_14323,N_14103);
or U14789 (N_14789,N_13943,N_14341);
and U14790 (N_14790,N_13933,N_14253);
nand U14791 (N_14791,N_14326,N_13764);
and U14792 (N_14792,N_14157,N_13781);
nand U14793 (N_14793,N_14066,N_14114);
xnor U14794 (N_14794,N_13786,N_14330);
xnor U14795 (N_14795,N_14225,N_13751);
or U14796 (N_14796,N_13780,N_14076);
nor U14797 (N_14797,N_14152,N_13943);
and U14798 (N_14798,N_14354,N_14257);
nand U14799 (N_14799,N_14314,N_14345);
xnor U14800 (N_14800,N_14103,N_13832);
nand U14801 (N_14801,N_13943,N_14136);
nand U14802 (N_14802,N_14262,N_14038);
xnor U14803 (N_14803,N_13866,N_14313);
xor U14804 (N_14804,N_13807,N_14311);
nor U14805 (N_14805,N_14050,N_13914);
nor U14806 (N_14806,N_13843,N_13959);
xor U14807 (N_14807,N_13780,N_13806);
or U14808 (N_14808,N_14325,N_14361);
or U14809 (N_14809,N_13985,N_13770);
and U14810 (N_14810,N_14342,N_14152);
and U14811 (N_14811,N_14052,N_14233);
nand U14812 (N_14812,N_13882,N_13978);
or U14813 (N_14813,N_14141,N_14202);
nand U14814 (N_14814,N_14119,N_13973);
xnor U14815 (N_14815,N_14259,N_13764);
nand U14816 (N_14816,N_13995,N_14248);
or U14817 (N_14817,N_13800,N_14252);
nand U14818 (N_14818,N_14091,N_14122);
or U14819 (N_14819,N_14051,N_14230);
nand U14820 (N_14820,N_14046,N_14116);
and U14821 (N_14821,N_13757,N_13793);
nor U14822 (N_14822,N_14311,N_14058);
or U14823 (N_14823,N_14130,N_13939);
and U14824 (N_14824,N_13994,N_14125);
nor U14825 (N_14825,N_14046,N_14025);
nor U14826 (N_14826,N_14098,N_14170);
or U14827 (N_14827,N_14079,N_14082);
nor U14828 (N_14828,N_13949,N_14203);
xor U14829 (N_14829,N_13797,N_14351);
nand U14830 (N_14830,N_14013,N_13883);
and U14831 (N_14831,N_13835,N_13942);
or U14832 (N_14832,N_14146,N_14126);
xor U14833 (N_14833,N_14194,N_13872);
nand U14834 (N_14834,N_13874,N_14090);
xnor U14835 (N_14835,N_14332,N_14009);
nor U14836 (N_14836,N_14040,N_13773);
and U14837 (N_14837,N_14038,N_13994);
and U14838 (N_14838,N_14048,N_14190);
nand U14839 (N_14839,N_14068,N_14178);
nand U14840 (N_14840,N_13915,N_14256);
or U14841 (N_14841,N_14258,N_14129);
or U14842 (N_14842,N_13823,N_14079);
nor U14843 (N_14843,N_14134,N_13796);
and U14844 (N_14844,N_13871,N_14053);
xor U14845 (N_14845,N_13908,N_13947);
and U14846 (N_14846,N_14109,N_13926);
and U14847 (N_14847,N_13950,N_13844);
nor U14848 (N_14848,N_13988,N_14042);
nor U14849 (N_14849,N_14072,N_13794);
and U14850 (N_14850,N_14209,N_13835);
or U14851 (N_14851,N_14001,N_14269);
and U14852 (N_14852,N_13941,N_14330);
nand U14853 (N_14853,N_14212,N_13993);
xnor U14854 (N_14854,N_14325,N_13814);
nand U14855 (N_14855,N_14094,N_13885);
or U14856 (N_14856,N_14041,N_14294);
xnor U14857 (N_14857,N_13977,N_14021);
xor U14858 (N_14858,N_14099,N_13826);
xnor U14859 (N_14859,N_13778,N_14126);
nor U14860 (N_14860,N_13801,N_14225);
or U14861 (N_14861,N_14050,N_13936);
xnor U14862 (N_14862,N_14163,N_14279);
nor U14863 (N_14863,N_13905,N_14334);
or U14864 (N_14864,N_13906,N_14135);
nor U14865 (N_14865,N_14316,N_13861);
nor U14866 (N_14866,N_13993,N_14369);
xor U14867 (N_14867,N_14249,N_13815);
xor U14868 (N_14868,N_14094,N_13903);
xor U14869 (N_14869,N_13788,N_13817);
nand U14870 (N_14870,N_14311,N_14299);
and U14871 (N_14871,N_13990,N_13776);
or U14872 (N_14872,N_14333,N_14188);
xnor U14873 (N_14873,N_13870,N_13858);
xnor U14874 (N_14874,N_14092,N_14077);
or U14875 (N_14875,N_13936,N_14005);
xnor U14876 (N_14876,N_14165,N_13909);
and U14877 (N_14877,N_13970,N_14072);
and U14878 (N_14878,N_13849,N_14297);
or U14879 (N_14879,N_14364,N_13761);
and U14880 (N_14880,N_13949,N_13981);
nor U14881 (N_14881,N_14325,N_14210);
nor U14882 (N_14882,N_13774,N_14134);
nand U14883 (N_14883,N_13876,N_14044);
xnor U14884 (N_14884,N_14021,N_14189);
xnor U14885 (N_14885,N_13863,N_14136);
nand U14886 (N_14886,N_14224,N_14131);
nand U14887 (N_14887,N_13920,N_14033);
or U14888 (N_14888,N_14248,N_13823);
nand U14889 (N_14889,N_14358,N_14360);
nor U14890 (N_14890,N_13768,N_13946);
or U14891 (N_14891,N_14075,N_14035);
nand U14892 (N_14892,N_14292,N_14236);
xor U14893 (N_14893,N_14020,N_13912);
nand U14894 (N_14894,N_13789,N_14181);
nand U14895 (N_14895,N_13774,N_14348);
nand U14896 (N_14896,N_14216,N_14322);
nand U14897 (N_14897,N_13916,N_14030);
xnor U14898 (N_14898,N_13797,N_13891);
nor U14899 (N_14899,N_14231,N_13939);
nand U14900 (N_14900,N_14073,N_14287);
and U14901 (N_14901,N_13906,N_13880);
nand U14902 (N_14902,N_14257,N_13839);
xnor U14903 (N_14903,N_14275,N_14310);
and U14904 (N_14904,N_13800,N_13793);
and U14905 (N_14905,N_13962,N_13862);
and U14906 (N_14906,N_14211,N_14041);
xnor U14907 (N_14907,N_14256,N_14296);
xnor U14908 (N_14908,N_13907,N_14129);
and U14909 (N_14909,N_13923,N_13760);
nor U14910 (N_14910,N_14202,N_13907);
and U14911 (N_14911,N_13895,N_14065);
nand U14912 (N_14912,N_13832,N_14253);
nand U14913 (N_14913,N_14374,N_14268);
nor U14914 (N_14914,N_13884,N_14149);
or U14915 (N_14915,N_14051,N_14358);
and U14916 (N_14916,N_13877,N_13846);
xor U14917 (N_14917,N_13810,N_14110);
xnor U14918 (N_14918,N_14246,N_14079);
xor U14919 (N_14919,N_13781,N_14227);
xnor U14920 (N_14920,N_13835,N_14196);
nor U14921 (N_14921,N_14181,N_14080);
or U14922 (N_14922,N_14172,N_14297);
nand U14923 (N_14923,N_14146,N_13772);
nor U14924 (N_14924,N_13777,N_14061);
and U14925 (N_14925,N_14108,N_14107);
or U14926 (N_14926,N_14252,N_14353);
xor U14927 (N_14927,N_14246,N_14289);
nor U14928 (N_14928,N_14042,N_13905);
nand U14929 (N_14929,N_14248,N_14143);
and U14930 (N_14930,N_13963,N_14357);
nand U14931 (N_14931,N_13976,N_14288);
and U14932 (N_14932,N_14363,N_14309);
and U14933 (N_14933,N_14186,N_13764);
and U14934 (N_14934,N_13886,N_14151);
and U14935 (N_14935,N_14233,N_14024);
nand U14936 (N_14936,N_14182,N_14243);
xnor U14937 (N_14937,N_14177,N_14274);
xor U14938 (N_14938,N_13806,N_13864);
nor U14939 (N_14939,N_13844,N_13845);
nor U14940 (N_14940,N_13922,N_14002);
and U14941 (N_14941,N_13952,N_14136);
and U14942 (N_14942,N_14244,N_14191);
nor U14943 (N_14943,N_14025,N_14290);
nor U14944 (N_14944,N_14203,N_14332);
or U14945 (N_14945,N_14075,N_13978);
xnor U14946 (N_14946,N_13765,N_14042);
nand U14947 (N_14947,N_14052,N_14308);
and U14948 (N_14948,N_13804,N_14191);
xor U14949 (N_14949,N_13911,N_14145);
xor U14950 (N_14950,N_13763,N_14073);
nor U14951 (N_14951,N_13877,N_13792);
nor U14952 (N_14952,N_14076,N_14016);
xor U14953 (N_14953,N_14150,N_13909);
nand U14954 (N_14954,N_14063,N_13933);
or U14955 (N_14955,N_14055,N_14040);
nor U14956 (N_14956,N_13906,N_13883);
or U14957 (N_14957,N_13832,N_14178);
and U14958 (N_14958,N_14210,N_14009);
nor U14959 (N_14959,N_13806,N_13829);
xnor U14960 (N_14960,N_14061,N_14306);
and U14961 (N_14961,N_14303,N_14171);
xor U14962 (N_14962,N_14193,N_14265);
xor U14963 (N_14963,N_13913,N_14321);
nor U14964 (N_14964,N_14082,N_14039);
nor U14965 (N_14965,N_13936,N_14264);
nor U14966 (N_14966,N_14229,N_14151);
nor U14967 (N_14967,N_14202,N_14230);
nor U14968 (N_14968,N_14068,N_14065);
xor U14969 (N_14969,N_14066,N_14336);
nand U14970 (N_14970,N_14288,N_14245);
nor U14971 (N_14971,N_13756,N_13999);
xor U14972 (N_14972,N_14115,N_13920);
and U14973 (N_14973,N_13759,N_14270);
nand U14974 (N_14974,N_13767,N_14126);
nand U14975 (N_14975,N_13819,N_14084);
and U14976 (N_14976,N_14271,N_13840);
nand U14977 (N_14977,N_14202,N_14371);
or U14978 (N_14978,N_14073,N_13958);
xor U14979 (N_14979,N_13983,N_13962);
xnor U14980 (N_14980,N_14125,N_13900);
and U14981 (N_14981,N_14214,N_14166);
and U14982 (N_14982,N_14239,N_13971);
and U14983 (N_14983,N_14072,N_14155);
xor U14984 (N_14984,N_14374,N_13837);
xor U14985 (N_14985,N_13820,N_14111);
nand U14986 (N_14986,N_14106,N_14311);
and U14987 (N_14987,N_13856,N_13852);
xnor U14988 (N_14988,N_14044,N_13857);
xnor U14989 (N_14989,N_14258,N_14126);
xor U14990 (N_14990,N_13771,N_13989);
xor U14991 (N_14991,N_14185,N_13849);
xor U14992 (N_14992,N_14208,N_14072);
or U14993 (N_14993,N_14151,N_13920);
xnor U14994 (N_14994,N_14033,N_14105);
nand U14995 (N_14995,N_14223,N_14102);
or U14996 (N_14996,N_14241,N_13853);
nand U14997 (N_14997,N_14169,N_13784);
and U14998 (N_14998,N_14261,N_14319);
nand U14999 (N_14999,N_14280,N_13896);
nand U15000 (N_15000,N_14865,N_14840);
nor U15001 (N_15001,N_14503,N_14803);
xnor U15002 (N_15002,N_14686,N_14455);
and U15003 (N_15003,N_14627,N_14843);
or U15004 (N_15004,N_14544,N_14827);
or U15005 (N_15005,N_14716,N_14641);
and U15006 (N_15006,N_14480,N_14941);
nand U15007 (N_15007,N_14910,N_14674);
or U15008 (N_15008,N_14412,N_14610);
and U15009 (N_15009,N_14731,N_14599);
xnor U15010 (N_15010,N_14977,N_14856);
nand U15011 (N_15011,N_14402,N_14978);
xor U15012 (N_15012,N_14702,N_14457);
xnor U15013 (N_15013,N_14450,N_14617);
or U15014 (N_15014,N_14399,N_14701);
nor U15015 (N_15015,N_14646,N_14597);
nand U15016 (N_15016,N_14768,N_14979);
xor U15017 (N_15017,N_14394,N_14870);
nor U15018 (N_15018,N_14476,N_14628);
nand U15019 (N_15019,N_14560,N_14633);
xor U15020 (N_15020,N_14595,N_14911);
nand U15021 (N_15021,N_14728,N_14386);
xnor U15022 (N_15022,N_14539,N_14789);
nor U15023 (N_15023,N_14389,N_14917);
nand U15024 (N_15024,N_14378,N_14837);
xor U15025 (N_15025,N_14593,N_14900);
nor U15026 (N_15026,N_14821,N_14393);
and U15027 (N_15027,N_14452,N_14937);
and U15028 (N_15028,N_14835,N_14944);
and U15029 (N_15029,N_14903,N_14715);
or U15030 (N_15030,N_14523,N_14462);
nor U15031 (N_15031,N_14665,N_14783);
xnor U15032 (N_15032,N_14976,N_14406);
nand U15033 (N_15033,N_14822,N_14380);
nor U15034 (N_15034,N_14514,N_14765);
or U15035 (N_15035,N_14990,N_14551);
nor U15036 (N_15036,N_14606,N_14634);
nor U15037 (N_15037,N_14586,N_14692);
xor U15038 (N_15038,N_14531,N_14517);
xnor U15039 (N_15039,N_14582,N_14748);
xnor U15040 (N_15040,N_14687,N_14534);
and U15041 (N_15041,N_14693,N_14823);
xor U15042 (N_15042,N_14567,N_14949);
xor U15043 (N_15043,N_14738,N_14994);
or U15044 (N_15044,N_14711,N_14968);
nor U15045 (N_15045,N_14395,N_14791);
nand U15046 (N_15046,N_14490,N_14905);
nand U15047 (N_15047,N_14709,N_14706);
nor U15048 (N_15048,N_14809,N_14779);
or U15049 (N_15049,N_14722,N_14578);
or U15050 (N_15050,N_14881,N_14461);
or U15051 (N_15051,N_14598,N_14594);
or U15052 (N_15052,N_14472,N_14961);
xnor U15053 (N_15053,N_14880,N_14828);
and U15054 (N_15054,N_14463,N_14605);
and U15055 (N_15055,N_14494,N_14908);
nor U15056 (N_15056,N_14985,N_14761);
nor U15057 (N_15057,N_14799,N_14888);
xnor U15058 (N_15058,N_14815,N_14755);
xor U15059 (N_15059,N_14564,N_14671);
or U15060 (N_15060,N_14580,N_14714);
or U15061 (N_15061,N_14964,N_14973);
or U15062 (N_15062,N_14410,N_14679);
and U15063 (N_15063,N_14683,N_14915);
nor U15064 (N_15064,N_14928,N_14611);
xnor U15065 (N_15065,N_14723,N_14591);
or U15066 (N_15066,N_14689,N_14474);
nand U15067 (N_15067,N_14848,N_14736);
and U15068 (N_15068,N_14688,N_14607);
or U15069 (N_15069,N_14705,N_14533);
nand U15070 (N_15070,N_14955,N_14696);
and U15071 (N_15071,N_14887,N_14566);
and U15072 (N_15072,N_14862,N_14588);
xnor U15073 (N_15073,N_14382,N_14868);
and U15074 (N_15074,N_14666,N_14802);
and U15075 (N_15075,N_14804,N_14397);
xor U15076 (N_15076,N_14651,N_14746);
nand U15077 (N_15077,N_14574,N_14506);
nand U15078 (N_15078,N_14409,N_14855);
nand U15079 (N_15079,N_14882,N_14999);
nor U15080 (N_15080,N_14925,N_14690);
or U15081 (N_15081,N_14869,N_14966);
xnor U15082 (N_15082,N_14430,N_14515);
xor U15083 (N_15083,N_14800,N_14730);
or U15084 (N_15084,N_14613,N_14647);
or U15085 (N_15085,N_14625,N_14744);
nor U15086 (N_15086,N_14739,N_14732);
or U15087 (N_15087,N_14993,N_14411);
or U15088 (N_15088,N_14839,N_14975);
nand U15089 (N_15089,N_14581,N_14519);
or U15090 (N_15090,N_14831,N_14918);
xnor U15091 (N_15091,N_14913,N_14773);
xnor U15092 (N_15092,N_14540,N_14429);
xor U15093 (N_15093,N_14826,N_14643);
or U15094 (N_15094,N_14554,N_14616);
xnor U15095 (N_15095,N_14547,N_14619);
or U15096 (N_15096,N_14682,N_14752);
or U15097 (N_15097,N_14872,N_14885);
nor U15098 (N_15098,N_14477,N_14431);
or U15099 (N_15099,N_14454,N_14650);
nor U15100 (N_15100,N_14559,N_14974);
xor U15101 (N_15101,N_14767,N_14672);
xor U15102 (N_15102,N_14659,N_14830);
or U15103 (N_15103,N_14640,N_14493);
nand U15104 (N_15104,N_14938,N_14914);
xor U15105 (N_15105,N_14878,N_14927);
nand U15106 (N_15106,N_14957,N_14642);
and U15107 (N_15107,N_14981,N_14573);
and U15108 (N_15108,N_14727,N_14829);
nor U15109 (N_15109,N_14898,N_14632);
and U15110 (N_15110,N_14897,N_14469);
xnor U15111 (N_15111,N_14618,N_14425);
nand U15112 (N_15112,N_14700,N_14959);
nor U15113 (N_15113,N_14453,N_14987);
and U15114 (N_15114,N_14838,N_14807);
nand U15115 (N_15115,N_14496,N_14526);
nor U15116 (N_15116,N_14423,N_14576);
or U15117 (N_15117,N_14583,N_14636);
nor U15118 (N_15118,N_14766,N_14909);
nand U15119 (N_15119,N_14537,N_14753);
nand U15120 (N_15120,N_14546,N_14670);
and U15121 (N_15121,N_14524,N_14675);
or U15122 (N_15122,N_14420,N_14720);
or U15123 (N_15123,N_14568,N_14798);
xnor U15124 (N_15124,N_14663,N_14895);
or U15125 (N_15125,N_14991,N_14572);
xnor U15126 (N_15126,N_14449,N_14518);
xor U15127 (N_15127,N_14933,N_14626);
xor U15128 (N_15128,N_14417,N_14456);
xor U15129 (N_15129,N_14784,N_14851);
xor U15130 (N_15130,N_14592,N_14879);
nor U15131 (N_15131,N_14601,N_14414);
and U15132 (N_15132,N_14710,N_14513);
and U15133 (N_15133,N_14875,N_14460);
nor U15134 (N_15134,N_14747,N_14522);
and U15135 (N_15135,N_14448,N_14892);
and U15136 (N_15136,N_14770,N_14762);
or U15137 (N_15137,N_14814,N_14734);
or U15138 (N_15138,N_14434,N_14407);
xor U15139 (N_15139,N_14510,N_14750);
or U15140 (N_15140,N_14653,N_14459);
nand U15141 (N_15141,N_14704,N_14561);
and U15142 (N_15142,N_14737,N_14408);
xnor U15143 (N_15143,N_14729,N_14956);
or U15144 (N_15144,N_14388,N_14891);
or U15145 (N_15145,N_14530,N_14585);
nand U15146 (N_15146,N_14781,N_14899);
nand U15147 (N_15147,N_14437,N_14970);
and U15148 (N_15148,N_14621,N_14889);
or U15149 (N_15149,N_14986,N_14376);
or U15150 (N_15150,N_14836,N_14971);
nor U15151 (N_15151,N_14805,N_14769);
xnor U15152 (N_15152,N_14669,N_14782);
or U15153 (N_15153,N_14849,N_14565);
or U15154 (N_15154,N_14624,N_14525);
and U15155 (N_15155,N_14404,N_14932);
nand U15156 (N_15156,N_14631,N_14439);
and U15157 (N_15157,N_14857,N_14542);
xnor U15158 (N_15158,N_14569,N_14742);
nor U15159 (N_15159,N_14777,N_14963);
xnor U15160 (N_15160,N_14906,N_14778);
nand U15161 (N_15161,N_14801,N_14620);
nand U15162 (N_15162,N_14751,N_14912);
nand U15163 (N_15163,N_14475,N_14396);
nor U15164 (N_15164,N_14708,N_14890);
nor U15165 (N_15165,N_14614,N_14931);
xnor U15166 (N_15166,N_14749,N_14864);
xnor U15167 (N_15167,N_14383,N_14527);
nand U15168 (N_15168,N_14577,N_14953);
nor U15169 (N_15169,N_14844,N_14668);
or U15170 (N_15170,N_14451,N_14441);
nand U15171 (N_15171,N_14458,N_14733);
nor U15172 (N_15172,N_14743,N_14507);
nor U15173 (N_15173,N_14965,N_14657);
or U15174 (N_15174,N_14645,N_14652);
nor U15175 (N_15175,N_14923,N_14866);
or U15176 (N_15176,N_14511,N_14757);
xnor U15177 (N_15177,N_14379,N_14609);
nor U15178 (N_15178,N_14886,N_14724);
and U15179 (N_15179,N_14995,N_14387);
or U15180 (N_15180,N_14992,N_14658);
xnor U15181 (N_15181,N_14982,N_14629);
or U15182 (N_15182,N_14557,N_14983);
nand U15183 (N_15183,N_14902,N_14392);
or U15184 (N_15184,N_14413,N_14442);
or U15185 (N_15185,N_14501,N_14787);
xor U15186 (N_15186,N_14754,N_14951);
or U15187 (N_15187,N_14936,N_14685);
nand U15188 (N_15188,N_14579,N_14471);
nor U15189 (N_15189,N_14846,N_14764);
and U15190 (N_15190,N_14400,N_14681);
and U15191 (N_15191,N_14589,N_14924);
xnor U15192 (N_15192,N_14958,N_14930);
xor U15193 (N_15193,N_14529,N_14435);
or U15194 (N_15194,N_14398,N_14418);
and U15195 (N_15195,N_14952,N_14945);
xor U15196 (N_15196,N_14859,N_14824);
nor U15197 (N_15197,N_14385,N_14896);
xnor U15198 (N_15198,N_14447,N_14570);
nand U15199 (N_15199,N_14445,N_14793);
and U15200 (N_15200,N_14488,N_14997);
xor U15201 (N_15201,N_14390,N_14863);
nor U15202 (N_15202,N_14502,N_14760);
or U15203 (N_15203,N_14818,N_14649);
and U15204 (N_15204,N_14813,N_14549);
and U15205 (N_15205,N_14491,N_14939);
nor U15206 (N_15206,N_14479,N_14639);
nor U15207 (N_15207,N_14419,N_14726);
or U15208 (N_15208,N_14998,N_14446);
nor U15209 (N_15209,N_14725,N_14416);
xnor U15210 (N_15210,N_14622,N_14548);
xnor U15211 (N_15211,N_14972,N_14482);
and U15212 (N_15212,N_14543,N_14984);
or U15213 (N_15213,N_14604,N_14916);
xor U15214 (N_15214,N_14630,N_14440);
nor U15215 (N_15215,N_14432,N_14771);
and U15216 (N_15216,N_14988,N_14788);
or U15217 (N_15217,N_14512,N_14426);
nor U15218 (N_15218,N_14558,N_14942);
or U15219 (N_15219,N_14673,N_14883);
nor U15220 (N_15220,N_14684,N_14536);
xor U15221 (N_15221,N_14528,N_14841);
xor U15222 (N_15222,N_14497,N_14735);
or U15223 (N_15223,N_14660,N_14858);
nand U15224 (N_15224,N_14817,N_14508);
or U15225 (N_15225,N_14719,N_14873);
xnor U15226 (N_15226,N_14648,N_14465);
and U15227 (N_15227,N_14545,N_14509);
xor U15228 (N_15228,N_14854,N_14467);
or U15229 (N_15229,N_14667,N_14877);
nand U15230 (N_15230,N_14820,N_14842);
or U15231 (N_15231,N_14833,N_14483);
or U15232 (N_15232,N_14785,N_14795);
and U15233 (N_15233,N_14960,N_14717);
nor U15234 (N_15234,N_14780,N_14521);
xor U15235 (N_15235,N_14834,N_14563);
or U15236 (N_15236,N_14384,N_14806);
nor U15237 (N_15237,N_14847,N_14444);
nor U15238 (N_15238,N_14405,N_14871);
nand U15239 (N_15239,N_14741,N_14421);
or U15240 (N_15240,N_14946,N_14495);
nand U15241 (N_15241,N_14662,N_14904);
xor U15242 (N_15242,N_14608,N_14943);
nand U15243 (N_15243,N_14699,N_14377);
and U15244 (N_15244,N_14600,N_14954);
xnor U15245 (N_15245,N_14562,N_14484);
nand U15246 (N_15246,N_14694,N_14745);
or U15247 (N_15247,N_14740,N_14989);
nand U15248 (N_15248,N_14721,N_14893);
or U15249 (N_15249,N_14424,N_14940);
xor U15250 (N_15250,N_14466,N_14401);
nor U15251 (N_15251,N_14676,N_14615);
xnor U15252 (N_15252,N_14655,N_14758);
or U15253 (N_15253,N_14464,N_14678);
or U15254 (N_15254,N_14926,N_14661);
nor U15255 (N_15255,N_14492,N_14861);
nand U15256 (N_15256,N_14555,N_14894);
and U15257 (N_15257,N_14697,N_14756);
xnor U15258 (N_15258,N_14920,N_14575);
or U15259 (N_15259,N_14935,N_14532);
nor U15260 (N_15260,N_14516,N_14695);
xor U15261 (N_15261,N_14481,N_14443);
and U15262 (N_15262,N_14929,N_14680);
nor U15263 (N_15263,N_14486,N_14656);
xnor U15264 (N_15264,N_14919,N_14612);
nor U15265 (N_15265,N_14500,N_14811);
nor U15266 (N_15266,N_14774,N_14853);
and U15267 (N_15267,N_14812,N_14677);
and U15268 (N_15268,N_14422,N_14470);
nor U15269 (N_15269,N_14552,N_14550);
nand U15270 (N_15270,N_14776,N_14884);
or U15271 (N_15271,N_14775,N_14796);
and U15272 (N_15272,N_14786,N_14571);
nand U15273 (N_15273,N_14556,N_14375);
xor U15274 (N_15274,N_14772,N_14438);
xnor U15275 (N_15275,N_14541,N_14934);
xnor U15276 (N_15276,N_14845,N_14901);
xor U15277 (N_15277,N_14948,N_14584);
and U15278 (N_15278,N_14602,N_14969);
or U15279 (N_15279,N_14980,N_14763);
and U15280 (N_15280,N_14644,N_14850);
and U15281 (N_15281,N_14874,N_14478);
nand U15282 (N_15282,N_14436,N_14499);
nand U15283 (N_15283,N_14415,N_14962);
or U15284 (N_15284,N_14712,N_14921);
nand U15285 (N_15285,N_14816,N_14759);
or U15286 (N_15286,N_14520,N_14950);
and U15287 (N_15287,N_14810,N_14587);
and U15288 (N_15288,N_14485,N_14867);
nand U15289 (N_15289,N_14596,N_14403);
or U15290 (N_15290,N_14468,N_14797);
or U15291 (N_15291,N_14473,N_14590);
nand U15292 (N_15292,N_14637,N_14967);
xor U15293 (N_15293,N_14691,N_14947);
nor U15294 (N_15294,N_14819,N_14876);
or U15295 (N_15295,N_14538,N_14654);
nor U15296 (N_15296,N_14498,N_14794);
nand U15297 (N_15297,N_14489,N_14718);
xnor U15298 (N_15298,N_14703,N_14433);
xnor U15299 (N_15299,N_14635,N_14623);
or U15300 (N_15300,N_14664,N_14638);
xnor U15301 (N_15301,N_14428,N_14603);
xor U15302 (N_15302,N_14487,N_14713);
xor U15303 (N_15303,N_14698,N_14922);
nor U15304 (N_15304,N_14792,N_14553);
nor U15305 (N_15305,N_14808,N_14391);
and U15306 (N_15306,N_14381,N_14707);
or U15307 (N_15307,N_14790,N_14825);
or U15308 (N_15308,N_14852,N_14832);
xnor U15309 (N_15309,N_14996,N_14505);
nor U15310 (N_15310,N_14907,N_14535);
nand U15311 (N_15311,N_14860,N_14504);
nor U15312 (N_15312,N_14427,N_14806);
nor U15313 (N_15313,N_14678,N_14679);
or U15314 (N_15314,N_14833,N_14718);
nand U15315 (N_15315,N_14888,N_14698);
and U15316 (N_15316,N_14847,N_14589);
or U15317 (N_15317,N_14965,N_14433);
nand U15318 (N_15318,N_14491,N_14480);
nor U15319 (N_15319,N_14950,N_14668);
or U15320 (N_15320,N_14887,N_14427);
xor U15321 (N_15321,N_14926,N_14845);
xnor U15322 (N_15322,N_14576,N_14480);
nor U15323 (N_15323,N_14963,N_14759);
or U15324 (N_15324,N_14873,N_14612);
and U15325 (N_15325,N_14388,N_14746);
and U15326 (N_15326,N_14389,N_14413);
nor U15327 (N_15327,N_14757,N_14817);
nand U15328 (N_15328,N_14969,N_14671);
nand U15329 (N_15329,N_14966,N_14479);
and U15330 (N_15330,N_14793,N_14993);
nand U15331 (N_15331,N_14777,N_14672);
or U15332 (N_15332,N_14468,N_14498);
xor U15333 (N_15333,N_14491,N_14552);
or U15334 (N_15334,N_14483,N_14606);
xnor U15335 (N_15335,N_14481,N_14438);
and U15336 (N_15336,N_14772,N_14956);
or U15337 (N_15337,N_14601,N_14548);
xnor U15338 (N_15338,N_14712,N_14849);
nand U15339 (N_15339,N_14706,N_14618);
or U15340 (N_15340,N_14826,N_14629);
or U15341 (N_15341,N_14956,N_14442);
or U15342 (N_15342,N_14927,N_14941);
nor U15343 (N_15343,N_14384,N_14780);
nor U15344 (N_15344,N_14381,N_14919);
or U15345 (N_15345,N_14687,N_14953);
and U15346 (N_15346,N_14544,N_14828);
nand U15347 (N_15347,N_14734,N_14904);
xor U15348 (N_15348,N_14687,N_14403);
xnor U15349 (N_15349,N_14536,N_14411);
xnor U15350 (N_15350,N_14878,N_14999);
nor U15351 (N_15351,N_14845,N_14636);
or U15352 (N_15352,N_14875,N_14851);
and U15353 (N_15353,N_14828,N_14745);
nand U15354 (N_15354,N_14804,N_14930);
xnor U15355 (N_15355,N_14863,N_14919);
xnor U15356 (N_15356,N_14390,N_14964);
and U15357 (N_15357,N_14858,N_14449);
nand U15358 (N_15358,N_14415,N_14744);
nand U15359 (N_15359,N_14589,N_14385);
or U15360 (N_15360,N_14409,N_14594);
nand U15361 (N_15361,N_14507,N_14681);
nor U15362 (N_15362,N_14656,N_14395);
xnor U15363 (N_15363,N_14634,N_14769);
and U15364 (N_15364,N_14464,N_14763);
xnor U15365 (N_15365,N_14994,N_14721);
xor U15366 (N_15366,N_14971,N_14812);
and U15367 (N_15367,N_14644,N_14947);
xor U15368 (N_15368,N_14451,N_14676);
nor U15369 (N_15369,N_14828,N_14800);
nor U15370 (N_15370,N_14407,N_14726);
and U15371 (N_15371,N_14748,N_14667);
nand U15372 (N_15372,N_14617,N_14671);
nor U15373 (N_15373,N_14694,N_14876);
xnor U15374 (N_15374,N_14580,N_14612);
and U15375 (N_15375,N_14823,N_14555);
xnor U15376 (N_15376,N_14823,N_14972);
xor U15377 (N_15377,N_14971,N_14646);
and U15378 (N_15378,N_14715,N_14616);
and U15379 (N_15379,N_14458,N_14972);
or U15380 (N_15380,N_14611,N_14464);
nor U15381 (N_15381,N_14906,N_14799);
and U15382 (N_15382,N_14870,N_14959);
and U15383 (N_15383,N_14947,N_14627);
and U15384 (N_15384,N_14899,N_14636);
nor U15385 (N_15385,N_14635,N_14533);
xnor U15386 (N_15386,N_14904,N_14933);
or U15387 (N_15387,N_14911,N_14946);
nor U15388 (N_15388,N_14497,N_14919);
and U15389 (N_15389,N_14390,N_14955);
nand U15390 (N_15390,N_14523,N_14826);
nor U15391 (N_15391,N_14614,N_14578);
or U15392 (N_15392,N_14907,N_14396);
nor U15393 (N_15393,N_14761,N_14917);
nor U15394 (N_15394,N_14879,N_14795);
or U15395 (N_15395,N_14722,N_14960);
nand U15396 (N_15396,N_14727,N_14934);
nand U15397 (N_15397,N_14528,N_14682);
or U15398 (N_15398,N_14782,N_14454);
and U15399 (N_15399,N_14963,N_14425);
and U15400 (N_15400,N_14725,N_14596);
nor U15401 (N_15401,N_14521,N_14427);
nand U15402 (N_15402,N_14467,N_14961);
or U15403 (N_15403,N_14779,N_14784);
and U15404 (N_15404,N_14449,N_14477);
nand U15405 (N_15405,N_14457,N_14713);
nand U15406 (N_15406,N_14922,N_14389);
and U15407 (N_15407,N_14905,N_14414);
nor U15408 (N_15408,N_14774,N_14593);
nor U15409 (N_15409,N_14741,N_14584);
nor U15410 (N_15410,N_14792,N_14725);
and U15411 (N_15411,N_14501,N_14606);
nand U15412 (N_15412,N_14517,N_14961);
or U15413 (N_15413,N_14751,N_14519);
nand U15414 (N_15414,N_14718,N_14654);
nand U15415 (N_15415,N_14754,N_14472);
or U15416 (N_15416,N_14550,N_14814);
nor U15417 (N_15417,N_14860,N_14571);
or U15418 (N_15418,N_14879,N_14601);
nand U15419 (N_15419,N_14815,N_14779);
nand U15420 (N_15420,N_14822,N_14763);
xor U15421 (N_15421,N_14937,N_14380);
nand U15422 (N_15422,N_14762,N_14717);
or U15423 (N_15423,N_14604,N_14720);
nor U15424 (N_15424,N_14845,N_14454);
nor U15425 (N_15425,N_14921,N_14549);
nand U15426 (N_15426,N_14959,N_14889);
and U15427 (N_15427,N_14692,N_14735);
nor U15428 (N_15428,N_14678,N_14542);
xnor U15429 (N_15429,N_14837,N_14431);
nor U15430 (N_15430,N_14818,N_14704);
and U15431 (N_15431,N_14660,N_14480);
or U15432 (N_15432,N_14597,N_14541);
nor U15433 (N_15433,N_14751,N_14399);
or U15434 (N_15434,N_14518,N_14423);
and U15435 (N_15435,N_14535,N_14745);
or U15436 (N_15436,N_14736,N_14830);
or U15437 (N_15437,N_14390,N_14944);
or U15438 (N_15438,N_14991,N_14986);
nor U15439 (N_15439,N_14917,N_14605);
nand U15440 (N_15440,N_14499,N_14709);
or U15441 (N_15441,N_14822,N_14935);
and U15442 (N_15442,N_14512,N_14591);
and U15443 (N_15443,N_14586,N_14828);
and U15444 (N_15444,N_14880,N_14845);
xnor U15445 (N_15445,N_14633,N_14745);
nor U15446 (N_15446,N_14672,N_14576);
xor U15447 (N_15447,N_14841,N_14931);
nand U15448 (N_15448,N_14450,N_14998);
xor U15449 (N_15449,N_14715,N_14706);
nor U15450 (N_15450,N_14763,N_14992);
nand U15451 (N_15451,N_14709,N_14442);
and U15452 (N_15452,N_14763,N_14562);
xnor U15453 (N_15453,N_14643,N_14574);
and U15454 (N_15454,N_14434,N_14879);
xnor U15455 (N_15455,N_14747,N_14680);
xnor U15456 (N_15456,N_14942,N_14468);
nand U15457 (N_15457,N_14688,N_14831);
nor U15458 (N_15458,N_14695,N_14585);
xor U15459 (N_15459,N_14484,N_14490);
nor U15460 (N_15460,N_14531,N_14846);
and U15461 (N_15461,N_14768,N_14980);
nand U15462 (N_15462,N_14862,N_14453);
nor U15463 (N_15463,N_14415,N_14877);
nor U15464 (N_15464,N_14564,N_14554);
or U15465 (N_15465,N_14408,N_14383);
nor U15466 (N_15466,N_14698,N_14645);
nand U15467 (N_15467,N_14644,N_14971);
xor U15468 (N_15468,N_14787,N_14591);
nand U15469 (N_15469,N_14593,N_14875);
and U15470 (N_15470,N_14755,N_14850);
or U15471 (N_15471,N_14555,N_14583);
xor U15472 (N_15472,N_14451,N_14536);
nor U15473 (N_15473,N_14533,N_14647);
nor U15474 (N_15474,N_14408,N_14398);
nand U15475 (N_15475,N_14568,N_14982);
xor U15476 (N_15476,N_14779,N_14685);
nand U15477 (N_15477,N_14403,N_14393);
nor U15478 (N_15478,N_14434,N_14892);
xor U15479 (N_15479,N_14892,N_14637);
xor U15480 (N_15480,N_14805,N_14549);
xnor U15481 (N_15481,N_14496,N_14477);
xor U15482 (N_15482,N_14384,N_14859);
xnor U15483 (N_15483,N_14778,N_14753);
nand U15484 (N_15484,N_14494,N_14924);
xor U15485 (N_15485,N_14688,N_14899);
xnor U15486 (N_15486,N_14608,N_14429);
and U15487 (N_15487,N_14410,N_14719);
nand U15488 (N_15488,N_14917,N_14658);
xor U15489 (N_15489,N_14988,N_14622);
nand U15490 (N_15490,N_14637,N_14643);
nor U15491 (N_15491,N_14699,N_14404);
nor U15492 (N_15492,N_14816,N_14778);
or U15493 (N_15493,N_14756,N_14978);
xor U15494 (N_15494,N_14974,N_14574);
xor U15495 (N_15495,N_14827,N_14497);
nand U15496 (N_15496,N_14797,N_14573);
xnor U15497 (N_15497,N_14641,N_14436);
nor U15498 (N_15498,N_14706,N_14525);
nand U15499 (N_15499,N_14658,N_14692);
nor U15500 (N_15500,N_14495,N_14655);
or U15501 (N_15501,N_14739,N_14665);
and U15502 (N_15502,N_14782,N_14668);
xor U15503 (N_15503,N_14820,N_14505);
xor U15504 (N_15504,N_14424,N_14993);
nor U15505 (N_15505,N_14568,N_14557);
or U15506 (N_15506,N_14675,N_14827);
nand U15507 (N_15507,N_14847,N_14898);
xor U15508 (N_15508,N_14500,N_14720);
or U15509 (N_15509,N_14559,N_14940);
nor U15510 (N_15510,N_14924,N_14917);
and U15511 (N_15511,N_14536,N_14401);
nor U15512 (N_15512,N_14545,N_14736);
xnor U15513 (N_15513,N_14603,N_14996);
nand U15514 (N_15514,N_14558,N_14712);
xor U15515 (N_15515,N_14799,N_14610);
xor U15516 (N_15516,N_14982,N_14917);
nor U15517 (N_15517,N_14957,N_14976);
or U15518 (N_15518,N_14716,N_14714);
and U15519 (N_15519,N_14950,N_14634);
nand U15520 (N_15520,N_14617,N_14750);
xor U15521 (N_15521,N_14747,N_14793);
xnor U15522 (N_15522,N_14898,N_14991);
xnor U15523 (N_15523,N_14818,N_14942);
nor U15524 (N_15524,N_14935,N_14781);
xor U15525 (N_15525,N_14558,N_14905);
nor U15526 (N_15526,N_14396,N_14681);
xnor U15527 (N_15527,N_14435,N_14993);
or U15528 (N_15528,N_14494,N_14960);
xor U15529 (N_15529,N_14665,N_14928);
xor U15530 (N_15530,N_14466,N_14381);
or U15531 (N_15531,N_14787,N_14459);
nand U15532 (N_15532,N_14893,N_14996);
and U15533 (N_15533,N_14602,N_14438);
or U15534 (N_15534,N_14759,N_14459);
nand U15535 (N_15535,N_14956,N_14706);
nand U15536 (N_15536,N_14819,N_14867);
nor U15537 (N_15537,N_14629,N_14622);
nand U15538 (N_15538,N_14925,N_14411);
and U15539 (N_15539,N_14734,N_14721);
and U15540 (N_15540,N_14690,N_14759);
and U15541 (N_15541,N_14475,N_14455);
nand U15542 (N_15542,N_14468,N_14419);
and U15543 (N_15543,N_14710,N_14629);
and U15544 (N_15544,N_14495,N_14669);
or U15545 (N_15545,N_14645,N_14765);
and U15546 (N_15546,N_14743,N_14495);
nor U15547 (N_15547,N_14931,N_14513);
or U15548 (N_15548,N_14747,N_14812);
and U15549 (N_15549,N_14535,N_14886);
or U15550 (N_15550,N_14615,N_14698);
or U15551 (N_15551,N_14818,N_14434);
or U15552 (N_15552,N_14631,N_14432);
xor U15553 (N_15553,N_14909,N_14413);
xnor U15554 (N_15554,N_14528,N_14935);
nand U15555 (N_15555,N_14673,N_14585);
nor U15556 (N_15556,N_14891,N_14671);
xnor U15557 (N_15557,N_14839,N_14652);
or U15558 (N_15558,N_14765,N_14625);
or U15559 (N_15559,N_14383,N_14767);
nand U15560 (N_15560,N_14696,N_14726);
xor U15561 (N_15561,N_14878,N_14920);
nand U15562 (N_15562,N_14376,N_14553);
or U15563 (N_15563,N_14440,N_14910);
xor U15564 (N_15564,N_14614,N_14883);
nand U15565 (N_15565,N_14933,N_14798);
and U15566 (N_15566,N_14912,N_14946);
or U15567 (N_15567,N_14383,N_14999);
and U15568 (N_15568,N_14890,N_14450);
xor U15569 (N_15569,N_14573,N_14631);
or U15570 (N_15570,N_14566,N_14748);
or U15571 (N_15571,N_14695,N_14451);
or U15572 (N_15572,N_14720,N_14562);
xnor U15573 (N_15573,N_14470,N_14877);
and U15574 (N_15574,N_14824,N_14423);
nand U15575 (N_15575,N_14774,N_14589);
xnor U15576 (N_15576,N_14475,N_14596);
nor U15577 (N_15577,N_14792,N_14945);
nand U15578 (N_15578,N_14407,N_14967);
xor U15579 (N_15579,N_14695,N_14849);
nor U15580 (N_15580,N_14509,N_14529);
and U15581 (N_15581,N_14762,N_14870);
and U15582 (N_15582,N_14672,N_14600);
nor U15583 (N_15583,N_14773,N_14701);
xor U15584 (N_15584,N_14851,N_14662);
xnor U15585 (N_15585,N_14932,N_14840);
nor U15586 (N_15586,N_14607,N_14767);
or U15587 (N_15587,N_14730,N_14954);
nand U15588 (N_15588,N_14573,N_14822);
nor U15589 (N_15589,N_14582,N_14605);
and U15590 (N_15590,N_14518,N_14917);
and U15591 (N_15591,N_14639,N_14676);
xnor U15592 (N_15592,N_14562,N_14393);
or U15593 (N_15593,N_14995,N_14704);
nand U15594 (N_15594,N_14718,N_14749);
and U15595 (N_15595,N_14984,N_14899);
nor U15596 (N_15596,N_14601,N_14487);
and U15597 (N_15597,N_14609,N_14691);
nor U15598 (N_15598,N_14751,N_14932);
nor U15599 (N_15599,N_14459,N_14954);
nand U15600 (N_15600,N_14979,N_14862);
nor U15601 (N_15601,N_14625,N_14984);
xnor U15602 (N_15602,N_14502,N_14829);
or U15603 (N_15603,N_14421,N_14479);
or U15604 (N_15604,N_14851,N_14611);
or U15605 (N_15605,N_14443,N_14381);
xnor U15606 (N_15606,N_14636,N_14376);
and U15607 (N_15607,N_14555,N_14728);
xor U15608 (N_15608,N_14506,N_14385);
nand U15609 (N_15609,N_14712,N_14432);
nand U15610 (N_15610,N_14665,N_14533);
or U15611 (N_15611,N_14920,N_14765);
or U15612 (N_15612,N_14934,N_14868);
or U15613 (N_15613,N_14646,N_14907);
nor U15614 (N_15614,N_14612,N_14766);
nor U15615 (N_15615,N_14620,N_14791);
nand U15616 (N_15616,N_14673,N_14696);
or U15617 (N_15617,N_14511,N_14648);
xnor U15618 (N_15618,N_14449,N_14640);
nand U15619 (N_15619,N_14552,N_14700);
or U15620 (N_15620,N_14965,N_14795);
xor U15621 (N_15621,N_14663,N_14816);
nand U15622 (N_15622,N_14620,N_14382);
nor U15623 (N_15623,N_14725,N_14491);
and U15624 (N_15624,N_14750,N_14572);
or U15625 (N_15625,N_15186,N_15457);
or U15626 (N_15626,N_15237,N_15328);
nand U15627 (N_15627,N_15319,N_15573);
xor U15628 (N_15628,N_15274,N_15444);
nand U15629 (N_15629,N_15144,N_15620);
nand U15630 (N_15630,N_15165,N_15018);
or U15631 (N_15631,N_15502,N_15490);
and U15632 (N_15632,N_15406,N_15145);
and U15633 (N_15633,N_15437,N_15324);
or U15634 (N_15634,N_15570,N_15006);
or U15635 (N_15635,N_15407,N_15501);
nor U15636 (N_15636,N_15472,N_15529);
xnor U15637 (N_15637,N_15446,N_15424);
and U15638 (N_15638,N_15057,N_15089);
nand U15639 (N_15639,N_15038,N_15115);
nand U15640 (N_15640,N_15409,N_15378);
xnor U15641 (N_15641,N_15366,N_15345);
nor U15642 (N_15642,N_15010,N_15303);
xor U15643 (N_15643,N_15403,N_15429);
nor U15644 (N_15644,N_15385,N_15491);
nor U15645 (N_15645,N_15558,N_15216);
or U15646 (N_15646,N_15100,N_15272);
xor U15647 (N_15647,N_15141,N_15454);
nand U15648 (N_15648,N_15563,N_15344);
xnor U15649 (N_15649,N_15126,N_15221);
nor U15650 (N_15650,N_15252,N_15200);
xor U15651 (N_15651,N_15325,N_15542);
xor U15652 (N_15652,N_15393,N_15477);
xor U15653 (N_15653,N_15132,N_15594);
xor U15654 (N_15654,N_15220,N_15508);
nand U15655 (N_15655,N_15230,N_15586);
and U15656 (N_15656,N_15166,N_15014);
nor U15657 (N_15657,N_15205,N_15447);
or U15658 (N_15658,N_15381,N_15597);
or U15659 (N_15659,N_15269,N_15267);
or U15660 (N_15660,N_15142,N_15521);
nand U15661 (N_15661,N_15131,N_15282);
or U15662 (N_15662,N_15510,N_15468);
nor U15663 (N_15663,N_15579,N_15334);
and U15664 (N_15664,N_15149,N_15375);
and U15665 (N_15665,N_15261,N_15493);
xor U15666 (N_15666,N_15433,N_15607);
and U15667 (N_15667,N_15610,N_15555);
nor U15668 (N_15668,N_15313,N_15562);
and U15669 (N_15669,N_15075,N_15373);
or U15670 (N_15670,N_15288,N_15096);
nor U15671 (N_15671,N_15157,N_15609);
nor U15672 (N_15672,N_15362,N_15600);
or U15673 (N_15673,N_15330,N_15370);
and U15674 (N_15674,N_15449,N_15314);
nand U15675 (N_15675,N_15538,N_15257);
or U15676 (N_15676,N_15582,N_15440);
nor U15677 (N_15677,N_15369,N_15549);
or U15678 (N_15678,N_15537,N_15540);
or U15679 (N_15679,N_15411,N_15172);
nor U15680 (N_15680,N_15225,N_15063);
or U15681 (N_15681,N_15129,N_15123);
and U15682 (N_15682,N_15333,N_15422);
nor U15683 (N_15683,N_15169,N_15599);
nor U15684 (N_15684,N_15109,N_15470);
or U15685 (N_15685,N_15374,N_15467);
or U15686 (N_15686,N_15613,N_15178);
or U15687 (N_15687,N_15404,N_15488);
or U15688 (N_15688,N_15384,N_15232);
nand U15689 (N_15689,N_15419,N_15055);
nor U15690 (N_15690,N_15133,N_15320);
nor U15691 (N_15691,N_15280,N_15505);
nor U15692 (N_15692,N_15294,N_15368);
xor U15693 (N_15693,N_15536,N_15532);
nand U15694 (N_15694,N_15047,N_15509);
nor U15695 (N_15695,N_15341,N_15154);
nand U15696 (N_15696,N_15098,N_15606);
nand U15697 (N_15697,N_15545,N_15360);
nor U15698 (N_15698,N_15079,N_15060);
or U15699 (N_15699,N_15116,N_15326);
or U15700 (N_15700,N_15571,N_15371);
xnor U15701 (N_15701,N_15179,N_15605);
nand U15702 (N_15702,N_15355,N_15199);
nor U15703 (N_15703,N_15574,N_15059);
and U15704 (N_15704,N_15614,N_15399);
and U15705 (N_15705,N_15479,N_15158);
nand U15706 (N_15706,N_15162,N_15560);
nor U15707 (N_15707,N_15364,N_15164);
nand U15708 (N_15708,N_15548,N_15443);
and U15709 (N_15709,N_15386,N_15522);
and U15710 (N_15710,N_15417,N_15050);
or U15711 (N_15711,N_15475,N_15283);
xnor U15712 (N_15712,N_15593,N_15278);
and U15713 (N_15713,N_15256,N_15530);
nand U15714 (N_15714,N_15321,N_15234);
or U15715 (N_15715,N_15284,N_15361);
xor U15716 (N_15716,N_15260,N_15622);
nand U15717 (N_15717,N_15596,N_15617);
and U15718 (N_15718,N_15623,N_15027);
nor U15719 (N_15719,N_15161,N_15524);
xnor U15720 (N_15720,N_15238,N_15483);
nand U15721 (N_15721,N_15557,N_15058);
and U15722 (N_15722,N_15020,N_15365);
xor U15723 (N_15723,N_15022,N_15621);
xnor U15724 (N_15724,N_15580,N_15137);
and U15725 (N_15725,N_15194,N_15004);
xor U15726 (N_15726,N_15598,N_15347);
or U15727 (N_15727,N_15286,N_15421);
or U15728 (N_15728,N_15255,N_15601);
nor U15729 (N_15729,N_15130,N_15181);
and U15730 (N_15730,N_15413,N_15327);
or U15731 (N_15731,N_15308,N_15067);
nor U15732 (N_15732,N_15412,N_15212);
and U15733 (N_15733,N_15478,N_15352);
or U15734 (N_15734,N_15246,N_15235);
nor U15735 (N_15735,N_15595,N_15189);
xnor U15736 (N_15736,N_15624,N_15346);
and U15737 (N_15737,N_15223,N_15083);
nand U15738 (N_15738,N_15460,N_15340);
nand U15739 (N_15739,N_15143,N_15489);
nand U15740 (N_15740,N_15188,N_15008);
and U15741 (N_15741,N_15439,N_15233);
nor U15742 (N_15742,N_15052,N_15054);
xor U15743 (N_15743,N_15480,N_15611);
or U15744 (N_15744,N_15565,N_15302);
and U15745 (N_15745,N_15315,N_15011);
or U15746 (N_15746,N_15306,N_15295);
xor U15747 (N_15747,N_15250,N_15281);
nand U15748 (N_15748,N_15533,N_15300);
xor U15749 (N_15749,N_15547,N_15243);
or U15750 (N_15750,N_15113,N_15608);
nand U15751 (N_15751,N_15139,N_15202);
nand U15752 (N_15752,N_15183,N_15318);
nor U15753 (N_15753,N_15253,N_15061);
nor U15754 (N_15754,N_15190,N_15591);
xor U15755 (N_15755,N_15270,N_15400);
nand U15756 (N_15756,N_15170,N_15209);
xor U15757 (N_15757,N_15051,N_15358);
and U15758 (N_15758,N_15031,N_15575);
or U15759 (N_15759,N_15535,N_15092);
nand U15760 (N_15760,N_15239,N_15019);
xnor U15761 (N_15761,N_15392,N_15367);
and U15762 (N_15762,N_15275,N_15523);
nor U15763 (N_15763,N_15091,N_15588);
and U15764 (N_15764,N_15329,N_15081);
or U15765 (N_15765,N_15394,N_15021);
nor U15766 (N_15766,N_15040,N_15507);
nand U15767 (N_15767,N_15331,N_15312);
and U15768 (N_15768,N_15003,N_15397);
xor U15769 (N_15769,N_15526,N_15259);
and U15770 (N_15770,N_15175,N_15520);
nand U15771 (N_15771,N_15258,N_15531);
or U15772 (N_15772,N_15553,N_15567);
and U15773 (N_15773,N_15583,N_15121);
and U15774 (N_15774,N_15114,N_15168);
or U15775 (N_15775,N_15527,N_15076);
nand U15776 (N_15776,N_15568,N_15110);
nor U15777 (N_15777,N_15512,N_15180);
xor U15778 (N_15778,N_15482,N_15388);
or U15779 (N_15779,N_15140,N_15117);
or U15780 (N_15780,N_15077,N_15576);
nor U15781 (N_15781,N_15518,N_15391);
or U15782 (N_15782,N_15556,N_15049);
and U15783 (N_15783,N_15002,N_15101);
or U15784 (N_15784,N_15438,N_15000);
nor U15785 (N_15785,N_15351,N_15338);
or U15786 (N_15786,N_15465,N_15078);
xor U15787 (N_15787,N_15554,N_15435);
nor U15788 (N_15788,N_15273,N_15147);
xnor U15789 (N_15789,N_15163,N_15012);
xor U15790 (N_15790,N_15276,N_15013);
and U15791 (N_15791,N_15396,N_15456);
or U15792 (N_15792,N_15289,N_15085);
or U15793 (N_15793,N_15036,N_15498);
nor U15794 (N_15794,N_15587,N_15032);
xnor U15795 (N_15795,N_15156,N_15105);
and U15796 (N_15796,N_15197,N_15087);
xor U15797 (N_15797,N_15108,N_15310);
xor U15798 (N_15798,N_15492,N_15048);
and U15799 (N_15799,N_15263,N_15045);
or U15800 (N_15800,N_15160,N_15128);
or U15801 (N_15801,N_15453,N_15213);
xor U15802 (N_15802,N_15569,N_15543);
and U15803 (N_15803,N_15578,N_15211);
nor U15804 (N_15804,N_15566,N_15309);
and U15805 (N_15805,N_15222,N_15187);
xor U15806 (N_15806,N_15317,N_15427);
or U15807 (N_15807,N_15219,N_15146);
xnor U15808 (N_15808,N_15033,N_15174);
and U15809 (N_15809,N_15009,N_15466);
and U15810 (N_15810,N_15217,N_15119);
and U15811 (N_15811,N_15451,N_15247);
nor U15812 (N_15812,N_15041,N_15441);
xnor U15813 (N_15813,N_15177,N_15240);
or U15814 (N_15814,N_15511,N_15426);
or U15815 (N_15815,N_15065,N_15503);
nor U15816 (N_15816,N_15215,N_15462);
nor U15817 (N_15817,N_15185,N_15514);
nand U15818 (N_15818,N_15420,N_15134);
xor U15819 (N_15819,N_15390,N_15432);
nor U15820 (N_15820,N_15589,N_15398);
and U15821 (N_15821,N_15459,N_15264);
nand U15822 (N_15822,N_15572,N_15069);
and U15823 (N_15823,N_15208,N_15042);
or U15824 (N_15824,N_15402,N_15332);
and U15825 (N_15825,N_15546,N_15350);
nor U15826 (N_15826,N_15266,N_15410);
and U15827 (N_15827,N_15292,N_15118);
nor U15828 (N_15828,N_15207,N_15618);
or U15829 (N_15829,N_15301,N_15495);
and U15830 (N_15830,N_15425,N_15044);
nor U15831 (N_15831,N_15463,N_15201);
nor U15832 (N_15832,N_15029,N_15564);
and U15833 (N_15833,N_15372,N_15182);
and U15834 (N_15834,N_15592,N_15070);
nand U15835 (N_15835,N_15349,N_15226);
nand U15836 (N_15836,N_15228,N_15290);
and U15837 (N_15837,N_15448,N_15389);
nand U15838 (N_15838,N_15436,N_15025);
or U15839 (N_15839,N_15363,N_15550);
and U15840 (N_15840,N_15107,N_15210);
or U15841 (N_15841,N_15464,N_15539);
or U15842 (N_15842,N_15559,N_15423);
nor U15843 (N_15843,N_15030,N_15103);
nor U15844 (N_15844,N_15171,N_15516);
or U15845 (N_15845,N_15016,N_15007);
nor U15846 (N_15846,N_15336,N_15307);
xor U15847 (N_15847,N_15619,N_15053);
and U15848 (N_15848,N_15153,N_15073);
and U15849 (N_15849,N_15254,N_15528);
and U15850 (N_15850,N_15001,N_15106);
nand U15851 (N_15851,N_15377,N_15244);
nand U15852 (N_15852,N_15487,N_15515);
nand U15853 (N_15853,N_15484,N_15469);
xnor U15854 (N_15854,N_15544,N_15176);
nand U15855 (N_15855,N_15311,N_15279);
or U15856 (N_15856,N_15037,N_15024);
and U15857 (N_15857,N_15428,N_15612);
and U15858 (N_15858,N_15015,N_15474);
nor U15859 (N_15859,N_15602,N_15494);
or U15860 (N_15860,N_15414,N_15080);
nor U15861 (N_15861,N_15120,N_15471);
xor U15862 (N_15862,N_15473,N_15072);
and U15863 (N_15863,N_15353,N_15506);
nor U15864 (N_15864,N_15585,N_15271);
nor U15865 (N_15865,N_15039,N_15615);
xor U15866 (N_15866,N_15481,N_15227);
xor U15867 (N_15867,N_15245,N_15342);
nor U15868 (N_15868,N_15616,N_15499);
or U15869 (N_15869,N_15450,N_15525);
and U15870 (N_15870,N_15339,N_15343);
nand U15871 (N_15871,N_15084,N_15517);
nand U15872 (N_15872,N_15066,N_15094);
xnor U15873 (N_15873,N_15150,N_15104);
nor U15874 (N_15874,N_15151,N_15214);
nor U15875 (N_15875,N_15354,N_15504);
nand U15876 (N_15876,N_15348,N_15095);
or U15877 (N_15877,N_15305,N_15102);
nor U15878 (N_15878,N_15125,N_15005);
xnor U15879 (N_15879,N_15383,N_15046);
nand U15880 (N_15880,N_15452,N_15249);
or U15881 (N_15881,N_15159,N_15395);
xnor U15882 (N_15882,N_15017,N_15229);
or U15883 (N_15883,N_15299,N_15122);
xor U15884 (N_15884,N_15382,N_15405);
and U15885 (N_15885,N_15380,N_15043);
xnor U15886 (N_15886,N_15298,N_15088);
or U15887 (N_15887,N_15124,N_15359);
and U15888 (N_15888,N_15248,N_15316);
nor U15889 (N_15889,N_15431,N_15192);
and U15890 (N_15890,N_15590,N_15379);
and U15891 (N_15891,N_15028,N_15026);
nand U15892 (N_15892,N_15430,N_15357);
xnor U15893 (N_15893,N_15111,N_15552);
and U15894 (N_15894,N_15082,N_15191);
and U15895 (N_15895,N_15236,N_15138);
nor U15896 (N_15896,N_15519,N_15241);
xnor U15897 (N_15897,N_15218,N_15496);
and U15898 (N_15898,N_15173,N_15086);
xor U15899 (N_15899,N_15513,N_15265);
or U15900 (N_15900,N_15034,N_15604);
xnor U15901 (N_15901,N_15155,N_15304);
nor U15902 (N_15902,N_15323,N_15062);
xor U15903 (N_15903,N_15064,N_15476);
and U15904 (N_15904,N_15203,N_15434);
nor U15905 (N_15905,N_15418,N_15603);
nand U15906 (N_15906,N_15297,N_15068);
or U15907 (N_15907,N_15416,N_15322);
nor U15908 (N_15908,N_15127,N_15277);
nand U15909 (N_15909,N_15486,N_15485);
nor U15910 (N_15910,N_15195,N_15458);
nand U15911 (N_15911,N_15136,N_15231);
nand U15912 (N_15912,N_15262,N_15287);
nand U15913 (N_15913,N_15056,N_15356);
nor U15914 (N_15914,N_15090,N_15500);
nand U15915 (N_15915,N_15184,N_15071);
nor U15916 (N_15916,N_15285,N_15534);
or U15917 (N_15917,N_15581,N_15561);
nand U15918 (N_15918,N_15442,N_15251);
and U15919 (N_15919,N_15577,N_15415);
and U15920 (N_15920,N_15167,N_15152);
or U15921 (N_15921,N_15206,N_15455);
and U15922 (N_15922,N_15242,N_15224);
or U15923 (N_15923,N_15196,N_15204);
nand U15924 (N_15924,N_15551,N_15387);
nand U15925 (N_15925,N_15337,N_15293);
nor U15926 (N_15926,N_15135,N_15497);
and U15927 (N_15927,N_15296,N_15376);
nand U15928 (N_15928,N_15445,N_15408);
xnor U15929 (N_15929,N_15148,N_15023);
xor U15930 (N_15930,N_15401,N_15268);
and U15931 (N_15931,N_15035,N_15097);
nand U15932 (N_15932,N_15112,N_15335);
xor U15933 (N_15933,N_15584,N_15291);
nand U15934 (N_15934,N_15461,N_15193);
or U15935 (N_15935,N_15541,N_15099);
or U15936 (N_15936,N_15198,N_15074);
xor U15937 (N_15937,N_15093,N_15604);
xor U15938 (N_15938,N_15389,N_15610);
nand U15939 (N_15939,N_15042,N_15284);
and U15940 (N_15940,N_15330,N_15203);
xor U15941 (N_15941,N_15299,N_15003);
nand U15942 (N_15942,N_15194,N_15310);
xnor U15943 (N_15943,N_15430,N_15112);
and U15944 (N_15944,N_15370,N_15439);
nor U15945 (N_15945,N_15389,N_15605);
xor U15946 (N_15946,N_15519,N_15165);
and U15947 (N_15947,N_15258,N_15059);
or U15948 (N_15948,N_15314,N_15539);
and U15949 (N_15949,N_15311,N_15132);
xor U15950 (N_15950,N_15311,N_15191);
nor U15951 (N_15951,N_15304,N_15195);
nand U15952 (N_15952,N_15048,N_15264);
or U15953 (N_15953,N_15199,N_15018);
or U15954 (N_15954,N_15316,N_15067);
or U15955 (N_15955,N_15615,N_15490);
or U15956 (N_15956,N_15423,N_15361);
nor U15957 (N_15957,N_15523,N_15115);
nor U15958 (N_15958,N_15308,N_15322);
xnor U15959 (N_15959,N_15216,N_15404);
and U15960 (N_15960,N_15231,N_15200);
nand U15961 (N_15961,N_15569,N_15554);
xnor U15962 (N_15962,N_15472,N_15339);
or U15963 (N_15963,N_15084,N_15543);
nor U15964 (N_15964,N_15575,N_15420);
nor U15965 (N_15965,N_15209,N_15003);
and U15966 (N_15966,N_15305,N_15558);
nor U15967 (N_15967,N_15468,N_15120);
nand U15968 (N_15968,N_15266,N_15571);
xor U15969 (N_15969,N_15267,N_15526);
and U15970 (N_15970,N_15495,N_15202);
xor U15971 (N_15971,N_15325,N_15100);
nand U15972 (N_15972,N_15276,N_15587);
or U15973 (N_15973,N_15387,N_15421);
xnor U15974 (N_15974,N_15355,N_15397);
xor U15975 (N_15975,N_15225,N_15490);
nand U15976 (N_15976,N_15020,N_15401);
or U15977 (N_15977,N_15581,N_15407);
and U15978 (N_15978,N_15368,N_15413);
nor U15979 (N_15979,N_15237,N_15475);
nor U15980 (N_15980,N_15468,N_15239);
nand U15981 (N_15981,N_15317,N_15460);
or U15982 (N_15982,N_15561,N_15153);
and U15983 (N_15983,N_15050,N_15232);
nand U15984 (N_15984,N_15441,N_15596);
or U15985 (N_15985,N_15404,N_15609);
xor U15986 (N_15986,N_15227,N_15435);
xor U15987 (N_15987,N_15292,N_15300);
and U15988 (N_15988,N_15574,N_15310);
nor U15989 (N_15989,N_15226,N_15543);
nor U15990 (N_15990,N_15485,N_15211);
and U15991 (N_15991,N_15259,N_15407);
nand U15992 (N_15992,N_15043,N_15187);
or U15993 (N_15993,N_15575,N_15234);
xor U15994 (N_15994,N_15304,N_15224);
or U15995 (N_15995,N_15026,N_15039);
nor U15996 (N_15996,N_15225,N_15497);
nor U15997 (N_15997,N_15039,N_15250);
nor U15998 (N_15998,N_15470,N_15287);
or U15999 (N_15999,N_15461,N_15207);
and U16000 (N_16000,N_15201,N_15370);
and U16001 (N_16001,N_15188,N_15135);
and U16002 (N_16002,N_15123,N_15176);
xnor U16003 (N_16003,N_15177,N_15278);
and U16004 (N_16004,N_15434,N_15345);
or U16005 (N_16005,N_15580,N_15179);
and U16006 (N_16006,N_15395,N_15595);
nand U16007 (N_16007,N_15083,N_15024);
and U16008 (N_16008,N_15282,N_15250);
xor U16009 (N_16009,N_15255,N_15367);
xnor U16010 (N_16010,N_15123,N_15442);
nor U16011 (N_16011,N_15252,N_15557);
nor U16012 (N_16012,N_15136,N_15554);
or U16013 (N_16013,N_15113,N_15251);
nor U16014 (N_16014,N_15096,N_15518);
and U16015 (N_16015,N_15175,N_15458);
xor U16016 (N_16016,N_15087,N_15174);
and U16017 (N_16017,N_15123,N_15515);
or U16018 (N_16018,N_15054,N_15308);
nor U16019 (N_16019,N_15582,N_15240);
or U16020 (N_16020,N_15247,N_15193);
or U16021 (N_16021,N_15426,N_15489);
nand U16022 (N_16022,N_15163,N_15482);
or U16023 (N_16023,N_15420,N_15299);
or U16024 (N_16024,N_15146,N_15151);
nand U16025 (N_16025,N_15318,N_15506);
nand U16026 (N_16026,N_15215,N_15348);
nor U16027 (N_16027,N_15169,N_15520);
xor U16028 (N_16028,N_15562,N_15005);
and U16029 (N_16029,N_15411,N_15149);
and U16030 (N_16030,N_15137,N_15442);
xor U16031 (N_16031,N_15128,N_15580);
xor U16032 (N_16032,N_15601,N_15411);
and U16033 (N_16033,N_15486,N_15377);
or U16034 (N_16034,N_15479,N_15568);
nor U16035 (N_16035,N_15269,N_15155);
xnor U16036 (N_16036,N_15307,N_15242);
nand U16037 (N_16037,N_15442,N_15353);
xnor U16038 (N_16038,N_15454,N_15567);
nand U16039 (N_16039,N_15403,N_15353);
xor U16040 (N_16040,N_15407,N_15226);
and U16041 (N_16041,N_15367,N_15307);
and U16042 (N_16042,N_15131,N_15305);
and U16043 (N_16043,N_15518,N_15353);
and U16044 (N_16044,N_15192,N_15153);
and U16045 (N_16045,N_15072,N_15272);
nand U16046 (N_16046,N_15442,N_15403);
and U16047 (N_16047,N_15134,N_15435);
or U16048 (N_16048,N_15516,N_15007);
and U16049 (N_16049,N_15017,N_15053);
xor U16050 (N_16050,N_15107,N_15163);
or U16051 (N_16051,N_15178,N_15486);
or U16052 (N_16052,N_15362,N_15095);
nand U16053 (N_16053,N_15001,N_15339);
and U16054 (N_16054,N_15103,N_15207);
xor U16055 (N_16055,N_15174,N_15555);
xor U16056 (N_16056,N_15283,N_15489);
nand U16057 (N_16057,N_15059,N_15140);
nor U16058 (N_16058,N_15029,N_15165);
or U16059 (N_16059,N_15204,N_15424);
and U16060 (N_16060,N_15472,N_15191);
and U16061 (N_16061,N_15255,N_15574);
nor U16062 (N_16062,N_15432,N_15521);
nor U16063 (N_16063,N_15124,N_15295);
nor U16064 (N_16064,N_15046,N_15288);
or U16065 (N_16065,N_15408,N_15174);
xnor U16066 (N_16066,N_15135,N_15548);
and U16067 (N_16067,N_15256,N_15507);
nand U16068 (N_16068,N_15561,N_15054);
or U16069 (N_16069,N_15204,N_15065);
nand U16070 (N_16070,N_15247,N_15522);
and U16071 (N_16071,N_15580,N_15473);
nand U16072 (N_16072,N_15564,N_15520);
and U16073 (N_16073,N_15588,N_15379);
xor U16074 (N_16074,N_15013,N_15166);
xnor U16075 (N_16075,N_15063,N_15372);
xor U16076 (N_16076,N_15031,N_15467);
nand U16077 (N_16077,N_15330,N_15016);
nand U16078 (N_16078,N_15402,N_15415);
nor U16079 (N_16079,N_15110,N_15586);
nor U16080 (N_16080,N_15502,N_15246);
nand U16081 (N_16081,N_15619,N_15020);
or U16082 (N_16082,N_15528,N_15320);
and U16083 (N_16083,N_15381,N_15437);
or U16084 (N_16084,N_15581,N_15431);
and U16085 (N_16085,N_15365,N_15222);
and U16086 (N_16086,N_15090,N_15418);
nor U16087 (N_16087,N_15308,N_15301);
nand U16088 (N_16088,N_15269,N_15305);
or U16089 (N_16089,N_15384,N_15154);
xnor U16090 (N_16090,N_15115,N_15321);
xor U16091 (N_16091,N_15417,N_15056);
nand U16092 (N_16092,N_15510,N_15174);
or U16093 (N_16093,N_15352,N_15417);
xnor U16094 (N_16094,N_15223,N_15240);
xor U16095 (N_16095,N_15083,N_15360);
or U16096 (N_16096,N_15624,N_15416);
and U16097 (N_16097,N_15191,N_15151);
xor U16098 (N_16098,N_15471,N_15404);
nand U16099 (N_16099,N_15417,N_15147);
and U16100 (N_16100,N_15238,N_15602);
xnor U16101 (N_16101,N_15521,N_15418);
or U16102 (N_16102,N_15325,N_15126);
xnor U16103 (N_16103,N_15577,N_15189);
nor U16104 (N_16104,N_15100,N_15022);
nand U16105 (N_16105,N_15363,N_15228);
nor U16106 (N_16106,N_15437,N_15060);
xnor U16107 (N_16107,N_15277,N_15106);
xnor U16108 (N_16108,N_15531,N_15472);
or U16109 (N_16109,N_15393,N_15536);
nand U16110 (N_16110,N_15042,N_15168);
and U16111 (N_16111,N_15426,N_15091);
and U16112 (N_16112,N_15049,N_15600);
nor U16113 (N_16113,N_15364,N_15582);
and U16114 (N_16114,N_15262,N_15417);
and U16115 (N_16115,N_15407,N_15595);
nor U16116 (N_16116,N_15551,N_15243);
nor U16117 (N_16117,N_15020,N_15428);
nor U16118 (N_16118,N_15438,N_15340);
nand U16119 (N_16119,N_15305,N_15006);
and U16120 (N_16120,N_15411,N_15511);
nor U16121 (N_16121,N_15127,N_15089);
and U16122 (N_16122,N_15103,N_15419);
and U16123 (N_16123,N_15042,N_15364);
nand U16124 (N_16124,N_15369,N_15429);
and U16125 (N_16125,N_15241,N_15369);
nand U16126 (N_16126,N_15559,N_15143);
xnor U16127 (N_16127,N_15185,N_15336);
and U16128 (N_16128,N_15068,N_15528);
nor U16129 (N_16129,N_15318,N_15251);
nand U16130 (N_16130,N_15595,N_15284);
nor U16131 (N_16131,N_15196,N_15316);
or U16132 (N_16132,N_15577,N_15518);
nor U16133 (N_16133,N_15439,N_15452);
xor U16134 (N_16134,N_15389,N_15565);
xnor U16135 (N_16135,N_15398,N_15421);
xnor U16136 (N_16136,N_15322,N_15035);
xnor U16137 (N_16137,N_15271,N_15145);
xnor U16138 (N_16138,N_15096,N_15380);
or U16139 (N_16139,N_15116,N_15061);
xor U16140 (N_16140,N_15383,N_15367);
nand U16141 (N_16141,N_15504,N_15524);
and U16142 (N_16142,N_15276,N_15107);
and U16143 (N_16143,N_15033,N_15173);
nand U16144 (N_16144,N_15352,N_15474);
xor U16145 (N_16145,N_15502,N_15489);
and U16146 (N_16146,N_15378,N_15396);
nor U16147 (N_16147,N_15580,N_15166);
nand U16148 (N_16148,N_15083,N_15267);
or U16149 (N_16149,N_15517,N_15293);
and U16150 (N_16150,N_15166,N_15594);
nor U16151 (N_16151,N_15265,N_15249);
and U16152 (N_16152,N_15351,N_15055);
nand U16153 (N_16153,N_15020,N_15056);
nor U16154 (N_16154,N_15135,N_15078);
and U16155 (N_16155,N_15276,N_15325);
or U16156 (N_16156,N_15072,N_15202);
nor U16157 (N_16157,N_15031,N_15624);
or U16158 (N_16158,N_15274,N_15579);
or U16159 (N_16159,N_15090,N_15383);
or U16160 (N_16160,N_15381,N_15559);
xnor U16161 (N_16161,N_15243,N_15602);
nor U16162 (N_16162,N_15513,N_15539);
nand U16163 (N_16163,N_15436,N_15213);
nand U16164 (N_16164,N_15322,N_15481);
nor U16165 (N_16165,N_15180,N_15562);
xnor U16166 (N_16166,N_15190,N_15362);
or U16167 (N_16167,N_15057,N_15249);
nor U16168 (N_16168,N_15006,N_15000);
and U16169 (N_16169,N_15402,N_15333);
xor U16170 (N_16170,N_15479,N_15201);
or U16171 (N_16171,N_15601,N_15308);
and U16172 (N_16172,N_15008,N_15174);
and U16173 (N_16173,N_15127,N_15514);
and U16174 (N_16174,N_15204,N_15369);
nand U16175 (N_16175,N_15393,N_15047);
or U16176 (N_16176,N_15041,N_15252);
and U16177 (N_16177,N_15250,N_15323);
or U16178 (N_16178,N_15202,N_15090);
xnor U16179 (N_16179,N_15480,N_15151);
xnor U16180 (N_16180,N_15547,N_15419);
nand U16181 (N_16181,N_15404,N_15493);
nor U16182 (N_16182,N_15013,N_15535);
nor U16183 (N_16183,N_15140,N_15381);
and U16184 (N_16184,N_15283,N_15296);
nand U16185 (N_16185,N_15098,N_15398);
nand U16186 (N_16186,N_15113,N_15152);
xnor U16187 (N_16187,N_15145,N_15297);
or U16188 (N_16188,N_15176,N_15060);
and U16189 (N_16189,N_15254,N_15118);
nor U16190 (N_16190,N_15587,N_15430);
xnor U16191 (N_16191,N_15601,N_15584);
nor U16192 (N_16192,N_15257,N_15104);
xor U16193 (N_16193,N_15614,N_15141);
xnor U16194 (N_16194,N_15095,N_15215);
nand U16195 (N_16195,N_15005,N_15156);
and U16196 (N_16196,N_15218,N_15254);
xor U16197 (N_16197,N_15472,N_15582);
xor U16198 (N_16198,N_15155,N_15358);
nand U16199 (N_16199,N_15208,N_15095);
nand U16200 (N_16200,N_15124,N_15106);
and U16201 (N_16201,N_15046,N_15031);
and U16202 (N_16202,N_15150,N_15377);
nand U16203 (N_16203,N_15229,N_15282);
nand U16204 (N_16204,N_15226,N_15175);
or U16205 (N_16205,N_15239,N_15473);
or U16206 (N_16206,N_15504,N_15237);
xnor U16207 (N_16207,N_15199,N_15527);
and U16208 (N_16208,N_15364,N_15493);
or U16209 (N_16209,N_15053,N_15393);
nand U16210 (N_16210,N_15055,N_15096);
and U16211 (N_16211,N_15413,N_15372);
nand U16212 (N_16212,N_15131,N_15537);
or U16213 (N_16213,N_15086,N_15541);
nand U16214 (N_16214,N_15236,N_15081);
nand U16215 (N_16215,N_15167,N_15374);
xor U16216 (N_16216,N_15450,N_15617);
or U16217 (N_16217,N_15316,N_15235);
and U16218 (N_16218,N_15126,N_15180);
xnor U16219 (N_16219,N_15034,N_15085);
xnor U16220 (N_16220,N_15007,N_15082);
nand U16221 (N_16221,N_15516,N_15164);
and U16222 (N_16222,N_15189,N_15378);
xor U16223 (N_16223,N_15495,N_15061);
or U16224 (N_16224,N_15310,N_15460);
nand U16225 (N_16225,N_15446,N_15160);
nand U16226 (N_16226,N_15294,N_15478);
or U16227 (N_16227,N_15557,N_15180);
and U16228 (N_16228,N_15302,N_15394);
xnor U16229 (N_16229,N_15357,N_15159);
and U16230 (N_16230,N_15333,N_15080);
nor U16231 (N_16231,N_15411,N_15145);
nor U16232 (N_16232,N_15217,N_15387);
or U16233 (N_16233,N_15129,N_15410);
and U16234 (N_16234,N_15124,N_15340);
or U16235 (N_16235,N_15413,N_15387);
xnor U16236 (N_16236,N_15561,N_15291);
and U16237 (N_16237,N_15472,N_15019);
and U16238 (N_16238,N_15473,N_15249);
and U16239 (N_16239,N_15258,N_15072);
nand U16240 (N_16240,N_15021,N_15411);
nor U16241 (N_16241,N_15553,N_15604);
xor U16242 (N_16242,N_15080,N_15348);
and U16243 (N_16243,N_15353,N_15515);
nor U16244 (N_16244,N_15262,N_15248);
and U16245 (N_16245,N_15184,N_15605);
or U16246 (N_16246,N_15044,N_15439);
xor U16247 (N_16247,N_15143,N_15072);
or U16248 (N_16248,N_15558,N_15490);
and U16249 (N_16249,N_15222,N_15072);
or U16250 (N_16250,N_16246,N_16108);
xor U16251 (N_16251,N_15847,N_16040);
or U16252 (N_16252,N_16195,N_15689);
xor U16253 (N_16253,N_15661,N_15741);
nor U16254 (N_16254,N_16215,N_16048);
and U16255 (N_16255,N_15869,N_15817);
nand U16256 (N_16256,N_15764,N_15800);
nand U16257 (N_16257,N_15819,N_15825);
nand U16258 (N_16258,N_16103,N_15791);
or U16259 (N_16259,N_15796,N_16110);
xnor U16260 (N_16260,N_15953,N_15842);
nand U16261 (N_16261,N_15839,N_16087);
xnor U16262 (N_16262,N_16165,N_15650);
nor U16263 (N_16263,N_15743,N_15895);
nor U16264 (N_16264,N_15705,N_16141);
xnor U16265 (N_16265,N_16187,N_16129);
nor U16266 (N_16266,N_16027,N_16009);
xor U16267 (N_16267,N_15632,N_15754);
nand U16268 (N_16268,N_15722,N_15983);
or U16269 (N_16269,N_15643,N_16095);
or U16270 (N_16270,N_15836,N_16072);
or U16271 (N_16271,N_16153,N_15674);
nor U16272 (N_16272,N_16163,N_16014);
or U16273 (N_16273,N_15845,N_15816);
nand U16274 (N_16274,N_15980,N_15948);
xnor U16275 (N_16275,N_16006,N_16058);
nor U16276 (N_16276,N_15725,N_15659);
nor U16277 (N_16277,N_15849,N_15850);
nor U16278 (N_16278,N_16241,N_16065);
or U16279 (N_16279,N_15731,N_15959);
and U16280 (N_16280,N_15843,N_15729);
and U16281 (N_16281,N_16075,N_15846);
or U16282 (N_16282,N_15943,N_16081);
nand U16283 (N_16283,N_15631,N_16015);
and U16284 (N_16284,N_16212,N_15768);
xor U16285 (N_16285,N_15781,N_16231);
nor U16286 (N_16286,N_15734,N_16148);
nor U16287 (N_16287,N_15914,N_16074);
or U16288 (N_16288,N_16184,N_15930);
or U16289 (N_16289,N_16094,N_15804);
nor U16290 (N_16290,N_15883,N_15999);
or U16291 (N_16291,N_16042,N_16107);
nand U16292 (N_16292,N_16076,N_15958);
nor U16293 (N_16293,N_15657,N_15864);
xor U16294 (N_16294,N_16023,N_16104);
or U16295 (N_16295,N_15684,N_15831);
and U16296 (N_16296,N_16240,N_16209);
and U16297 (N_16297,N_15759,N_15991);
xor U16298 (N_16298,N_15784,N_15704);
nor U16299 (N_16299,N_16106,N_16233);
nor U16300 (N_16300,N_15848,N_15637);
nor U16301 (N_16301,N_15712,N_16125);
or U16302 (N_16302,N_15979,N_15665);
xor U16303 (N_16303,N_15949,N_15968);
and U16304 (N_16304,N_15899,N_15802);
nor U16305 (N_16305,N_15931,N_15870);
nor U16306 (N_16306,N_15940,N_15862);
nand U16307 (N_16307,N_16071,N_16045);
and U16308 (N_16308,N_16002,N_15830);
xor U16309 (N_16309,N_15765,N_16057);
nand U16310 (N_16310,N_16208,N_15746);
or U16311 (N_16311,N_16176,N_15717);
or U16312 (N_16312,N_15801,N_15651);
or U16313 (N_16313,N_15767,N_15710);
or U16314 (N_16314,N_16008,N_16211);
or U16315 (N_16315,N_15766,N_15866);
xor U16316 (N_16316,N_16235,N_16224);
and U16317 (N_16317,N_15779,N_15835);
or U16318 (N_16318,N_16016,N_15805);
nor U16319 (N_16319,N_16080,N_16068);
nand U16320 (N_16320,N_16193,N_15673);
nand U16321 (N_16321,N_15906,N_15871);
or U16322 (N_16322,N_15957,N_16144);
and U16323 (N_16323,N_15737,N_15880);
nor U16324 (N_16324,N_15910,N_15857);
or U16325 (N_16325,N_16160,N_15660);
or U16326 (N_16326,N_15723,N_15955);
and U16327 (N_16327,N_15820,N_15882);
xor U16328 (N_16328,N_16205,N_16177);
nand U16329 (N_16329,N_15769,N_16118);
or U16330 (N_16330,N_15993,N_16122);
or U16331 (N_16331,N_15989,N_15954);
xor U16332 (N_16332,N_16194,N_16063);
nand U16333 (N_16333,N_15709,N_15797);
nand U16334 (N_16334,N_15821,N_15966);
and U16335 (N_16335,N_15916,N_15985);
nor U16336 (N_16336,N_15942,N_16159);
nor U16337 (N_16337,N_16239,N_15923);
nor U16338 (N_16338,N_15788,N_15630);
xnor U16339 (N_16339,N_15655,N_16003);
nand U16340 (N_16340,N_15828,N_15860);
xor U16341 (N_16341,N_15858,N_15794);
xor U16342 (N_16342,N_15834,N_16025);
nand U16343 (N_16343,N_15833,N_16226);
and U16344 (N_16344,N_15720,N_15711);
nand U16345 (N_16345,N_16225,N_15981);
nor U16346 (N_16346,N_16112,N_15738);
or U16347 (N_16347,N_15898,N_16090);
nand U16348 (N_16348,N_15702,N_16079);
or U16349 (N_16349,N_15918,N_15971);
nand U16350 (N_16350,N_15874,N_15680);
xor U16351 (N_16351,N_15907,N_16117);
nand U16352 (N_16352,N_15822,N_15676);
or U16353 (N_16353,N_15811,N_16030);
nand U16354 (N_16354,N_16020,N_15771);
or U16355 (N_16355,N_15787,N_16183);
xor U16356 (N_16356,N_15658,N_16060);
nand U16357 (N_16357,N_15698,N_16073);
or U16358 (N_16358,N_15855,N_15678);
nor U16359 (N_16359,N_16032,N_15877);
xor U16360 (N_16360,N_15716,N_15947);
and U16361 (N_16361,N_15629,N_15750);
and U16362 (N_16362,N_15917,N_16138);
nor U16363 (N_16363,N_16085,N_16132);
nand U16364 (N_16364,N_16078,N_15903);
or U16365 (N_16365,N_16036,N_15932);
and U16366 (N_16366,N_15925,N_15776);
nor U16367 (N_16367,N_16244,N_15688);
nor U16368 (N_16368,N_15886,N_16067);
and U16369 (N_16369,N_16134,N_15964);
xnor U16370 (N_16370,N_16230,N_15675);
nor U16371 (N_16371,N_15793,N_15815);
or U16372 (N_16372,N_15946,N_15915);
nand U16373 (N_16373,N_16082,N_15854);
or U16374 (N_16374,N_15736,N_15703);
or U16375 (N_16375,N_16083,N_16221);
xor U16376 (N_16376,N_15856,N_15863);
or U16377 (N_16377,N_16242,N_16105);
xnor U16378 (N_16378,N_16156,N_15721);
xor U16379 (N_16379,N_15708,N_16001);
nor U16380 (N_16380,N_15975,N_16100);
nand U16381 (N_16381,N_15978,N_15992);
xor U16382 (N_16382,N_16007,N_16114);
or U16383 (N_16383,N_15639,N_15653);
xor U16384 (N_16384,N_15982,N_16228);
or U16385 (N_16385,N_15691,N_16111);
or U16386 (N_16386,N_15945,N_16054);
xor U16387 (N_16387,N_15837,N_16140);
nor U16388 (N_16388,N_16031,N_15645);
xnor U16389 (N_16389,N_16227,N_15933);
xnor U16390 (N_16390,N_15818,N_15640);
and U16391 (N_16391,N_16180,N_15666);
or U16392 (N_16392,N_16084,N_16147);
nor U16393 (N_16393,N_15715,N_16202);
and U16394 (N_16394,N_15777,N_15697);
nand U16395 (N_16395,N_16029,N_15726);
and U16396 (N_16396,N_15668,N_16102);
xnor U16397 (N_16397,N_15696,N_15881);
nor U16398 (N_16398,N_16167,N_15662);
nand U16399 (N_16399,N_16249,N_15841);
or U16400 (N_16400,N_15900,N_15969);
xnor U16401 (N_16401,N_16052,N_16070);
and U16402 (N_16402,N_16088,N_15913);
xnor U16403 (N_16403,N_15656,N_15664);
nor U16404 (N_16404,N_15799,N_16200);
nand U16405 (N_16405,N_15713,N_15692);
nor U16406 (N_16406,N_16237,N_15681);
and U16407 (N_16407,N_16017,N_15924);
nand U16408 (N_16408,N_15896,N_15757);
or U16409 (N_16409,N_15685,N_15865);
nor U16410 (N_16410,N_16028,N_15648);
nor U16411 (N_16411,N_15634,N_15908);
or U16412 (N_16412,N_15770,N_15827);
nor U16413 (N_16413,N_16019,N_16039);
or U16414 (N_16414,N_16203,N_15707);
and U16415 (N_16415,N_15967,N_16044);
nor U16416 (N_16416,N_16086,N_15751);
nor U16417 (N_16417,N_15937,N_16005);
and U16418 (N_16418,N_16201,N_15778);
xor U16419 (N_16419,N_15625,N_15838);
nor U16420 (N_16420,N_15956,N_15944);
nand U16421 (N_16421,N_15927,N_15986);
xor U16422 (N_16422,N_16043,N_16155);
nand U16423 (N_16423,N_15739,N_15928);
or U16424 (N_16424,N_15683,N_16116);
xor U16425 (N_16425,N_16055,N_15667);
and U16426 (N_16426,N_16164,N_15939);
nor U16427 (N_16427,N_15994,N_15852);
and U16428 (N_16428,N_15627,N_15642);
or U16429 (N_16429,N_15965,N_16053);
xnor U16430 (N_16430,N_15829,N_15891);
xor U16431 (N_16431,N_16022,N_15761);
nand U16432 (N_16432,N_15961,N_15844);
and U16433 (N_16433,N_16247,N_15744);
nor U16434 (N_16434,N_15868,N_16109);
xnor U16435 (N_16435,N_15654,N_15652);
xnor U16436 (N_16436,N_16050,N_16124);
nand U16437 (N_16437,N_15694,N_15693);
nand U16438 (N_16438,N_16185,N_16064);
xor U16439 (N_16439,N_15878,N_15887);
nor U16440 (N_16440,N_15687,N_16161);
nand U16441 (N_16441,N_15872,N_15789);
or U16442 (N_16442,N_15941,N_16168);
xnor U16443 (N_16443,N_16190,N_16131);
and U16444 (N_16444,N_16169,N_15775);
nand U16445 (N_16445,N_16136,N_16013);
nor U16446 (N_16446,N_16216,N_16232);
or U16447 (N_16447,N_15889,N_16097);
xnor U16448 (N_16448,N_16222,N_16145);
nand U16449 (N_16449,N_15879,N_15774);
or U16450 (N_16450,N_15984,N_15671);
nand U16451 (N_16451,N_16018,N_15669);
nand U16452 (N_16452,N_16098,N_16192);
and U16453 (N_16453,N_16171,N_16004);
nor U16454 (N_16454,N_15686,N_15748);
xnor U16455 (N_16455,N_15792,N_15960);
xnor U16456 (N_16456,N_15756,N_16234);
and U16457 (N_16457,N_16077,N_15682);
nor U16458 (N_16458,N_16198,N_15990);
nor U16459 (N_16459,N_16170,N_16038);
nand U16460 (N_16460,N_15803,N_15859);
and U16461 (N_16461,N_15772,N_15890);
nand U16462 (N_16462,N_15644,N_15635);
nor U16463 (N_16463,N_15782,N_15763);
and U16464 (N_16464,N_15998,N_15884);
and U16465 (N_16465,N_15695,N_15780);
and U16466 (N_16466,N_16223,N_15892);
and U16467 (N_16467,N_16149,N_15783);
and U16468 (N_16468,N_15876,N_15851);
nand U16469 (N_16469,N_15626,N_16173);
nor U16470 (N_16470,N_15718,N_15745);
or U16471 (N_16471,N_15976,N_16069);
or U16472 (N_16472,N_15790,N_15952);
nor U16473 (N_16473,N_16172,N_15824);
nand U16474 (N_16474,N_15996,N_16120);
or U16475 (N_16475,N_16062,N_15912);
nand U16476 (N_16476,N_16047,N_16126);
xnor U16477 (N_16477,N_15742,N_15638);
nand U16478 (N_16478,N_15911,N_16158);
nand U16479 (N_16479,N_16012,N_16174);
or U16480 (N_16480,N_16000,N_15646);
nand U16481 (N_16481,N_16142,N_15809);
and U16482 (N_16482,N_15970,N_15755);
or U16483 (N_16483,N_16096,N_16181);
or U16484 (N_16484,N_15810,N_16139);
or U16485 (N_16485,N_16146,N_15901);
and U16486 (N_16486,N_15875,N_15706);
or U16487 (N_16487,N_16189,N_15728);
xnor U16488 (N_16488,N_16123,N_15919);
nor U16489 (N_16489,N_15735,N_15786);
xnor U16490 (N_16490,N_15840,N_16207);
xor U16491 (N_16491,N_15988,N_16220);
and U16492 (N_16492,N_15987,N_15773);
xnor U16493 (N_16493,N_15758,N_16011);
or U16494 (N_16494,N_16204,N_15647);
nor U16495 (N_16495,N_16214,N_15853);
xor U16496 (N_16496,N_15808,N_16197);
nor U16497 (N_16497,N_16137,N_15813);
nand U16498 (N_16498,N_15740,N_15893);
or U16499 (N_16499,N_16059,N_16101);
or U16500 (N_16500,N_15641,N_15873);
and U16501 (N_16501,N_16037,N_16061);
or U16502 (N_16502,N_15867,N_16099);
and U16503 (N_16503,N_15905,N_16026);
nand U16504 (N_16504,N_16121,N_16179);
or U16505 (N_16505,N_15663,N_16046);
and U16506 (N_16506,N_16093,N_16182);
and U16507 (N_16507,N_16162,N_16135);
or U16508 (N_16508,N_16178,N_16119);
nand U16509 (N_16509,N_16245,N_15785);
nor U16510 (N_16510,N_15938,N_15700);
nand U16511 (N_16511,N_16188,N_16033);
and U16512 (N_16512,N_15894,N_15814);
or U16513 (N_16513,N_15935,N_16217);
nand U16514 (N_16514,N_15861,N_15973);
xnor U16515 (N_16515,N_16219,N_16248);
nor U16516 (N_16516,N_15730,N_16066);
or U16517 (N_16517,N_16151,N_15727);
or U16518 (N_16518,N_15732,N_16154);
and U16519 (N_16519,N_16089,N_16152);
nand U16520 (N_16520,N_15690,N_16133);
and U16521 (N_16521,N_15950,N_16034);
nand U16522 (N_16522,N_16035,N_15926);
or U16523 (N_16523,N_15922,N_16127);
nand U16524 (N_16524,N_15762,N_15752);
xnor U16525 (N_16525,N_15963,N_16128);
and U16526 (N_16526,N_15714,N_16213);
or U16527 (N_16527,N_16092,N_15672);
nand U16528 (N_16528,N_16130,N_16196);
and U16529 (N_16529,N_15628,N_16157);
or U16530 (N_16530,N_15972,N_16199);
nand U16531 (N_16531,N_15724,N_15753);
nand U16532 (N_16532,N_16218,N_16206);
nand U16533 (N_16533,N_15997,N_15951);
or U16534 (N_16534,N_15812,N_16238);
and U16535 (N_16535,N_15888,N_15902);
nand U16536 (N_16536,N_16051,N_16115);
xor U16537 (N_16537,N_15677,N_15929);
nand U16538 (N_16538,N_15921,N_16186);
and U16539 (N_16539,N_15806,N_16024);
or U16540 (N_16540,N_16243,N_16010);
nand U16541 (N_16541,N_15909,N_15807);
or U16542 (N_16542,N_15649,N_15934);
xor U16543 (N_16543,N_16056,N_16041);
or U16544 (N_16544,N_15733,N_15798);
nor U16545 (N_16545,N_16049,N_15670);
nand U16546 (N_16546,N_15904,N_15760);
xnor U16547 (N_16547,N_15974,N_15936);
and U16548 (N_16548,N_15832,N_16229);
and U16549 (N_16549,N_15747,N_15679);
nor U16550 (N_16550,N_15995,N_16143);
nand U16551 (N_16551,N_15885,N_15823);
nand U16552 (N_16552,N_16210,N_16175);
xor U16553 (N_16553,N_15636,N_15749);
nor U16554 (N_16554,N_16150,N_15977);
nor U16555 (N_16555,N_16166,N_16236);
nand U16556 (N_16556,N_15897,N_15920);
or U16557 (N_16557,N_16113,N_15701);
or U16558 (N_16558,N_16021,N_16191);
or U16559 (N_16559,N_15699,N_16091);
xor U16560 (N_16560,N_15826,N_15962);
xor U16561 (N_16561,N_15795,N_15633);
and U16562 (N_16562,N_15719,N_16154);
xnor U16563 (N_16563,N_16192,N_16114);
nor U16564 (N_16564,N_16052,N_16003);
nand U16565 (N_16565,N_15988,N_15937);
or U16566 (N_16566,N_15705,N_15699);
nor U16567 (N_16567,N_15813,N_15838);
nor U16568 (N_16568,N_15703,N_16102);
nand U16569 (N_16569,N_15769,N_15841);
and U16570 (N_16570,N_15912,N_15723);
xnor U16571 (N_16571,N_15999,N_15654);
nor U16572 (N_16572,N_16136,N_15978);
nor U16573 (N_16573,N_15783,N_15814);
or U16574 (N_16574,N_15717,N_16142);
or U16575 (N_16575,N_15867,N_15635);
and U16576 (N_16576,N_16072,N_15807);
nor U16577 (N_16577,N_15729,N_15672);
nor U16578 (N_16578,N_16233,N_15687);
xnor U16579 (N_16579,N_15808,N_15849);
and U16580 (N_16580,N_16212,N_16180);
or U16581 (N_16581,N_15771,N_15797);
or U16582 (N_16582,N_16098,N_16142);
and U16583 (N_16583,N_15985,N_16066);
nor U16584 (N_16584,N_15640,N_15895);
xnor U16585 (N_16585,N_15678,N_16112);
nand U16586 (N_16586,N_15866,N_15911);
and U16587 (N_16587,N_16097,N_16232);
nand U16588 (N_16588,N_15795,N_16091);
nand U16589 (N_16589,N_16216,N_15684);
nor U16590 (N_16590,N_16045,N_15733);
nor U16591 (N_16591,N_15684,N_15919);
and U16592 (N_16592,N_15983,N_15918);
and U16593 (N_16593,N_16160,N_15798);
xor U16594 (N_16594,N_15780,N_15799);
xor U16595 (N_16595,N_15783,N_15642);
or U16596 (N_16596,N_15865,N_16117);
nand U16597 (N_16597,N_15842,N_16022);
and U16598 (N_16598,N_16115,N_15667);
nand U16599 (N_16599,N_15688,N_15796);
xor U16600 (N_16600,N_15910,N_16016);
xnor U16601 (N_16601,N_15884,N_16166);
nand U16602 (N_16602,N_15881,N_15931);
nor U16603 (N_16603,N_15900,N_15651);
xnor U16604 (N_16604,N_16180,N_15794);
nand U16605 (N_16605,N_15890,N_15963);
and U16606 (N_16606,N_15896,N_16151);
or U16607 (N_16607,N_15959,N_16106);
nor U16608 (N_16608,N_15652,N_16021);
and U16609 (N_16609,N_16122,N_15782);
nand U16610 (N_16610,N_15770,N_15758);
nand U16611 (N_16611,N_16126,N_15741);
nor U16612 (N_16612,N_16192,N_15878);
xnor U16613 (N_16613,N_16137,N_16164);
nand U16614 (N_16614,N_15977,N_16156);
and U16615 (N_16615,N_15836,N_16212);
or U16616 (N_16616,N_15676,N_16194);
nand U16617 (N_16617,N_15992,N_15635);
xnor U16618 (N_16618,N_15977,N_15918);
xor U16619 (N_16619,N_16205,N_15687);
nand U16620 (N_16620,N_15738,N_15958);
nor U16621 (N_16621,N_16245,N_15859);
or U16622 (N_16622,N_16058,N_15702);
or U16623 (N_16623,N_15817,N_15845);
and U16624 (N_16624,N_16068,N_16021);
xor U16625 (N_16625,N_15754,N_15637);
and U16626 (N_16626,N_16198,N_16035);
and U16627 (N_16627,N_15985,N_15718);
or U16628 (N_16628,N_15978,N_16060);
and U16629 (N_16629,N_15646,N_16215);
xnor U16630 (N_16630,N_16157,N_16186);
and U16631 (N_16631,N_15647,N_15992);
and U16632 (N_16632,N_15945,N_15839);
nand U16633 (N_16633,N_15851,N_15701);
nor U16634 (N_16634,N_15743,N_16154);
xor U16635 (N_16635,N_15654,N_15758);
nor U16636 (N_16636,N_15705,N_15683);
xnor U16637 (N_16637,N_15910,N_15637);
or U16638 (N_16638,N_15714,N_15807);
and U16639 (N_16639,N_16125,N_16231);
nor U16640 (N_16640,N_16036,N_15816);
xor U16641 (N_16641,N_15973,N_15955);
nor U16642 (N_16642,N_16148,N_15952);
or U16643 (N_16643,N_15822,N_15783);
nand U16644 (N_16644,N_16164,N_16185);
or U16645 (N_16645,N_15665,N_15805);
nand U16646 (N_16646,N_15645,N_16198);
and U16647 (N_16647,N_15981,N_15698);
or U16648 (N_16648,N_15625,N_15654);
nand U16649 (N_16649,N_16226,N_15721);
nand U16650 (N_16650,N_16063,N_15925);
nor U16651 (N_16651,N_15773,N_15902);
xor U16652 (N_16652,N_16229,N_15750);
xor U16653 (N_16653,N_16132,N_16026);
nand U16654 (N_16654,N_15626,N_16245);
nand U16655 (N_16655,N_16095,N_15928);
and U16656 (N_16656,N_16238,N_15847);
nor U16657 (N_16657,N_15707,N_15925);
or U16658 (N_16658,N_15970,N_16145);
nor U16659 (N_16659,N_15738,N_15740);
or U16660 (N_16660,N_15826,N_15782);
or U16661 (N_16661,N_15890,N_15751);
or U16662 (N_16662,N_15658,N_16246);
or U16663 (N_16663,N_15763,N_15647);
or U16664 (N_16664,N_15659,N_15877);
nor U16665 (N_16665,N_15974,N_15832);
and U16666 (N_16666,N_15728,N_16220);
nor U16667 (N_16667,N_16049,N_15871);
and U16668 (N_16668,N_16191,N_15940);
xnor U16669 (N_16669,N_15885,N_15888);
xor U16670 (N_16670,N_15727,N_16095);
and U16671 (N_16671,N_15996,N_15681);
nor U16672 (N_16672,N_15824,N_16108);
and U16673 (N_16673,N_15766,N_15988);
nor U16674 (N_16674,N_16136,N_15934);
nor U16675 (N_16675,N_15698,N_15960);
nor U16676 (N_16676,N_16161,N_16175);
and U16677 (N_16677,N_15913,N_15734);
or U16678 (N_16678,N_15812,N_15941);
nand U16679 (N_16679,N_15924,N_15827);
nand U16680 (N_16680,N_15856,N_16077);
nor U16681 (N_16681,N_15903,N_15770);
xnor U16682 (N_16682,N_15910,N_15758);
or U16683 (N_16683,N_15836,N_15849);
xor U16684 (N_16684,N_15661,N_15715);
nand U16685 (N_16685,N_16036,N_15796);
or U16686 (N_16686,N_15931,N_15670);
and U16687 (N_16687,N_16221,N_16019);
xnor U16688 (N_16688,N_15871,N_15851);
and U16689 (N_16689,N_16006,N_15982);
nor U16690 (N_16690,N_15764,N_15973);
nand U16691 (N_16691,N_16008,N_15982);
or U16692 (N_16692,N_15668,N_16009);
and U16693 (N_16693,N_16152,N_15655);
or U16694 (N_16694,N_15717,N_15693);
or U16695 (N_16695,N_16005,N_15646);
nor U16696 (N_16696,N_15755,N_15866);
and U16697 (N_16697,N_15739,N_16039);
nand U16698 (N_16698,N_16234,N_16058);
or U16699 (N_16699,N_15888,N_15720);
xor U16700 (N_16700,N_15865,N_16083);
xor U16701 (N_16701,N_15676,N_15686);
nand U16702 (N_16702,N_15925,N_16206);
nand U16703 (N_16703,N_16194,N_15748);
nand U16704 (N_16704,N_15916,N_16049);
nor U16705 (N_16705,N_16173,N_15629);
nor U16706 (N_16706,N_15955,N_15913);
nand U16707 (N_16707,N_15970,N_15657);
and U16708 (N_16708,N_16060,N_15805);
or U16709 (N_16709,N_16125,N_15928);
and U16710 (N_16710,N_15639,N_15943);
and U16711 (N_16711,N_16009,N_15711);
and U16712 (N_16712,N_15668,N_15686);
and U16713 (N_16713,N_15876,N_15924);
or U16714 (N_16714,N_15871,N_16180);
and U16715 (N_16715,N_15883,N_15804);
nand U16716 (N_16716,N_15933,N_16098);
or U16717 (N_16717,N_16077,N_15772);
and U16718 (N_16718,N_16205,N_15926);
nand U16719 (N_16719,N_15671,N_16155);
xor U16720 (N_16720,N_15771,N_15862);
nor U16721 (N_16721,N_15625,N_15729);
xnor U16722 (N_16722,N_15741,N_16125);
nand U16723 (N_16723,N_15646,N_15995);
xor U16724 (N_16724,N_16028,N_15830);
nor U16725 (N_16725,N_15669,N_15809);
or U16726 (N_16726,N_15774,N_15657);
or U16727 (N_16727,N_16065,N_15693);
and U16728 (N_16728,N_15935,N_16214);
or U16729 (N_16729,N_15716,N_15961);
nor U16730 (N_16730,N_16229,N_16045);
and U16731 (N_16731,N_16094,N_16008);
xnor U16732 (N_16732,N_16073,N_15720);
or U16733 (N_16733,N_15974,N_16098);
nand U16734 (N_16734,N_16008,N_15894);
nor U16735 (N_16735,N_15646,N_16094);
nor U16736 (N_16736,N_16071,N_15894);
xor U16737 (N_16737,N_15700,N_15780);
nand U16738 (N_16738,N_15935,N_16168);
nand U16739 (N_16739,N_16085,N_16029);
nand U16740 (N_16740,N_16089,N_15870);
or U16741 (N_16741,N_16042,N_15895);
and U16742 (N_16742,N_16046,N_15666);
and U16743 (N_16743,N_15802,N_16210);
nand U16744 (N_16744,N_16018,N_15718);
and U16745 (N_16745,N_15672,N_15821);
and U16746 (N_16746,N_15833,N_15724);
nand U16747 (N_16747,N_16110,N_15983);
nand U16748 (N_16748,N_15629,N_16134);
or U16749 (N_16749,N_15647,N_15754);
nor U16750 (N_16750,N_16173,N_16191);
and U16751 (N_16751,N_15954,N_15640);
xor U16752 (N_16752,N_16064,N_15996);
xor U16753 (N_16753,N_16237,N_16128);
and U16754 (N_16754,N_16046,N_15792);
and U16755 (N_16755,N_16063,N_16196);
xor U16756 (N_16756,N_15828,N_16043);
nand U16757 (N_16757,N_16007,N_16076);
nor U16758 (N_16758,N_15918,N_16109);
and U16759 (N_16759,N_15864,N_16136);
or U16760 (N_16760,N_16210,N_16109);
and U16761 (N_16761,N_16047,N_15868);
and U16762 (N_16762,N_15666,N_15701);
nor U16763 (N_16763,N_16182,N_16068);
and U16764 (N_16764,N_15719,N_15661);
xnor U16765 (N_16765,N_15879,N_15711);
nand U16766 (N_16766,N_16105,N_15980);
and U16767 (N_16767,N_15912,N_16004);
or U16768 (N_16768,N_15655,N_16007);
or U16769 (N_16769,N_15854,N_16201);
or U16770 (N_16770,N_16024,N_16228);
or U16771 (N_16771,N_16047,N_15627);
xor U16772 (N_16772,N_15825,N_15733);
nor U16773 (N_16773,N_15877,N_15645);
nor U16774 (N_16774,N_16083,N_15946);
xor U16775 (N_16775,N_15829,N_15889);
and U16776 (N_16776,N_16221,N_16219);
nor U16777 (N_16777,N_15995,N_15805);
nand U16778 (N_16778,N_15658,N_15833);
nor U16779 (N_16779,N_16036,N_15770);
xor U16780 (N_16780,N_15690,N_15768);
and U16781 (N_16781,N_15820,N_15767);
and U16782 (N_16782,N_15931,N_16019);
xnor U16783 (N_16783,N_16236,N_16157);
nor U16784 (N_16784,N_15890,N_15815);
xnor U16785 (N_16785,N_16124,N_16081);
and U16786 (N_16786,N_16161,N_16019);
or U16787 (N_16787,N_15908,N_15659);
and U16788 (N_16788,N_15859,N_15833);
nor U16789 (N_16789,N_15709,N_15872);
xnor U16790 (N_16790,N_15893,N_15927);
nand U16791 (N_16791,N_15928,N_16239);
nor U16792 (N_16792,N_16103,N_15753);
xnor U16793 (N_16793,N_15652,N_16221);
and U16794 (N_16794,N_16151,N_15777);
xnor U16795 (N_16795,N_16089,N_16165);
nor U16796 (N_16796,N_16139,N_15880);
or U16797 (N_16797,N_15633,N_15948);
nand U16798 (N_16798,N_16032,N_16238);
nand U16799 (N_16799,N_16021,N_16215);
or U16800 (N_16800,N_16000,N_15975);
nand U16801 (N_16801,N_16022,N_15801);
nand U16802 (N_16802,N_15770,N_16011);
nand U16803 (N_16803,N_16188,N_16083);
or U16804 (N_16804,N_16157,N_16179);
nand U16805 (N_16805,N_16039,N_16075);
nand U16806 (N_16806,N_15757,N_16058);
xnor U16807 (N_16807,N_16199,N_16158);
and U16808 (N_16808,N_16127,N_15834);
and U16809 (N_16809,N_15749,N_15798);
nor U16810 (N_16810,N_15783,N_15852);
nand U16811 (N_16811,N_15998,N_15781);
and U16812 (N_16812,N_16236,N_15990);
or U16813 (N_16813,N_16240,N_16109);
nor U16814 (N_16814,N_15822,N_15746);
nand U16815 (N_16815,N_15650,N_15950);
nor U16816 (N_16816,N_15909,N_15865);
xor U16817 (N_16817,N_16220,N_15646);
nor U16818 (N_16818,N_15941,N_15904);
xor U16819 (N_16819,N_15748,N_16085);
nand U16820 (N_16820,N_15642,N_16075);
xnor U16821 (N_16821,N_15947,N_15698);
xnor U16822 (N_16822,N_16105,N_16082);
xnor U16823 (N_16823,N_15697,N_15628);
and U16824 (N_16824,N_15649,N_16249);
nor U16825 (N_16825,N_16138,N_15970);
and U16826 (N_16826,N_15700,N_16027);
or U16827 (N_16827,N_16244,N_15986);
or U16828 (N_16828,N_15751,N_16021);
nor U16829 (N_16829,N_16197,N_15695);
nor U16830 (N_16830,N_16061,N_15997);
xor U16831 (N_16831,N_15701,N_15673);
xor U16832 (N_16832,N_15700,N_15833);
or U16833 (N_16833,N_15994,N_15876);
xnor U16834 (N_16834,N_16008,N_16129);
nand U16835 (N_16835,N_15832,N_16084);
or U16836 (N_16836,N_15748,N_15862);
xnor U16837 (N_16837,N_15743,N_15811);
nor U16838 (N_16838,N_16070,N_15785);
nor U16839 (N_16839,N_15898,N_15934);
and U16840 (N_16840,N_16244,N_15931);
and U16841 (N_16841,N_16074,N_16142);
or U16842 (N_16842,N_16168,N_15955);
xnor U16843 (N_16843,N_15765,N_15961);
nor U16844 (N_16844,N_16030,N_15983);
xnor U16845 (N_16845,N_15927,N_15720);
nand U16846 (N_16846,N_15844,N_16136);
nand U16847 (N_16847,N_16240,N_15961);
nor U16848 (N_16848,N_16248,N_16247);
xnor U16849 (N_16849,N_15702,N_15740);
xor U16850 (N_16850,N_15747,N_15730);
nand U16851 (N_16851,N_15769,N_16048);
or U16852 (N_16852,N_16203,N_15632);
and U16853 (N_16853,N_15685,N_15839);
nand U16854 (N_16854,N_16150,N_15689);
or U16855 (N_16855,N_15696,N_16088);
nor U16856 (N_16856,N_16012,N_16093);
or U16857 (N_16857,N_15798,N_15801);
or U16858 (N_16858,N_16054,N_15662);
nand U16859 (N_16859,N_16025,N_15852);
and U16860 (N_16860,N_16046,N_15722);
nand U16861 (N_16861,N_15722,N_16163);
and U16862 (N_16862,N_15884,N_15722);
nand U16863 (N_16863,N_16168,N_15960);
or U16864 (N_16864,N_15632,N_15859);
nand U16865 (N_16865,N_16202,N_16057);
xor U16866 (N_16866,N_16230,N_16053);
and U16867 (N_16867,N_15927,N_16098);
xnor U16868 (N_16868,N_15870,N_16099);
xor U16869 (N_16869,N_15725,N_16058);
xor U16870 (N_16870,N_16180,N_15961);
or U16871 (N_16871,N_16035,N_16239);
xor U16872 (N_16872,N_16237,N_15988);
nor U16873 (N_16873,N_15888,N_15799);
xnor U16874 (N_16874,N_15922,N_15933);
xnor U16875 (N_16875,N_16651,N_16761);
and U16876 (N_16876,N_16434,N_16496);
xnor U16877 (N_16877,N_16757,N_16563);
xnor U16878 (N_16878,N_16424,N_16273);
and U16879 (N_16879,N_16281,N_16792);
nor U16880 (N_16880,N_16607,N_16663);
nand U16881 (N_16881,N_16411,N_16858);
or U16882 (N_16882,N_16445,N_16597);
xnor U16883 (N_16883,N_16861,N_16730);
xnor U16884 (N_16884,N_16564,N_16364);
nor U16885 (N_16885,N_16749,N_16259);
xor U16886 (N_16886,N_16303,N_16536);
or U16887 (N_16887,N_16280,N_16801);
nand U16888 (N_16888,N_16726,N_16793);
nor U16889 (N_16889,N_16475,N_16823);
nor U16890 (N_16890,N_16418,N_16457);
nor U16891 (N_16891,N_16746,N_16282);
xor U16892 (N_16892,N_16745,N_16656);
and U16893 (N_16893,N_16449,N_16350);
or U16894 (N_16894,N_16738,N_16531);
and U16895 (N_16895,N_16441,N_16501);
or U16896 (N_16896,N_16308,N_16348);
xor U16897 (N_16897,N_16355,N_16453);
or U16898 (N_16898,N_16603,N_16648);
and U16899 (N_16899,N_16809,N_16483);
nand U16900 (N_16900,N_16312,N_16758);
nor U16901 (N_16901,N_16268,N_16686);
nor U16902 (N_16902,N_16313,N_16406);
and U16903 (N_16903,N_16345,N_16669);
and U16904 (N_16904,N_16495,N_16407);
or U16905 (N_16905,N_16720,N_16650);
nor U16906 (N_16906,N_16714,N_16609);
and U16907 (N_16907,N_16602,N_16431);
and U16908 (N_16908,N_16599,N_16291);
nor U16909 (N_16909,N_16815,N_16567);
or U16910 (N_16910,N_16554,N_16575);
or U16911 (N_16911,N_16665,N_16551);
and U16912 (N_16912,N_16808,N_16822);
nor U16913 (N_16913,N_16293,N_16865);
xor U16914 (N_16914,N_16849,N_16391);
xnor U16915 (N_16915,N_16344,N_16356);
nand U16916 (N_16916,N_16487,N_16836);
or U16917 (N_16917,N_16477,N_16335);
nor U16918 (N_16918,N_16872,N_16634);
and U16919 (N_16919,N_16598,N_16804);
nand U16920 (N_16920,N_16645,N_16400);
nand U16921 (N_16921,N_16416,N_16777);
nand U16922 (N_16922,N_16253,N_16397);
and U16923 (N_16923,N_16640,N_16276);
nor U16924 (N_16924,N_16586,N_16744);
nor U16925 (N_16925,N_16351,N_16835);
nand U16926 (N_16926,N_16322,N_16780);
nand U16927 (N_16927,N_16731,N_16805);
and U16928 (N_16928,N_16543,N_16393);
xnor U16929 (N_16929,N_16839,N_16723);
nand U16930 (N_16930,N_16638,N_16257);
nand U16931 (N_16931,N_16250,N_16300);
or U16932 (N_16932,N_16410,N_16833);
xor U16933 (N_16933,N_16621,N_16334);
and U16934 (N_16934,N_16526,N_16628);
xnor U16935 (N_16935,N_16811,N_16552);
nor U16936 (N_16936,N_16314,N_16261);
nor U16937 (N_16937,N_16736,N_16519);
nand U16938 (N_16938,N_16381,N_16388);
nand U16939 (N_16939,N_16830,N_16613);
and U16940 (N_16940,N_16256,N_16409);
nand U16941 (N_16941,N_16729,N_16820);
and U16942 (N_16942,N_16685,N_16265);
xor U16943 (N_16943,N_16376,N_16759);
and U16944 (N_16944,N_16641,N_16318);
nand U16945 (N_16945,N_16688,N_16587);
and U16946 (N_16946,N_16592,N_16724);
and U16947 (N_16947,N_16392,N_16333);
nor U16948 (N_16948,N_16399,N_16639);
nor U16949 (N_16949,N_16689,N_16432);
nand U16950 (N_16950,N_16420,N_16748);
or U16951 (N_16951,N_16324,N_16684);
or U16952 (N_16952,N_16525,N_16306);
nand U16953 (N_16953,N_16384,N_16845);
or U16954 (N_16954,N_16368,N_16571);
xor U16955 (N_16955,N_16838,N_16427);
or U16956 (N_16956,N_16659,N_16576);
nor U16957 (N_16957,N_16874,N_16817);
nor U16958 (N_16958,N_16498,N_16497);
nand U16959 (N_16959,N_16649,N_16798);
nor U16960 (N_16960,N_16795,N_16588);
xnor U16961 (N_16961,N_16537,N_16462);
xor U16962 (N_16962,N_16664,N_16784);
nand U16963 (N_16963,N_16700,N_16474);
xor U16964 (N_16964,N_16605,N_16678);
or U16965 (N_16965,N_16271,N_16841);
nor U16966 (N_16966,N_16850,N_16661);
and U16967 (N_16967,N_16781,N_16524);
or U16968 (N_16968,N_16658,N_16620);
or U16969 (N_16969,N_16360,N_16252);
nand U16970 (N_16970,N_16553,N_16787);
nor U16971 (N_16971,N_16535,N_16718);
xor U16972 (N_16972,N_16488,N_16298);
xor U16973 (N_16973,N_16354,N_16414);
or U16974 (N_16974,N_16561,N_16471);
or U16975 (N_16975,N_16819,N_16813);
and U16976 (N_16976,N_16452,N_16717);
nand U16977 (N_16977,N_16579,N_16546);
nand U16978 (N_16978,N_16654,N_16617);
xor U16979 (N_16979,N_16466,N_16657);
nor U16980 (N_16980,N_16721,N_16490);
nand U16981 (N_16981,N_16679,N_16572);
xor U16982 (N_16982,N_16556,N_16295);
or U16983 (N_16983,N_16646,N_16251);
nand U16984 (N_16984,N_16387,N_16596);
nand U16985 (N_16985,N_16606,N_16705);
xnor U16986 (N_16986,N_16622,N_16816);
nand U16987 (N_16987,N_16735,N_16425);
and U16988 (N_16988,N_16283,N_16515);
or U16989 (N_16989,N_16800,N_16755);
nor U16990 (N_16990,N_16570,N_16618);
or U16991 (N_16991,N_16328,N_16520);
and U16992 (N_16992,N_16331,N_16713);
nand U16993 (N_16993,N_16568,N_16402);
or U16994 (N_16994,N_16644,N_16437);
xor U16995 (N_16995,N_16267,N_16762);
nor U16996 (N_16996,N_16357,N_16873);
or U16997 (N_16997,N_16869,N_16767);
xor U16998 (N_16998,N_16580,N_16595);
nor U16999 (N_16999,N_16843,N_16523);
and U17000 (N_17000,N_16484,N_16538);
and U17001 (N_17001,N_16851,N_16734);
or U17002 (N_17002,N_16372,N_16503);
or U17003 (N_17003,N_16367,N_16739);
xnor U17004 (N_17004,N_16547,N_16712);
xnor U17005 (N_17005,N_16701,N_16751);
and U17006 (N_17006,N_16770,N_16481);
or U17007 (N_17007,N_16840,N_16773);
nand U17008 (N_17008,N_16539,N_16301);
or U17009 (N_17009,N_16337,N_16396);
nand U17010 (N_17010,N_16383,N_16534);
xor U17011 (N_17011,N_16390,N_16677);
or U17012 (N_17012,N_16829,N_16860);
xor U17013 (N_17013,N_16470,N_16545);
xnor U17014 (N_17014,N_16302,N_16855);
and U17015 (N_17015,N_16783,N_16670);
nor U17016 (N_17016,N_16785,N_16429);
or U17017 (N_17017,N_16447,N_16662);
or U17018 (N_17018,N_16386,N_16451);
xnor U17019 (N_17019,N_16435,N_16803);
and U17020 (N_17020,N_16741,N_16653);
nor U17021 (N_17021,N_16710,N_16864);
and U17022 (N_17022,N_16455,N_16269);
nor U17023 (N_17023,N_16775,N_16442);
xor U17024 (N_17024,N_16422,N_16696);
nand U17025 (N_17025,N_16491,N_16789);
nor U17026 (N_17026,N_16352,N_16668);
xnor U17027 (N_17027,N_16358,N_16857);
and U17028 (N_17028,N_16325,N_16389);
or U17029 (N_17029,N_16541,N_16275);
and U17030 (N_17030,N_16807,N_16395);
nand U17031 (N_17031,N_16492,N_16310);
xor U17032 (N_17032,N_16788,N_16467);
nor U17033 (N_17033,N_16676,N_16270);
xor U17034 (N_17034,N_16593,N_16272);
xor U17035 (N_17035,N_16405,N_16332);
xor U17036 (N_17036,N_16377,N_16747);
or U17037 (N_17037,N_16725,N_16732);
nand U17038 (N_17038,N_16737,N_16786);
nor U17039 (N_17039,N_16585,N_16608);
and U17040 (N_17040,N_16562,N_16502);
or U17041 (N_17041,N_16320,N_16382);
nand U17042 (N_17042,N_16459,N_16419);
or U17043 (N_17043,N_16278,N_16702);
and U17044 (N_17044,N_16577,N_16507);
or U17045 (N_17045,N_16548,N_16286);
nand U17046 (N_17046,N_16415,N_16366);
or U17047 (N_17047,N_16660,N_16363);
nor U17048 (N_17048,N_16615,N_16589);
xnor U17049 (N_17049,N_16461,N_16408);
nand U17050 (N_17050,N_16549,N_16500);
nor U17051 (N_17051,N_16818,N_16307);
xor U17052 (N_17052,N_16258,N_16870);
xor U17053 (N_17053,N_16473,N_16292);
nand U17054 (N_17054,N_16478,N_16578);
and U17055 (N_17055,N_16590,N_16633);
and U17056 (N_17056,N_16687,N_16378);
xnor U17057 (N_17057,N_16530,N_16297);
and U17058 (N_17058,N_16752,N_16610);
nor U17059 (N_17059,N_16706,N_16594);
and U17060 (N_17060,N_16769,N_16672);
or U17061 (N_17061,N_16288,N_16458);
nor U17062 (N_17062,N_16683,N_16439);
nand U17063 (N_17063,N_16814,N_16834);
or U17064 (N_17064,N_16740,N_16790);
nand U17065 (N_17065,N_16369,N_16326);
nand U17066 (N_17066,N_16772,N_16476);
and U17067 (N_17067,N_16796,N_16768);
or U17068 (N_17068,N_16707,N_16379);
or U17069 (N_17069,N_16330,N_16719);
nor U17070 (N_17070,N_16697,N_16844);
and U17071 (N_17071,N_16339,N_16557);
or U17072 (N_17072,N_16299,N_16279);
nor U17073 (N_17073,N_16509,N_16401);
and U17074 (N_17074,N_16479,N_16489);
nand U17075 (N_17075,N_16652,N_16647);
or U17076 (N_17076,N_16438,N_16550);
nor U17077 (N_17077,N_16722,N_16763);
or U17078 (N_17078,N_16616,N_16499);
xor U17079 (N_17079,N_16573,N_16806);
or U17080 (N_17080,N_16756,N_16682);
or U17081 (N_17081,N_16454,N_16255);
xor U17082 (N_17082,N_16847,N_16626);
xnor U17083 (N_17083,N_16512,N_16493);
nor U17084 (N_17084,N_16304,N_16285);
nand U17085 (N_17085,N_16655,N_16340);
nor U17086 (N_17086,N_16863,N_16623);
and U17087 (N_17087,N_16266,N_16812);
xnor U17088 (N_17088,N_16778,N_16637);
xor U17089 (N_17089,N_16604,N_16558);
nor U17090 (N_17090,N_16398,N_16456);
nor U17091 (N_17091,N_16837,N_16574);
nor U17092 (N_17092,N_16284,N_16824);
xor U17093 (N_17093,N_16359,N_16450);
nand U17094 (N_17094,N_16412,N_16264);
or U17095 (N_17095,N_16635,N_16516);
xnor U17096 (N_17096,N_16533,N_16370);
xor U17097 (N_17097,N_16627,N_16518);
xor U17098 (N_17098,N_16867,N_16315);
xnor U17099 (N_17099,N_16540,N_16263);
nand U17100 (N_17100,N_16465,N_16342);
xor U17101 (N_17101,N_16582,N_16583);
xor U17102 (N_17102,N_16698,N_16373);
or U17103 (N_17103,N_16305,N_16742);
and U17104 (N_17104,N_16522,N_16630);
xnor U17105 (N_17105,N_16394,N_16528);
nand U17106 (N_17106,N_16560,N_16614);
nor U17107 (N_17107,N_16826,N_16591);
and U17108 (N_17108,N_16517,N_16694);
xor U17109 (N_17109,N_16827,N_16317);
nand U17110 (N_17110,N_16692,N_16703);
or U17111 (N_17111,N_16619,N_16868);
nor U17112 (N_17112,N_16289,N_16529);
nor U17113 (N_17113,N_16862,N_16629);
xnor U17114 (N_17114,N_16711,N_16631);
nor U17115 (N_17115,N_16294,N_16277);
nand U17116 (N_17116,N_16510,N_16385);
xor U17117 (N_17117,N_16504,N_16680);
and U17118 (N_17118,N_16754,N_16346);
nor U17119 (N_17119,N_16433,N_16667);
nand U17120 (N_17120,N_16675,N_16374);
nand U17121 (N_17121,N_16715,N_16632);
and U17122 (N_17122,N_16513,N_16274);
xnor U17123 (N_17123,N_16810,N_16309);
nor U17124 (N_17124,N_16600,N_16779);
xnor U17125 (N_17125,N_16353,N_16423);
and U17126 (N_17126,N_16428,N_16771);
nor U17127 (N_17127,N_16750,N_16709);
or U17128 (N_17128,N_16776,N_16327);
xnor U17129 (N_17129,N_16316,N_16468);
nand U17130 (N_17130,N_16336,N_16791);
or U17131 (N_17131,N_16403,N_16254);
xnor U17132 (N_17132,N_16674,N_16821);
nor U17133 (N_17133,N_16569,N_16404);
nor U17134 (N_17134,N_16691,N_16601);
nor U17135 (N_17135,N_16774,N_16371);
or U17136 (N_17136,N_16642,N_16361);
or U17137 (N_17137,N_16733,N_16704);
xnor U17138 (N_17138,N_16311,N_16321);
nor U17139 (N_17139,N_16542,N_16584);
xnor U17140 (N_17140,N_16413,N_16469);
or U17141 (N_17141,N_16693,N_16765);
or U17142 (N_17142,N_16699,N_16766);
nand U17143 (N_17143,N_16794,N_16581);
nor U17144 (N_17144,N_16559,N_16430);
and U17145 (N_17145,N_16728,N_16831);
and U17146 (N_17146,N_16625,N_16362);
and U17147 (N_17147,N_16421,N_16443);
and U17148 (N_17148,N_16482,N_16532);
nor U17149 (N_17149,N_16486,N_16480);
xnor U17150 (N_17150,N_16681,N_16505);
xor U17151 (N_17151,N_16566,N_16859);
nand U17152 (N_17152,N_16262,N_16508);
and U17153 (N_17153,N_16764,N_16472);
nand U17154 (N_17154,N_16565,N_16832);
or U17155 (N_17155,N_16329,N_16666);
nand U17156 (N_17156,N_16828,N_16871);
nor U17157 (N_17157,N_16612,N_16463);
or U17158 (N_17158,N_16611,N_16695);
or U17159 (N_17159,N_16347,N_16743);
nand U17160 (N_17160,N_16446,N_16287);
and U17161 (N_17161,N_16636,N_16290);
or U17162 (N_17162,N_16506,N_16799);
xnor U17163 (N_17163,N_16866,N_16341);
or U17164 (N_17164,N_16797,N_16782);
xnor U17165 (N_17165,N_16319,N_16464);
or U17166 (N_17166,N_16426,N_16521);
or U17167 (N_17167,N_16544,N_16485);
xnor U17168 (N_17168,N_16440,N_16753);
nor U17169 (N_17169,N_16380,N_16527);
xnor U17170 (N_17170,N_16448,N_16727);
and U17171 (N_17171,N_16856,N_16343);
or U17172 (N_17172,N_16854,N_16444);
and U17173 (N_17173,N_16624,N_16260);
nand U17174 (N_17174,N_16716,N_16673);
nor U17175 (N_17175,N_16825,N_16852);
nand U17176 (N_17176,N_16514,N_16760);
nand U17177 (N_17177,N_16802,N_16436);
or U17178 (N_17178,N_16643,N_16511);
and U17179 (N_17179,N_16349,N_16296);
xor U17180 (N_17180,N_16842,N_16853);
xor U17181 (N_17181,N_16338,N_16417);
nand U17182 (N_17182,N_16671,N_16708);
nor U17183 (N_17183,N_16690,N_16375);
nand U17184 (N_17184,N_16460,N_16555);
or U17185 (N_17185,N_16365,N_16494);
xor U17186 (N_17186,N_16846,N_16323);
nor U17187 (N_17187,N_16848,N_16802);
or U17188 (N_17188,N_16366,N_16825);
and U17189 (N_17189,N_16628,N_16319);
nor U17190 (N_17190,N_16543,N_16631);
or U17191 (N_17191,N_16427,N_16283);
nand U17192 (N_17192,N_16586,N_16788);
xor U17193 (N_17193,N_16424,N_16491);
and U17194 (N_17194,N_16640,N_16721);
xor U17195 (N_17195,N_16536,N_16803);
nand U17196 (N_17196,N_16356,N_16482);
xor U17197 (N_17197,N_16677,N_16444);
or U17198 (N_17198,N_16279,N_16645);
nand U17199 (N_17199,N_16379,N_16490);
and U17200 (N_17200,N_16672,N_16598);
or U17201 (N_17201,N_16419,N_16755);
nand U17202 (N_17202,N_16260,N_16495);
xnor U17203 (N_17203,N_16562,N_16848);
and U17204 (N_17204,N_16804,N_16768);
or U17205 (N_17205,N_16811,N_16349);
nand U17206 (N_17206,N_16725,N_16319);
xor U17207 (N_17207,N_16700,N_16809);
nand U17208 (N_17208,N_16749,N_16483);
xor U17209 (N_17209,N_16469,N_16691);
nand U17210 (N_17210,N_16428,N_16311);
nand U17211 (N_17211,N_16367,N_16523);
xor U17212 (N_17212,N_16869,N_16603);
nor U17213 (N_17213,N_16660,N_16328);
and U17214 (N_17214,N_16600,N_16277);
nand U17215 (N_17215,N_16726,N_16258);
xor U17216 (N_17216,N_16403,N_16748);
nor U17217 (N_17217,N_16819,N_16799);
nand U17218 (N_17218,N_16573,N_16712);
and U17219 (N_17219,N_16407,N_16512);
xor U17220 (N_17220,N_16505,N_16348);
xnor U17221 (N_17221,N_16551,N_16847);
or U17222 (N_17222,N_16406,N_16862);
and U17223 (N_17223,N_16734,N_16327);
nand U17224 (N_17224,N_16866,N_16629);
nor U17225 (N_17225,N_16857,N_16796);
or U17226 (N_17226,N_16749,N_16613);
xnor U17227 (N_17227,N_16447,N_16472);
nand U17228 (N_17228,N_16534,N_16747);
nand U17229 (N_17229,N_16560,N_16578);
nand U17230 (N_17230,N_16296,N_16506);
or U17231 (N_17231,N_16693,N_16712);
and U17232 (N_17232,N_16696,N_16839);
or U17233 (N_17233,N_16468,N_16627);
and U17234 (N_17234,N_16665,N_16350);
or U17235 (N_17235,N_16354,N_16655);
and U17236 (N_17236,N_16355,N_16732);
or U17237 (N_17237,N_16870,N_16853);
or U17238 (N_17238,N_16435,N_16535);
nand U17239 (N_17239,N_16650,N_16417);
nand U17240 (N_17240,N_16345,N_16391);
xor U17241 (N_17241,N_16470,N_16715);
nor U17242 (N_17242,N_16353,N_16387);
nor U17243 (N_17243,N_16530,N_16342);
or U17244 (N_17244,N_16307,N_16551);
nand U17245 (N_17245,N_16463,N_16425);
nand U17246 (N_17246,N_16314,N_16807);
nand U17247 (N_17247,N_16720,N_16519);
xnor U17248 (N_17248,N_16287,N_16283);
xor U17249 (N_17249,N_16641,N_16291);
nand U17250 (N_17250,N_16807,N_16707);
and U17251 (N_17251,N_16722,N_16621);
or U17252 (N_17252,N_16830,N_16486);
and U17253 (N_17253,N_16725,N_16320);
xor U17254 (N_17254,N_16361,N_16840);
or U17255 (N_17255,N_16661,N_16269);
nor U17256 (N_17256,N_16549,N_16724);
xnor U17257 (N_17257,N_16634,N_16478);
or U17258 (N_17258,N_16412,N_16753);
and U17259 (N_17259,N_16257,N_16342);
nor U17260 (N_17260,N_16291,N_16728);
nand U17261 (N_17261,N_16530,N_16771);
nand U17262 (N_17262,N_16395,N_16487);
nor U17263 (N_17263,N_16273,N_16455);
or U17264 (N_17264,N_16323,N_16745);
nor U17265 (N_17265,N_16312,N_16480);
or U17266 (N_17266,N_16662,N_16542);
nand U17267 (N_17267,N_16865,N_16327);
xor U17268 (N_17268,N_16428,N_16722);
and U17269 (N_17269,N_16761,N_16332);
or U17270 (N_17270,N_16618,N_16624);
nand U17271 (N_17271,N_16704,N_16724);
nor U17272 (N_17272,N_16581,N_16314);
xor U17273 (N_17273,N_16829,N_16506);
and U17274 (N_17274,N_16755,N_16843);
or U17275 (N_17275,N_16778,N_16856);
nand U17276 (N_17276,N_16824,N_16589);
nor U17277 (N_17277,N_16266,N_16328);
nor U17278 (N_17278,N_16653,N_16280);
xnor U17279 (N_17279,N_16273,N_16383);
nand U17280 (N_17280,N_16672,N_16341);
xnor U17281 (N_17281,N_16330,N_16840);
xnor U17282 (N_17282,N_16373,N_16307);
nand U17283 (N_17283,N_16520,N_16871);
xor U17284 (N_17284,N_16633,N_16558);
xnor U17285 (N_17285,N_16712,N_16364);
nor U17286 (N_17286,N_16344,N_16394);
nand U17287 (N_17287,N_16646,N_16379);
and U17288 (N_17288,N_16336,N_16693);
and U17289 (N_17289,N_16622,N_16449);
nor U17290 (N_17290,N_16560,N_16682);
nand U17291 (N_17291,N_16633,N_16257);
xnor U17292 (N_17292,N_16657,N_16254);
nand U17293 (N_17293,N_16711,N_16650);
and U17294 (N_17294,N_16763,N_16346);
nor U17295 (N_17295,N_16742,N_16668);
nor U17296 (N_17296,N_16380,N_16721);
nor U17297 (N_17297,N_16524,N_16874);
xor U17298 (N_17298,N_16846,N_16855);
nand U17299 (N_17299,N_16400,N_16451);
nand U17300 (N_17300,N_16555,N_16327);
nand U17301 (N_17301,N_16652,N_16830);
nor U17302 (N_17302,N_16357,N_16615);
and U17303 (N_17303,N_16443,N_16372);
nand U17304 (N_17304,N_16638,N_16730);
or U17305 (N_17305,N_16575,N_16711);
nor U17306 (N_17306,N_16645,N_16708);
xnor U17307 (N_17307,N_16417,N_16646);
nor U17308 (N_17308,N_16821,N_16349);
nor U17309 (N_17309,N_16775,N_16765);
nand U17310 (N_17310,N_16280,N_16680);
or U17311 (N_17311,N_16272,N_16730);
nand U17312 (N_17312,N_16322,N_16627);
nor U17313 (N_17313,N_16563,N_16443);
nor U17314 (N_17314,N_16753,N_16329);
nor U17315 (N_17315,N_16703,N_16292);
nand U17316 (N_17316,N_16694,N_16545);
and U17317 (N_17317,N_16681,N_16534);
nand U17318 (N_17318,N_16367,N_16428);
or U17319 (N_17319,N_16381,N_16252);
nand U17320 (N_17320,N_16486,N_16661);
nand U17321 (N_17321,N_16474,N_16551);
nor U17322 (N_17322,N_16723,N_16417);
nand U17323 (N_17323,N_16301,N_16811);
xnor U17324 (N_17324,N_16808,N_16500);
nand U17325 (N_17325,N_16789,N_16870);
and U17326 (N_17326,N_16666,N_16345);
nor U17327 (N_17327,N_16292,N_16276);
and U17328 (N_17328,N_16640,N_16560);
nand U17329 (N_17329,N_16440,N_16693);
or U17330 (N_17330,N_16670,N_16470);
and U17331 (N_17331,N_16634,N_16537);
nand U17332 (N_17332,N_16625,N_16310);
xnor U17333 (N_17333,N_16278,N_16692);
nand U17334 (N_17334,N_16866,N_16485);
or U17335 (N_17335,N_16370,N_16550);
nand U17336 (N_17336,N_16514,N_16681);
nor U17337 (N_17337,N_16538,N_16320);
xnor U17338 (N_17338,N_16742,N_16845);
nor U17339 (N_17339,N_16325,N_16841);
and U17340 (N_17340,N_16671,N_16318);
or U17341 (N_17341,N_16681,N_16718);
xnor U17342 (N_17342,N_16438,N_16720);
xor U17343 (N_17343,N_16514,N_16571);
nor U17344 (N_17344,N_16641,N_16425);
and U17345 (N_17345,N_16251,N_16467);
nor U17346 (N_17346,N_16852,N_16693);
and U17347 (N_17347,N_16533,N_16396);
nor U17348 (N_17348,N_16549,N_16352);
or U17349 (N_17349,N_16427,N_16760);
nand U17350 (N_17350,N_16821,N_16291);
and U17351 (N_17351,N_16560,N_16853);
and U17352 (N_17352,N_16499,N_16454);
and U17353 (N_17353,N_16766,N_16404);
nand U17354 (N_17354,N_16333,N_16461);
and U17355 (N_17355,N_16751,N_16546);
nor U17356 (N_17356,N_16781,N_16601);
and U17357 (N_17357,N_16601,N_16282);
xnor U17358 (N_17358,N_16394,N_16303);
nor U17359 (N_17359,N_16297,N_16318);
xnor U17360 (N_17360,N_16296,N_16865);
and U17361 (N_17361,N_16743,N_16514);
xor U17362 (N_17362,N_16647,N_16377);
xnor U17363 (N_17363,N_16470,N_16489);
nor U17364 (N_17364,N_16514,N_16857);
xor U17365 (N_17365,N_16784,N_16422);
nor U17366 (N_17366,N_16367,N_16352);
and U17367 (N_17367,N_16818,N_16577);
xnor U17368 (N_17368,N_16436,N_16582);
and U17369 (N_17369,N_16412,N_16282);
or U17370 (N_17370,N_16443,N_16449);
nand U17371 (N_17371,N_16274,N_16626);
xor U17372 (N_17372,N_16374,N_16814);
nand U17373 (N_17373,N_16871,N_16347);
nor U17374 (N_17374,N_16710,N_16309);
nor U17375 (N_17375,N_16588,N_16536);
nor U17376 (N_17376,N_16540,N_16437);
or U17377 (N_17377,N_16581,N_16619);
or U17378 (N_17378,N_16504,N_16319);
or U17379 (N_17379,N_16514,N_16348);
and U17380 (N_17380,N_16869,N_16798);
nor U17381 (N_17381,N_16838,N_16660);
nor U17382 (N_17382,N_16685,N_16492);
nand U17383 (N_17383,N_16440,N_16525);
nor U17384 (N_17384,N_16644,N_16529);
or U17385 (N_17385,N_16305,N_16370);
or U17386 (N_17386,N_16497,N_16737);
nand U17387 (N_17387,N_16697,N_16689);
or U17388 (N_17388,N_16833,N_16692);
nor U17389 (N_17389,N_16470,N_16730);
nor U17390 (N_17390,N_16340,N_16773);
and U17391 (N_17391,N_16369,N_16440);
xor U17392 (N_17392,N_16437,N_16804);
nand U17393 (N_17393,N_16457,N_16797);
nor U17394 (N_17394,N_16759,N_16383);
and U17395 (N_17395,N_16654,N_16252);
nand U17396 (N_17396,N_16307,N_16856);
or U17397 (N_17397,N_16825,N_16597);
and U17398 (N_17398,N_16713,N_16775);
or U17399 (N_17399,N_16398,N_16270);
or U17400 (N_17400,N_16765,N_16374);
nor U17401 (N_17401,N_16687,N_16482);
nand U17402 (N_17402,N_16420,N_16422);
or U17403 (N_17403,N_16261,N_16272);
nand U17404 (N_17404,N_16384,N_16506);
nor U17405 (N_17405,N_16541,N_16747);
xor U17406 (N_17406,N_16833,N_16625);
nand U17407 (N_17407,N_16764,N_16305);
and U17408 (N_17408,N_16764,N_16268);
nor U17409 (N_17409,N_16792,N_16486);
xnor U17410 (N_17410,N_16527,N_16736);
xnor U17411 (N_17411,N_16314,N_16791);
nor U17412 (N_17412,N_16526,N_16834);
nand U17413 (N_17413,N_16611,N_16660);
and U17414 (N_17414,N_16421,N_16366);
nor U17415 (N_17415,N_16437,N_16820);
xor U17416 (N_17416,N_16293,N_16619);
and U17417 (N_17417,N_16484,N_16733);
and U17418 (N_17418,N_16873,N_16332);
or U17419 (N_17419,N_16305,N_16316);
or U17420 (N_17420,N_16393,N_16369);
or U17421 (N_17421,N_16607,N_16793);
nand U17422 (N_17422,N_16413,N_16253);
nor U17423 (N_17423,N_16363,N_16871);
nor U17424 (N_17424,N_16679,N_16797);
nand U17425 (N_17425,N_16808,N_16503);
xor U17426 (N_17426,N_16703,N_16284);
and U17427 (N_17427,N_16778,N_16370);
nor U17428 (N_17428,N_16663,N_16710);
and U17429 (N_17429,N_16827,N_16425);
or U17430 (N_17430,N_16818,N_16736);
xor U17431 (N_17431,N_16713,N_16280);
or U17432 (N_17432,N_16841,N_16283);
nor U17433 (N_17433,N_16405,N_16865);
nand U17434 (N_17434,N_16847,N_16421);
or U17435 (N_17435,N_16751,N_16809);
nor U17436 (N_17436,N_16737,N_16535);
and U17437 (N_17437,N_16320,N_16676);
xnor U17438 (N_17438,N_16437,N_16407);
and U17439 (N_17439,N_16672,N_16431);
or U17440 (N_17440,N_16407,N_16827);
nand U17441 (N_17441,N_16331,N_16567);
and U17442 (N_17442,N_16599,N_16351);
or U17443 (N_17443,N_16475,N_16653);
nand U17444 (N_17444,N_16290,N_16345);
nand U17445 (N_17445,N_16729,N_16853);
xor U17446 (N_17446,N_16670,N_16334);
xnor U17447 (N_17447,N_16498,N_16331);
or U17448 (N_17448,N_16377,N_16733);
nand U17449 (N_17449,N_16397,N_16446);
and U17450 (N_17450,N_16470,N_16554);
nand U17451 (N_17451,N_16633,N_16358);
or U17452 (N_17452,N_16375,N_16327);
nor U17453 (N_17453,N_16864,N_16427);
or U17454 (N_17454,N_16756,N_16857);
nor U17455 (N_17455,N_16508,N_16761);
and U17456 (N_17456,N_16769,N_16408);
xor U17457 (N_17457,N_16465,N_16692);
and U17458 (N_17458,N_16258,N_16659);
nor U17459 (N_17459,N_16817,N_16614);
xor U17460 (N_17460,N_16415,N_16642);
nor U17461 (N_17461,N_16715,N_16594);
or U17462 (N_17462,N_16473,N_16764);
or U17463 (N_17463,N_16558,N_16262);
and U17464 (N_17464,N_16867,N_16629);
nand U17465 (N_17465,N_16308,N_16678);
xor U17466 (N_17466,N_16313,N_16809);
and U17467 (N_17467,N_16591,N_16290);
and U17468 (N_17468,N_16799,N_16385);
xnor U17469 (N_17469,N_16358,N_16545);
or U17470 (N_17470,N_16637,N_16752);
nand U17471 (N_17471,N_16593,N_16624);
nand U17472 (N_17472,N_16549,N_16268);
nor U17473 (N_17473,N_16855,N_16353);
and U17474 (N_17474,N_16636,N_16425);
nand U17475 (N_17475,N_16559,N_16446);
nor U17476 (N_17476,N_16656,N_16532);
or U17477 (N_17477,N_16410,N_16424);
nor U17478 (N_17478,N_16626,N_16420);
and U17479 (N_17479,N_16519,N_16381);
nor U17480 (N_17480,N_16686,N_16485);
xor U17481 (N_17481,N_16723,N_16409);
nor U17482 (N_17482,N_16828,N_16477);
nand U17483 (N_17483,N_16510,N_16532);
nand U17484 (N_17484,N_16507,N_16387);
nand U17485 (N_17485,N_16331,N_16661);
or U17486 (N_17486,N_16323,N_16360);
nor U17487 (N_17487,N_16676,N_16705);
or U17488 (N_17488,N_16639,N_16448);
or U17489 (N_17489,N_16854,N_16619);
nand U17490 (N_17490,N_16320,N_16271);
and U17491 (N_17491,N_16593,N_16810);
nor U17492 (N_17492,N_16498,N_16608);
nand U17493 (N_17493,N_16499,N_16636);
or U17494 (N_17494,N_16505,N_16639);
nand U17495 (N_17495,N_16752,N_16611);
nand U17496 (N_17496,N_16775,N_16515);
nor U17497 (N_17497,N_16671,N_16681);
xor U17498 (N_17498,N_16458,N_16764);
and U17499 (N_17499,N_16584,N_16337);
or U17500 (N_17500,N_17465,N_16905);
xor U17501 (N_17501,N_17148,N_17348);
and U17502 (N_17502,N_16935,N_16956);
or U17503 (N_17503,N_17046,N_17138);
nor U17504 (N_17504,N_17000,N_17087);
or U17505 (N_17505,N_17400,N_17399);
xnor U17506 (N_17506,N_16994,N_17214);
xor U17507 (N_17507,N_17357,N_17246);
and U17508 (N_17508,N_17055,N_17277);
and U17509 (N_17509,N_17198,N_17178);
or U17510 (N_17510,N_16911,N_17059);
and U17511 (N_17511,N_16974,N_17434);
and U17512 (N_17512,N_17019,N_17157);
xnor U17513 (N_17513,N_17469,N_17403);
or U17514 (N_17514,N_17407,N_16998);
xnor U17515 (N_17515,N_16936,N_17171);
xnor U17516 (N_17516,N_17075,N_17451);
xnor U17517 (N_17517,N_17231,N_17293);
nor U17518 (N_17518,N_17083,N_17464);
nand U17519 (N_17519,N_17385,N_16888);
nor U17520 (N_17520,N_16975,N_17350);
nor U17521 (N_17521,N_17209,N_17028);
xnor U17522 (N_17522,N_17474,N_17193);
xnor U17523 (N_17523,N_17227,N_17298);
nor U17524 (N_17524,N_16947,N_17127);
nor U17525 (N_17525,N_17174,N_16928);
nand U17526 (N_17526,N_17067,N_17307);
nor U17527 (N_17527,N_17487,N_17168);
nor U17528 (N_17528,N_17011,N_17191);
xnor U17529 (N_17529,N_17016,N_16977);
nand U17530 (N_17530,N_17339,N_17017);
and U17531 (N_17531,N_16913,N_16951);
xnor U17532 (N_17532,N_17404,N_17163);
or U17533 (N_17533,N_16976,N_17472);
or U17534 (N_17534,N_17423,N_17468);
nor U17535 (N_17535,N_17143,N_17386);
or U17536 (N_17536,N_17279,N_16941);
xnor U17537 (N_17537,N_17115,N_17485);
nand U17538 (N_17538,N_17327,N_16916);
and U17539 (N_17539,N_17460,N_17336);
nand U17540 (N_17540,N_17034,N_16980);
and U17541 (N_17541,N_16971,N_17160);
and U17542 (N_17542,N_17424,N_17475);
nand U17543 (N_17543,N_17065,N_17181);
and U17544 (N_17544,N_17388,N_17345);
and U17545 (N_17545,N_17090,N_17483);
xor U17546 (N_17546,N_16986,N_17054);
xor U17547 (N_17547,N_17351,N_17006);
and U17548 (N_17548,N_17128,N_17096);
nand U17549 (N_17549,N_17499,N_17481);
nor U17550 (N_17550,N_17377,N_17466);
xor U17551 (N_17551,N_17235,N_17108);
xnor U17552 (N_17552,N_17250,N_17050);
xnor U17553 (N_17553,N_17410,N_17306);
nand U17554 (N_17554,N_17333,N_17111);
xnor U17555 (N_17555,N_17442,N_16996);
nand U17556 (N_17556,N_17486,N_17176);
nand U17557 (N_17557,N_17249,N_17304);
or U17558 (N_17558,N_17383,N_17081);
nor U17559 (N_17559,N_17069,N_16981);
or U17560 (N_17560,N_17002,N_17353);
or U17561 (N_17561,N_17213,N_17370);
nand U17562 (N_17562,N_17489,N_17317);
and U17563 (N_17563,N_17030,N_17493);
or U17564 (N_17564,N_17195,N_17380);
nor U17565 (N_17565,N_17378,N_16995);
xnor U17566 (N_17566,N_17360,N_16906);
xnor U17567 (N_17567,N_17261,N_17420);
and U17568 (N_17568,N_17440,N_17478);
nor U17569 (N_17569,N_16959,N_17072);
xnor U17570 (N_17570,N_17484,N_17390);
or U17571 (N_17571,N_16880,N_17452);
nor U17572 (N_17572,N_16886,N_17431);
nor U17573 (N_17573,N_16918,N_17161);
xnor U17574 (N_17574,N_17189,N_17029);
and U17575 (N_17575,N_16964,N_17273);
xor U17576 (N_17576,N_16919,N_17256);
xor U17577 (N_17577,N_16982,N_16910);
or U17578 (N_17578,N_17435,N_16875);
nor U17579 (N_17579,N_17175,N_16883);
xnor U17580 (N_17580,N_17013,N_16926);
nor U17581 (N_17581,N_16940,N_17076);
nor U17582 (N_17582,N_17280,N_17276);
nand U17583 (N_17583,N_17457,N_17091);
xnor U17584 (N_17584,N_16907,N_17392);
and U17585 (N_17585,N_17286,N_17365);
xnor U17586 (N_17586,N_17254,N_16973);
nand U17587 (N_17587,N_17165,N_16927);
and U17588 (N_17588,N_16882,N_17459);
nor U17589 (N_17589,N_17239,N_17042);
xor U17590 (N_17590,N_17409,N_17375);
nand U17591 (N_17591,N_17238,N_17397);
xor U17592 (N_17592,N_17453,N_17344);
or U17593 (N_17593,N_17325,N_17288);
xnor U17594 (N_17594,N_17221,N_17234);
nand U17595 (N_17595,N_17335,N_17308);
nand U17596 (N_17596,N_17158,N_16988);
or U17597 (N_17597,N_17272,N_17122);
xor U17598 (N_17598,N_16889,N_17026);
and U17599 (N_17599,N_17057,N_17190);
xnor U17600 (N_17600,N_17425,N_16891);
and U17601 (N_17601,N_17018,N_16942);
or U17602 (N_17602,N_16970,N_17292);
or U17603 (N_17603,N_17264,N_16929);
nor U17604 (N_17604,N_16902,N_17008);
and U17605 (N_17605,N_17226,N_17462);
or U17606 (N_17606,N_16932,N_17043);
xnor U17607 (N_17607,N_17051,N_17166);
or U17608 (N_17608,N_17173,N_17172);
nor U17609 (N_17609,N_17156,N_17202);
xor U17610 (N_17610,N_17428,N_17114);
nand U17611 (N_17611,N_17224,N_16885);
or U17612 (N_17612,N_16992,N_17093);
or U17613 (N_17613,N_17498,N_16904);
or U17614 (N_17614,N_17020,N_17053);
or U17615 (N_17615,N_17123,N_17032);
nor U17616 (N_17616,N_17037,N_17334);
and U17617 (N_17617,N_16962,N_17041);
nand U17618 (N_17618,N_16949,N_16899);
nand U17619 (N_17619,N_16923,N_17346);
xor U17620 (N_17620,N_17140,N_17267);
or U17621 (N_17621,N_17117,N_17203);
nor U17622 (N_17622,N_16878,N_17355);
xnor U17623 (N_17623,N_17302,N_17027);
xnor U17624 (N_17624,N_16945,N_17154);
or U17625 (N_17625,N_16895,N_17066);
xor U17626 (N_17626,N_16997,N_17247);
nand U17627 (N_17627,N_16903,N_16963);
xnor U17628 (N_17628,N_17242,N_16985);
or U17629 (N_17629,N_17290,N_17147);
and U17630 (N_17630,N_17199,N_17401);
xnor U17631 (N_17631,N_17183,N_16967);
xnor U17632 (N_17632,N_17482,N_17294);
nand U17633 (N_17633,N_17271,N_17496);
and U17634 (N_17634,N_17303,N_16979);
and U17635 (N_17635,N_16917,N_17413);
nor U17636 (N_17636,N_17429,N_17391);
nor U17637 (N_17637,N_16983,N_17461);
or U17638 (N_17638,N_17121,N_17282);
nand U17639 (N_17639,N_17326,N_16989);
nor U17640 (N_17640,N_17206,N_16953);
xor U17641 (N_17641,N_17196,N_16897);
nor U17642 (N_17642,N_17291,N_17218);
xnor U17643 (N_17643,N_16987,N_17358);
or U17644 (N_17644,N_17044,N_17110);
or U17645 (N_17645,N_17359,N_17275);
nor U17646 (N_17646,N_17211,N_17124);
xor U17647 (N_17647,N_17185,N_17473);
or U17648 (N_17648,N_16914,N_17396);
nand U17649 (N_17649,N_16909,N_17118);
or U17650 (N_17650,N_17444,N_17217);
xor U17651 (N_17651,N_17314,N_17471);
xnor U17652 (N_17652,N_17343,N_16930);
xnor U17653 (N_17653,N_17039,N_17448);
nand U17654 (N_17654,N_17092,N_17463);
nand U17655 (N_17655,N_17438,N_17188);
xor U17656 (N_17656,N_17169,N_17480);
nand U17657 (N_17657,N_17036,N_17492);
nor U17658 (N_17658,N_17159,N_17103);
and U17659 (N_17659,N_16934,N_17330);
nand U17660 (N_17660,N_17406,N_17144);
xnor U17661 (N_17661,N_17058,N_17268);
xnor U17662 (N_17662,N_17412,N_16898);
or U17663 (N_17663,N_17073,N_17015);
or U17664 (N_17664,N_17419,N_17074);
or U17665 (N_17665,N_16968,N_16938);
nand U17666 (N_17666,N_17257,N_17329);
or U17667 (N_17667,N_17430,N_17299);
nand U17668 (N_17668,N_17338,N_17102);
and U17669 (N_17669,N_17088,N_17269);
or U17670 (N_17670,N_17236,N_17374);
xor U17671 (N_17671,N_17446,N_17497);
nor U17672 (N_17672,N_17152,N_17084);
nand U17673 (N_17673,N_17177,N_17426);
xor U17674 (N_17674,N_17225,N_17142);
and U17675 (N_17675,N_17322,N_16901);
xor U17676 (N_17676,N_17321,N_17099);
xor U17677 (N_17677,N_16944,N_17309);
xnor U17678 (N_17678,N_17427,N_17210);
and U17679 (N_17679,N_17048,N_17033);
or U17680 (N_17680,N_17184,N_17433);
or U17681 (N_17681,N_17164,N_16931);
or U17682 (N_17682,N_17205,N_16990);
nor U17683 (N_17683,N_17001,N_17323);
and U17684 (N_17684,N_17113,N_17207);
or U17685 (N_17685,N_16961,N_16965);
nand U17686 (N_17686,N_17216,N_17192);
and U17687 (N_17687,N_17415,N_17311);
nand U17688 (N_17688,N_17394,N_17296);
nand U17689 (N_17689,N_17182,N_17135);
nand U17690 (N_17690,N_16946,N_17204);
nand U17691 (N_17691,N_16915,N_16966);
or U17692 (N_17692,N_17405,N_16933);
or U17693 (N_17693,N_17106,N_17283);
nor U17694 (N_17694,N_17062,N_17031);
nor U17695 (N_17695,N_17445,N_17258);
xor U17696 (N_17696,N_17371,N_17432);
and U17697 (N_17697,N_17362,N_17316);
and U17698 (N_17698,N_17479,N_17363);
nand U17699 (N_17699,N_17477,N_17025);
and U17700 (N_17700,N_16892,N_17187);
or U17701 (N_17701,N_17418,N_17153);
and U17702 (N_17702,N_17449,N_17285);
and U17703 (N_17703,N_17393,N_17009);
and U17704 (N_17704,N_17134,N_17136);
nor U17705 (N_17705,N_17131,N_17060);
nor U17706 (N_17706,N_17082,N_17324);
nand U17707 (N_17707,N_17064,N_16960);
nor U17708 (N_17708,N_16972,N_17229);
nand U17709 (N_17709,N_17443,N_17310);
nand U17710 (N_17710,N_16884,N_17270);
nor U17711 (N_17711,N_16999,N_17130);
nand U17712 (N_17712,N_17274,N_17010);
and U17713 (N_17713,N_17259,N_17109);
and U17714 (N_17714,N_17056,N_16894);
or U17715 (N_17715,N_17450,N_17197);
and U17716 (N_17716,N_17494,N_17212);
nor U17717 (N_17717,N_17382,N_17266);
or U17718 (N_17718,N_17364,N_17023);
nand U17719 (N_17719,N_17422,N_17107);
xor U17720 (N_17720,N_16879,N_17414);
or U17721 (N_17721,N_17337,N_17003);
xnor U17722 (N_17722,N_16952,N_16937);
or U17723 (N_17723,N_17230,N_16969);
xnor U17724 (N_17724,N_16958,N_17495);
or U17725 (N_17725,N_17300,N_17328);
xnor U17726 (N_17726,N_17265,N_17395);
xor U17727 (N_17727,N_17305,N_17208);
or U17728 (N_17728,N_17233,N_16939);
nor U17729 (N_17729,N_17278,N_17070);
or U17730 (N_17730,N_17222,N_17180);
xnor U17731 (N_17731,N_17047,N_17488);
xor U17732 (N_17732,N_17421,N_17248);
and U17733 (N_17733,N_17170,N_17320);
xor U17734 (N_17734,N_17194,N_17253);
xor U17735 (N_17735,N_16978,N_17086);
xor U17736 (N_17736,N_17476,N_17078);
nand U17737 (N_17737,N_17155,N_17458);
nand U17738 (N_17738,N_17439,N_16993);
nand U17739 (N_17739,N_16984,N_17384);
and U17740 (N_17740,N_17347,N_16948);
or U17741 (N_17741,N_17139,N_17361);
nand U17742 (N_17742,N_17436,N_17366);
or U17743 (N_17743,N_17260,N_17437);
nand U17744 (N_17744,N_16920,N_17022);
xnor U17745 (N_17745,N_17342,N_17319);
and U17746 (N_17746,N_17417,N_17132);
xnor U17747 (N_17747,N_17079,N_17112);
or U17748 (N_17748,N_17098,N_17416);
or U17749 (N_17749,N_17376,N_17145);
or U17750 (N_17750,N_17455,N_17167);
or U17751 (N_17751,N_17295,N_17297);
xnor U17752 (N_17752,N_17241,N_16912);
or U17753 (N_17753,N_16877,N_17045);
xnor U17754 (N_17754,N_17315,N_17137);
nor U17755 (N_17755,N_17133,N_17237);
nor U17756 (N_17756,N_17332,N_17220);
xor U17757 (N_17757,N_17095,N_17387);
or U17758 (N_17758,N_17119,N_17367);
and U17759 (N_17759,N_17162,N_17245);
xnor U17760 (N_17760,N_17490,N_16896);
xnor U17761 (N_17761,N_17352,N_16957);
xnor U17762 (N_17762,N_17200,N_16908);
nor U17763 (N_17763,N_17116,N_17318);
and U17764 (N_17764,N_17186,N_17105);
nor U17765 (N_17765,N_17262,N_17240);
nand U17766 (N_17766,N_17408,N_17179);
nor U17767 (N_17767,N_17150,N_17369);
nor U17768 (N_17768,N_17005,N_17402);
nand U17769 (N_17769,N_17012,N_17052);
and U17770 (N_17770,N_17035,N_17125);
nor U17771 (N_17771,N_17441,N_17120);
nor U17772 (N_17772,N_17251,N_17372);
nor U17773 (N_17773,N_17071,N_17068);
nand U17774 (N_17774,N_17232,N_17381);
nor U17775 (N_17775,N_16925,N_17287);
nand U17776 (N_17776,N_17252,N_17063);
and U17777 (N_17777,N_17411,N_17014);
and U17778 (N_17778,N_17356,N_17223);
or U17779 (N_17779,N_17097,N_16887);
xor U17780 (N_17780,N_17141,N_17061);
and U17781 (N_17781,N_16900,N_17313);
nor U17782 (N_17782,N_17024,N_17126);
nor U17783 (N_17783,N_17094,N_16943);
or U17784 (N_17784,N_17349,N_17215);
and U17785 (N_17785,N_17243,N_17049);
nor U17786 (N_17786,N_17219,N_17040);
xor U17787 (N_17787,N_17470,N_17341);
and U17788 (N_17788,N_16893,N_17398);
nand U17789 (N_17789,N_17077,N_17089);
and U17790 (N_17790,N_17447,N_17101);
nor U17791 (N_17791,N_17201,N_17021);
xor U17792 (N_17792,N_16924,N_16954);
nor U17793 (N_17793,N_17301,N_17085);
nand U17794 (N_17794,N_17080,N_17312);
xor U17795 (N_17795,N_17007,N_16922);
and U17796 (N_17796,N_17289,N_16991);
nand U17797 (N_17797,N_17149,N_17263);
or U17798 (N_17798,N_17244,N_16955);
nor U17799 (N_17799,N_17354,N_17331);
and U17800 (N_17800,N_17467,N_17281);
and U17801 (N_17801,N_16876,N_17373);
xnor U17802 (N_17802,N_17146,N_17228);
or U17803 (N_17803,N_17368,N_17129);
nand U17804 (N_17804,N_17100,N_17454);
and U17805 (N_17805,N_16921,N_17340);
xnor U17806 (N_17806,N_17491,N_17004);
nor U17807 (N_17807,N_17456,N_16950);
and U17808 (N_17808,N_17284,N_16890);
xor U17809 (N_17809,N_17389,N_17151);
nand U17810 (N_17810,N_17379,N_17104);
nand U17811 (N_17811,N_17255,N_16881);
xor U17812 (N_17812,N_17038,N_17378);
or U17813 (N_17813,N_17394,N_17419);
nand U17814 (N_17814,N_16921,N_17194);
nor U17815 (N_17815,N_17021,N_17031);
or U17816 (N_17816,N_17186,N_17412);
nor U17817 (N_17817,N_16922,N_17033);
and U17818 (N_17818,N_17034,N_16923);
nand U17819 (N_17819,N_17177,N_17474);
nand U17820 (N_17820,N_17433,N_17087);
nand U17821 (N_17821,N_17037,N_17032);
nand U17822 (N_17822,N_17094,N_17116);
or U17823 (N_17823,N_16982,N_17173);
nand U17824 (N_17824,N_17205,N_17295);
or U17825 (N_17825,N_17432,N_17253);
and U17826 (N_17826,N_17430,N_17336);
xor U17827 (N_17827,N_17318,N_17236);
nor U17828 (N_17828,N_17004,N_17339);
xor U17829 (N_17829,N_17489,N_17440);
nand U17830 (N_17830,N_17383,N_17348);
and U17831 (N_17831,N_16984,N_17219);
and U17832 (N_17832,N_17201,N_17193);
xnor U17833 (N_17833,N_16929,N_17429);
and U17834 (N_17834,N_17213,N_17104);
xnor U17835 (N_17835,N_17241,N_17398);
and U17836 (N_17836,N_17102,N_17149);
nor U17837 (N_17837,N_17159,N_16968);
and U17838 (N_17838,N_17168,N_17208);
or U17839 (N_17839,N_17101,N_17445);
or U17840 (N_17840,N_17231,N_17120);
xor U17841 (N_17841,N_17051,N_17041);
or U17842 (N_17842,N_17329,N_16923);
nor U17843 (N_17843,N_17409,N_16921);
nand U17844 (N_17844,N_17351,N_17219);
nor U17845 (N_17845,N_17264,N_17391);
and U17846 (N_17846,N_17487,N_17104);
and U17847 (N_17847,N_17358,N_17246);
nand U17848 (N_17848,N_17005,N_17311);
and U17849 (N_17849,N_17450,N_17390);
nor U17850 (N_17850,N_17413,N_16957);
nand U17851 (N_17851,N_16977,N_16927);
or U17852 (N_17852,N_17337,N_16904);
or U17853 (N_17853,N_17448,N_17371);
nand U17854 (N_17854,N_17013,N_17046);
or U17855 (N_17855,N_17440,N_17474);
or U17856 (N_17856,N_16893,N_17224);
and U17857 (N_17857,N_17042,N_17133);
or U17858 (N_17858,N_16899,N_17474);
nand U17859 (N_17859,N_17433,N_17348);
nor U17860 (N_17860,N_16886,N_17086);
nor U17861 (N_17861,N_17357,N_16988);
and U17862 (N_17862,N_16990,N_17389);
xor U17863 (N_17863,N_17466,N_16982);
nor U17864 (N_17864,N_17297,N_16900);
nand U17865 (N_17865,N_17416,N_17147);
and U17866 (N_17866,N_17360,N_16963);
or U17867 (N_17867,N_17020,N_17065);
and U17868 (N_17868,N_17054,N_17228);
nor U17869 (N_17869,N_17386,N_17343);
or U17870 (N_17870,N_17071,N_17097);
xnor U17871 (N_17871,N_17371,N_17143);
or U17872 (N_17872,N_17480,N_17286);
xnor U17873 (N_17873,N_16921,N_17291);
and U17874 (N_17874,N_17468,N_17409);
nand U17875 (N_17875,N_17310,N_17272);
xnor U17876 (N_17876,N_17450,N_17470);
nor U17877 (N_17877,N_17057,N_16891);
or U17878 (N_17878,N_16969,N_17428);
or U17879 (N_17879,N_17372,N_17199);
nand U17880 (N_17880,N_17123,N_16899);
or U17881 (N_17881,N_17067,N_17487);
nor U17882 (N_17882,N_17369,N_17452);
nand U17883 (N_17883,N_17138,N_17441);
nand U17884 (N_17884,N_17456,N_16958);
nand U17885 (N_17885,N_17386,N_17078);
nand U17886 (N_17886,N_17165,N_17394);
nor U17887 (N_17887,N_16893,N_16878);
xor U17888 (N_17888,N_17132,N_17090);
xnor U17889 (N_17889,N_17289,N_17188);
nor U17890 (N_17890,N_17003,N_17469);
nor U17891 (N_17891,N_17427,N_17436);
and U17892 (N_17892,N_17292,N_17487);
xnor U17893 (N_17893,N_17072,N_16957);
or U17894 (N_17894,N_17252,N_17289);
or U17895 (N_17895,N_17185,N_17191);
nand U17896 (N_17896,N_17124,N_17463);
nor U17897 (N_17897,N_17075,N_16939);
nand U17898 (N_17898,N_17236,N_16891);
and U17899 (N_17899,N_17388,N_16947);
nor U17900 (N_17900,N_17333,N_17217);
or U17901 (N_17901,N_17220,N_17196);
or U17902 (N_17902,N_17042,N_16934);
nand U17903 (N_17903,N_17146,N_17221);
xor U17904 (N_17904,N_17481,N_16993);
nor U17905 (N_17905,N_17304,N_17375);
or U17906 (N_17906,N_16892,N_17298);
or U17907 (N_17907,N_17464,N_17438);
xnor U17908 (N_17908,N_17247,N_17408);
or U17909 (N_17909,N_17021,N_17353);
and U17910 (N_17910,N_17304,N_17119);
xor U17911 (N_17911,N_17106,N_17020);
or U17912 (N_17912,N_17425,N_17446);
nand U17913 (N_17913,N_16931,N_17276);
or U17914 (N_17914,N_16890,N_17222);
nand U17915 (N_17915,N_16879,N_17083);
and U17916 (N_17916,N_17491,N_17071);
nand U17917 (N_17917,N_17064,N_17250);
nand U17918 (N_17918,N_17402,N_17299);
xor U17919 (N_17919,N_17491,N_17295);
or U17920 (N_17920,N_17498,N_17247);
or U17921 (N_17921,N_17382,N_17012);
nand U17922 (N_17922,N_16900,N_17352);
nor U17923 (N_17923,N_17433,N_17143);
and U17924 (N_17924,N_17369,N_17314);
nand U17925 (N_17925,N_17194,N_17077);
and U17926 (N_17926,N_17015,N_17270);
nor U17927 (N_17927,N_16984,N_17187);
nand U17928 (N_17928,N_17324,N_17074);
xor U17929 (N_17929,N_17009,N_17378);
nor U17930 (N_17930,N_17418,N_17266);
nand U17931 (N_17931,N_16895,N_17378);
or U17932 (N_17932,N_17499,N_16928);
nor U17933 (N_17933,N_17293,N_16987);
and U17934 (N_17934,N_17344,N_17318);
nand U17935 (N_17935,N_17222,N_17232);
or U17936 (N_17936,N_16939,N_16975);
nand U17937 (N_17937,N_17429,N_17348);
nand U17938 (N_17938,N_17156,N_16951);
nor U17939 (N_17939,N_16994,N_17376);
and U17940 (N_17940,N_17042,N_17142);
nor U17941 (N_17941,N_17088,N_17363);
or U17942 (N_17942,N_17351,N_17019);
nand U17943 (N_17943,N_17345,N_16956);
xor U17944 (N_17944,N_17239,N_17160);
nor U17945 (N_17945,N_17456,N_17246);
xor U17946 (N_17946,N_16977,N_17342);
or U17947 (N_17947,N_16992,N_16916);
or U17948 (N_17948,N_17195,N_17356);
xnor U17949 (N_17949,N_17144,N_17152);
and U17950 (N_17950,N_17202,N_17200);
nand U17951 (N_17951,N_16915,N_17084);
xnor U17952 (N_17952,N_17372,N_17407);
nor U17953 (N_17953,N_16879,N_16904);
xor U17954 (N_17954,N_17482,N_17486);
and U17955 (N_17955,N_17409,N_17322);
nand U17956 (N_17956,N_16891,N_17023);
nand U17957 (N_17957,N_17214,N_16924);
nand U17958 (N_17958,N_17452,N_17246);
nand U17959 (N_17959,N_17266,N_17070);
or U17960 (N_17960,N_17060,N_17494);
xnor U17961 (N_17961,N_17212,N_17384);
or U17962 (N_17962,N_17245,N_17106);
and U17963 (N_17963,N_16997,N_16914);
nor U17964 (N_17964,N_17174,N_17350);
nand U17965 (N_17965,N_17193,N_17019);
or U17966 (N_17966,N_17275,N_17358);
nor U17967 (N_17967,N_17455,N_17371);
and U17968 (N_17968,N_16898,N_17065);
or U17969 (N_17969,N_16886,N_17267);
or U17970 (N_17970,N_17244,N_17207);
or U17971 (N_17971,N_16885,N_17040);
nor U17972 (N_17972,N_16972,N_17391);
xor U17973 (N_17973,N_16924,N_17240);
xnor U17974 (N_17974,N_17374,N_17378);
nand U17975 (N_17975,N_17428,N_17394);
and U17976 (N_17976,N_16924,N_16908);
nand U17977 (N_17977,N_17242,N_17002);
nand U17978 (N_17978,N_16884,N_17217);
nor U17979 (N_17979,N_17199,N_16983);
nor U17980 (N_17980,N_17429,N_17208);
or U17981 (N_17981,N_16938,N_17022);
or U17982 (N_17982,N_17144,N_17136);
nor U17983 (N_17983,N_17023,N_16997);
nand U17984 (N_17984,N_17081,N_17075);
xor U17985 (N_17985,N_17162,N_17229);
and U17986 (N_17986,N_16918,N_17028);
nand U17987 (N_17987,N_17387,N_16913);
and U17988 (N_17988,N_17455,N_16930);
and U17989 (N_17989,N_17169,N_17018);
and U17990 (N_17990,N_17296,N_16920);
and U17991 (N_17991,N_16911,N_17114);
and U17992 (N_17992,N_17022,N_17492);
nor U17993 (N_17993,N_16965,N_17218);
nand U17994 (N_17994,N_17481,N_17389);
nor U17995 (N_17995,N_17398,N_17056);
or U17996 (N_17996,N_17413,N_17227);
nand U17997 (N_17997,N_16974,N_17315);
nor U17998 (N_17998,N_17320,N_17166);
xor U17999 (N_17999,N_16902,N_16946);
and U18000 (N_18000,N_17164,N_17369);
nor U18001 (N_18001,N_17120,N_17488);
or U18002 (N_18002,N_17001,N_17229);
or U18003 (N_18003,N_16888,N_17169);
or U18004 (N_18004,N_17183,N_16937);
xnor U18005 (N_18005,N_16905,N_17407);
or U18006 (N_18006,N_17460,N_17275);
and U18007 (N_18007,N_17350,N_17090);
nand U18008 (N_18008,N_17113,N_17422);
or U18009 (N_18009,N_16981,N_17063);
and U18010 (N_18010,N_17268,N_17022);
nor U18011 (N_18011,N_17340,N_17123);
nand U18012 (N_18012,N_17085,N_16879);
and U18013 (N_18013,N_17166,N_17182);
nor U18014 (N_18014,N_16935,N_17318);
nand U18015 (N_18015,N_17355,N_17257);
or U18016 (N_18016,N_17345,N_17245);
or U18017 (N_18017,N_17034,N_16951);
or U18018 (N_18018,N_17436,N_17032);
xnor U18019 (N_18019,N_17154,N_17066);
xor U18020 (N_18020,N_17181,N_17069);
or U18021 (N_18021,N_16935,N_17229);
nand U18022 (N_18022,N_17300,N_17263);
xnor U18023 (N_18023,N_17065,N_17494);
and U18024 (N_18024,N_16956,N_17267);
or U18025 (N_18025,N_17411,N_17218);
nand U18026 (N_18026,N_16989,N_17369);
or U18027 (N_18027,N_17028,N_16932);
and U18028 (N_18028,N_17230,N_16992);
and U18029 (N_18029,N_17346,N_16927);
and U18030 (N_18030,N_17161,N_17215);
and U18031 (N_18031,N_17328,N_17265);
nand U18032 (N_18032,N_17118,N_17363);
or U18033 (N_18033,N_17137,N_16909);
and U18034 (N_18034,N_16921,N_17341);
xnor U18035 (N_18035,N_17442,N_17094);
nor U18036 (N_18036,N_17094,N_17326);
or U18037 (N_18037,N_17364,N_16941);
and U18038 (N_18038,N_17401,N_17299);
nor U18039 (N_18039,N_16912,N_17024);
nand U18040 (N_18040,N_17120,N_17201);
or U18041 (N_18041,N_17002,N_16983);
nand U18042 (N_18042,N_17046,N_17317);
or U18043 (N_18043,N_17386,N_17414);
and U18044 (N_18044,N_17061,N_17267);
nor U18045 (N_18045,N_17329,N_17256);
or U18046 (N_18046,N_17419,N_16968);
nand U18047 (N_18047,N_17315,N_17473);
nor U18048 (N_18048,N_17039,N_17105);
or U18049 (N_18049,N_17358,N_17203);
or U18050 (N_18050,N_16962,N_16957);
nand U18051 (N_18051,N_17312,N_17400);
nand U18052 (N_18052,N_17038,N_16925);
nand U18053 (N_18053,N_17378,N_17309);
nand U18054 (N_18054,N_16950,N_17471);
nand U18055 (N_18055,N_17179,N_17328);
nand U18056 (N_18056,N_17064,N_17277);
or U18057 (N_18057,N_17404,N_16985);
or U18058 (N_18058,N_17486,N_17143);
and U18059 (N_18059,N_17181,N_17015);
nor U18060 (N_18060,N_17213,N_17383);
nor U18061 (N_18061,N_17357,N_17347);
nand U18062 (N_18062,N_17215,N_17122);
nand U18063 (N_18063,N_17333,N_17316);
nor U18064 (N_18064,N_16979,N_17392);
nor U18065 (N_18065,N_17451,N_17114);
and U18066 (N_18066,N_17368,N_17053);
and U18067 (N_18067,N_16991,N_17452);
and U18068 (N_18068,N_16930,N_17449);
and U18069 (N_18069,N_17488,N_17101);
or U18070 (N_18070,N_17272,N_17018);
nand U18071 (N_18071,N_16948,N_16888);
or U18072 (N_18072,N_17417,N_17064);
and U18073 (N_18073,N_17066,N_17491);
or U18074 (N_18074,N_17495,N_17425);
nor U18075 (N_18075,N_16972,N_16884);
or U18076 (N_18076,N_16946,N_17039);
xnor U18077 (N_18077,N_17264,N_17064);
nor U18078 (N_18078,N_17382,N_17491);
nor U18079 (N_18079,N_16929,N_16931);
nor U18080 (N_18080,N_17272,N_17044);
and U18081 (N_18081,N_17283,N_17488);
xor U18082 (N_18082,N_17451,N_16898);
nand U18083 (N_18083,N_17351,N_17138);
or U18084 (N_18084,N_17291,N_17492);
and U18085 (N_18085,N_17395,N_17118);
nor U18086 (N_18086,N_17090,N_17410);
and U18087 (N_18087,N_17160,N_17046);
nand U18088 (N_18088,N_17156,N_17250);
xor U18089 (N_18089,N_17484,N_17007);
and U18090 (N_18090,N_17216,N_17088);
and U18091 (N_18091,N_16999,N_17296);
and U18092 (N_18092,N_17275,N_17111);
and U18093 (N_18093,N_17468,N_17342);
and U18094 (N_18094,N_17135,N_17329);
nor U18095 (N_18095,N_17196,N_16963);
nor U18096 (N_18096,N_17221,N_17131);
or U18097 (N_18097,N_17175,N_17022);
nor U18098 (N_18098,N_17308,N_17044);
or U18099 (N_18099,N_17376,N_17078);
or U18100 (N_18100,N_17245,N_17113);
or U18101 (N_18101,N_17169,N_17113);
and U18102 (N_18102,N_17095,N_17478);
xor U18103 (N_18103,N_17055,N_17136);
nor U18104 (N_18104,N_17008,N_17328);
nor U18105 (N_18105,N_17008,N_16880);
or U18106 (N_18106,N_17043,N_17268);
nor U18107 (N_18107,N_17024,N_17287);
xor U18108 (N_18108,N_17220,N_17431);
xnor U18109 (N_18109,N_17311,N_16977);
nor U18110 (N_18110,N_17049,N_17472);
xor U18111 (N_18111,N_17466,N_16959);
and U18112 (N_18112,N_17332,N_17149);
or U18113 (N_18113,N_17159,N_17278);
or U18114 (N_18114,N_17405,N_17395);
and U18115 (N_18115,N_17471,N_17165);
or U18116 (N_18116,N_16905,N_16996);
and U18117 (N_18117,N_17194,N_16886);
nand U18118 (N_18118,N_17269,N_16911);
or U18119 (N_18119,N_17476,N_17146);
or U18120 (N_18120,N_17120,N_17082);
xor U18121 (N_18121,N_17118,N_17227);
nor U18122 (N_18122,N_17016,N_16918);
and U18123 (N_18123,N_16946,N_17373);
nand U18124 (N_18124,N_16991,N_17152);
and U18125 (N_18125,N_17557,N_17836);
xnor U18126 (N_18126,N_17908,N_17930);
xnor U18127 (N_18127,N_17970,N_17582);
nand U18128 (N_18128,N_18091,N_17918);
and U18129 (N_18129,N_17821,N_17719);
nand U18130 (N_18130,N_17548,N_17617);
nand U18131 (N_18131,N_17656,N_17576);
nand U18132 (N_18132,N_17827,N_17929);
or U18133 (N_18133,N_17839,N_18029);
or U18134 (N_18134,N_17952,N_17990);
xnor U18135 (N_18135,N_17607,N_18115);
or U18136 (N_18136,N_17815,N_17636);
nand U18137 (N_18137,N_17530,N_17851);
and U18138 (N_18138,N_18035,N_18064);
nor U18139 (N_18139,N_17740,N_17692);
or U18140 (N_18140,N_17822,N_17893);
nand U18141 (N_18141,N_17599,N_17524);
and U18142 (N_18142,N_18004,N_17956);
xor U18143 (N_18143,N_17537,N_17872);
xor U18144 (N_18144,N_17529,N_17534);
or U18145 (N_18145,N_18097,N_17980);
nor U18146 (N_18146,N_18065,N_17566);
nand U18147 (N_18147,N_17921,N_17977);
xor U18148 (N_18148,N_17514,N_17632);
xnor U18149 (N_18149,N_17637,N_17809);
nor U18150 (N_18150,N_18015,N_17666);
and U18151 (N_18151,N_18075,N_17759);
and U18152 (N_18152,N_17650,N_18051);
and U18153 (N_18153,N_18063,N_18036);
nand U18154 (N_18154,N_17609,N_17782);
xnor U18155 (N_18155,N_18016,N_17832);
xnor U18156 (N_18156,N_17813,N_18095);
and U18157 (N_18157,N_17902,N_17628);
nand U18158 (N_18158,N_17506,N_17954);
nand U18159 (N_18159,N_17849,N_17772);
and U18160 (N_18160,N_17941,N_17885);
nor U18161 (N_18161,N_17794,N_18005);
or U18162 (N_18162,N_18041,N_18020);
nand U18163 (N_18163,N_17743,N_17861);
nand U18164 (N_18164,N_18000,N_17526);
nor U18165 (N_18165,N_17671,N_17659);
or U18166 (N_18166,N_17838,N_18014);
nor U18167 (N_18167,N_17716,N_17700);
and U18168 (N_18168,N_18072,N_18059);
and U18169 (N_18169,N_18050,N_17555);
xnor U18170 (N_18170,N_17604,N_17735);
nor U18171 (N_18171,N_17638,N_18113);
nor U18172 (N_18172,N_17586,N_18011);
nand U18173 (N_18173,N_17926,N_17748);
xnor U18174 (N_18174,N_18106,N_17799);
nor U18175 (N_18175,N_18066,N_17792);
nand U18176 (N_18176,N_17697,N_17855);
nor U18177 (N_18177,N_17718,N_17664);
nor U18178 (N_18178,N_18112,N_17767);
nor U18179 (N_18179,N_17684,N_17900);
nand U18180 (N_18180,N_18100,N_17592);
xnor U18181 (N_18181,N_17940,N_17979);
and U18182 (N_18182,N_17909,N_18105);
xor U18183 (N_18183,N_17906,N_17876);
nor U18184 (N_18184,N_17840,N_18068);
xor U18185 (N_18185,N_17711,N_17846);
nor U18186 (N_18186,N_17695,N_17841);
nor U18187 (N_18187,N_18027,N_18052);
or U18188 (N_18188,N_17866,N_17919);
nor U18189 (N_18189,N_17675,N_17608);
and U18190 (N_18190,N_18096,N_17795);
and U18191 (N_18191,N_17683,N_17696);
and U18192 (N_18192,N_17550,N_17913);
xor U18193 (N_18193,N_17594,N_17669);
xnor U18194 (N_18194,N_17646,N_18071);
xor U18195 (N_18195,N_18053,N_17976);
nor U18196 (N_18196,N_17710,N_17528);
or U18197 (N_18197,N_18006,N_17639);
and U18198 (N_18198,N_17925,N_17654);
xnor U18199 (N_18199,N_17867,N_18087);
xor U18200 (N_18200,N_17972,N_17706);
nand U18201 (N_18201,N_17641,N_17755);
and U18202 (N_18202,N_17691,N_18002);
nor U18203 (N_18203,N_17904,N_17510);
and U18204 (N_18204,N_17721,N_17613);
xnor U18205 (N_18205,N_17982,N_17801);
nand U18206 (N_18206,N_18108,N_17788);
nand U18207 (N_18207,N_17729,N_18069);
xnor U18208 (N_18208,N_17544,N_17583);
xnor U18209 (N_18209,N_17842,N_17648);
and U18210 (N_18210,N_17560,N_17702);
and U18211 (N_18211,N_17728,N_17730);
and U18212 (N_18212,N_17854,N_17917);
or U18213 (N_18213,N_17749,N_18062);
nand U18214 (N_18214,N_17516,N_17665);
xor U18215 (N_18215,N_17989,N_17525);
nand U18216 (N_18216,N_17533,N_17668);
and U18217 (N_18217,N_17810,N_17873);
or U18218 (N_18218,N_17717,N_17947);
nand U18219 (N_18219,N_17546,N_18093);
xor U18220 (N_18220,N_18074,N_17833);
and U18221 (N_18221,N_17674,N_18025);
or U18222 (N_18222,N_17737,N_17698);
or U18223 (N_18223,N_17511,N_18099);
and U18224 (N_18224,N_18111,N_17614);
nand U18225 (N_18225,N_17817,N_17657);
xnor U18226 (N_18226,N_17574,N_17722);
nor U18227 (N_18227,N_17881,N_17766);
or U18228 (N_18228,N_18120,N_17714);
nand U18229 (N_18229,N_17553,N_18049);
nand U18230 (N_18230,N_18008,N_17770);
and U18231 (N_18231,N_17741,N_17775);
nor U18232 (N_18232,N_17850,N_18023);
xnor U18233 (N_18233,N_17727,N_17967);
and U18234 (N_18234,N_17581,N_17680);
xor U18235 (N_18235,N_17959,N_17898);
nand U18236 (N_18236,N_17883,N_17603);
nor U18237 (N_18237,N_17595,N_18033);
xnor U18238 (N_18238,N_17814,N_17760);
or U18239 (N_18239,N_17720,N_17757);
xnor U18240 (N_18240,N_17862,N_17562);
nor U18241 (N_18241,N_17563,N_17658);
or U18242 (N_18242,N_18037,N_17521);
nand U18243 (N_18243,N_17573,N_17556);
or U18244 (N_18244,N_17865,N_18076);
xor U18245 (N_18245,N_17784,N_17914);
nor U18246 (N_18246,N_17884,N_17983);
xnor U18247 (N_18247,N_17903,N_17931);
or U18248 (N_18248,N_17723,N_17611);
nor U18249 (N_18249,N_17958,N_17783);
xnor U18250 (N_18250,N_18085,N_17747);
nand U18251 (N_18251,N_17762,N_18101);
nor U18252 (N_18252,N_17629,N_17523);
xnor U18253 (N_18253,N_17874,N_17540);
or U18254 (N_18254,N_17853,N_17732);
and U18255 (N_18255,N_17785,N_18084);
nand U18256 (N_18256,N_17974,N_17907);
or U18257 (N_18257,N_18047,N_18019);
and U18258 (N_18258,N_17942,N_17824);
nand U18259 (N_18259,N_17704,N_17751);
and U18260 (N_18260,N_17500,N_17960);
or U18261 (N_18261,N_18022,N_18104);
and U18262 (N_18262,N_17763,N_17912);
xor U18263 (N_18263,N_17645,N_17731);
or U18264 (N_18264,N_17996,N_17713);
nand U18265 (N_18265,N_17803,N_18092);
and U18266 (N_18266,N_18042,N_17891);
nand U18267 (N_18267,N_17619,N_17955);
nor U18268 (N_18268,N_17764,N_17975);
nand U18269 (N_18269,N_17808,N_17519);
nor U18270 (N_18270,N_18030,N_17936);
xnor U18271 (N_18271,N_17777,N_17937);
and U18272 (N_18272,N_18046,N_17834);
or U18273 (N_18273,N_18124,N_18078);
or U18274 (N_18274,N_17949,N_18054);
nor U18275 (N_18275,N_17831,N_18057);
or U18276 (N_18276,N_18056,N_18028);
nand U18277 (N_18277,N_17779,N_17640);
xor U18278 (N_18278,N_17991,N_17542);
or U18279 (N_18279,N_17590,N_17739);
nor U18280 (N_18280,N_17580,N_17651);
nand U18281 (N_18281,N_17986,N_17627);
nand U18282 (N_18282,N_17830,N_17559);
or U18283 (N_18283,N_18055,N_17998);
xnor U18284 (N_18284,N_18079,N_17642);
nor U18285 (N_18285,N_17859,N_17758);
nand U18286 (N_18286,N_17802,N_17950);
nor U18287 (N_18287,N_17899,N_17892);
and U18288 (N_18288,N_17826,N_17571);
or U18289 (N_18289,N_18012,N_17520);
and U18290 (N_18290,N_17857,N_17856);
nor U18291 (N_18291,N_17828,N_17987);
nand U18292 (N_18292,N_17752,N_17943);
xnor U18293 (N_18293,N_17558,N_17549);
or U18294 (N_18294,N_17633,N_17522);
or U18295 (N_18295,N_17791,N_18088);
and U18296 (N_18296,N_17561,N_17689);
and U18297 (N_18297,N_17649,N_17685);
nand U18298 (N_18298,N_17825,N_17660);
nand U18299 (N_18299,N_17835,N_17630);
nor U18300 (N_18300,N_17963,N_17682);
or U18301 (N_18301,N_17678,N_17786);
or U18302 (N_18302,N_18090,N_17769);
nor U18303 (N_18303,N_17591,N_18122);
xnor U18304 (N_18304,N_17733,N_18003);
xor U18305 (N_18305,N_17570,N_17602);
nand U18306 (N_18306,N_17889,N_17897);
nor U18307 (N_18307,N_17634,N_18089);
and U18308 (N_18308,N_17653,N_17806);
and U18309 (N_18309,N_17864,N_17596);
or U18310 (N_18310,N_17644,N_17616);
xor U18311 (N_18311,N_17667,N_17819);
and U18312 (N_18312,N_17858,N_17852);
and U18313 (N_18313,N_17672,N_17957);
or U18314 (N_18314,N_17652,N_17552);
nand U18315 (N_18315,N_18116,N_17501);
or U18316 (N_18316,N_17915,N_17539);
xor U18317 (N_18317,N_18048,N_18107);
xor U18318 (N_18318,N_17545,N_17860);
and U18319 (N_18319,N_17875,N_18094);
nor U18320 (N_18320,N_18018,N_17820);
xor U18321 (N_18321,N_17890,N_17527);
nand U18322 (N_18322,N_17938,N_17978);
xor U18323 (N_18323,N_18123,N_17910);
xor U18324 (N_18324,N_17575,N_17726);
and U18325 (N_18325,N_17886,N_17804);
nor U18326 (N_18326,N_17724,N_17536);
nand U18327 (N_18327,N_17997,N_17626);
or U18328 (N_18328,N_18017,N_17948);
and U18329 (N_18329,N_17871,N_17584);
nor U18330 (N_18330,N_17703,N_17934);
and U18331 (N_18331,N_17712,N_17631);
nor U18332 (N_18332,N_17935,N_17887);
nor U18333 (N_18333,N_17811,N_17756);
xor U18334 (N_18334,N_18032,N_18026);
and U18335 (N_18335,N_17916,N_18117);
nand U18336 (N_18336,N_17746,N_17734);
nor U18337 (N_18337,N_17961,N_18010);
xnor U18338 (N_18338,N_17964,N_17965);
or U18339 (N_18339,N_17688,N_17508);
nor U18340 (N_18340,N_17681,N_17988);
or U18341 (N_18341,N_17620,N_17993);
or U18342 (N_18342,N_17635,N_17715);
xor U18343 (N_18343,N_17612,N_17837);
xor U18344 (N_18344,N_17600,N_18083);
xor U18345 (N_18345,N_17781,N_17677);
or U18346 (N_18346,N_17823,N_17878);
or U18347 (N_18347,N_17554,N_17693);
and U18348 (N_18348,N_17798,N_18118);
nand U18349 (N_18349,N_17761,N_17572);
xnor U18350 (N_18350,N_17778,N_17922);
nor U18351 (N_18351,N_17610,N_18058);
nor U18352 (N_18352,N_17844,N_17984);
nor U18353 (N_18353,N_17962,N_17845);
nand U18354 (N_18354,N_17927,N_17694);
and U18355 (N_18355,N_17968,N_17622);
xnor U18356 (N_18356,N_17701,N_18110);
or U18357 (N_18357,N_17509,N_17789);
nor U18358 (N_18358,N_17992,N_17655);
nor U18359 (N_18359,N_17621,N_17805);
xnor U18360 (N_18360,N_17597,N_17933);
nor U18361 (N_18361,N_17971,N_17924);
xor U18362 (N_18362,N_17797,N_17848);
or U18363 (N_18363,N_18098,N_17870);
xor U18364 (N_18364,N_18103,N_17829);
and U18365 (N_18365,N_18102,N_17538);
and U18366 (N_18366,N_17565,N_17793);
xor U18367 (N_18367,N_17507,N_17882);
nand U18368 (N_18368,N_17880,N_17796);
or U18369 (N_18369,N_17615,N_17503);
or U18370 (N_18370,N_17624,N_18045);
and U18371 (N_18371,N_17547,N_18081);
nor U18372 (N_18372,N_17567,N_17946);
nor U18373 (N_18373,N_18060,N_17568);
nor U18374 (N_18374,N_17699,N_17773);
or U18375 (N_18375,N_17888,N_18001);
nand U18376 (N_18376,N_17995,N_18073);
nand U18377 (N_18377,N_17745,N_18119);
or U18378 (N_18378,N_17541,N_17593);
or U18379 (N_18379,N_17515,N_17736);
nor U18380 (N_18380,N_17939,N_17725);
xor U18381 (N_18381,N_17847,N_18077);
or U18382 (N_18382,N_17768,N_17589);
xor U18383 (N_18383,N_18007,N_18114);
nand U18384 (N_18384,N_17673,N_18040);
or U18385 (N_18385,N_17690,N_17800);
or U18386 (N_18386,N_17754,N_17843);
nand U18387 (N_18387,N_18034,N_17569);
xor U18388 (N_18388,N_17863,N_17807);
xor U18389 (N_18389,N_17738,N_17513);
nor U18390 (N_18390,N_17578,N_17894);
nand U18391 (N_18391,N_17517,N_17643);
nor U18392 (N_18392,N_17744,N_17812);
nor U18393 (N_18393,N_18013,N_17911);
nor U18394 (N_18394,N_18043,N_17901);
nand U18395 (N_18395,N_17750,N_18024);
nand U18396 (N_18396,N_17647,N_17780);
nor U18397 (N_18397,N_17869,N_17601);
nand U18398 (N_18398,N_17928,N_17535);
nand U18399 (N_18399,N_18044,N_17505);
and U18400 (N_18400,N_17709,N_17923);
nand U18401 (N_18401,N_17816,N_17588);
nand U18402 (N_18402,N_17905,N_17945);
nor U18403 (N_18403,N_17551,N_17504);
xor U18404 (N_18404,N_17973,N_17577);
nor U18405 (N_18405,N_17765,N_17896);
nand U18406 (N_18406,N_17679,N_17686);
or U18407 (N_18407,N_18109,N_17774);
and U18408 (N_18408,N_17502,N_17951);
nand U18409 (N_18409,N_17981,N_17787);
xor U18410 (N_18410,N_17985,N_17771);
or U18411 (N_18411,N_18080,N_17944);
nor U18412 (N_18412,N_17753,N_17868);
nor U18413 (N_18413,N_17687,N_18039);
xor U18414 (N_18414,N_18082,N_18070);
xor U18415 (N_18415,N_18031,N_17877);
and U18416 (N_18416,N_17623,N_17895);
and U18417 (N_18417,N_17966,N_17705);
nor U18418 (N_18418,N_18021,N_18061);
nor U18419 (N_18419,N_18121,N_17598);
nor U18420 (N_18420,N_17543,N_17776);
xor U18421 (N_18421,N_17625,N_17662);
or U18422 (N_18422,N_17707,N_17605);
xor U18423 (N_18423,N_17531,N_17670);
nand U18424 (N_18424,N_17994,N_17579);
xor U18425 (N_18425,N_17676,N_17618);
nand U18426 (N_18426,N_17518,N_17953);
or U18427 (N_18427,N_17790,N_17708);
xor U18428 (N_18428,N_17879,N_18038);
or U18429 (N_18429,N_18086,N_17564);
or U18430 (N_18430,N_17920,N_18067);
nor U18431 (N_18431,N_17663,N_17818);
nor U18432 (N_18432,N_17512,N_17532);
and U18433 (N_18433,N_18009,N_17587);
nor U18434 (N_18434,N_17606,N_17661);
and U18435 (N_18435,N_17999,N_17742);
nand U18436 (N_18436,N_17585,N_17932);
nand U18437 (N_18437,N_17969,N_17819);
xor U18438 (N_18438,N_17769,N_18026);
and U18439 (N_18439,N_17506,N_17592);
or U18440 (N_18440,N_18085,N_17711);
xor U18441 (N_18441,N_17899,N_18028);
xor U18442 (N_18442,N_17699,N_17805);
xor U18443 (N_18443,N_18104,N_18014);
and U18444 (N_18444,N_17837,N_17785);
or U18445 (N_18445,N_17933,N_18023);
and U18446 (N_18446,N_17564,N_17877);
xor U18447 (N_18447,N_18011,N_17592);
or U18448 (N_18448,N_18093,N_17717);
nor U18449 (N_18449,N_17611,N_18107);
and U18450 (N_18450,N_17813,N_18100);
nor U18451 (N_18451,N_17932,N_17870);
xnor U18452 (N_18452,N_18019,N_17837);
nand U18453 (N_18453,N_17734,N_17690);
nand U18454 (N_18454,N_18017,N_17666);
nor U18455 (N_18455,N_18055,N_17530);
and U18456 (N_18456,N_17785,N_17973);
and U18457 (N_18457,N_18106,N_17570);
nand U18458 (N_18458,N_17689,N_17669);
and U18459 (N_18459,N_17862,N_18004);
xnor U18460 (N_18460,N_17992,N_18017);
xor U18461 (N_18461,N_17630,N_17583);
and U18462 (N_18462,N_17604,N_17782);
or U18463 (N_18463,N_17822,N_17597);
and U18464 (N_18464,N_17904,N_18113);
nand U18465 (N_18465,N_18059,N_17879);
and U18466 (N_18466,N_17530,N_17777);
nand U18467 (N_18467,N_17630,N_17723);
or U18468 (N_18468,N_17974,N_17592);
nor U18469 (N_18469,N_17728,N_18055);
nand U18470 (N_18470,N_17643,N_17562);
or U18471 (N_18471,N_17867,N_17706);
nor U18472 (N_18472,N_17576,N_18089);
nand U18473 (N_18473,N_18016,N_17713);
nand U18474 (N_18474,N_17754,N_17547);
nor U18475 (N_18475,N_17647,N_18065);
nor U18476 (N_18476,N_17705,N_18080);
or U18477 (N_18477,N_17569,N_17974);
nor U18478 (N_18478,N_18029,N_17986);
xor U18479 (N_18479,N_17739,N_17832);
xor U18480 (N_18480,N_17959,N_17652);
or U18481 (N_18481,N_17760,N_17714);
or U18482 (N_18482,N_17975,N_17822);
xor U18483 (N_18483,N_17809,N_17939);
or U18484 (N_18484,N_17959,N_17631);
nand U18485 (N_18485,N_17824,N_17761);
nand U18486 (N_18486,N_17756,N_18032);
nand U18487 (N_18487,N_17823,N_17665);
nor U18488 (N_18488,N_17961,N_17571);
nand U18489 (N_18489,N_17545,N_17686);
xnor U18490 (N_18490,N_17557,N_17911);
xor U18491 (N_18491,N_17506,N_17719);
or U18492 (N_18492,N_18042,N_17626);
and U18493 (N_18493,N_17575,N_17584);
and U18494 (N_18494,N_17812,N_17786);
or U18495 (N_18495,N_18067,N_17645);
xor U18496 (N_18496,N_17983,N_17657);
and U18497 (N_18497,N_18115,N_17730);
nor U18498 (N_18498,N_17651,N_17819);
or U18499 (N_18499,N_17904,N_17564);
xor U18500 (N_18500,N_17959,N_18102);
nor U18501 (N_18501,N_17963,N_17529);
and U18502 (N_18502,N_17556,N_17895);
nor U18503 (N_18503,N_17990,N_17645);
and U18504 (N_18504,N_18057,N_17581);
or U18505 (N_18505,N_17953,N_18088);
or U18506 (N_18506,N_17907,N_18117);
xor U18507 (N_18507,N_17786,N_18120);
nor U18508 (N_18508,N_17733,N_17774);
or U18509 (N_18509,N_17796,N_17672);
nand U18510 (N_18510,N_18016,N_17981);
and U18511 (N_18511,N_17910,N_17618);
xor U18512 (N_18512,N_17515,N_17966);
nand U18513 (N_18513,N_17820,N_17537);
nor U18514 (N_18514,N_17938,N_17620);
xor U18515 (N_18515,N_17918,N_18096);
or U18516 (N_18516,N_17976,N_17588);
and U18517 (N_18517,N_17640,N_17937);
nor U18518 (N_18518,N_17620,N_18110);
xnor U18519 (N_18519,N_17680,N_17883);
or U18520 (N_18520,N_18020,N_18099);
xnor U18521 (N_18521,N_17847,N_18038);
nor U18522 (N_18522,N_17710,N_17825);
nor U18523 (N_18523,N_17535,N_17603);
and U18524 (N_18524,N_17567,N_17922);
xnor U18525 (N_18525,N_17925,N_17851);
nand U18526 (N_18526,N_18009,N_18015);
or U18527 (N_18527,N_17708,N_17548);
or U18528 (N_18528,N_17855,N_17545);
xor U18529 (N_18529,N_17704,N_17703);
nor U18530 (N_18530,N_17868,N_17919);
xnor U18531 (N_18531,N_17693,N_17742);
nor U18532 (N_18532,N_17558,N_17557);
and U18533 (N_18533,N_17734,N_18057);
xor U18534 (N_18534,N_17722,N_17956);
and U18535 (N_18535,N_17953,N_18032);
or U18536 (N_18536,N_18072,N_17697);
xnor U18537 (N_18537,N_17972,N_17746);
nand U18538 (N_18538,N_17806,N_17968);
and U18539 (N_18539,N_17696,N_18122);
nand U18540 (N_18540,N_17877,N_17857);
xnor U18541 (N_18541,N_18059,N_17947);
xnor U18542 (N_18542,N_17578,N_17954);
nor U18543 (N_18543,N_17946,N_17962);
nand U18544 (N_18544,N_17946,N_17600);
or U18545 (N_18545,N_17722,N_17616);
nand U18546 (N_18546,N_17577,N_18072);
and U18547 (N_18547,N_17708,N_17779);
nand U18548 (N_18548,N_17827,N_17683);
xor U18549 (N_18549,N_17985,N_17628);
and U18550 (N_18550,N_17789,N_18041);
or U18551 (N_18551,N_17963,N_17944);
or U18552 (N_18552,N_17862,N_17589);
nand U18553 (N_18553,N_17620,N_18094);
xnor U18554 (N_18554,N_17609,N_17924);
xnor U18555 (N_18555,N_17744,N_17642);
nand U18556 (N_18556,N_18094,N_18008);
xor U18557 (N_18557,N_17699,N_17520);
and U18558 (N_18558,N_17629,N_17502);
or U18559 (N_18559,N_17772,N_18074);
nand U18560 (N_18560,N_17529,N_18108);
or U18561 (N_18561,N_17985,N_17939);
and U18562 (N_18562,N_17761,N_17587);
nor U18563 (N_18563,N_17947,N_17626);
nor U18564 (N_18564,N_18051,N_17665);
nor U18565 (N_18565,N_17771,N_18070);
xor U18566 (N_18566,N_17812,N_17791);
or U18567 (N_18567,N_18063,N_17826);
nand U18568 (N_18568,N_17908,N_17517);
nor U18569 (N_18569,N_17514,N_18085);
xor U18570 (N_18570,N_17660,N_17880);
xnor U18571 (N_18571,N_17830,N_17999);
or U18572 (N_18572,N_17968,N_17765);
or U18573 (N_18573,N_17969,N_18046);
and U18574 (N_18574,N_17656,N_17626);
xor U18575 (N_18575,N_18034,N_17670);
and U18576 (N_18576,N_17522,N_17558);
nor U18577 (N_18577,N_17711,N_17940);
or U18578 (N_18578,N_17818,N_17737);
or U18579 (N_18579,N_17637,N_17568);
xnor U18580 (N_18580,N_17832,N_17638);
and U18581 (N_18581,N_18070,N_17559);
nor U18582 (N_18582,N_17658,N_17625);
nor U18583 (N_18583,N_17827,N_18085);
or U18584 (N_18584,N_17997,N_17893);
and U18585 (N_18585,N_17979,N_18031);
or U18586 (N_18586,N_17620,N_18074);
nand U18587 (N_18587,N_17838,N_17835);
nand U18588 (N_18588,N_18110,N_17902);
xnor U18589 (N_18589,N_17586,N_18053);
or U18590 (N_18590,N_17772,N_18107);
and U18591 (N_18591,N_17855,N_17563);
xor U18592 (N_18592,N_17547,N_18020);
and U18593 (N_18593,N_18083,N_17724);
and U18594 (N_18594,N_17577,N_17519);
xnor U18595 (N_18595,N_17785,N_17502);
nand U18596 (N_18596,N_17803,N_17585);
xnor U18597 (N_18597,N_17655,N_17616);
and U18598 (N_18598,N_17894,N_17674);
nor U18599 (N_18599,N_17923,N_17914);
or U18600 (N_18600,N_17999,N_17934);
nand U18601 (N_18601,N_17699,N_17659);
or U18602 (N_18602,N_17980,N_17831);
and U18603 (N_18603,N_17818,N_17725);
nor U18604 (N_18604,N_18028,N_17613);
xor U18605 (N_18605,N_17969,N_17703);
xnor U18606 (N_18606,N_17877,N_18052);
xor U18607 (N_18607,N_17823,N_17831);
nand U18608 (N_18608,N_17852,N_17889);
or U18609 (N_18609,N_17605,N_17803);
nand U18610 (N_18610,N_17576,N_18074);
or U18611 (N_18611,N_17546,N_18004);
nor U18612 (N_18612,N_17625,N_17708);
nor U18613 (N_18613,N_17649,N_17779);
xor U18614 (N_18614,N_17918,N_17562);
nand U18615 (N_18615,N_17601,N_17814);
nand U18616 (N_18616,N_17708,N_17566);
nor U18617 (N_18617,N_17593,N_17914);
or U18618 (N_18618,N_17772,N_17588);
and U18619 (N_18619,N_17752,N_17788);
xnor U18620 (N_18620,N_17675,N_18032);
nand U18621 (N_18621,N_18025,N_17976);
nor U18622 (N_18622,N_17884,N_17988);
or U18623 (N_18623,N_17873,N_17675);
xor U18624 (N_18624,N_17757,N_17996);
or U18625 (N_18625,N_17816,N_18004);
nand U18626 (N_18626,N_17540,N_17586);
or U18627 (N_18627,N_18070,N_17519);
xor U18628 (N_18628,N_17873,N_17620);
xor U18629 (N_18629,N_18071,N_17600);
and U18630 (N_18630,N_17975,N_17891);
nand U18631 (N_18631,N_17698,N_17748);
xnor U18632 (N_18632,N_18012,N_17685);
and U18633 (N_18633,N_17842,N_17660);
xnor U18634 (N_18634,N_17837,N_17712);
xnor U18635 (N_18635,N_17562,N_17682);
nand U18636 (N_18636,N_18027,N_18045);
nor U18637 (N_18637,N_18103,N_17555);
nand U18638 (N_18638,N_18078,N_17909);
nand U18639 (N_18639,N_17851,N_18114);
xor U18640 (N_18640,N_18070,N_17629);
or U18641 (N_18641,N_17578,N_17875);
xnor U18642 (N_18642,N_17680,N_17650);
or U18643 (N_18643,N_18085,N_17741);
or U18644 (N_18644,N_17638,N_17679);
or U18645 (N_18645,N_17763,N_17590);
and U18646 (N_18646,N_17948,N_17852);
or U18647 (N_18647,N_17518,N_17895);
nand U18648 (N_18648,N_17873,N_18012);
nor U18649 (N_18649,N_17763,N_17545);
nor U18650 (N_18650,N_18119,N_18040);
nor U18651 (N_18651,N_17776,N_18067);
xor U18652 (N_18652,N_17860,N_17573);
nor U18653 (N_18653,N_17877,N_18033);
or U18654 (N_18654,N_17510,N_18033);
nand U18655 (N_18655,N_17602,N_17556);
xnor U18656 (N_18656,N_18068,N_18015);
nand U18657 (N_18657,N_18010,N_17955);
nor U18658 (N_18658,N_17938,N_17864);
or U18659 (N_18659,N_17994,N_17684);
xnor U18660 (N_18660,N_17766,N_17508);
or U18661 (N_18661,N_17809,N_17842);
nand U18662 (N_18662,N_17598,N_17655);
nor U18663 (N_18663,N_17715,N_17796);
or U18664 (N_18664,N_18045,N_17607);
or U18665 (N_18665,N_17648,N_17613);
and U18666 (N_18666,N_17846,N_17814);
and U18667 (N_18667,N_17605,N_17945);
nand U18668 (N_18668,N_17684,N_17933);
or U18669 (N_18669,N_18047,N_17809);
and U18670 (N_18670,N_18044,N_17922);
xnor U18671 (N_18671,N_17786,N_17782);
and U18672 (N_18672,N_17825,N_17581);
nor U18673 (N_18673,N_17783,N_17725);
nand U18674 (N_18674,N_17636,N_18058);
or U18675 (N_18675,N_18088,N_17572);
and U18676 (N_18676,N_17865,N_17531);
nor U18677 (N_18677,N_18101,N_17656);
or U18678 (N_18678,N_17511,N_17858);
nor U18679 (N_18679,N_17691,N_17912);
nor U18680 (N_18680,N_17814,N_17658);
nor U18681 (N_18681,N_17804,N_17864);
or U18682 (N_18682,N_17842,N_18025);
nor U18683 (N_18683,N_17703,N_17780);
xnor U18684 (N_18684,N_17716,N_17991);
nor U18685 (N_18685,N_17987,N_17915);
and U18686 (N_18686,N_18120,N_17565);
xnor U18687 (N_18687,N_17546,N_17767);
and U18688 (N_18688,N_18045,N_17570);
nand U18689 (N_18689,N_17549,N_17647);
nor U18690 (N_18690,N_17894,N_18111);
nand U18691 (N_18691,N_18013,N_17774);
or U18692 (N_18692,N_17787,N_17829);
or U18693 (N_18693,N_17930,N_18100);
nand U18694 (N_18694,N_17836,N_17619);
xor U18695 (N_18695,N_17622,N_17601);
nand U18696 (N_18696,N_17950,N_17627);
xnor U18697 (N_18697,N_17801,N_17983);
nor U18698 (N_18698,N_17951,N_18106);
or U18699 (N_18699,N_17743,N_17841);
nand U18700 (N_18700,N_17972,N_17605);
or U18701 (N_18701,N_17735,N_17812);
nor U18702 (N_18702,N_17786,N_17642);
and U18703 (N_18703,N_17846,N_17610);
nor U18704 (N_18704,N_18055,N_17967);
or U18705 (N_18705,N_17895,N_17776);
xor U18706 (N_18706,N_17928,N_17670);
nand U18707 (N_18707,N_17530,N_18116);
and U18708 (N_18708,N_18013,N_17763);
xnor U18709 (N_18709,N_17546,N_18040);
nand U18710 (N_18710,N_18016,N_17653);
nor U18711 (N_18711,N_17599,N_17706);
xor U18712 (N_18712,N_18112,N_17926);
and U18713 (N_18713,N_17681,N_18034);
nor U18714 (N_18714,N_17758,N_17631);
or U18715 (N_18715,N_17503,N_17680);
and U18716 (N_18716,N_17566,N_17504);
or U18717 (N_18717,N_17974,N_17792);
nand U18718 (N_18718,N_17529,N_17807);
nand U18719 (N_18719,N_17937,N_17667);
nand U18720 (N_18720,N_17624,N_17979);
or U18721 (N_18721,N_17867,N_17556);
or U18722 (N_18722,N_17727,N_18032);
nor U18723 (N_18723,N_17532,N_17668);
or U18724 (N_18724,N_18000,N_17753);
nor U18725 (N_18725,N_17759,N_18124);
and U18726 (N_18726,N_17721,N_17757);
xnor U18727 (N_18727,N_17864,N_17628);
nand U18728 (N_18728,N_17714,N_17945);
xor U18729 (N_18729,N_17722,N_17914);
or U18730 (N_18730,N_17540,N_17918);
and U18731 (N_18731,N_17938,N_18104);
xor U18732 (N_18732,N_17810,N_17988);
or U18733 (N_18733,N_18115,N_17881);
and U18734 (N_18734,N_18059,N_18015);
or U18735 (N_18735,N_17824,N_17519);
or U18736 (N_18736,N_17991,N_18105);
nand U18737 (N_18737,N_17558,N_17897);
nor U18738 (N_18738,N_17872,N_18016);
and U18739 (N_18739,N_17619,N_17828);
or U18740 (N_18740,N_17896,N_17645);
nor U18741 (N_18741,N_18013,N_17507);
and U18742 (N_18742,N_17612,N_17624);
xnor U18743 (N_18743,N_17663,N_17830);
or U18744 (N_18744,N_17525,N_17511);
and U18745 (N_18745,N_18029,N_17964);
xnor U18746 (N_18746,N_17735,N_17792);
nand U18747 (N_18747,N_17581,N_17977);
nor U18748 (N_18748,N_17666,N_17880);
or U18749 (N_18749,N_17540,N_17807);
xnor U18750 (N_18750,N_18446,N_18306);
and U18751 (N_18751,N_18723,N_18683);
nor U18752 (N_18752,N_18496,N_18200);
nand U18753 (N_18753,N_18272,N_18587);
nand U18754 (N_18754,N_18583,N_18475);
or U18755 (N_18755,N_18418,N_18642);
nor U18756 (N_18756,N_18665,N_18623);
xnor U18757 (N_18757,N_18342,N_18182);
nand U18758 (N_18758,N_18327,N_18678);
xnor U18759 (N_18759,N_18749,N_18478);
xor U18760 (N_18760,N_18682,N_18740);
nor U18761 (N_18761,N_18181,N_18634);
or U18762 (N_18762,N_18132,N_18442);
nand U18763 (N_18763,N_18133,N_18258);
nor U18764 (N_18764,N_18491,N_18397);
xor U18765 (N_18765,N_18308,N_18325);
and U18766 (N_18766,N_18138,N_18169);
or U18767 (N_18767,N_18193,N_18404);
xnor U18768 (N_18768,N_18318,N_18298);
xor U18769 (N_18769,N_18350,N_18519);
nand U18770 (N_18770,N_18285,N_18690);
nor U18771 (N_18771,N_18620,N_18321);
xor U18772 (N_18772,N_18562,N_18507);
nor U18773 (N_18773,N_18431,N_18307);
and U18774 (N_18774,N_18376,N_18277);
xor U18775 (N_18775,N_18559,N_18425);
nor U18776 (N_18776,N_18159,N_18359);
or U18777 (N_18777,N_18379,N_18411);
nor U18778 (N_18778,N_18651,N_18636);
nor U18779 (N_18779,N_18432,N_18509);
nand U18780 (N_18780,N_18729,N_18282);
nand U18781 (N_18781,N_18203,N_18534);
nor U18782 (N_18782,N_18174,N_18545);
and U18783 (N_18783,N_18556,N_18443);
xor U18784 (N_18784,N_18485,N_18151);
xor U18785 (N_18785,N_18716,N_18275);
xor U18786 (N_18786,N_18353,N_18468);
nor U18787 (N_18787,N_18361,N_18453);
and U18788 (N_18788,N_18499,N_18211);
nor U18789 (N_18789,N_18252,N_18546);
nor U18790 (N_18790,N_18273,N_18595);
and U18791 (N_18791,N_18538,N_18558);
xor U18792 (N_18792,N_18675,N_18399);
xor U18793 (N_18793,N_18388,N_18560);
nor U18794 (N_18794,N_18234,N_18736);
xor U18795 (N_18795,N_18142,N_18419);
nor U18796 (N_18796,N_18511,N_18561);
xnor U18797 (N_18797,N_18661,N_18390);
nand U18798 (N_18798,N_18223,N_18673);
and U18799 (N_18799,N_18360,N_18548);
xor U18800 (N_18800,N_18549,N_18155);
and U18801 (N_18801,N_18704,N_18192);
and U18802 (N_18802,N_18482,N_18221);
xor U18803 (N_18803,N_18236,N_18702);
xnor U18804 (N_18804,N_18691,N_18245);
and U18805 (N_18805,N_18225,N_18185);
nand U18806 (N_18806,N_18590,N_18671);
xor U18807 (N_18807,N_18337,N_18429);
nor U18808 (N_18808,N_18341,N_18312);
nor U18809 (N_18809,N_18378,N_18190);
nand U18810 (N_18810,N_18125,N_18608);
nand U18811 (N_18811,N_18274,N_18730);
nand U18812 (N_18812,N_18264,N_18612);
xor U18813 (N_18813,N_18664,N_18160);
or U18814 (N_18814,N_18293,N_18450);
nand U18815 (N_18815,N_18156,N_18692);
and U18816 (N_18816,N_18317,N_18403);
nor U18817 (N_18817,N_18335,N_18618);
and U18818 (N_18818,N_18551,N_18638);
or U18819 (N_18819,N_18394,N_18235);
nor U18820 (N_18820,N_18314,N_18709);
xor U18821 (N_18821,N_18537,N_18448);
and U18822 (N_18822,N_18693,N_18153);
nor U18823 (N_18823,N_18139,N_18256);
nor U18824 (N_18824,N_18363,N_18462);
nor U18825 (N_18825,N_18512,N_18385);
or U18826 (N_18826,N_18148,N_18165);
or U18827 (N_18827,N_18689,N_18149);
or U18828 (N_18828,N_18247,N_18492);
and U18829 (N_18829,N_18616,N_18703);
xnor U18830 (N_18830,N_18714,N_18470);
nor U18831 (N_18831,N_18533,N_18624);
and U18832 (N_18832,N_18416,N_18246);
nand U18833 (N_18833,N_18348,N_18295);
and U18834 (N_18834,N_18393,N_18488);
and U18835 (N_18835,N_18180,N_18594);
xnor U18836 (N_18836,N_18739,N_18748);
and U18837 (N_18837,N_18224,N_18652);
nand U18838 (N_18838,N_18424,N_18451);
and U18839 (N_18839,N_18194,N_18564);
and U18840 (N_18840,N_18212,N_18710);
xnor U18841 (N_18841,N_18720,N_18309);
xnor U18842 (N_18842,N_18251,N_18198);
and U18843 (N_18843,N_18323,N_18480);
nand U18844 (N_18844,N_18574,N_18576);
nor U18845 (N_18845,N_18553,N_18366);
or U18846 (N_18846,N_18345,N_18286);
xor U18847 (N_18847,N_18179,N_18655);
or U18848 (N_18848,N_18728,N_18554);
nor U18849 (N_18849,N_18137,N_18172);
nand U18850 (N_18850,N_18573,N_18715);
xor U18851 (N_18851,N_18498,N_18644);
and U18852 (N_18852,N_18228,N_18296);
and U18853 (N_18853,N_18501,N_18186);
xor U18854 (N_18854,N_18128,N_18303);
or U18855 (N_18855,N_18222,N_18628);
nor U18856 (N_18856,N_18745,N_18591);
nor U18857 (N_18857,N_18449,N_18542);
xnor U18858 (N_18858,N_18288,N_18197);
and U18859 (N_18859,N_18268,N_18412);
or U18860 (N_18860,N_18371,N_18183);
xnor U18861 (N_18861,N_18281,N_18271);
nand U18862 (N_18862,N_18402,N_18505);
nor U18863 (N_18863,N_18469,N_18544);
or U18864 (N_18864,N_18486,N_18218);
and U18865 (N_18865,N_18134,N_18520);
xor U18866 (N_18866,N_18580,N_18334);
and U18867 (N_18867,N_18530,N_18528);
nand U18868 (N_18868,N_18632,N_18706);
nor U18869 (N_18869,N_18602,N_18435);
nor U18870 (N_18870,N_18414,N_18428);
nor U18871 (N_18871,N_18267,N_18744);
nand U18872 (N_18872,N_18467,N_18539);
xnor U18873 (N_18873,N_18438,N_18255);
nor U18874 (N_18874,N_18143,N_18369);
xnor U18875 (N_18875,N_18582,N_18726);
or U18876 (N_18876,N_18625,N_18357);
nor U18877 (N_18877,N_18515,N_18188);
nand U18878 (N_18878,N_18202,N_18208);
nor U18879 (N_18879,N_18521,N_18619);
and U18880 (N_18880,N_18565,N_18698);
xnor U18881 (N_18881,N_18621,N_18687);
xor U18882 (N_18882,N_18171,N_18526);
and U18883 (N_18883,N_18215,N_18130);
and U18884 (N_18884,N_18217,N_18260);
or U18885 (N_18885,N_18238,N_18654);
and U18886 (N_18886,N_18466,N_18207);
or U18887 (N_18887,N_18204,N_18173);
or U18888 (N_18888,N_18490,N_18206);
and U18889 (N_18889,N_18504,N_18170);
and U18890 (N_18890,N_18658,N_18647);
nand U18891 (N_18891,N_18524,N_18472);
or U18892 (N_18892,N_18452,N_18413);
nor U18893 (N_18893,N_18331,N_18679);
xnor U18894 (N_18894,N_18610,N_18510);
or U18895 (N_18895,N_18579,N_18734);
and U18896 (N_18896,N_18484,N_18588);
nor U18897 (N_18897,N_18604,N_18343);
or U18898 (N_18898,N_18494,N_18316);
xnor U18899 (N_18899,N_18550,N_18543);
nor U18900 (N_18900,N_18313,N_18301);
and U18901 (N_18901,N_18291,N_18351);
xnor U18902 (N_18902,N_18708,N_18199);
xnor U18903 (N_18903,N_18522,N_18427);
and U18904 (N_18904,N_18639,N_18700);
and U18905 (N_18905,N_18210,N_18458);
xnor U18906 (N_18906,N_18441,N_18253);
and U18907 (N_18907,N_18731,N_18471);
and U18908 (N_18908,N_18146,N_18436);
nor U18909 (N_18909,N_18555,N_18575);
nand U18910 (N_18910,N_18384,N_18685);
and U18911 (N_18911,N_18220,N_18479);
nor U18912 (N_18912,N_18358,N_18297);
xnor U18913 (N_18913,N_18699,N_18493);
and U18914 (N_18914,N_18166,N_18677);
nand U18915 (N_18915,N_18231,N_18536);
and U18916 (N_18916,N_18392,N_18289);
nand U18917 (N_18917,N_18606,N_18355);
xor U18918 (N_18918,N_18569,N_18649);
or U18919 (N_18919,N_18311,N_18696);
nand U18920 (N_18920,N_18326,N_18667);
nand U18921 (N_18921,N_18571,N_18417);
nor U18922 (N_18922,N_18167,N_18670);
nand U18923 (N_18923,N_18514,N_18630);
nand U18924 (N_18924,N_18241,N_18684);
nor U18925 (N_18925,N_18315,N_18324);
nor U18926 (N_18926,N_18680,N_18426);
and U18927 (N_18927,N_18237,N_18532);
nand U18928 (N_18928,N_18398,N_18410);
xnor U18929 (N_18929,N_18263,N_18158);
and U18930 (N_18930,N_18535,N_18287);
and U18931 (N_18931,N_18660,N_18592);
xor U18932 (N_18932,N_18147,N_18136);
nor U18933 (N_18933,N_18746,N_18395);
and U18934 (N_18934,N_18456,N_18645);
xor U18935 (N_18935,N_18336,N_18219);
or U18936 (N_18936,N_18129,N_18354);
and U18937 (N_18937,N_18659,N_18668);
nand U18938 (N_18938,N_18141,N_18567);
or U18939 (N_18939,N_18455,N_18257);
xnor U18940 (N_18940,N_18266,N_18681);
nor U18941 (N_18941,N_18254,N_18641);
nand U18942 (N_18942,N_18711,N_18319);
xnor U18943 (N_18943,N_18572,N_18408);
nand U18944 (N_18944,N_18674,N_18598);
or U18945 (N_18945,N_18695,N_18196);
xnor U18946 (N_18946,N_18205,N_18135);
nor U18947 (N_18947,N_18742,N_18459);
or U18948 (N_18948,N_18332,N_18292);
or U18949 (N_18949,N_18581,N_18214);
nand U18950 (N_18950,N_18523,N_18557);
or U18951 (N_18951,N_18547,N_18421);
xnor U18952 (N_18952,N_18676,N_18629);
and U18953 (N_18953,N_18304,N_18725);
nand U18954 (N_18954,N_18525,N_18503);
and U18955 (N_18955,N_18387,N_18662);
and U18956 (N_18956,N_18631,N_18440);
and U18957 (N_18957,N_18747,N_18226);
or U18958 (N_18958,N_18259,N_18191);
or U18959 (N_18959,N_18603,N_18433);
or U18960 (N_18960,N_18338,N_18447);
nor U18961 (N_18961,N_18294,N_18473);
or U18962 (N_18962,N_18409,N_18340);
nor U18963 (N_18963,N_18540,N_18373);
nor U18964 (N_18964,N_18465,N_18474);
nor U18965 (N_18965,N_18701,N_18401);
nand U18966 (N_18966,N_18423,N_18502);
nand U18967 (N_18967,N_18280,N_18389);
or U18968 (N_18968,N_18707,N_18383);
xor U18969 (N_18969,N_18157,N_18614);
and U18970 (N_18970,N_18733,N_18650);
nor U18971 (N_18971,N_18420,N_18721);
nand U18972 (N_18972,N_18497,N_18600);
and U18973 (N_18973,N_18593,N_18643);
xor U18974 (N_18974,N_18232,N_18305);
xor U18975 (N_18975,N_18364,N_18666);
and U18976 (N_18976,N_18195,N_18622);
nand U18977 (N_18977,N_18741,N_18601);
or U18978 (N_18978,N_18239,N_18265);
and U18979 (N_18979,N_18300,N_18518);
or U18980 (N_18980,N_18405,N_18362);
nor U18981 (N_18981,N_18635,N_18227);
nand U18982 (N_18982,N_18717,N_18483);
nor U18983 (N_18983,N_18476,N_18249);
nor U18984 (N_18984,N_18640,N_18500);
nor U18985 (N_18985,N_18463,N_18611);
xnor U18986 (N_18986,N_18365,N_18377);
nor U18987 (N_18987,N_18517,N_18299);
and U18988 (N_18988,N_18250,N_18140);
or U18989 (N_18989,N_18656,N_18585);
or U18990 (N_18990,N_18302,N_18184);
and U18991 (N_18991,N_18460,N_18162);
xnor U18992 (N_18992,N_18552,N_18131);
and U18993 (N_18993,N_18310,N_18516);
and U18994 (N_18994,N_18400,N_18722);
and U18995 (N_18995,N_18617,N_18627);
and U18996 (N_18996,N_18596,N_18607);
xor U18997 (N_18997,N_18737,N_18344);
nor U18998 (N_18998,N_18657,N_18589);
nor U18999 (N_18999,N_18374,N_18481);
nor U19000 (N_19000,N_18577,N_18279);
xor U19001 (N_19001,N_18609,N_18445);
xnor U19002 (N_19002,N_18270,N_18461);
nor U19003 (N_19003,N_18372,N_18176);
nand U19004 (N_19004,N_18697,N_18144);
nand U19005 (N_19005,N_18407,N_18527);
nand U19006 (N_19006,N_18244,N_18669);
nor U19007 (N_19007,N_18391,N_18339);
or U19008 (N_19008,N_18381,N_18349);
and U19009 (N_19009,N_18563,N_18724);
or U19010 (N_19010,N_18175,N_18663);
and U19011 (N_19011,N_18370,N_18346);
nor U19012 (N_19012,N_18686,N_18615);
xor U19013 (N_19013,N_18477,N_18487);
xor U19014 (N_19014,N_18328,N_18727);
and U19015 (N_19015,N_18329,N_18127);
or U19016 (N_19016,N_18489,N_18230);
and U19017 (N_19017,N_18283,N_18168);
nor U19018 (N_19018,N_18672,N_18269);
nor U19019 (N_19019,N_18648,N_18613);
xnor U19020 (N_19020,N_18382,N_18599);
or U19021 (N_19021,N_18347,N_18578);
xor U19022 (N_19022,N_18368,N_18444);
nor U19023 (N_19023,N_18126,N_18566);
and U19024 (N_19024,N_18178,N_18718);
and U19025 (N_19025,N_18333,N_18597);
xnor U19026 (N_19026,N_18261,N_18434);
nor U19027 (N_19027,N_18352,N_18570);
and U19028 (N_19028,N_18705,N_18508);
and U19029 (N_19029,N_18262,N_18464);
or U19030 (N_19030,N_18240,N_18322);
and U19031 (N_19031,N_18568,N_18145);
nand U19032 (N_19032,N_18177,N_18367);
nand U19033 (N_19033,N_18738,N_18164);
nor U19034 (N_19034,N_18422,N_18229);
nor U19035 (N_19035,N_18320,N_18284);
and U19036 (N_19036,N_18150,N_18529);
and U19037 (N_19037,N_18633,N_18375);
or U19038 (N_19038,N_18732,N_18276);
nor U19039 (N_19039,N_18531,N_18584);
nor U19040 (N_19040,N_18213,N_18454);
xnor U19041 (N_19041,N_18161,N_18637);
xnor U19042 (N_19042,N_18396,N_18646);
xor U19043 (N_19043,N_18290,N_18415);
or U19044 (N_19044,N_18278,N_18719);
xor U19045 (N_19045,N_18187,N_18189);
and U19046 (N_19046,N_18495,N_18216);
or U19047 (N_19047,N_18653,N_18605);
and U19048 (N_19048,N_18688,N_18506);
nand U19049 (N_19049,N_18713,N_18330);
and U19050 (N_19050,N_18694,N_18152);
and U19051 (N_19051,N_18437,N_18242);
or U19052 (N_19052,N_18380,N_18586);
or U19053 (N_19053,N_18626,N_18712);
nor U19054 (N_19054,N_18243,N_18513);
nand U19055 (N_19055,N_18201,N_18439);
and U19056 (N_19056,N_18386,N_18163);
xor U19057 (N_19057,N_18457,N_18154);
nand U19058 (N_19058,N_18743,N_18735);
and U19059 (N_19059,N_18248,N_18233);
xor U19060 (N_19060,N_18209,N_18356);
nand U19061 (N_19061,N_18430,N_18406);
nor U19062 (N_19062,N_18541,N_18324);
or U19063 (N_19063,N_18553,N_18535);
nor U19064 (N_19064,N_18483,N_18668);
and U19065 (N_19065,N_18272,N_18459);
nor U19066 (N_19066,N_18265,N_18295);
nand U19067 (N_19067,N_18503,N_18147);
nand U19068 (N_19068,N_18668,N_18684);
nor U19069 (N_19069,N_18263,N_18310);
nor U19070 (N_19070,N_18695,N_18401);
xnor U19071 (N_19071,N_18218,N_18541);
xnor U19072 (N_19072,N_18235,N_18259);
or U19073 (N_19073,N_18746,N_18169);
xnor U19074 (N_19074,N_18345,N_18299);
and U19075 (N_19075,N_18747,N_18353);
and U19076 (N_19076,N_18517,N_18494);
or U19077 (N_19077,N_18633,N_18267);
and U19078 (N_19078,N_18134,N_18517);
nor U19079 (N_19079,N_18538,N_18712);
nand U19080 (N_19080,N_18202,N_18157);
nand U19081 (N_19081,N_18137,N_18136);
or U19082 (N_19082,N_18206,N_18685);
nor U19083 (N_19083,N_18265,N_18677);
xnor U19084 (N_19084,N_18666,N_18729);
and U19085 (N_19085,N_18141,N_18306);
xor U19086 (N_19086,N_18527,N_18584);
and U19087 (N_19087,N_18383,N_18548);
or U19088 (N_19088,N_18410,N_18445);
xor U19089 (N_19089,N_18156,N_18428);
nand U19090 (N_19090,N_18231,N_18593);
nand U19091 (N_19091,N_18724,N_18364);
xor U19092 (N_19092,N_18569,N_18140);
xor U19093 (N_19093,N_18430,N_18696);
or U19094 (N_19094,N_18458,N_18231);
and U19095 (N_19095,N_18483,N_18350);
nor U19096 (N_19096,N_18351,N_18161);
nor U19097 (N_19097,N_18702,N_18516);
nor U19098 (N_19098,N_18543,N_18707);
or U19099 (N_19099,N_18471,N_18273);
xor U19100 (N_19100,N_18591,N_18492);
nor U19101 (N_19101,N_18420,N_18444);
nor U19102 (N_19102,N_18457,N_18536);
xnor U19103 (N_19103,N_18363,N_18205);
or U19104 (N_19104,N_18611,N_18541);
or U19105 (N_19105,N_18437,N_18175);
or U19106 (N_19106,N_18229,N_18402);
or U19107 (N_19107,N_18500,N_18509);
or U19108 (N_19108,N_18260,N_18334);
nand U19109 (N_19109,N_18745,N_18611);
nor U19110 (N_19110,N_18742,N_18253);
and U19111 (N_19111,N_18247,N_18267);
and U19112 (N_19112,N_18549,N_18389);
nor U19113 (N_19113,N_18436,N_18516);
or U19114 (N_19114,N_18718,N_18692);
or U19115 (N_19115,N_18221,N_18465);
nor U19116 (N_19116,N_18712,N_18671);
xor U19117 (N_19117,N_18254,N_18709);
nand U19118 (N_19118,N_18371,N_18226);
xnor U19119 (N_19119,N_18244,N_18136);
nor U19120 (N_19120,N_18436,N_18402);
xor U19121 (N_19121,N_18187,N_18539);
and U19122 (N_19122,N_18724,N_18623);
and U19123 (N_19123,N_18449,N_18628);
nor U19124 (N_19124,N_18295,N_18649);
or U19125 (N_19125,N_18520,N_18132);
nand U19126 (N_19126,N_18594,N_18668);
xor U19127 (N_19127,N_18663,N_18467);
nand U19128 (N_19128,N_18517,N_18430);
or U19129 (N_19129,N_18411,N_18160);
nand U19130 (N_19130,N_18355,N_18469);
and U19131 (N_19131,N_18623,N_18632);
xor U19132 (N_19132,N_18716,N_18351);
and U19133 (N_19133,N_18471,N_18304);
nand U19134 (N_19134,N_18695,N_18578);
nor U19135 (N_19135,N_18710,N_18563);
xnor U19136 (N_19136,N_18509,N_18381);
and U19137 (N_19137,N_18606,N_18167);
and U19138 (N_19138,N_18632,N_18479);
and U19139 (N_19139,N_18706,N_18483);
nand U19140 (N_19140,N_18625,N_18450);
xor U19141 (N_19141,N_18638,N_18148);
nand U19142 (N_19142,N_18425,N_18381);
nor U19143 (N_19143,N_18250,N_18620);
and U19144 (N_19144,N_18564,N_18317);
xor U19145 (N_19145,N_18648,N_18632);
or U19146 (N_19146,N_18187,N_18304);
nor U19147 (N_19147,N_18179,N_18507);
and U19148 (N_19148,N_18344,N_18349);
nor U19149 (N_19149,N_18182,N_18239);
nor U19150 (N_19150,N_18732,N_18475);
nor U19151 (N_19151,N_18240,N_18349);
and U19152 (N_19152,N_18288,N_18564);
and U19153 (N_19153,N_18391,N_18666);
or U19154 (N_19154,N_18495,N_18162);
and U19155 (N_19155,N_18745,N_18270);
and U19156 (N_19156,N_18549,N_18378);
and U19157 (N_19157,N_18201,N_18254);
or U19158 (N_19158,N_18675,N_18182);
nor U19159 (N_19159,N_18467,N_18294);
nand U19160 (N_19160,N_18736,N_18496);
and U19161 (N_19161,N_18281,N_18357);
or U19162 (N_19162,N_18606,N_18548);
nor U19163 (N_19163,N_18677,N_18457);
nor U19164 (N_19164,N_18534,N_18652);
and U19165 (N_19165,N_18676,N_18306);
xnor U19166 (N_19166,N_18204,N_18619);
and U19167 (N_19167,N_18699,N_18308);
and U19168 (N_19168,N_18631,N_18606);
and U19169 (N_19169,N_18461,N_18658);
nor U19170 (N_19170,N_18468,N_18233);
or U19171 (N_19171,N_18457,N_18688);
xor U19172 (N_19172,N_18713,N_18126);
nor U19173 (N_19173,N_18442,N_18738);
xor U19174 (N_19174,N_18199,N_18139);
nand U19175 (N_19175,N_18568,N_18181);
nand U19176 (N_19176,N_18720,N_18373);
nand U19177 (N_19177,N_18549,N_18382);
and U19178 (N_19178,N_18329,N_18241);
and U19179 (N_19179,N_18409,N_18566);
xnor U19180 (N_19180,N_18550,N_18567);
and U19181 (N_19181,N_18208,N_18292);
and U19182 (N_19182,N_18175,N_18479);
and U19183 (N_19183,N_18635,N_18614);
nand U19184 (N_19184,N_18578,N_18234);
nand U19185 (N_19185,N_18379,N_18512);
or U19186 (N_19186,N_18180,N_18644);
nand U19187 (N_19187,N_18253,N_18537);
or U19188 (N_19188,N_18634,N_18479);
xnor U19189 (N_19189,N_18216,N_18302);
and U19190 (N_19190,N_18543,N_18150);
nand U19191 (N_19191,N_18576,N_18699);
or U19192 (N_19192,N_18562,N_18706);
and U19193 (N_19193,N_18300,N_18648);
nand U19194 (N_19194,N_18138,N_18292);
nand U19195 (N_19195,N_18673,N_18547);
or U19196 (N_19196,N_18630,N_18471);
or U19197 (N_19197,N_18409,N_18323);
xor U19198 (N_19198,N_18509,N_18598);
or U19199 (N_19199,N_18378,N_18192);
xnor U19200 (N_19200,N_18234,N_18489);
and U19201 (N_19201,N_18548,N_18596);
xor U19202 (N_19202,N_18717,N_18677);
nand U19203 (N_19203,N_18320,N_18183);
nand U19204 (N_19204,N_18549,N_18359);
and U19205 (N_19205,N_18160,N_18713);
nand U19206 (N_19206,N_18457,N_18666);
nor U19207 (N_19207,N_18344,N_18511);
nand U19208 (N_19208,N_18180,N_18185);
or U19209 (N_19209,N_18227,N_18188);
or U19210 (N_19210,N_18509,N_18643);
nand U19211 (N_19211,N_18313,N_18704);
nand U19212 (N_19212,N_18533,N_18409);
xor U19213 (N_19213,N_18128,N_18497);
or U19214 (N_19214,N_18226,N_18234);
nand U19215 (N_19215,N_18743,N_18606);
nor U19216 (N_19216,N_18677,N_18167);
nor U19217 (N_19217,N_18163,N_18645);
xnor U19218 (N_19218,N_18556,N_18202);
and U19219 (N_19219,N_18612,N_18296);
and U19220 (N_19220,N_18642,N_18215);
and U19221 (N_19221,N_18529,N_18436);
nor U19222 (N_19222,N_18553,N_18303);
xor U19223 (N_19223,N_18281,N_18594);
xor U19224 (N_19224,N_18209,N_18396);
nor U19225 (N_19225,N_18469,N_18240);
nor U19226 (N_19226,N_18366,N_18322);
nand U19227 (N_19227,N_18324,N_18390);
or U19228 (N_19228,N_18359,N_18565);
and U19229 (N_19229,N_18749,N_18201);
nand U19230 (N_19230,N_18345,N_18194);
and U19231 (N_19231,N_18608,N_18507);
nand U19232 (N_19232,N_18320,N_18158);
xnor U19233 (N_19233,N_18418,N_18623);
nor U19234 (N_19234,N_18744,N_18483);
nand U19235 (N_19235,N_18177,N_18372);
and U19236 (N_19236,N_18133,N_18329);
or U19237 (N_19237,N_18606,N_18411);
or U19238 (N_19238,N_18401,N_18524);
and U19239 (N_19239,N_18181,N_18504);
nor U19240 (N_19240,N_18493,N_18694);
nor U19241 (N_19241,N_18513,N_18125);
nand U19242 (N_19242,N_18681,N_18487);
nor U19243 (N_19243,N_18210,N_18133);
nor U19244 (N_19244,N_18133,N_18160);
and U19245 (N_19245,N_18265,N_18127);
nor U19246 (N_19246,N_18243,N_18517);
nor U19247 (N_19247,N_18147,N_18708);
nand U19248 (N_19248,N_18432,N_18636);
or U19249 (N_19249,N_18144,N_18309);
xnor U19250 (N_19250,N_18255,N_18565);
and U19251 (N_19251,N_18227,N_18379);
nor U19252 (N_19252,N_18303,N_18487);
nor U19253 (N_19253,N_18406,N_18384);
nand U19254 (N_19254,N_18147,N_18434);
nand U19255 (N_19255,N_18668,N_18359);
xnor U19256 (N_19256,N_18610,N_18658);
and U19257 (N_19257,N_18574,N_18407);
nand U19258 (N_19258,N_18579,N_18570);
nor U19259 (N_19259,N_18467,N_18277);
nand U19260 (N_19260,N_18634,N_18619);
or U19261 (N_19261,N_18137,N_18287);
or U19262 (N_19262,N_18434,N_18230);
nor U19263 (N_19263,N_18479,N_18648);
nand U19264 (N_19264,N_18675,N_18673);
and U19265 (N_19265,N_18708,N_18524);
nor U19266 (N_19266,N_18434,N_18429);
nand U19267 (N_19267,N_18452,N_18299);
nor U19268 (N_19268,N_18243,N_18349);
and U19269 (N_19269,N_18322,N_18309);
or U19270 (N_19270,N_18594,N_18397);
xor U19271 (N_19271,N_18220,N_18267);
nand U19272 (N_19272,N_18262,N_18238);
nor U19273 (N_19273,N_18481,N_18696);
or U19274 (N_19274,N_18314,N_18214);
nand U19275 (N_19275,N_18399,N_18517);
and U19276 (N_19276,N_18627,N_18468);
xor U19277 (N_19277,N_18674,N_18665);
and U19278 (N_19278,N_18164,N_18319);
or U19279 (N_19279,N_18296,N_18389);
xnor U19280 (N_19280,N_18466,N_18403);
or U19281 (N_19281,N_18412,N_18463);
or U19282 (N_19282,N_18214,N_18674);
and U19283 (N_19283,N_18248,N_18266);
and U19284 (N_19284,N_18173,N_18369);
xor U19285 (N_19285,N_18371,N_18665);
or U19286 (N_19286,N_18734,N_18200);
xor U19287 (N_19287,N_18210,N_18555);
and U19288 (N_19288,N_18614,N_18127);
xnor U19289 (N_19289,N_18140,N_18402);
or U19290 (N_19290,N_18174,N_18240);
nand U19291 (N_19291,N_18686,N_18296);
nand U19292 (N_19292,N_18433,N_18618);
and U19293 (N_19293,N_18278,N_18675);
and U19294 (N_19294,N_18558,N_18217);
xor U19295 (N_19295,N_18515,N_18575);
xor U19296 (N_19296,N_18354,N_18131);
nand U19297 (N_19297,N_18132,N_18398);
and U19298 (N_19298,N_18157,N_18225);
nand U19299 (N_19299,N_18448,N_18133);
and U19300 (N_19300,N_18744,N_18749);
and U19301 (N_19301,N_18649,N_18724);
nor U19302 (N_19302,N_18209,N_18507);
or U19303 (N_19303,N_18351,N_18247);
xnor U19304 (N_19304,N_18462,N_18528);
nand U19305 (N_19305,N_18556,N_18389);
or U19306 (N_19306,N_18200,N_18347);
nand U19307 (N_19307,N_18202,N_18590);
xor U19308 (N_19308,N_18528,N_18352);
or U19309 (N_19309,N_18301,N_18147);
or U19310 (N_19310,N_18656,N_18216);
and U19311 (N_19311,N_18402,N_18656);
and U19312 (N_19312,N_18584,N_18126);
or U19313 (N_19313,N_18386,N_18713);
nand U19314 (N_19314,N_18700,N_18283);
and U19315 (N_19315,N_18301,N_18519);
nor U19316 (N_19316,N_18459,N_18166);
nand U19317 (N_19317,N_18216,N_18344);
nor U19318 (N_19318,N_18537,N_18533);
or U19319 (N_19319,N_18707,N_18282);
and U19320 (N_19320,N_18201,N_18491);
nand U19321 (N_19321,N_18394,N_18631);
and U19322 (N_19322,N_18413,N_18407);
xor U19323 (N_19323,N_18723,N_18493);
or U19324 (N_19324,N_18684,N_18373);
nor U19325 (N_19325,N_18326,N_18356);
xor U19326 (N_19326,N_18388,N_18163);
xnor U19327 (N_19327,N_18748,N_18645);
xor U19328 (N_19328,N_18451,N_18674);
or U19329 (N_19329,N_18223,N_18482);
and U19330 (N_19330,N_18432,N_18554);
or U19331 (N_19331,N_18214,N_18321);
nand U19332 (N_19332,N_18334,N_18251);
xnor U19333 (N_19333,N_18301,N_18419);
nand U19334 (N_19334,N_18450,N_18456);
nand U19335 (N_19335,N_18253,N_18440);
or U19336 (N_19336,N_18500,N_18260);
or U19337 (N_19337,N_18334,N_18234);
nor U19338 (N_19338,N_18673,N_18213);
nand U19339 (N_19339,N_18642,N_18486);
nand U19340 (N_19340,N_18350,N_18412);
xnor U19341 (N_19341,N_18744,N_18256);
or U19342 (N_19342,N_18635,N_18553);
and U19343 (N_19343,N_18678,N_18506);
nand U19344 (N_19344,N_18649,N_18217);
xor U19345 (N_19345,N_18288,N_18504);
nor U19346 (N_19346,N_18192,N_18595);
xnor U19347 (N_19347,N_18612,N_18235);
nand U19348 (N_19348,N_18201,N_18324);
nor U19349 (N_19349,N_18640,N_18460);
and U19350 (N_19350,N_18718,N_18294);
nand U19351 (N_19351,N_18177,N_18396);
xor U19352 (N_19352,N_18142,N_18211);
nand U19353 (N_19353,N_18500,N_18730);
or U19354 (N_19354,N_18332,N_18458);
or U19355 (N_19355,N_18481,N_18422);
or U19356 (N_19356,N_18285,N_18680);
or U19357 (N_19357,N_18699,N_18377);
nand U19358 (N_19358,N_18444,N_18713);
xor U19359 (N_19359,N_18127,N_18258);
nor U19360 (N_19360,N_18562,N_18214);
nor U19361 (N_19361,N_18602,N_18198);
or U19362 (N_19362,N_18485,N_18420);
or U19363 (N_19363,N_18549,N_18138);
nand U19364 (N_19364,N_18143,N_18128);
nand U19365 (N_19365,N_18383,N_18352);
nand U19366 (N_19366,N_18228,N_18182);
and U19367 (N_19367,N_18521,N_18668);
nor U19368 (N_19368,N_18237,N_18535);
nand U19369 (N_19369,N_18617,N_18340);
or U19370 (N_19370,N_18148,N_18295);
nand U19371 (N_19371,N_18482,N_18383);
and U19372 (N_19372,N_18423,N_18206);
or U19373 (N_19373,N_18563,N_18211);
nand U19374 (N_19374,N_18414,N_18300);
and U19375 (N_19375,N_18788,N_19222);
nand U19376 (N_19376,N_19063,N_19165);
nand U19377 (N_19377,N_19031,N_19114);
nor U19378 (N_19378,N_18867,N_19081);
nand U19379 (N_19379,N_18989,N_18937);
nand U19380 (N_19380,N_19070,N_18962);
and U19381 (N_19381,N_19197,N_18791);
xor U19382 (N_19382,N_19060,N_19011);
xor U19383 (N_19383,N_18979,N_19178);
or U19384 (N_19384,N_18930,N_19168);
or U19385 (N_19385,N_18983,N_19030);
or U19386 (N_19386,N_18778,N_18811);
nor U19387 (N_19387,N_19048,N_18925);
nand U19388 (N_19388,N_18908,N_18942);
xnor U19389 (N_19389,N_18934,N_18870);
xor U19390 (N_19390,N_19200,N_19280);
xnor U19391 (N_19391,N_18768,N_19170);
nor U19392 (N_19392,N_18765,N_18862);
xor U19393 (N_19393,N_18893,N_18885);
nor U19394 (N_19394,N_19020,N_19198);
xnor U19395 (N_19395,N_19265,N_19318);
or U19396 (N_19396,N_18807,N_19314);
or U19397 (N_19397,N_19151,N_18803);
and U19398 (N_19398,N_19327,N_18894);
and U19399 (N_19399,N_19321,N_19342);
nand U19400 (N_19400,N_18907,N_18875);
nand U19401 (N_19401,N_18993,N_19305);
nor U19402 (N_19402,N_19279,N_18816);
nand U19403 (N_19403,N_19336,N_19079);
nor U19404 (N_19404,N_19303,N_19106);
nor U19405 (N_19405,N_19053,N_18964);
nand U19406 (N_19406,N_19292,N_19082);
nor U19407 (N_19407,N_18767,N_19115);
nand U19408 (N_19408,N_19025,N_19135);
nor U19409 (N_19409,N_18770,N_19185);
xor U19410 (N_19410,N_19267,N_18773);
nand U19411 (N_19411,N_19354,N_18923);
or U19412 (N_19412,N_18986,N_19364);
nor U19413 (N_19413,N_19270,N_18882);
or U19414 (N_19414,N_19100,N_19138);
nor U19415 (N_19415,N_19144,N_19158);
and U19416 (N_19416,N_18782,N_19365);
or U19417 (N_19417,N_19174,N_19210);
nor U19418 (N_19418,N_18779,N_18864);
nand U19419 (N_19419,N_19110,N_19142);
xor U19420 (N_19420,N_19171,N_18752);
nor U19421 (N_19421,N_18881,N_18769);
xor U19422 (N_19422,N_19050,N_18860);
nand U19423 (N_19423,N_18785,N_19074);
or U19424 (N_19424,N_18975,N_19231);
xnor U19425 (N_19425,N_18815,N_19049);
nor U19426 (N_19426,N_19213,N_18884);
or U19427 (N_19427,N_19004,N_19224);
or U19428 (N_19428,N_19358,N_19322);
or U19429 (N_19429,N_19104,N_19090);
xor U19430 (N_19430,N_18776,N_19067);
and U19431 (N_19431,N_18903,N_19304);
nor U19432 (N_19432,N_18780,N_19337);
and U19433 (N_19433,N_18910,N_18957);
xnor U19434 (N_19434,N_19083,N_19014);
xnor U19435 (N_19435,N_19355,N_18754);
xnor U19436 (N_19436,N_18758,N_19299);
nand U19437 (N_19437,N_19340,N_19162);
nand U19438 (N_19438,N_19109,N_19236);
xnor U19439 (N_19439,N_19061,N_18997);
nor U19440 (N_19440,N_19320,N_18980);
nor U19441 (N_19441,N_19002,N_18996);
nor U19442 (N_19442,N_19080,N_19042);
or U19443 (N_19443,N_18947,N_19140);
nand U19444 (N_19444,N_19127,N_18771);
nand U19445 (N_19445,N_19278,N_18931);
xnor U19446 (N_19446,N_19290,N_19017);
nor U19447 (N_19447,N_18866,N_18981);
and U19448 (N_19448,N_19244,N_19214);
nor U19449 (N_19449,N_19264,N_19359);
or U19450 (N_19450,N_18914,N_19262);
nor U19451 (N_19451,N_18918,N_19289);
or U19452 (N_19452,N_18959,N_19208);
nand U19453 (N_19453,N_19247,N_19124);
nand U19454 (N_19454,N_18974,N_19297);
xnor U19455 (N_19455,N_19033,N_19350);
and U19456 (N_19456,N_18880,N_18821);
or U19457 (N_19457,N_19096,N_18802);
and U19458 (N_19458,N_18793,N_19223);
nand U19459 (N_19459,N_19179,N_19040);
or U19460 (N_19460,N_18965,N_19065);
and U19461 (N_19461,N_18854,N_18865);
nand U19462 (N_19462,N_19075,N_18820);
and U19463 (N_19463,N_19362,N_18840);
nor U19464 (N_19464,N_19284,N_19054);
nor U19465 (N_19465,N_18805,N_19023);
nand U19466 (N_19466,N_19332,N_18834);
or U19467 (N_19467,N_19041,N_18789);
and U19468 (N_19468,N_19245,N_18833);
or U19469 (N_19469,N_19206,N_19293);
and U19470 (N_19470,N_19175,N_18909);
nand U19471 (N_19471,N_18762,N_19274);
xor U19472 (N_19472,N_18929,N_18944);
nor U19473 (N_19473,N_19351,N_19077);
xnor U19474 (N_19474,N_18863,N_18960);
xnor U19475 (N_19475,N_19008,N_19013);
nor U19476 (N_19476,N_19037,N_18756);
nor U19477 (N_19477,N_18890,N_18935);
and U19478 (N_19478,N_19333,N_19016);
and U19479 (N_19479,N_19182,N_19241);
or U19480 (N_19480,N_19216,N_18963);
or U19481 (N_19481,N_19329,N_19131);
and U19482 (N_19482,N_19349,N_19370);
nor U19483 (N_19483,N_19312,N_18850);
nand U19484 (N_19484,N_18796,N_18859);
xor U19485 (N_19485,N_19301,N_18915);
and U19486 (N_19486,N_19219,N_19258);
nand U19487 (N_19487,N_19188,N_19027);
and U19488 (N_19488,N_19192,N_19311);
xor U19489 (N_19489,N_18783,N_18861);
nor U19490 (N_19490,N_19325,N_19288);
nand U19491 (N_19491,N_19072,N_19323);
nor U19492 (N_19492,N_18972,N_18943);
nor U19493 (N_19493,N_18795,N_19345);
nor U19494 (N_19494,N_19007,N_19024);
and U19495 (N_19495,N_19112,N_19137);
nor U19496 (N_19496,N_19058,N_19328);
nand U19497 (N_19497,N_18982,N_19134);
nor U19498 (N_19498,N_18899,N_18829);
and U19499 (N_19499,N_19240,N_19266);
nand U19500 (N_19500,N_18940,N_18971);
or U19501 (N_19501,N_18938,N_18878);
nor U19502 (N_19502,N_18764,N_19164);
xnor U19503 (N_19503,N_18818,N_18766);
xor U19504 (N_19504,N_18990,N_18921);
xnor U19505 (N_19505,N_18868,N_18933);
or U19506 (N_19506,N_18988,N_19071);
xnor U19507 (N_19507,N_19028,N_18994);
nand U19508 (N_19508,N_19268,N_19120);
and U19509 (N_19509,N_18750,N_19069);
or U19510 (N_19510,N_18876,N_19009);
and U19511 (N_19511,N_19018,N_19116);
nor U19512 (N_19512,N_18948,N_18753);
xor U19513 (N_19513,N_18917,N_19205);
or U19514 (N_19514,N_19043,N_18777);
or U19515 (N_19515,N_19105,N_19287);
nor U19516 (N_19516,N_18872,N_19209);
or U19517 (N_19517,N_19035,N_19285);
nor U19518 (N_19518,N_18912,N_18845);
xnor U19519 (N_19519,N_19253,N_19225);
xor U19520 (N_19520,N_18759,N_18800);
or U19521 (N_19521,N_18836,N_19338);
nor U19522 (N_19522,N_18945,N_19226);
and U19523 (N_19523,N_19026,N_19038);
and U19524 (N_19524,N_18784,N_19233);
xor U19525 (N_19525,N_18904,N_19057);
nor U19526 (N_19526,N_19126,N_18801);
or U19527 (N_19527,N_19235,N_19125);
nor U19528 (N_19528,N_19294,N_18920);
xnor U19529 (N_19529,N_18823,N_18887);
or U19530 (N_19530,N_19036,N_19194);
and U19531 (N_19531,N_19005,N_19203);
nor U19532 (N_19532,N_19146,N_18855);
xor U19533 (N_19533,N_19101,N_18774);
nand U19534 (N_19534,N_19257,N_19298);
xor U19535 (N_19535,N_19207,N_19121);
nor U19536 (N_19536,N_18911,N_18900);
xnor U19537 (N_19537,N_19357,N_18831);
or U19538 (N_19538,N_19148,N_18772);
nand U19539 (N_19539,N_18763,N_19360);
and U19540 (N_19540,N_19186,N_19335);
nand U19541 (N_19541,N_19220,N_19029);
or U19542 (N_19542,N_19324,N_18794);
and U19543 (N_19543,N_19097,N_19059);
nor U19544 (N_19544,N_19184,N_19353);
or U19545 (N_19545,N_18961,N_19147);
xor U19546 (N_19546,N_18761,N_19202);
xnor U19547 (N_19547,N_19319,N_18891);
xor U19548 (N_19548,N_18852,N_19150);
nand U19549 (N_19549,N_18838,N_19128);
and U19550 (N_19550,N_18985,N_18842);
nor U19551 (N_19551,N_19176,N_18927);
and U19552 (N_19552,N_19143,N_18792);
and U19553 (N_19553,N_18926,N_19102);
nand U19554 (N_19554,N_19313,N_19371);
nor U19555 (N_19555,N_19092,N_18919);
or U19556 (N_19556,N_18873,N_18819);
nand U19557 (N_19557,N_18760,N_19308);
nor U19558 (N_19558,N_18968,N_19085);
or U19559 (N_19559,N_19275,N_18822);
and U19560 (N_19560,N_18847,N_19177);
nand U19561 (N_19561,N_18949,N_19089);
nor U19562 (N_19562,N_19094,N_18956);
nand U19563 (N_19563,N_18992,N_18955);
xor U19564 (N_19564,N_18827,N_19339);
nor U19565 (N_19565,N_19086,N_19196);
or U19566 (N_19566,N_18906,N_19046);
or U19567 (N_19567,N_19249,N_19256);
xnor U19568 (N_19568,N_19238,N_19347);
or U19569 (N_19569,N_18998,N_19242);
and U19570 (N_19570,N_19276,N_18916);
xor U19571 (N_19571,N_19103,N_18809);
xnor U19572 (N_19572,N_19368,N_19001);
xnor U19573 (N_19573,N_19118,N_19088);
nor U19574 (N_19574,N_18999,N_19263);
nand U19575 (N_19575,N_18889,N_19123);
or U19576 (N_19576,N_19145,N_19052);
and U19577 (N_19577,N_19095,N_19056);
and U19578 (N_19578,N_18950,N_19260);
and U19579 (N_19579,N_18913,N_19309);
or U19580 (N_19580,N_19155,N_19167);
nand U19581 (N_19581,N_18835,N_19366);
xnor U19582 (N_19582,N_19129,N_18939);
or U19583 (N_19583,N_19169,N_19141);
xor U19584 (N_19584,N_18858,N_19295);
and U19585 (N_19585,N_19315,N_18976);
and U19586 (N_19586,N_19372,N_19283);
nor U19587 (N_19587,N_19254,N_19078);
xor U19588 (N_19588,N_19201,N_19068);
or U19589 (N_19589,N_18857,N_19239);
nand U19590 (N_19590,N_18987,N_19361);
nor U19591 (N_19591,N_19229,N_19087);
xor U19592 (N_19592,N_19000,N_18869);
or U19593 (N_19593,N_18828,N_19136);
or U19594 (N_19594,N_19291,N_19012);
nand U19595 (N_19595,N_19271,N_19373);
and U19596 (N_19596,N_18922,N_19152);
nor U19597 (N_19597,N_18902,N_19367);
xor U19598 (N_19598,N_18825,N_19187);
nor U19599 (N_19599,N_19193,N_18966);
nor U19600 (N_19600,N_18888,N_19084);
or U19601 (N_19601,N_18898,N_19132);
xnor U19602 (N_19602,N_19246,N_18808);
or U19603 (N_19603,N_19228,N_19204);
nand U19604 (N_19604,N_19006,N_18849);
nor U19605 (N_19605,N_18799,N_19232);
and U19606 (N_19606,N_18895,N_18941);
nor U19607 (N_19607,N_19099,N_19032);
xor U19608 (N_19608,N_18841,N_19255);
xnor U19609 (N_19609,N_19215,N_19363);
or U19610 (N_19610,N_19076,N_18952);
and U19611 (N_19611,N_19021,N_19051);
and U19612 (N_19612,N_19093,N_18843);
and U19613 (N_19613,N_18946,N_19133);
or U19614 (N_19614,N_18879,N_19066);
or U19615 (N_19615,N_19252,N_19212);
nand U19616 (N_19616,N_18897,N_19108);
nand U19617 (N_19617,N_18932,N_19166);
or U19618 (N_19618,N_18928,N_18991);
nand U19619 (N_19619,N_19190,N_18877);
or U19620 (N_19620,N_19243,N_18832);
nand U19621 (N_19621,N_19044,N_19282);
or U19622 (N_19622,N_19352,N_19119);
nor U19623 (N_19623,N_19163,N_19227);
xor U19624 (N_19624,N_18837,N_18830);
nor U19625 (N_19625,N_19374,N_19111);
or U19626 (N_19626,N_19159,N_19334);
nor U19627 (N_19627,N_18969,N_18797);
and U19628 (N_19628,N_18786,N_18851);
and U19629 (N_19629,N_18970,N_18839);
nand U19630 (N_19630,N_18810,N_18787);
or U19631 (N_19631,N_19172,N_19181);
xor U19632 (N_19632,N_19348,N_18886);
nor U19633 (N_19633,N_19230,N_19300);
xor U19634 (N_19634,N_19064,N_18804);
nand U19635 (N_19635,N_19149,N_19369);
and U19636 (N_19636,N_19269,N_18826);
or U19637 (N_19637,N_19317,N_19062);
and U19638 (N_19638,N_18846,N_19055);
or U19639 (N_19639,N_19307,N_19296);
and U19640 (N_19640,N_18958,N_19330);
or U19641 (N_19641,N_19191,N_19356);
nand U19642 (N_19642,N_18848,N_19341);
nand U19643 (N_19643,N_18853,N_19195);
and U19644 (N_19644,N_19154,N_18973);
nor U19645 (N_19645,N_19281,N_18901);
nand U19646 (N_19646,N_18883,N_18790);
nand U19647 (N_19647,N_19019,N_19261);
and U19648 (N_19648,N_19039,N_18951);
or U19649 (N_19649,N_19045,N_18984);
nand U19650 (N_19650,N_19221,N_18924);
and U19651 (N_19651,N_18892,N_19022);
or U19652 (N_19652,N_19237,N_19250);
nor U19653 (N_19653,N_18751,N_18755);
and U19654 (N_19654,N_18775,N_18954);
nand U19655 (N_19655,N_19286,N_18812);
xor U19656 (N_19656,N_19113,N_19277);
nand U19657 (N_19657,N_18967,N_18824);
nand U19658 (N_19658,N_19173,N_18817);
xnor U19659 (N_19659,N_19091,N_19306);
nor U19660 (N_19660,N_19273,N_19117);
and U19661 (N_19661,N_19160,N_19211);
and U19662 (N_19662,N_19153,N_19015);
nor U19663 (N_19663,N_19139,N_19047);
xor U19664 (N_19664,N_18781,N_18874);
xnor U19665 (N_19665,N_19310,N_18871);
or U19666 (N_19666,N_19234,N_19272);
and U19667 (N_19667,N_19316,N_18798);
and U19668 (N_19668,N_19003,N_19199);
or U19669 (N_19669,N_19259,N_19180);
or U19670 (N_19670,N_19346,N_19161);
nor U19671 (N_19671,N_18844,N_19010);
nor U19672 (N_19672,N_18905,N_19034);
and U19673 (N_19673,N_19326,N_19248);
and U19674 (N_19674,N_19098,N_18814);
xnor U19675 (N_19675,N_19107,N_18813);
nor U19676 (N_19676,N_18978,N_18806);
xnor U19677 (N_19677,N_19157,N_19343);
xor U19678 (N_19678,N_19073,N_19251);
xnor U19679 (N_19679,N_18995,N_18896);
and U19680 (N_19680,N_19183,N_19156);
or U19681 (N_19681,N_19217,N_18977);
xor U19682 (N_19682,N_18936,N_19344);
nand U19683 (N_19683,N_19302,N_18757);
nand U19684 (N_19684,N_18856,N_19331);
xor U19685 (N_19685,N_19218,N_18953);
nor U19686 (N_19686,N_19130,N_19122);
nand U19687 (N_19687,N_19189,N_18974);
and U19688 (N_19688,N_19314,N_19069);
nand U19689 (N_19689,N_19277,N_18898);
xnor U19690 (N_19690,N_19273,N_19131);
nand U19691 (N_19691,N_18790,N_19260);
or U19692 (N_19692,N_19062,N_18840);
or U19693 (N_19693,N_19192,N_18848);
xor U19694 (N_19694,N_19122,N_19199);
and U19695 (N_19695,N_19239,N_19059);
nand U19696 (N_19696,N_19033,N_18979);
nor U19697 (N_19697,N_19113,N_18868);
or U19698 (N_19698,N_19046,N_19246);
xor U19699 (N_19699,N_18851,N_19163);
and U19700 (N_19700,N_19053,N_19180);
and U19701 (N_19701,N_18912,N_19082);
xor U19702 (N_19702,N_19131,N_19066);
xnor U19703 (N_19703,N_19254,N_19031);
nand U19704 (N_19704,N_19251,N_18954);
nand U19705 (N_19705,N_18763,N_18942);
nand U19706 (N_19706,N_19020,N_18924);
nand U19707 (N_19707,N_18887,N_19268);
or U19708 (N_19708,N_19310,N_18976);
nor U19709 (N_19709,N_19006,N_19274);
or U19710 (N_19710,N_19197,N_19175);
nor U19711 (N_19711,N_19103,N_19208);
or U19712 (N_19712,N_18888,N_19117);
or U19713 (N_19713,N_19172,N_19164);
nand U19714 (N_19714,N_19082,N_19353);
nand U19715 (N_19715,N_19208,N_19325);
xor U19716 (N_19716,N_18823,N_19150);
nor U19717 (N_19717,N_18847,N_19109);
and U19718 (N_19718,N_18983,N_19190);
nor U19719 (N_19719,N_18848,N_19172);
and U19720 (N_19720,N_19205,N_19124);
and U19721 (N_19721,N_19316,N_18902);
nor U19722 (N_19722,N_19014,N_19148);
or U19723 (N_19723,N_18973,N_19273);
or U19724 (N_19724,N_19360,N_19134);
xnor U19725 (N_19725,N_19345,N_19230);
or U19726 (N_19726,N_18937,N_19233);
and U19727 (N_19727,N_18986,N_19328);
or U19728 (N_19728,N_18916,N_19239);
nand U19729 (N_19729,N_19189,N_19235);
xnor U19730 (N_19730,N_18960,N_19284);
xor U19731 (N_19731,N_19093,N_18806);
and U19732 (N_19732,N_19178,N_18962);
and U19733 (N_19733,N_19183,N_18909);
nor U19734 (N_19734,N_19209,N_18801);
and U19735 (N_19735,N_18890,N_19007);
or U19736 (N_19736,N_18760,N_18930);
xnor U19737 (N_19737,N_18980,N_18804);
and U19738 (N_19738,N_18769,N_19198);
or U19739 (N_19739,N_19047,N_18972);
and U19740 (N_19740,N_18884,N_18969);
and U19741 (N_19741,N_18919,N_19137);
or U19742 (N_19742,N_19187,N_19161);
and U19743 (N_19743,N_19130,N_19038);
nand U19744 (N_19744,N_18992,N_18903);
nor U19745 (N_19745,N_18989,N_19027);
xnor U19746 (N_19746,N_19002,N_18957);
or U19747 (N_19747,N_19331,N_19325);
nor U19748 (N_19748,N_19211,N_18933);
or U19749 (N_19749,N_19149,N_18927);
or U19750 (N_19750,N_19177,N_19336);
xnor U19751 (N_19751,N_19157,N_19242);
and U19752 (N_19752,N_19147,N_19007);
nand U19753 (N_19753,N_18920,N_19078);
or U19754 (N_19754,N_19203,N_19109);
or U19755 (N_19755,N_18889,N_19017);
and U19756 (N_19756,N_18925,N_18990);
and U19757 (N_19757,N_19018,N_18893);
and U19758 (N_19758,N_18836,N_18755);
and U19759 (N_19759,N_19246,N_18846);
and U19760 (N_19760,N_18873,N_18856);
nor U19761 (N_19761,N_18761,N_19247);
xnor U19762 (N_19762,N_19021,N_19133);
nand U19763 (N_19763,N_18895,N_19172);
or U19764 (N_19764,N_19195,N_18890);
and U19765 (N_19765,N_18986,N_18846);
nand U19766 (N_19766,N_19082,N_18900);
xnor U19767 (N_19767,N_19036,N_19124);
nand U19768 (N_19768,N_19161,N_18775);
xnor U19769 (N_19769,N_19286,N_18873);
or U19770 (N_19770,N_18937,N_19008);
xor U19771 (N_19771,N_19037,N_18861);
nor U19772 (N_19772,N_18889,N_18938);
nor U19773 (N_19773,N_18884,N_19281);
nor U19774 (N_19774,N_19184,N_19083);
nand U19775 (N_19775,N_19231,N_18836);
xnor U19776 (N_19776,N_18810,N_18917);
nor U19777 (N_19777,N_18941,N_18810);
and U19778 (N_19778,N_19147,N_19306);
xor U19779 (N_19779,N_19173,N_18764);
nor U19780 (N_19780,N_19123,N_19233);
nor U19781 (N_19781,N_19314,N_19145);
nor U19782 (N_19782,N_19331,N_19162);
nand U19783 (N_19783,N_18884,N_19233);
and U19784 (N_19784,N_19305,N_19318);
and U19785 (N_19785,N_19190,N_19312);
nor U19786 (N_19786,N_18855,N_18922);
xnor U19787 (N_19787,N_19241,N_18902);
nand U19788 (N_19788,N_19356,N_18981);
nor U19789 (N_19789,N_18937,N_18837);
xnor U19790 (N_19790,N_18927,N_19162);
and U19791 (N_19791,N_18823,N_18964);
nor U19792 (N_19792,N_18955,N_18958);
xor U19793 (N_19793,N_18967,N_19180);
xnor U19794 (N_19794,N_19121,N_18844);
nand U19795 (N_19795,N_19033,N_19021);
xor U19796 (N_19796,N_18793,N_19225);
or U19797 (N_19797,N_18752,N_19274);
xor U19798 (N_19798,N_19343,N_19151);
or U19799 (N_19799,N_19108,N_18935);
xnor U19800 (N_19800,N_18964,N_18893);
nand U19801 (N_19801,N_19108,N_18895);
xor U19802 (N_19802,N_18873,N_18822);
or U19803 (N_19803,N_18750,N_19359);
xor U19804 (N_19804,N_19199,N_18771);
nor U19805 (N_19805,N_19196,N_18777);
and U19806 (N_19806,N_18757,N_18904);
and U19807 (N_19807,N_18879,N_18816);
and U19808 (N_19808,N_18770,N_18839);
xor U19809 (N_19809,N_19105,N_19249);
nand U19810 (N_19810,N_19170,N_19203);
and U19811 (N_19811,N_18774,N_19265);
or U19812 (N_19812,N_19308,N_19169);
nor U19813 (N_19813,N_18977,N_19193);
xnor U19814 (N_19814,N_18847,N_19298);
xnor U19815 (N_19815,N_18863,N_19160);
xnor U19816 (N_19816,N_18782,N_19201);
nor U19817 (N_19817,N_19353,N_18865);
or U19818 (N_19818,N_18876,N_19239);
nand U19819 (N_19819,N_19229,N_18904);
or U19820 (N_19820,N_19266,N_19364);
xnor U19821 (N_19821,N_19269,N_19352);
nor U19822 (N_19822,N_19045,N_19199);
nor U19823 (N_19823,N_19299,N_18773);
xnor U19824 (N_19824,N_18774,N_19070);
xor U19825 (N_19825,N_19070,N_18949);
nor U19826 (N_19826,N_19074,N_18783);
nor U19827 (N_19827,N_18894,N_18999);
or U19828 (N_19828,N_18916,N_18893);
nor U19829 (N_19829,N_18897,N_19101);
and U19830 (N_19830,N_19052,N_19183);
nand U19831 (N_19831,N_19078,N_19276);
or U19832 (N_19832,N_18808,N_18857);
xnor U19833 (N_19833,N_19106,N_19091);
nor U19834 (N_19834,N_19217,N_19011);
or U19835 (N_19835,N_19245,N_19304);
or U19836 (N_19836,N_19007,N_18981);
and U19837 (N_19837,N_19035,N_19247);
or U19838 (N_19838,N_18890,N_19163);
xnor U19839 (N_19839,N_19366,N_18859);
nor U19840 (N_19840,N_19287,N_19124);
nor U19841 (N_19841,N_19022,N_19038);
nor U19842 (N_19842,N_19049,N_19007);
xnor U19843 (N_19843,N_19203,N_18939);
and U19844 (N_19844,N_18984,N_19027);
and U19845 (N_19845,N_18989,N_18829);
nand U19846 (N_19846,N_19080,N_19074);
nand U19847 (N_19847,N_19373,N_18932);
nor U19848 (N_19848,N_19371,N_18866);
nand U19849 (N_19849,N_18795,N_18903);
nand U19850 (N_19850,N_18944,N_18935);
and U19851 (N_19851,N_19329,N_19116);
or U19852 (N_19852,N_18861,N_18933);
nor U19853 (N_19853,N_19293,N_18810);
or U19854 (N_19854,N_19034,N_19033);
or U19855 (N_19855,N_19074,N_19331);
xor U19856 (N_19856,N_18907,N_18996);
and U19857 (N_19857,N_18801,N_19367);
or U19858 (N_19858,N_19085,N_19010);
and U19859 (N_19859,N_18844,N_18956);
and U19860 (N_19860,N_18906,N_19372);
nor U19861 (N_19861,N_19074,N_19329);
and U19862 (N_19862,N_18836,N_19070);
and U19863 (N_19863,N_18981,N_19275);
or U19864 (N_19864,N_19231,N_19046);
nor U19865 (N_19865,N_19256,N_19329);
or U19866 (N_19866,N_19212,N_19356);
xor U19867 (N_19867,N_19331,N_19372);
nand U19868 (N_19868,N_19113,N_19099);
and U19869 (N_19869,N_18964,N_18941);
or U19870 (N_19870,N_19084,N_18776);
xnor U19871 (N_19871,N_18835,N_18795);
nand U19872 (N_19872,N_19067,N_18845);
nor U19873 (N_19873,N_19352,N_18934);
xor U19874 (N_19874,N_19343,N_19112);
and U19875 (N_19875,N_19207,N_19374);
nor U19876 (N_19876,N_19021,N_18913);
xnor U19877 (N_19877,N_18756,N_18881);
xnor U19878 (N_19878,N_19080,N_19159);
nor U19879 (N_19879,N_19110,N_19254);
or U19880 (N_19880,N_18865,N_18999);
xor U19881 (N_19881,N_19318,N_18876);
nand U19882 (N_19882,N_19071,N_19024);
nor U19883 (N_19883,N_19231,N_19279);
and U19884 (N_19884,N_19295,N_18944);
and U19885 (N_19885,N_19367,N_19255);
nand U19886 (N_19886,N_18944,N_18934);
xor U19887 (N_19887,N_19297,N_19150);
nand U19888 (N_19888,N_19061,N_19114);
or U19889 (N_19889,N_19033,N_19068);
nor U19890 (N_19890,N_19107,N_18917);
nor U19891 (N_19891,N_19255,N_18791);
xnor U19892 (N_19892,N_19361,N_19257);
nor U19893 (N_19893,N_18805,N_18924);
nor U19894 (N_19894,N_18939,N_19177);
nor U19895 (N_19895,N_18791,N_19009);
xor U19896 (N_19896,N_19208,N_19159);
nor U19897 (N_19897,N_19113,N_18892);
or U19898 (N_19898,N_18820,N_19132);
or U19899 (N_19899,N_18829,N_19050);
and U19900 (N_19900,N_19239,N_18993);
nand U19901 (N_19901,N_19231,N_18951);
nand U19902 (N_19902,N_18785,N_19022);
and U19903 (N_19903,N_19064,N_19259);
xor U19904 (N_19904,N_18868,N_19193);
nand U19905 (N_19905,N_18917,N_19217);
and U19906 (N_19906,N_19173,N_18843);
xor U19907 (N_19907,N_18855,N_19017);
nand U19908 (N_19908,N_19078,N_18935);
nor U19909 (N_19909,N_19299,N_19166);
or U19910 (N_19910,N_18822,N_18996);
xnor U19911 (N_19911,N_18786,N_19347);
xor U19912 (N_19912,N_18857,N_19103);
nand U19913 (N_19913,N_19035,N_19082);
xnor U19914 (N_19914,N_19274,N_19063);
and U19915 (N_19915,N_19053,N_19070);
nor U19916 (N_19916,N_18930,N_19372);
nand U19917 (N_19917,N_19279,N_18831);
nand U19918 (N_19918,N_19369,N_18808);
and U19919 (N_19919,N_19372,N_18909);
and U19920 (N_19920,N_19266,N_19270);
xor U19921 (N_19921,N_19366,N_19220);
and U19922 (N_19922,N_19038,N_19088);
xnor U19923 (N_19923,N_19371,N_19149);
nand U19924 (N_19924,N_19324,N_18830);
nor U19925 (N_19925,N_19316,N_19029);
nand U19926 (N_19926,N_18799,N_19326);
or U19927 (N_19927,N_19192,N_19066);
nor U19928 (N_19928,N_19033,N_18902);
nor U19929 (N_19929,N_18904,N_19146);
nand U19930 (N_19930,N_19056,N_19009);
and U19931 (N_19931,N_19195,N_18815);
and U19932 (N_19932,N_19003,N_18827);
nand U19933 (N_19933,N_19114,N_19204);
nor U19934 (N_19934,N_19142,N_18768);
nand U19935 (N_19935,N_19274,N_18804);
or U19936 (N_19936,N_19231,N_18783);
and U19937 (N_19937,N_19315,N_19043);
nor U19938 (N_19938,N_18763,N_19183);
xor U19939 (N_19939,N_19221,N_18948);
nand U19940 (N_19940,N_19204,N_19091);
and U19941 (N_19941,N_19072,N_19000);
nand U19942 (N_19942,N_18848,N_19260);
and U19943 (N_19943,N_18772,N_18883);
xnor U19944 (N_19944,N_18952,N_18769);
nor U19945 (N_19945,N_18794,N_19267);
nor U19946 (N_19946,N_19199,N_19154);
xnor U19947 (N_19947,N_18903,N_19088);
and U19948 (N_19948,N_19253,N_18873);
nor U19949 (N_19949,N_19128,N_18819);
or U19950 (N_19950,N_18863,N_19274);
xnor U19951 (N_19951,N_18907,N_19268);
or U19952 (N_19952,N_19059,N_19350);
and U19953 (N_19953,N_19075,N_19224);
nand U19954 (N_19954,N_18769,N_19216);
nand U19955 (N_19955,N_19128,N_19134);
nor U19956 (N_19956,N_19173,N_19324);
or U19957 (N_19957,N_18808,N_19201);
or U19958 (N_19958,N_19053,N_19269);
nand U19959 (N_19959,N_19166,N_19123);
or U19960 (N_19960,N_19111,N_19101);
and U19961 (N_19961,N_18915,N_18889);
or U19962 (N_19962,N_18899,N_18880);
nand U19963 (N_19963,N_19204,N_18930);
nand U19964 (N_19964,N_18801,N_18981);
or U19965 (N_19965,N_19214,N_19046);
xnor U19966 (N_19966,N_19062,N_19158);
xor U19967 (N_19967,N_19086,N_19057);
and U19968 (N_19968,N_19047,N_19258);
and U19969 (N_19969,N_19201,N_19341);
nand U19970 (N_19970,N_18776,N_19245);
nand U19971 (N_19971,N_19037,N_19229);
and U19972 (N_19972,N_18756,N_18934);
nand U19973 (N_19973,N_18864,N_19244);
and U19974 (N_19974,N_18797,N_19165);
xnor U19975 (N_19975,N_19228,N_18857);
xnor U19976 (N_19976,N_18949,N_18796);
and U19977 (N_19977,N_19214,N_19027);
xor U19978 (N_19978,N_18794,N_19244);
xor U19979 (N_19979,N_19350,N_18991);
xnor U19980 (N_19980,N_18945,N_19274);
or U19981 (N_19981,N_19228,N_18877);
xnor U19982 (N_19982,N_18879,N_18890);
xnor U19983 (N_19983,N_19148,N_19080);
nand U19984 (N_19984,N_18945,N_19102);
xnor U19985 (N_19985,N_19247,N_19278);
nand U19986 (N_19986,N_18760,N_19131);
nor U19987 (N_19987,N_18966,N_19162);
nand U19988 (N_19988,N_19213,N_18898);
nor U19989 (N_19989,N_18950,N_19301);
or U19990 (N_19990,N_19191,N_19300);
nor U19991 (N_19991,N_19011,N_18891);
xnor U19992 (N_19992,N_19146,N_18895);
or U19993 (N_19993,N_19341,N_19335);
xnor U19994 (N_19994,N_18839,N_19222);
nor U19995 (N_19995,N_18751,N_18974);
xnor U19996 (N_19996,N_19241,N_18906);
nor U19997 (N_19997,N_19213,N_18808);
nor U19998 (N_19998,N_18787,N_19124);
xnor U19999 (N_19999,N_19197,N_19319);
and U20000 (N_20000,N_19651,N_19870);
nor U20001 (N_20001,N_19965,N_19503);
and U20002 (N_20002,N_19936,N_19866);
nand U20003 (N_20003,N_19874,N_19898);
xnor U20004 (N_20004,N_19468,N_19706);
and U20005 (N_20005,N_19774,N_19384);
nand U20006 (N_20006,N_19598,N_19457);
nor U20007 (N_20007,N_19765,N_19612);
nor U20008 (N_20008,N_19982,N_19822);
or U20009 (N_20009,N_19692,N_19970);
nor U20010 (N_20010,N_19516,N_19449);
xor U20011 (N_20011,N_19740,N_19672);
and U20012 (N_20012,N_19572,N_19865);
nor U20013 (N_20013,N_19742,N_19971);
xnor U20014 (N_20014,N_19677,N_19434);
and U20015 (N_20015,N_19416,N_19981);
nand U20016 (N_20016,N_19633,N_19940);
or U20017 (N_20017,N_19423,N_19404);
or U20018 (N_20018,N_19979,N_19844);
or U20019 (N_20019,N_19479,N_19688);
nor U20020 (N_20020,N_19925,N_19494);
and U20021 (N_20021,N_19796,N_19816);
nand U20022 (N_20022,N_19665,N_19858);
and U20023 (N_20023,N_19725,N_19535);
or U20024 (N_20024,N_19775,N_19689);
nand U20025 (N_20025,N_19398,N_19393);
nand U20026 (N_20026,N_19795,N_19698);
or U20027 (N_20027,N_19712,N_19838);
and U20028 (N_20028,N_19442,N_19536);
or U20029 (N_20029,N_19653,N_19949);
nand U20030 (N_20030,N_19426,N_19611);
nor U20031 (N_20031,N_19475,N_19744);
nor U20032 (N_20032,N_19815,N_19854);
nor U20033 (N_20033,N_19730,N_19837);
nor U20034 (N_20034,N_19827,N_19558);
or U20035 (N_20035,N_19380,N_19548);
or U20036 (N_20036,N_19968,N_19717);
and U20037 (N_20037,N_19962,N_19711);
or U20038 (N_20038,N_19439,N_19552);
and U20039 (N_20039,N_19853,N_19509);
or U20040 (N_20040,N_19731,N_19459);
or U20041 (N_20041,N_19763,N_19986);
nor U20042 (N_20042,N_19451,N_19830);
nand U20043 (N_20043,N_19504,N_19570);
nor U20044 (N_20044,N_19780,N_19669);
nand U20045 (N_20045,N_19998,N_19578);
nor U20046 (N_20046,N_19583,N_19424);
and U20047 (N_20047,N_19593,N_19631);
nand U20048 (N_20048,N_19691,N_19828);
or U20049 (N_20049,N_19544,N_19462);
xor U20050 (N_20050,N_19739,N_19464);
or U20051 (N_20051,N_19630,N_19715);
or U20052 (N_20052,N_19762,N_19794);
xnor U20053 (N_20053,N_19819,N_19681);
and U20054 (N_20054,N_19871,N_19522);
xor U20055 (N_20055,N_19834,N_19879);
nand U20056 (N_20056,N_19953,N_19663);
nand U20057 (N_20057,N_19541,N_19802);
or U20058 (N_20058,N_19679,N_19942);
and U20059 (N_20059,N_19957,N_19642);
nand U20060 (N_20060,N_19619,N_19496);
and U20061 (N_20061,N_19980,N_19594);
nor U20062 (N_20062,N_19894,N_19841);
nand U20063 (N_20063,N_19845,N_19421);
or U20064 (N_20064,N_19564,N_19389);
and U20065 (N_20065,N_19502,N_19429);
nand U20066 (N_20066,N_19403,N_19568);
or U20067 (N_20067,N_19883,N_19929);
and U20068 (N_20068,N_19718,N_19878);
nand U20069 (N_20069,N_19961,N_19420);
nand U20070 (N_20070,N_19767,N_19835);
nand U20071 (N_20071,N_19667,N_19895);
nand U20072 (N_20072,N_19450,N_19397);
and U20073 (N_20073,N_19527,N_19388);
or U20074 (N_20074,N_19955,N_19406);
and U20075 (N_20075,N_19662,N_19812);
nor U20076 (N_20076,N_19484,N_19738);
and U20077 (N_20077,N_19620,N_19799);
and U20078 (N_20078,N_19975,N_19480);
xor U20079 (N_20079,N_19753,N_19410);
xor U20080 (N_20080,N_19614,N_19787);
xnor U20081 (N_20081,N_19576,N_19749);
or U20082 (N_20082,N_19560,N_19921);
nor U20083 (N_20083,N_19400,N_19624);
xor U20084 (N_20084,N_19716,N_19719);
and U20085 (N_20085,N_19656,N_19847);
xnor U20086 (N_20086,N_19638,N_19938);
or U20087 (N_20087,N_19991,N_19820);
and U20088 (N_20088,N_19566,N_19987);
xnor U20089 (N_20089,N_19481,N_19513);
and U20090 (N_20090,N_19759,N_19413);
nand U20091 (N_20091,N_19990,N_19761);
and U20092 (N_20092,N_19944,N_19732);
xor U20093 (N_20093,N_19563,N_19747);
nand U20094 (N_20094,N_19632,N_19924);
and U20095 (N_20095,N_19378,N_19618);
xnor U20096 (N_20096,N_19432,N_19546);
xor U20097 (N_20097,N_19797,N_19456);
and U20098 (N_20098,N_19628,N_19993);
and U20099 (N_20099,N_19776,N_19728);
nand U20100 (N_20100,N_19913,N_19448);
and U20101 (N_20101,N_19860,N_19491);
or U20102 (N_20102,N_19801,N_19682);
nor U20103 (N_20103,N_19673,N_19495);
nand U20104 (N_20104,N_19466,N_19512);
or U20105 (N_20105,N_19863,N_19402);
nand U20106 (N_20106,N_19637,N_19640);
xnor U20107 (N_20107,N_19909,N_19528);
xnor U20108 (N_20108,N_19600,N_19463);
nor U20109 (N_20109,N_19997,N_19989);
xor U20110 (N_20110,N_19999,N_19994);
or U20111 (N_20111,N_19721,N_19707);
or U20112 (N_20112,N_19789,N_19649);
or U20113 (N_20113,N_19607,N_19983);
nor U20114 (N_20114,N_19606,N_19533);
nand U20115 (N_20115,N_19967,N_19788);
nand U20116 (N_20116,N_19490,N_19394);
nor U20117 (N_20117,N_19574,N_19786);
xnor U20118 (N_20118,N_19823,N_19557);
xnor U20119 (N_20119,N_19538,N_19727);
nor U20120 (N_20120,N_19671,N_19508);
nand U20121 (N_20121,N_19932,N_19948);
nand U20122 (N_20122,N_19554,N_19696);
and U20123 (N_20123,N_19960,N_19793);
and U20124 (N_20124,N_19876,N_19903);
and U20125 (N_20125,N_19390,N_19811);
nand U20126 (N_20126,N_19680,N_19455);
xor U20127 (N_20127,N_19585,N_19708);
nand U20128 (N_20128,N_19399,N_19922);
or U20129 (N_20129,N_19988,N_19567);
nor U20130 (N_20130,N_19805,N_19613);
and U20131 (N_20131,N_19750,N_19650);
nor U20132 (N_20132,N_19754,N_19984);
and U20133 (N_20133,N_19777,N_19526);
and U20134 (N_20134,N_19447,N_19918);
xor U20135 (N_20135,N_19724,N_19621);
nor U20136 (N_20136,N_19843,N_19935);
nor U20137 (N_20137,N_19800,N_19829);
nor U20138 (N_20138,N_19849,N_19422);
nor U20139 (N_20139,N_19617,N_19969);
nor U20140 (N_20140,N_19582,N_19931);
nand U20141 (N_20141,N_19722,N_19684);
and U20142 (N_20142,N_19460,N_19781);
or U20143 (N_20143,N_19930,N_19972);
or U20144 (N_20144,N_19499,N_19493);
nand U20145 (N_20145,N_19911,N_19872);
xnor U20146 (N_20146,N_19419,N_19427);
nor U20147 (N_20147,N_19756,N_19889);
xnor U20148 (N_20148,N_19498,N_19483);
nor U20149 (N_20149,N_19588,N_19927);
nor U20150 (N_20150,N_19565,N_19492);
nor U20151 (N_20151,N_19609,N_19531);
nand U20152 (N_20152,N_19610,N_19848);
nor U20153 (N_20153,N_19881,N_19386);
and U20154 (N_20154,N_19454,N_19584);
or U20155 (N_20155,N_19379,N_19412);
xnor U20156 (N_20156,N_19446,N_19652);
or U20157 (N_20157,N_19912,N_19720);
and U20158 (N_20158,N_19813,N_19791);
or U20159 (N_20159,N_19690,N_19868);
nor U20160 (N_20160,N_19603,N_19798);
nor U20161 (N_20161,N_19933,N_19745);
and U20162 (N_20162,N_19452,N_19976);
and U20163 (N_20163,N_19519,N_19615);
and U20164 (N_20164,N_19375,N_19657);
nand U20165 (N_20165,N_19809,N_19770);
nor U20166 (N_20166,N_19861,N_19532);
nor U20167 (N_20167,N_19697,N_19401);
xor U20168 (N_20168,N_19445,N_19807);
nand U20169 (N_20169,N_19573,N_19951);
and U20170 (N_20170,N_19947,N_19840);
nor U20171 (N_20171,N_19857,N_19596);
nor U20172 (N_20172,N_19977,N_19501);
xnor U20173 (N_20173,N_19973,N_19907);
and U20174 (N_20174,N_19595,N_19525);
and U20175 (N_20175,N_19824,N_19952);
nand U20176 (N_20176,N_19832,N_19647);
and U20177 (N_20177,N_19411,N_19443);
and U20178 (N_20178,N_19623,N_19683);
xnor U20179 (N_20179,N_19655,N_19906);
nand U20180 (N_20180,N_19597,N_19592);
nor U20181 (N_20181,N_19414,N_19897);
xnor U20182 (N_20182,N_19937,N_19555);
nand U20183 (N_20183,N_19441,N_19709);
nor U20184 (N_20184,N_19825,N_19985);
nor U20185 (N_20185,N_19859,N_19629);
or U20186 (N_20186,N_19852,N_19729);
nand U20187 (N_20187,N_19392,N_19641);
nand U20188 (N_20188,N_19836,N_19458);
xnor U20189 (N_20189,N_19575,N_19757);
xor U20190 (N_20190,N_19995,N_19896);
nor U20191 (N_20191,N_19507,N_19383);
or U20192 (N_20192,N_19687,N_19648);
or U20193 (N_20193,N_19864,N_19635);
nand U20194 (N_20194,N_19803,N_19486);
nor U20195 (N_20195,N_19685,N_19645);
nand U20196 (N_20196,N_19417,N_19471);
nor U20197 (N_20197,N_19856,N_19407);
and U20198 (N_20198,N_19437,N_19601);
or U20199 (N_20199,N_19833,N_19892);
nand U20200 (N_20200,N_19808,N_19875);
nor U20201 (N_20201,N_19425,N_19473);
and U20202 (N_20202,N_19551,N_19659);
nand U20203 (N_20203,N_19626,N_19604);
nand U20204 (N_20204,N_19428,N_19752);
xnor U20205 (N_20205,N_19511,N_19764);
xnor U20206 (N_20206,N_19549,N_19939);
and U20207 (N_20207,N_19545,N_19735);
or U20208 (N_20208,N_19751,N_19608);
and U20209 (N_20209,N_19950,N_19550);
and U20210 (N_20210,N_19839,N_19736);
nor U20211 (N_20211,N_19644,N_19470);
nor U20212 (N_20212,N_19435,N_19755);
nor U20213 (N_20213,N_19943,N_19477);
and U20214 (N_20214,N_19666,N_19946);
nor U20215 (N_20215,N_19902,N_19636);
and U20216 (N_20216,N_19766,N_19415);
xor U20217 (N_20217,N_19701,N_19916);
xnor U20218 (N_20218,N_19467,N_19846);
or U20219 (N_20219,N_19743,N_19395);
and U20220 (N_20220,N_19885,N_19867);
or U20221 (N_20221,N_19873,N_19431);
and U20222 (N_20222,N_19627,N_19489);
nand U20223 (N_20223,N_19444,N_19625);
nor U20224 (N_20224,N_19741,N_19804);
and U20225 (N_20225,N_19882,N_19562);
xor U20226 (N_20226,N_19855,N_19810);
and U20227 (N_20227,N_19524,N_19919);
or U20228 (N_20228,N_19561,N_19699);
nor U20229 (N_20229,N_19643,N_19616);
nand U20230 (N_20230,N_19577,N_19487);
and U20231 (N_20231,N_19886,N_19478);
nor U20232 (N_20232,N_19862,N_19978);
xnor U20233 (N_20233,N_19959,N_19587);
and U20234 (N_20234,N_19469,N_19589);
xor U20235 (N_20235,N_19992,N_19580);
and U20236 (N_20236,N_19704,N_19530);
nand U20237 (N_20237,N_19826,N_19778);
nor U20238 (N_20238,N_19670,N_19482);
nor U20239 (N_20239,N_19851,N_19784);
or U20240 (N_20240,N_19668,N_19622);
or U20241 (N_20241,N_19387,N_19382);
and U20242 (N_20242,N_19817,N_19880);
and U20243 (N_20243,N_19945,N_19887);
or U20244 (N_20244,N_19510,N_19433);
nor U20245 (N_20245,N_19996,N_19639);
or U20246 (N_20246,N_19539,N_19914);
xor U20247 (N_20247,N_19408,N_19806);
nand U20248 (N_20248,N_19705,N_19385);
nand U20249 (N_20249,N_19694,N_19377);
and U20250 (N_20250,N_19405,N_19904);
nor U20251 (N_20251,N_19605,N_19954);
nor U20252 (N_20252,N_19569,N_19773);
nor U20253 (N_20253,N_19521,N_19440);
nand U20254 (N_20254,N_19702,N_19520);
and U20255 (N_20255,N_19461,N_19831);
or U20256 (N_20256,N_19540,N_19926);
xor U20257 (N_20257,N_19488,N_19418);
and U20258 (N_20258,N_19964,N_19381);
and U20259 (N_20259,N_19695,N_19658);
nor U20260 (N_20260,N_19453,N_19686);
xor U20261 (N_20261,N_19726,N_19664);
nor U20262 (N_20262,N_19771,N_19910);
xnor U20263 (N_20263,N_19571,N_19915);
xnor U20264 (N_20264,N_19529,N_19966);
or U20265 (N_20265,N_19772,N_19714);
nor U20266 (N_20266,N_19900,N_19893);
and U20267 (N_20267,N_19505,N_19792);
nand U20268 (N_20268,N_19591,N_19586);
xnor U20269 (N_20269,N_19737,N_19901);
nand U20270 (N_20270,N_19506,N_19654);
nor U20271 (N_20271,N_19941,N_19537);
nand U20272 (N_20272,N_19884,N_19472);
and U20273 (N_20273,N_19465,N_19923);
and U20274 (N_20274,N_19917,N_19409);
and U20275 (N_20275,N_19850,N_19928);
nand U20276 (N_20276,N_19474,N_19559);
nor U20277 (N_20277,N_19890,N_19678);
nand U20278 (N_20278,N_19703,N_19783);
and U20279 (N_20279,N_19700,N_19877);
nand U20280 (N_20280,N_19956,N_19391);
xnor U20281 (N_20281,N_19869,N_19818);
nor U20282 (N_20282,N_19590,N_19634);
nor U20283 (N_20283,N_19599,N_19674);
nand U20284 (N_20284,N_19543,N_19891);
and U20285 (N_20285,N_19779,N_19958);
or U20286 (N_20286,N_19842,N_19710);
and U20287 (N_20287,N_19888,N_19769);
or U20288 (N_20288,N_19693,N_19790);
xor U20289 (N_20289,N_19396,N_19734);
xor U20290 (N_20290,N_19514,N_19713);
or U20291 (N_20291,N_19547,N_19733);
xor U20292 (N_20292,N_19785,N_19661);
nor U20293 (N_20293,N_19542,N_19646);
and U20294 (N_20294,N_19515,N_19963);
and U20295 (N_20295,N_19518,N_19556);
nor U20296 (N_20296,N_19602,N_19934);
nor U20297 (N_20297,N_19746,N_19758);
or U20298 (N_20298,N_19523,N_19974);
and U20299 (N_20299,N_19814,N_19760);
or U20300 (N_20300,N_19920,N_19748);
nand U20301 (N_20301,N_19821,N_19782);
or U20302 (N_20302,N_19436,N_19376);
or U20303 (N_20303,N_19534,N_19485);
xor U20304 (N_20304,N_19553,N_19908);
or U20305 (N_20305,N_19676,N_19438);
nor U20306 (N_20306,N_19675,N_19899);
nor U20307 (N_20307,N_19517,N_19905);
and U20308 (N_20308,N_19430,N_19500);
or U20309 (N_20309,N_19581,N_19497);
and U20310 (N_20310,N_19660,N_19579);
nand U20311 (N_20311,N_19476,N_19723);
nand U20312 (N_20312,N_19768,N_19847);
nand U20313 (N_20313,N_19954,N_19434);
xnor U20314 (N_20314,N_19737,N_19888);
xor U20315 (N_20315,N_19535,N_19915);
xor U20316 (N_20316,N_19913,N_19813);
or U20317 (N_20317,N_19832,N_19998);
nand U20318 (N_20318,N_19851,N_19835);
nor U20319 (N_20319,N_19468,N_19498);
or U20320 (N_20320,N_19788,N_19428);
nor U20321 (N_20321,N_19594,N_19505);
and U20322 (N_20322,N_19722,N_19889);
nand U20323 (N_20323,N_19609,N_19398);
and U20324 (N_20324,N_19865,N_19906);
nor U20325 (N_20325,N_19567,N_19549);
and U20326 (N_20326,N_19843,N_19691);
or U20327 (N_20327,N_19547,N_19411);
or U20328 (N_20328,N_19747,N_19542);
nand U20329 (N_20329,N_19765,N_19820);
nand U20330 (N_20330,N_19621,N_19604);
and U20331 (N_20331,N_19802,N_19971);
and U20332 (N_20332,N_19443,N_19855);
nor U20333 (N_20333,N_19582,N_19972);
or U20334 (N_20334,N_19530,N_19941);
or U20335 (N_20335,N_19395,N_19907);
xnor U20336 (N_20336,N_19864,N_19731);
nor U20337 (N_20337,N_19825,N_19411);
or U20338 (N_20338,N_19483,N_19793);
or U20339 (N_20339,N_19468,N_19787);
xor U20340 (N_20340,N_19645,N_19583);
nand U20341 (N_20341,N_19412,N_19986);
xnor U20342 (N_20342,N_19943,N_19584);
nand U20343 (N_20343,N_19525,N_19964);
nor U20344 (N_20344,N_19502,N_19645);
xnor U20345 (N_20345,N_19676,N_19904);
xor U20346 (N_20346,N_19401,N_19985);
nor U20347 (N_20347,N_19957,N_19849);
and U20348 (N_20348,N_19990,N_19661);
xor U20349 (N_20349,N_19561,N_19851);
xnor U20350 (N_20350,N_19778,N_19389);
nand U20351 (N_20351,N_19969,N_19392);
and U20352 (N_20352,N_19777,N_19898);
nor U20353 (N_20353,N_19912,N_19468);
nand U20354 (N_20354,N_19739,N_19579);
xnor U20355 (N_20355,N_19601,N_19452);
or U20356 (N_20356,N_19683,N_19914);
or U20357 (N_20357,N_19852,N_19411);
or U20358 (N_20358,N_19733,N_19499);
and U20359 (N_20359,N_19661,N_19544);
nand U20360 (N_20360,N_19706,N_19818);
or U20361 (N_20361,N_19854,N_19510);
xor U20362 (N_20362,N_19927,N_19590);
and U20363 (N_20363,N_19939,N_19614);
and U20364 (N_20364,N_19512,N_19856);
xor U20365 (N_20365,N_19706,N_19709);
or U20366 (N_20366,N_19574,N_19604);
and U20367 (N_20367,N_19528,N_19833);
nand U20368 (N_20368,N_19427,N_19437);
xnor U20369 (N_20369,N_19561,N_19999);
or U20370 (N_20370,N_19618,N_19572);
nor U20371 (N_20371,N_19571,N_19413);
or U20372 (N_20372,N_19493,N_19706);
nor U20373 (N_20373,N_19540,N_19997);
or U20374 (N_20374,N_19446,N_19630);
or U20375 (N_20375,N_19575,N_19570);
nor U20376 (N_20376,N_19637,N_19721);
nand U20377 (N_20377,N_19583,N_19436);
or U20378 (N_20378,N_19889,N_19501);
or U20379 (N_20379,N_19491,N_19390);
nand U20380 (N_20380,N_19753,N_19500);
and U20381 (N_20381,N_19711,N_19579);
nor U20382 (N_20382,N_19948,N_19584);
nor U20383 (N_20383,N_19480,N_19643);
or U20384 (N_20384,N_19381,N_19987);
xor U20385 (N_20385,N_19745,N_19627);
and U20386 (N_20386,N_19999,N_19453);
xor U20387 (N_20387,N_19686,N_19884);
nand U20388 (N_20388,N_19733,N_19697);
or U20389 (N_20389,N_19632,N_19936);
and U20390 (N_20390,N_19464,N_19719);
or U20391 (N_20391,N_19557,N_19710);
or U20392 (N_20392,N_19818,N_19816);
nand U20393 (N_20393,N_19972,N_19875);
or U20394 (N_20394,N_19832,N_19683);
nand U20395 (N_20395,N_19420,N_19564);
nor U20396 (N_20396,N_19767,N_19868);
nor U20397 (N_20397,N_19903,N_19591);
xnor U20398 (N_20398,N_19791,N_19899);
xor U20399 (N_20399,N_19914,N_19933);
nand U20400 (N_20400,N_19996,N_19610);
xnor U20401 (N_20401,N_19569,N_19411);
and U20402 (N_20402,N_19681,N_19487);
nor U20403 (N_20403,N_19520,N_19565);
nand U20404 (N_20404,N_19958,N_19830);
or U20405 (N_20405,N_19959,N_19508);
nand U20406 (N_20406,N_19574,N_19547);
and U20407 (N_20407,N_19886,N_19888);
xor U20408 (N_20408,N_19987,N_19837);
xnor U20409 (N_20409,N_19814,N_19396);
and U20410 (N_20410,N_19428,N_19815);
or U20411 (N_20411,N_19652,N_19920);
xor U20412 (N_20412,N_19779,N_19816);
nor U20413 (N_20413,N_19465,N_19955);
or U20414 (N_20414,N_19789,N_19414);
nor U20415 (N_20415,N_19543,N_19508);
and U20416 (N_20416,N_19950,N_19642);
nand U20417 (N_20417,N_19808,N_19440);
and U20418 (N_20418,N_19529,N_19645);
or U20419 (N_20419,N_19692,N_19407);
nor U20420 (N_20420,N_19626,N_19407);
or U20421 (N_20421,N_19758,N_19629);
nand U20422 (N_20422,N_19552,N_19618);
nand U20423 (N_20423,N_19401,N_19594);
xor U20424 (N_20424,N_19491,N_19978);
or U20425 (N_20425,N_19622,N_19579);
xor U20426 (N_20426,N_19538,N_19890);
nand U20427 (N_20427,N_19957,N_19610);
nor U20428 (N_20428,N_19554,N_19832);
nor U20429 (N_20429,N_19964,N_19766);
or U20430 (N_20430,N_19660,N_19941);
nor U20431 (N_20431,N_19408,N_19386);
or U20432 (N_20432,N_19695,N_19725);
or U20433 (N_20433,N_19380,N_19427);
and U20434 (N_20434,N_19860,N_19919);
xnor U20435 (N_20435,N_19672,N_19546);
and U20436 (N_20436,N_19720,N_19635);
xor U20437 (N_20437,N_19707,N_19898);
nand U20438 (N_20438,N_19553,N_19925);
and U20439 (N_20439,N_19481,N_19384);
or U20440 (N_20440,N_19692,N_19845);
and U20441 (N_20441,N_19997,N_19650);
or U20442 (N_20442,N_19825,N_19693);
xor U20443 (N_20443,N_19636,N_19607);
nor U20444 (N_20444,N_19859,N_19615);
xnor U20445 (N_20445,N_19488,N_19811);
or U20446 (N_20446,N_19931,N_19405);
nor U20447 (N_20447,N_19531,N_19731);
and U20448 (N_20448,N_19782,N_19577);
nor U20449 (N_20449,N_19994,N_19538);
and U20450 (N_20450,N_19427,N_19544);
or U20451 (N_20451,N_19797,N_19851);
or U20452 (N_20452,N_19609,N_19675);
or U20453 (N_20453,N_19569,N_19606);
nand U20454 (N_20454,N_19450,N_19572);
nor U20455 (N_20455,N_19735,N_19489);
nor U20456 (N_20456,N_19551,N_19453);
xor U20457 (N_20457,N_19876,N_19606);
nand U20458 (N_20458,N_19728,N_19798);
or U20459 (N_20459,N_19974,N_19940);
or U20460 (N_20460,N_19760,N_19422);
nand U20461 (N_20461,N_19723,N_19735);
nand U20462 (N_20462,N_19590,N_19434);
xor U20463 (N_20463,N_19740,N_19810);
nor U20464 (N_20464,N_19476,N_19584);
or U20465 (N_20465,N_19866,N_19803);
nand U20466 (N_20466,N_19619,N_19841);
nor U20467 (N_20467,N_19708,N_19946);
nor U20468 (N_20468,N_19610,N_19968);
nor U20469 (N_20469,N_19928,N_19826);
or U20470 (N_20470,N_19688,N_19875);
xor U20471 (N_20471,N_19476,N_19605);
or U20472 (N_20472,N_19401,N_19417);
xnor U20473 (N_20473,N_19696,N_19551);
or U20474 (N_20474,N_19460,N_19539);
nor U20475 (N_20475,N_19682,N_19456);
and U20476 (N_20476,N_19946,N_19673);
and U20477 (N_20477,N_19711,N_19837);
nand U20478 (N_20478,N_19613,N_19435);
nor U20479 (N_20479,N_19553,N_19769);
or U20480 (N_20480,N_19650,N_19393);
or U20481 (N_20481,N_19825,N_19848);
xor U20482 (N_20482,N_19920,N_19534);
and U20483 (N_20483,N_19829,N_19742);
nor U20484 (N_20484,N_19420,N_19723);
or U20485 (N_20485,N_19706,N_19986);
nand U20486 (N_20486,N_19506,N_19520);
xnor U20487 (N_20487,N_19712,N_19476);
and U20488 (N_20488,N_19660,N_19868);
nand U20489 (N_20489,N_19795,N_19771);
or U20490 (N_20490,N_19982,N_19680);
nand U20491 (N_20491,N_19713,N_19843);
or U20492 (N_20492,N_19886,N_19718);
nand U20493 (N_20493,N_19481,N_19709);
or U20494 (N_20494,N_19607,N_19810);
and U20495 (N_20495,N_19447,N_19409);
nor U20496 (N_20496,N_19747,N_19582);
or U20497 (N_20497,N_19453,N_19414);
or U20498 (N_20498,N_19926,N_19438);
or U20499 (N_20499,N_19388,N_19720);
xnor U20500 (N_20500,N_19563,N_19746);
nor U20501 (N_20501,N_19513,N_19852);
nor U20502 (N_20502,N_19729,N_19643);
and U20503 (N_20503,N_19531,N_19689);
xnor U20504 (N_20504,N_19484,N_19546);
or U20505 (N_20505,N_19616,N_19627);
nor U20506 (N_20506,N_19410,N_19394);
xor U20507 (N_20507,N_19555,N_19465);
nor U20508 (N_20508,N_19400,N_19687);
and U20509 (N_20509,N_19469,N_19381);
and U20510 (N_20510,N_19560,N_19766);
xor U20511 (N_20511,N_19683,N_19900);
or U20512 (N_20512,N_19891,N_19791);
xnor U20513 (N_20513,N_19459,N_19888);
nor U20514 (N_20514,N_19536,N_19690);
nand U20515 (N_20515,N_19440,N_19591);
xnor U20516 (N_20516,N_19964,N_19436);
or U20517 (N_20517,N_19491,N_19891);
xor U20518 (N_20518,N_19907,N_19614);
xor U20519 (N_20519,N_19651,N_19956);
xor U20520 (N_20520,N_19794,N_19442);
and U20521 (N_20521,N_19394,N_19609);
nor U20522 (N_20522,N_19869,N_19682);
nor U20523 (N_20523,N_19845,N_19635);
and U20524 (N_20524,N_19649,N_19804);
nor U20525 (N_20525,N_19545,N_19849);
xnor U20526 (N_20526,N_19568,N_19480);
nor U20527 (N_20527,N_19947,N_19903);
and U20528 (N_20528,N_19381,N_19509);
and U20529 (N_20529,N_19728,N_19669);
xnor U20530 (N_20530,N_19613,N_19472);
nor U20531 (N_20531,N_19439,N_19996);
nand U20532 (N_20532,N_19764,N_19388);
xnor U20533 (N_20533,N_19843,N_19994);
xnor U20534 (N_20534,N_19672,N_19948);
nand U20535 (N_20535,N_19787,N_19418);
and U20536 (N_20536,N_19423,N_19878);
nor U20537 (N_20537,N_19820,N_19621);
or U20538 (N_20538,N_19758,N_19908);
nor U20539 (N_20539,N_19802,N_19931);
nand U20540 (N_20540,N_19760,N_19603);
nand U20541 (N_20541,N_19508,N_19737);
and U20542 (N_20542,N_19593,N_19420);
xnor U20543 (N_20543,N_19948,N_19902);
xor U20544 (N_20544,N_19633,N_19836);
or U20545 (N_20545,N_19981,N_19516);
and U20546 (N_20546,N_19869,N_19879);
or U20547 (N_20547,N_19758,N_19666);
and U20548 (N_20548,N_19434,N_19772);
or U20549 (N_20549,N_19724,N_19516);
nor U20550 (N_20550,N_19552,N_19443);
or U20551 (N_20551,N_19608,N_19510);
or U20552 (N_20552,N_19983,N_19616);
nand U20553 (N_20553,N_19899,N_19852);
or U20554 (N_20554,N_19895,N_19512);
nor U20555 (N_20555,N_19672,N_19645);
or U20556 (N_20556,N_19503,N_19859);
nand U20557 (N_20557,N_19522,N_19648);
or U20558 (N_20558,N_19999,N_19775);
nand U20559 (N_20559,N_19653,N_19655);
and U20560 (N_20560,N_19486,N_19466);
and U20561 (N_20561,N_19777,N_19378);
xnor U20562 (N_20562,N_19656,N_19774);
nor U20563 (N_20563,N_19757,N_19687);
and U20564 (N_20564,N_19986,N_19703);
xnor U20565 (N_20565,N_19380,N_19927);
xor U20566 (N_20566,N_19384,N_19879);
xnor U20567 (N_20567,N_19904,N_19508);
and U20568 (N_20568,N_19452,N_19837);
nand U20569 (N_20569,N_19955,N_19447);
or U20570 (N_20570,N_19889,N_19580);
or U20571 (N_20571,N_19799,N_19378);
and U20572 (N_20572,N_19972,N_19831);
or U20573 (N_20573,N_19433,N_19453);
nor U20574 (N_20574,N_19724,N_19570);
or U20575 (N_20575,N_19801,N_19850);
or U20576 (N_20576,N_19549,N_19632);
nor U20577 (N_20577,N_19798,N_19453);
nand U20578 (N_20578,N_19803,N_19440);
or U20579 (N_20579,N_19995,N_19410);
nand U20580 (N_20580,N_19989,N_19414);
nor U20581 (N_20581,N_19765,N_19408);
or U20582 (N_20582,N_19656,N_19949);
nand U20583 (N_20583,N_19706,N_19685);
nand U20584 (N_20584,N_19807,N_19684);
and U20585 (N_20585,N_19450,N_19885);
xnor U20586 (N_20586,N_19785,N_19777);
nor U20587 (N_20587,N_19889,N_19863);
and U20588 (N_20588,N_19496,N_19723);
or U20589 (N_20589,N_19625,N_19384);
and U20590 (N_20590,N_19897,N_19637);
nor U20591 (N_20591,N_19959,N_19652);
and U20592 (N_20592,N_19597,N_19751);
or U20593 (N_20593,N_19481,N_19395);
nor U20594 (N_20594,N_19539,N_19789);
xor U20595 (N_20595,N_19818,N_19534);
nor U20596 (N_20596,N_19698,N_19460);
and U20597 (N_20597,N_19480,N_19586);
and U20598 (N_20598,N_19684,N_19982);
nand U20599 (N_20599,N_19856,N_19668);
nand U20600 (N_20600,N_19697,N_19958);
or U20601 (N_20601,N_19744,N_19627);
and U20602 (N_20602,N_19778,N_19508);
nand U20603 (N_20603,N_19907,N_19866);
xnor U20604 (N_20604,N_19415,N_19412);
nand U20605 (N_20605,N_19523,N_19861);
and U20606 (N_20606,N_19909,N_19848);
xnor U20607 (N_20607,N_19724,N_19640);
nand U20608 (N_20608,N_19394,N_19517);
and U20609 (N_20609,N_19571,N_19655);
or U20610 (N_20610,N_19840,N_19902);
and U20611 (N_20611,N_19877,N_19644);
or U20612 (N_20612,N_19738,N_19953);
nor U20613 (N_20613,N_19852,N_19600);
or U20614 (N_20614,N_19631,N_19485);
and U20615 (N_20615,N_19380,N_19624);
nand U20616 (N_20616,N_19490,N_19674);
nor U20617 (N_20617,N_19733,N_19984);
or U20618 (N_20618,N_19379,N_19998);
or U20619 (N_20619,N_19798,N_19444);
and U20620 (N_20620,N_19802,N_19595);
xor U20621 (N_20621,N_19741,N_19863);
nand U20622 (N_20622,N_19503,N_19799);
nand U20623 (N_20623,N_19796,N_19519);
and U20624 (N_20624,N_19794,N_19980);
nand U20625 (N_20625,N_20081,N_20582);
or U20626 (N_20626,N_20165,N_20158);
and U20627 (N_20627,N_20012,N_20524);
or U20628 (N_20628,N_20440,N_20494);
nand U20629 (N_20629,N_20557,N_20079);
nor U20630 (N_20630,N_20003,N_20608);
or U20631 (N_20631,N_20229,N_20269);
xnor U20632 (N_20632,N_20225,N_20106);
nor U20633 (N_20633,N_20196,N_20025);
nor U20634 (N_20634,N_20323,N_20104);
nor U20635 (N_20635,N_20147,N_20171);
and U20636 (N_20636,N_20359,N_20004);
nand U20637 (N_20637,N_20318,N_20372);
nor U20638 (N_20638,N_20390,N_20342);
or U20639 (N_20639,N_20271,N_20449);
and U20640 (N_20640,N_20045,N_20437);
nand U20641 (N_20641,N_20534,N_20419);
and U20642 (N_20642,N_20255,N_20009);
or U20643 (N_20643,N_20547,N_20264);
or U20644 (N_20644,N_20388,N_20102);
or U20645 (N_20645,N_20083,N_20175);
nor U20646 (N_20646,N_20493,N_20191);
or U20647 (N_20647,N_20461,N_20065);
xnor U20648 (N_20648,N_20606,N_20377);
xnor U20649 (N_20649,N_20263,N_20221);
or U20650 (N_20650,N_20595,N_20412);
and U20651 (N_20651,N_20089,N_20035);
nand U20652 (N_20652,N_20140,N_20274);
and U20653 (N_20653,N_20513,N_20570);
xnor U20654 (N_20654,N_20261,N_20369);
nor U20655 (N_20655,N_20001,N_20093);
nor U20656 (N_20656,N_20098,N_20566);
nor U20657 (N_20657,N_20476,N_20549);
xor U20658 (N_20658,N_20074,N_20242);
nand U20659 (N_20659,N_20523,N_20135);
or U20660 (N_20660,N_20039,N_20022);
xor U20661 (N_20661,N_20542,N_20017);
nor U20662 (N_20662,N_20087,N_20061);
or U20663 (N_20663,N_20545,N_20115);
nor U20664 (N_20664,N_20238,N_20525);
xor U20665 (N_20665,N_20294,N_20601);
xnor U20666 (N_20666,N_20468,N_20210);
nand U20667 (N_20667,N_20163,N_20179);
nand U20668 (N_20668,N_20042,N_20550);
and U20669 (N_20669,N_20145,N_20485);
and U20670 (N_20670,N_20455,N_20162);
or U20671 (N_20671,N_20190,N_20603);
xnor U20672 (N_20672,N_20467,N_20330);
nand U20673 (N_20673,N_20075,N_20002);
nand U20674 (N_20674,N_20405,N_20030);
or U20675 (N_20675,N_20232,N_20054);
xor U20676 (N_20676,N_20077,N_20354);
xor U20677 (N_20677,N_20483,N_20118);
nand U20678 (N_20678,N_20548,N_20040);
nand U20679 (N_20679,N_20230,N_20464);
or U20680 (N_20680,N_20010,N_20267);
nor U20681 (N_20681,N_20346,N_20178);
nor U20682 (N_20682,N_20599,N_20117);
xnor U20683 (N_20683,N_20568,N_20151);
nand U20684 (N_20684,N_20362,N_20224);
nand U20685 (N_20685,N_20302,N_20306);
nor U20686 (N_20686,N_20182,N_20373);
xnor U20687 (N_20687,N_20382,N_20265);
and U20688 (N_20688,N_20516,N_20291);
xor U20689 (N_20689,N_20514,N_20421);
nor U20690 (N_20690,N_20028,N_20082);
xnor U20691 (N_20691,N_20212,N_20143);
or U20692 (N_20692,N_20452,N_20319);
nor U20693 (N_20693,N_20586,N_20157);
xor U20694 (N_20694,N_20048,N_20097);
nor U20695 (N_20695,N_20005,N_20403);
nand U20696 (N_20696,N_20609,N_20007);
and U20697 (N_20697,N_20283,N_20192);
and U20698 (N_20698,N_20357,N_20553);
and U20699 (N_20699,N_20019,N_20481);
nand U20700 (N_20700,N_20521,N_20059);
and U20701 (N_20701,N_20617,N_20571);
nor U20702 (N_20702,N_20398,N_20307);
nand U20703 (N_20703,N_20458,N_20141);
nand U20704 (N_20704,N_20374,N_20051);
nor U20705 (N_20705,N_20310,N_20465);
and U20706 (N_20706,N_20137,N_20590);
xor U20707 (N_20707,N_20000,N_20278);
or U20708 (N_20708,N_20084,N_20486);
xnor U20709 (N_20709,N_20327,N_20287);
nand U20710 (N_20710,N_20340,N_20088);
and U20711 (N_20711,N_20155,N_20574);
nand U20712 (N_20712,N_20298,N_20381);
nor U20713 (N_20713,N_20144,N_20047);
and U20714 (N_20714,N_20125,N_20069);
or U20715 (N_20715,N_20236,N_20320);
xnor U20716 (N_20716,N_20326,N_20462);
and U20717 (N_20717,N_20161,N_20413);
and U20718 (N_20718,N_20539,N_20506);
and U20719 (N_20719,N_20138,N_20100);
and U20720 (N_20720,N_20597,N_20253);
nand U20721 (N_20721,N_20598,N_20480);
and U20722 (N_20722,N_20428,N_20111);
nor U20723 (N_20723,N_20049,N_20376);
nand U20724 (N_20724,N_20173,N_20168);
nand U20725 (N_20725,N_20361,N_20197);
nand U20726 (N_20726,N_20488,N_20510);
xor U20727 (N_20727,N_20367,N_20114);
xor U20728 (N_20728,N_20492,N_20529);
nor U20729 (N_20729,N_20363,N_20136);
xor U20730 (N_20730,N_20573,N_20420);
and U20731 (N_20731,N_20406,N_20233);
nor U20732 (N_20732,N_20371,N_20551);
xor U20733 (N_20733,N_20418,N_20482);
xor U20734 (N_20734,N_20335,N_20073);
or U20735 (N_20735,N_20415,N_20579);
xnor U20736 (N_20736,N_20129,N_20497);
xor U20737 (N_20737,N_20613,N_20396);
nand U20738 (N_20738,N_20247,N_20299);
nand U20739 (N_20739,N_20459,N_20411);
nor U20740 (N_20740,N_20260,N_20495);
and U20741 (N_20741,N_20202,N_20123);
or U20742 (N_20742,N_20214,N_20066);
or U20743 (N_20743,N_20441,N_20543);
or U20744 (N_20744,N_20502,N_20394);
nor U20745 (N_20745,N_20471,N_20474);
xnor U20746 (N_20746,N_20531,N_20107);
nand U20747 (N_20747,N_20174,N_20316);
and U20748 (N_20748,N_20037,N_20344);
or U20749 (N_20749,N_20222,N_20275);
or U20750 (N_20750,N_20353,N_20209);
and U20751 (N_20751,N_20332,N_20023);
nor U20752 (N_20752,N_20305,N_20600);
xnor U20753 (N_20753,N_20577,N_20149);
and U20754 (N_20754,N_20569,N_20333);
xor U20755 (N_20755,N_20504,N_20228);
nor U20756 (N_20756,N_20400,N_20619);
nand U20757 (N_20757,N_20578,N_20554);
or U20758 (N_20758,N_20544,N_20248);
and U20759 (N_20759,N_20068,N_20234);
nor U20760 (N_20760,N_20142,N_20176);
xor U20761 (N_20761,N_20303,N_20257);
xnor U20762 (N_20762,N_20610,N_20169);
nand U20763 (N_20763,N_20477,N_20041);
nor U20764 (N_20764,N_20127,N_20385);
nor U20765 (N_20765,N_20245,N_20511);
nor U20766 (N_20766,N_20116,N_20220);
or U20767 (N_20767,N_20195,N_20226);
and U20768 (N_20768,N_20311,N_20383);
xnor U20769 (N_20769,N_20067,N_20063);
nor U20770 (N_20770,N_20526,N_20172);
nor U20771 (N_20771,N_20080,N_20094);
xor U20772 (N_20772,N_20499,N_20139);
nand U20773 (N_20773,N_20046,N_20512);
and U20774 (N_20774,N_20090,N_20515);
xnor U20775 (N_20775,N_20343,N_20113);
or U20776 (N_20776,N_20008,N_20108);
nand U20777 (N_20777,N_20487,N_20062);
nor U20778 (N_20778,N_20128,N_20223);
xor U20779 (N_20779,N_20297,N_20289);
or U20780 (N_20780,N_20414,N_20496);
xor U20781 (N_20781,N_20126,N_20038);
nor U20782 (N_20782,N_20285,N_20053);
and U20783 (N_20783,N_20375,N_20188);
nor U20784 (N_20784,N_20517,N_20624);
xor U20785 (N_20785,N_20313,N_20470);
nand U20786 (N_20786,N_20270,N_20575);
or U20787 (N_20787,N_20201,N_20044);
or U20788 (N_20788,N_20432,N_20286);
and U20789 (N_20789,N_20607,N_20200);
and U20790 (N_20790,N_20364,N_20594);
nand U20791 (N_20791,N_20021,N_20535);
xor U20792 (N_20792,N_20217,N_20015);
nor U20793 (N_20793,N_20519,N_20614);
xnor U20794 (N_20794,N_20295,N_20150);
and U20795 (N_20795,N_20266,N_20300);
or U20796 (N_20796,N_20556,N_20057);
xor U20797 (N_20797,N_20086,N_20427);
nand U20798 (N_20798,N_20448,N_20078);
nand U20799 (N_20799,N_20564,N_20541);
xnor U20800 (N_20800,N_20309,N_20589);
xnor U20801 (N_20801,N_20215,N_20130);
xor U20802 (N_20802,N_20058,N_20186);
or U20803 (N_20803,N_20424,N_20160);
nor U20804 (N_20804,N_20429,N_20532);
and U20805 (N_20805,N_20387,N_20254);
nand U20806 (N_20806,N_20076,N_20153);
xor U20807 (N_20807,N_20356,N_20416);
and U20808 (N_20808,N_20463,N_20407);
or U20809 (N_20809,N_20146,N_20583);
and U20810 (N_20810,N_20132,N_20218);
nand U20811 (N_20811,N_20325,N_20091);
nor U20812 (N_20812,N_20443,N_20050);
nor U20813 (N_20813,N_20378,N_20425);
xor U20814 (N_20814,N_20592,N_20092);
xnor U20815 (N_20815,N_20211,N_20436);
and U20816 (N_20816,N_20540,N_20337);
nor U20817 (N_20817,N_20011,N_20164);
or U20818 (N_20818,N_20249,N_20240);
or U20819 (N_20819,N_20239,N_20189);
and U20820 (N_20820,N_20446,N_20293);
or U20821 (N_20821,N_20386,N_20308);
nand U20822 (N_20822,N_20622,N_20351);
nand U20823 (N_20823,N_20006,N_20032);
and U20824 (N_20824,N_20304,N_20024);
nand U20825 (N_20825,N_20417,N_20321);
nor U20826 (N_20826,N_20454,N_20134);
nor U20827 (N_20827,N_20101,N_20029);
or U20828 (N_20828,N_20591,N_20281);
or U20829 (N_20829,N_20013,N_20623);
and U20830 (N_20830,N_20558,N_20280);
xnor U20831 (N_20831,N_20014,N_20241);
nor U20832 (N_20832,N_20208,N_20479);
xor U20833 (N_20833,N_20256,N_20433);
and U20834 (N_20834,N_20530,N_20020);
or U20835 (N_20835,N_20018,N_20434);
and U20836 (N_20836,N_20352,N_20404);
nand U20837 (N_20837,N_20576,N_20154);
and U20838 (N_20838,N_20565,N_20183);
nor U20839 (N_20839,N_20581,N_20027);
or U20840 (N_20840,N_20508,N_20537);
nand U20841 (N_20841,N_20314,N_20096);
nand U20842 (N_20842,N_20453,N_20099);
xor U20843 (N_20843,N_20505,N_20276);
nor U20844 (N_20844,N_20070,N_20445);
and U20845 (N_20845,N_20219,N_20469);
nand U20846 (N_20846,N_20166,N_20365);
or U20847 (N_20847,N_20052,N_20277);
or U20848 (N_20848,N_20207,N_20426);
and U20849 (N_20849,N_20472,N_20456);
nand U20850 (N_20850,N_20243,N_20447);
or U20851 (N_20851,N_20284,N_20442);
xor U20852 (N_20852,N_20338,N_20339);
nand U20853 (N_20853,N_20273,N_20334);
nand U20854 (N_20854,N_20290,N_20205);
nand U20855 (N_20855,N_20203,N_20272);
xor U20856 (N_20856,N_20397,N_20588);
nor U20857 (N_20857,N_20324,N_20509);
nand U20858 (N_20858,N_20252,N_20312);
nand U20859 (N_20859,N_20621,N_20408);
nand U20860 (N_20860,N_20016,N_20615);
xor U20861 (N_20861,N_20131,N_20602);
and U20862 (N_20862,N_20122,N_20555);
xor U20863 (N_20863,N_20246,N_20235);
and U20864 (N_20864,N_20187,N_20301);
nand U20865 (N_20865,N_20216,N_20444);
nor U20866 (N_20866,N_20064,N_20501);
or U20867 (N_20867,N_20536,N_20036);
or U20868 (N_20868,N_20349,N_20292);
or U20869 (N_20869,N_20237,N_20056);
nand U20870 (N_20870,N_20152,N_20500);
nor U20871 (N_20871,N_20604,N_20401);
or U20872 (N_20872,N_20395,N_20350);
nand U20873 (N_20873,N_20498,N_20559);
xor U20874 (N_20874,N_20194,N_20593);
nor U20875 (N_20875,N_20180,N_20331);
and U20876 (N_20876,N_20616,N_20206);
nor U20877 (N_20877,N_20296,N_20204);
nand U20878 (N_20878,N_20584,N_20409);
nor U20879 (N_20879,N_20288,N_20360);
nand U20880 (N_20880,N_20489,N_20193);
or U20881 (N_20881,N_20198,N_20244);
nand U20882 (N_20882,N_20055,N_20355);
nand U20883 (N_20883,N_20156,N_20105);
or U20884 (N_20884,N_20391,N_20358);
nor U20885 (N_20885,N_20345,N_20250);
nor U20886 (N_20886,N_20177,N_20181);
or U20887 (N_20887,N_20438,N_20562);
nor U20888 (N_20888,N_20620,N_20466);
nor U20889 (N_20889,N_20533,N_20384);
and U20890 (N_20890,N_20430,N_20560);
nor U20891 (N_20891,N_20612,N_20034);
and U20892 (N_20892,N_20347,N_20348);
and U20893 (N_20893,N_20518,N_20085);
xnor U20894 (N_20894,N_20328,N_20133);
or U20895 (N_20895,N_20341,N_20185);
xor U20896 (N_20896,N_20431,N_20507);
or U20897 (N_20897,N_20259,N_20460);
nand U20898 (N_20898,N_20563,N_20528);
nand U20899 (N_20899,N_20213,N_20370);
nand U20900 (N_20900,N_20435,N_20043);
nand U20901 (N_20901,N_20120,N_20439);
and U20902 (N_20902,N_20315,N_20184);
xor U20903 (N_20903,N_20605,N_20478);
or U20904 (N_20904,N_20410,N_20572);
nand U20905 (N_20905,N_20112,N_20121);
and U20906 (N_20906,N_20587,N_20329);
nand U20907 (N_20907,N_20268,N_20336);
and U20908 (N_20908,N_20317,N_20561);
or U20909 (N_20909,N_20033,N_20322);
or U20910 (N_20910,N_20148,N_20072);
nand U20911 (N_20911,N_20251,N_20473);
and U20912 (N_20912,N_20484,N_20124);
or U20913 (N_20913,N_20546,N_20393);
xor U20914 (N_20914,N_20368,N_20031);
nor U20915 (N_20915,N_20380,N_20392);
and U20916 (N_20916,N_20167,N_20450);
nand U20917 (N_20917,N_20503,N_20119);
and U20918 (N_20918,N_20399,N_20522);
or U20919 (N_20919,N_20282,N_20618);
and U20920 (N_20920,N_20258,N_20103);
nor U20921 (N_20921,N_20389,N_20231);
and U20922 (N_20922,N_20423,N_20071);
nand U20923 (N_20923,N_20611,N_20110);
and U20924 (N_20924,N_20199,N_20596);
nand U20925 (N_20925,N_20060,N_20527);
and U20926 (N_20926,N_20227,N_20475);
nor U20927 (N_20927,N_20451,N_20580);
nand U20928 (N_20928,N_20279,N_20490);
or U20929 (N_20929,N_20491,N_20170);
and U20930 (N_20930,N_20366,N_20567);
xnor U20931 (N_20931,N_20109,N_20402);
and U20932 (N_20932,N_20262,N_20538);
or U20933 (N_20933,N_20095,N_20026);
and U20934 (N_20934,N_20159,N_20552);
nor U20935 (N_20935,N_20585,N_20422);
xnor U20936 (N_20936,N_20457,N_20379);
and U20937 (N_20937,N_20520,N_20056);
nor U20938 (N_20938,N_20224,N_20333);
and U20939 (N_20939,N_20485,N_20016);
and U20940 (N_20940,N_20338,N_20153);
or U20941 (N_20941,N_20071,N_20104);
nand U20942 (N_20942,N_20003,N_20567);
or U20943 (N_20943,N_20442,N_20425);
or U20944 (N_20944,N_20584,N_20204);
and U20945 (N_20945,N_20064,N_20431);
nand U20946 (N_20946,N_20338,N_20196);
nor U20947 (N_20947,N_20624,N_20212);
nand U20948 (N_20948,N_20051,N_20368);
or U20949 (N_20949,N_20389,N_20136);
nand U20950 (N_20950,N_20264,N_20011);
nand U20951 (N_20951,N_20227,N_20363);
or U20952 (N_20952,N_20212,N_20352);
nor U20953 (N_20953,N_20359,N_20097);
xor U20954 (N_20954,N_20343,N_20203);
nor U20955 (N_20955,N_20593,N_20410);
nor U20956 (N_20956,N_20067,N_20292);
and U20957 (N_20957,N_20248,N_20435);
nor U20958 (N_20958,N_20285,N_20246);
nand U20959 (N_20959,N_20556,N_20120);
nor U20960 (N_20960,N_20276,N_20537);
xnor U20961 (N_20961,N_20516,N_20450);
nand U20962 (N_20962,N_20338,N_20618);
or U20963 (N_20963,N_20169,N_20186);
and U20964 (N_20964,N_20187,N_20527);
nand U20965 (N_20965,N_20604,N_20088);
and U20966 (N_20966,N_20495,N_20404);
nand U20967 (N_20967,N_20437,N_20041);
nor U20968 (N_20968,N_20438,N_20454);
xnor U20969 (N_20969,N_20540,N_20577);
nand U20970 (N_20970,N_20432,N_20153);
nand U20971 (N_20971,N_20181,N_20364);
or U20972 (N_20972,N_20067,N_20116);
nand U20973 (N_20973,N_20166,N_20616);
xnor U20974 (N_20974,N_20392,N_20296);
and U20975 (N_20975,N_20164,N_20530);
nand U20976 (N_20976,N_20399,N_20528);
nor U20977 (N_20977,N_20345,N_20461);
and U20978 (N_20978,N_20343,N_20450);
xnor U20979 (N_20979,N_20046,N_20293);
and U20980 (N_20980,N_20377,N_20268);
and U20981 (N_20981,N_20268,N_20391);
or U20982 (N_20982,N_20436,N_20127);
nand U20983 (N_20983,N_20379,N_20484);
or U20984 (N_20984,N_20446,N_20012);
and U20985 (N_20985,N_20078,N_20065);
and U20986 (N_20986,N_20552,N_20169);
nor U20987 (N_20987,N_20394,N_20169);
or U20988 (N_20988,N_20289,N_20614);
or U20989 (N_20989,N_20310,N_20021);
nor U20990 (N_20990,N_20011,N_20051);
nor U20991 (N_20991,N_20122,N_20231);
nor U20992 (N_20992,N_20293,N_20547);
nand U20993 (N_20993,N_20276,N_20277);
or U20994 (N_20994,N_20380,N_20397);
xnor U20995 (N_20995,N_20326,N_20167);
or U20996 (N_20996,N_20611,N_20536);
nor U20997 (N_20997,N_20239,N_20327);
nand U20998 (N_20998,N_20251,N_20495);
and U20999 (N_20999,N_20291,N_20247);
and U21000 (N_21000,N_20348,N_20152);
nand U21001 (N_21001,N_20143,N_20156);
xor U21002 (N_21002,N_20084,N_20589);
or U21003 (N_21003,N_20051,N_20136);
nand U21004 (N_21004,N_20444,N_20415);
nor U21005 (N_21005,N_20345,N_20268);
nand U21006 (N_21006,N_20061,N_20197);
nand U21007 (N_21007,N_20427,N_20191);
or U21008 (N_21008,N_20562,N_20044);
or U21009 (N_21009,N_20254,N_20557);
xnor U21010 (N_21010,N_20442,N_20250);
and U21011 (N_21011,N_20103,N_20480);
and U21012 (N_21012,N_20358,N_20011);
or U21013 (N_21013,N_20279,N_20030);
nor U21014 (N_21014,N_20580,N_20387);
xnor U21015 (N_21015,N_20351,N_20209);
and U21016 (N_21016,N_20596,N_20247);
and U21017 (N_21017,N_20185,N_20383);
xnor U21018 (N_21018,N_20447,N_20322);
nor U21019 (N_21019,N_20345,N_20429);
nand U21020 (N_21020,N_20073,N_20008);
or U21021 (N_21021,N_20445,N_20245);
or U21022 (N_21022,N_20343,N_20622);
xor U21023 (N_21023,N_20207,N_20456);
xnor U21024 (N_21024,N_20589,N_20545);
xnor U21025 (N_21025,N_20299,N_20507);
xor U21026 (N_21026,N_20001,N_20164);
nor U21027 (N_21027,N_20178,N_20319);
or U21028 (N_21028,N_20118,N_20247);
or U21029 (N_21029,N_20440,N_20155);
nand U21030 (N_21030,N_20044,N_20307);
nor U21031 (N_21031,N_20257,N_20522);
and U21032 (N_21032,N_20618,N_20343);
or U21033 (N_21033,N_20116,N_20575);
nor U21034 (N_21034,N_20492,N_20562);
nand U21035 (N_21035,N_20080,N_20123);
and U21036 (N_21036,N_20516,N_20622);
and U21037 (N_21037,N_20220,N_20048);
or U21038 (N_21038,N_20234,N_20442);
and U21039 (N_21039,N_20525,N_20126);
nand U21040 (N_21040,N_20607,N_20488);
nor U21041 (N_21041,N_20554,N_20337);
nand U21042 (N_21042,N_20346,N_20373);
nor U21043 (N_21043,N_20292,N_20090);
xnor U21044 (N_21044,N_20326,N_20215);
or U21045 (N_21045,N_20541,N_20027);
nor U21046 (N_21046,N_20289,N_20546);
or U21047 (N_21047,N_20443,N_20154);
xor U21048 (N_21048,N_20417,N_20270);
xor U21049 (N_21049,N_20449,N_20419);
nor U21050 (N_21050,N_20074,N_20091);
or U21051 (N_21051,N_20454,N_20124);
nor U21052 (N_21052,N_20244,N_20270);
nor U21053 (N_21053,N_20308,N_20184);
nand U21054 (N_21054,N_20382,N_20055);
or U21055 (N_21055,N_20256,N_20278);
or U21056 (N_21056,N_20557,N_20585);
nor U21057 (N_21057,N_20484,N_20032);
nor U21058 (N_21058,N_20421,N_20181);
nand U21059 (N_21059,N_20263,N_20438);
nand U21060 (N_21060,N_20526,N_20349);
nor U21061 (N_21061,N_20069,N_20425);
nand U21062 (N_21062,N_20409,N_20510);
and U21063 (N_21063,N_20116,N_20214);
xor U21064 (N_21064,N_20081,N_20215);
xnor U21065 (N_21065,N_20609,N_20610);
xor U21066 (N_21066,N_20052,N_20041);
xor U21067 (N_21067,N_20414,N_20211);
or U21068 (N_21068,N_20462,N_20612);
nand U21069 (N_21069,N_20397,N_20026);
nor U21070 (N_21070,N_20061,N_20475);
xnor U21071 (N_21071,N_20224,N_20264);
xor U21072 (N_21072,N_20321,N_20086);
xnor U21073 (N_21073,N_20446,N_20121);
or U21074 (N_21074,N_20256,N_20281);
xor U21075 (N_21075,N_20155,N_20339);
nand U21076 (N_21076,N_20213,N_20023);
or U21077 (N_21077,N_20480,N_20544);
and U21078 (N_21078,N_20111,N_20131);
or U21079 (N_21079,N_20092,N_20059);
and U21080 (N_21080,N_20005,N_20231);
or U21081 (N_21081,N_20031,N_20354);
or U21082 (N_21082,N_20252,N_20470);
xnor U21083 (N_21083,N_20036,N_20543);
nand U21084 (N_21084,N_20597,N_20567);
or U21085 (N_21085,N_20140,N_20603);
or U21086 (N_21086,N_20270,N_20526);
nor U21087 (N_21087,N_20444,N_20581);
and U21088 (N_21088,N_20274,N_20076);
and U21089 (N_21089,N_20007,N_20598);
nand U21090 (N_21090,N_20028,N_20570);
and U21091 (N_21091,N_20064,N_20414);
and U21092 (N_21092,N_20308,N_20568);
and U21093 (N_21093,N_20069,N_20414);
and U21094 (N_21094,N_20223,N_20506);
xnor U21095 (N_21095,N_20126,N_20353);
nor U21096 (N_21096,N_20344,N_20332);
xor U21097 (N_21097,N_20453,N_20498);
nor U21098 (N_21098,N_20581,N_20591);
xnor U21099 (N_21099,N_20450,N_20402);
xnor U21100 (N_21100,N_20044,N_20275);
nand U21101 (N_21101,N_20264,N_20157);
xor U21102 (N_21102,N_20181,N_20577);
or U21103 (N_21103,N_20259,N_20129);
xnor U21104 (N_21104,N_20033,N_20126);
or U21105 (N_21105,N_20452,N_20179);
and U21106 (N_21106,N_20402,N_20437);
nor U21107 (N_21107,N_20367,N_20535);
and U21108 (N_21108,N_20111,N_20110);
or U21109 (N_21109,N_20481,N_20113);
and U21110 (N_21110,N_20398,N_20489);
and U21111 (N_21111,N_20163,N_20241);
nor U21112 (N_21112,N_20540,N_20106);
and U21113 (N_21113,N_20468,N_20600);
xor U21114 (N_21114,N_20412,N_20081);
xor U21115 (N_21115,N_20209,N_20589);
nor U21116 (N_21116,N_20527,N_20382);
nand U21117 (N_21117,N_20456,N_20229);
and U21118 (N_21118,N_20084,N_20043);
nor U21119 (N_21119,N_20208,N_20495);
and U21120 (N_21120,N_20006,N_20113);
nand U21121 (N_21121,N_20465,N_20336);
and U21122 (N_21122,N_20608,N_20574);
and U21123 (N_21123,N_20409,N_20161);
nor U21124 (N_21124,N_20529,N_20197);
and U21125 (N_21125,N_20188,N_20119);
xor U21126 (N_21126,N_20307,N_20236);
nand U21127 (N_21127,N_20077,N_20441);
and U21128 (N_21128,N_20148,N_20206);
nand U21129 (N_21129,N_20078,N_20591);
nand U21130 (N_21130,N_20589,N_20360);
xnor U21131 (N_21131,N_20095,N_20324);
and U21132 (N_21132,N_20351,N_20190);
and U21133 (N_21133,N_20164,N_20424);
xor U21134 (N_21134,N_20275,N_20021);
nor U21135 (N_21135,N_20454,N_20392);
and U21136 (N_21136,N_20047,N_20464);
nand U21137 (N_21137,N_20583,N_20391);
and U21138 (N_21138,N_20019,N_20291);
and U21139 (N_21139,N_20521,N_20525);
nand U21140 (N_21140,N_20328,N_20149);
or U21141 (N_21141,N_20394,N_20035);
or U21142 (N_21142,N_20472,N_20337);
nor U21143 (N_21143,N_20055,N_20204);
and U21144 (N_21144,N_20007,N_20404);
xor U21145 (N_21145,N_20544,N_20426);
and U21146 (N_21146,N_20135,N_20603);
or U21147 (N_21147,N_20570,N_20521);
or U21148 (N_21148,N_20383,N_20496);
xnor U21149 (N_21149,N_20495,N_20585);
nor U21150 (N_21150,N_20543,N_20526);
or U21151 (N_21151,N_20043,N_20039);
nor U21152 (N_21152,N_20071,N_20357);
nor U21153 (N_21153,N_20241,N_20081);
or U21154 (N_21154,N_20218,N_20045);
nand U21155 (N_21155,N_20079,N_20090);
nor U21156 (N_21156,N_20495,N_20079);
nand U21157 (N_21157,N_20043,N_20258);
nor U21158 (N_21158,N_20112,N_20454);
and U21159 (N_21159,N_20392,N_20021);
xor U21160 (N_21160,N_20516,N_20474);
and U21161 (N_21161,N_20609,N_20378);
and U21162 (N_21162,N_20357,N_20401);
xnor U21163 (N_21163,N_20450,N_20119);
and U21164 (N_21164,N_20488,N_20490);
and U21165 (N_21165,N_20020,N_20109);
nand U21166 (N_21166,N_20591,N_20199);
and U21167 (N_21167,N_20519,N_20511);
or U21168 (N_21168,N_20444,N_20599);
nand U21169 (N_21169,N_20257,N_20362);
and U21170 (N_21170,N_20165,N_20148);
and U21171 (N_21171,N_20461,N_20609);
or U21172 (N_21172,N_20574,N_20353);
nor U21173 (N_21173,N_20095,N_20161);
and U21174 (N_21174,N_20466,N_20317);
or U21175 (N_21175,N_20318,N_20341);
nor U21176 (N_21176,N_20309,N_20301);
and U21177 (N_21177,N_20487,N_20477);
or U21178 (N_21178,N_20058,N_20374);
xor U21179 (N_21179,N_20021,N_20095);
or U21180 (N_21180,N_20409,N_20027);
xor U21181 (N_21181,N_20428,N_20159);
and U21182 (N_21182,N_20213,N_20071);
and U21183 (N_21183,N_20287,N_20464);
nand U21184 (N_21184,N_20069,N_20039);
or U21185 (N_21185,N_20430,N_20613);
nand U21186 (N_21186,N_20615,N_20198);
or U21187 (N_21187,N_20022,N_20609);
xor U21188 (N_21188,N_20039,N_20173);
nand U21189 (N_21189,N_20238,N_20577);
or U21190 (N_21190,N_20283,N_20563);
xnor U21191 (N_21191,N_20390,N_20160);
xor U21192 (N_21192,N_20294,N_20480);
nor U21193 (N_21193,N_20254,N_20379);
nand U21194 (N_21194,N_20600,N_20500);
and U21195 (N_21195,N_20385,N_20167);
or U21196 (N_21196,N_20491,N_20031);
nand U21197 (N_21197,N_20150,N_20029);
nor U21198 (N_21198,N_20337,N_20505);
xnor U21199 (N_21199,N_20187,N_20217);
nor U21200 (N_21200,N_20377,N_20231);
xor U21201 (N_21201,N_20453,N_20617);
or U21202 (N_21202,N_20324,N_20455);
and U21203 (N_21203,N_20412,N_20002);
or U21204 (N_21204,N_20336,N_20243);
or U21205 (N_21205,N_20292,N_20145);
xnor U21206 (N_21206,N_20063,N_20617);
nor U21207 (N_21207,N_20000,N_20486);
or U21208 (N_21208,N_20329,N_20023);
nor U21209 (N_21209,N_20570,N_20335);
nor U21210 (N_21210,N_20204,N_20339);
nor U21211 (N_21211,N_20446,N_20353);
xor U21212 (N_21212,N_20180,N_20376);
or U21213 (N_21213,N_20133,N_20283);
nor U21214 (N_21214,N_20264,N_20569);
nor U21215 (N_21215,N_20077,N_20027);
nand U21216 (N_21216,N_20060,N_20613);
nor U21217 (N_21217,N_20002,N_20247);
xor U21218 (N_21218,N_20021,N_20505);
nand U21219 (N_21219,N_20134,N_20071);
nor U21220 (N_21220,N_20147,N_20314);
and U21221 (N_21221,N_20508,N_20404);
or U21222 (N_21222,N_20019,N_20506);
or U21223 (N_21223,N_20043,N_20013);
xor U21224 (N_21224,N_20331,N_20496);
xnor U21225 (N_21225,N_20594,N_20173);
nand U21226 (N_21226,N_20367,N_20458);
and U21227 (N_21227,N_20262,N_20467);
nand U21228 (N_21228,N_20548,N_20456);
nand U21229 (N_21229,N_20332,N_20276);
xor U21230 (N_21230,N_20275,N_20013);
and U21231 (N_21231,N_20503,N_20397);
nand U21232 (N_21232,N_20155,N_20531);
or U21233 (N_21233,N_20226,N_20163);
xor U21234 (N_21234,N_20457,N_20299);
and U21235 (N_21235,N_20601,N_20466);
nor U21236 (N_21236,N_20564,N_20602);
nand U21237 (N_21237,N_20551,N_20539);
nand U21238 (N_21238,N_20370,N_20313);
nand U21239 (N_21239,N_20318,N_20087);
or U21240 (N_21240,N_20267,N_20565);
nand U21241 (N_21241,N_20173,N_20599);
xnor U21242 (N_21242,N_20291,N_20515);
nand U21243 (N_21243,N_20023,N_20323);
and U21244 (N_21244,N_20500,N_20331);
nand U21245 (N_21245,N_20564,N_20061);
xnor U21246 (N_21246,N_20270,N_20160);
xor U21247 (N_21247,N_20565,N_20453);
nor U21248 (N_21248,N_20372,N_20058);
or U21249 (N_21249,N_20404,N_20428);
nor U21250 (N_21250,N_20696,N_21167);
or U21251 (N_21251,N_21232,N_20749);
xor U21252 (N_21252,N_21009,N_20771);
xor U21253 (N_21253,N_20675,N_21213);
nor U21254 (N_21254,N_20763,N_21031);
nor U21255 (N_21255,N_20667,N_20787);
xnor U21256 (N_21256,N_20789,N_21155);
or U21257 (N_21257,N_21141,N_21112);
nor U21258 (N_21258,N_21061,N_21073);
or U21259 (N_21259,N_20945,N_20698);
and U21260 (N_21260,N_20692,N_20855);
xor U21261 (N_21261,N_20985,N_20765);
or U21262 (N_21262,N_20753,N_20902);
xor U21263 (N_21263,N_20846,N_20861);
and U21264 (N_21264,N_20877,N_21018);
or U21265 (N_21265,N_20971,N_20874);
nand U21266 (N_21266,N_21199,N_20786);
xnor U21267 (N_21267,N_20873,N_21211);
nand U21268 (N_21268,N_21166,N_21131);
nand U21269 (N_21269,N_20734,N_20654);
nand U21270 (N_21270,N_20638,N_21045);
and U21271 (N_21271,N_21138,N_20705);
nand U21272 (N_21272,N_20837,N_20688);
xnor U21273 (N_21273,N_21176,N_21072);
xnor U21274 (N_21274,N_20921,N_20648);
and U21275 (N_21275,N_20870,N_21204);
nand U21276 (N_21276,N_20904,N_21066);
nand U21277 (N_21277,N_21084,N_20981);
and U21278 (N_21278,N_21212,N_20661);
nand U21279 (N_21279,N_20947,N_20650);
and U21280 (N_21280,N_21020,N_20948);
xor U21281 (N_21281,N_20956,N_20750);
nand U21282 (N_21282,N_21107,N_21001);
nor U21283 (N_21283,N_20911,N_20668);
xor U21284 (N_21284,N_20881,N_21185);
nand U21285 (N_21285,N_20728,N_20726);
nand U21286 (N_21286,N_21148,N_20989);
and U21287 (N_21287,N_20838,N_21218);
and U21288 (N_21288,N_21115,N_21075);
xnor U21289 (N_21289,N_20813,N_20653);
or U21290 (N_21290,N_20941,N_21026);
and U21291 (N_21291,N_21109,N_20931);
nor U21292 (N_21292,N_20903,N_21024);
nand U21293 (N_21293,N_20759,N_21043);
xor U21294 (N_21294,N_20633,N_20715);
nand U21295 (N_21295,N_20818,N_20984);
xor U21296 (N_21296,N_20965,N_21229);
xor U21297 (N_21297,N_20707,N_21231);
or U21298 (N_21298,N_20792,N_20731);
nand U21299 (N_21299,N_20997,N_20736);
and U21300 (N_21300,N_20784,N_20852);
nand U21301 (N_21301,N_21165,N_20991);
or U21302 (N_21302,N_20729,N_20889);
nand U21303 (N_21303,N_20915,N_20793);
or U21304 (N_21304,N_20848,N_20927);
and U21305 (N_21305,N_21140,N_20906);
and U21306 (N_21306,N_21007,N_21145);
nand U21307 (N_21307,N_20737,N_20944);
or U21308 (N_21308,N_20907,N_21106);
or U21309 (N_21309,N_20741,N_21198);
nor U21310 (N_21310,N_21130,N_20917);
and U21311 (N_21311,N_21224,N_21022);
nor U21312 (N_21312,N_21119,N_20842);
nand U21313 (N_21313,N_20628,N_20883);
nand U21314 (N_21314,N_20804,N_21027);
nor U21315 (N_21315,N_20890,N_20836);
or U21316 (N_21316,N_20651,N_21210);
nor U21317 (N_21317,N_21159,N_21032);
nand U21318 (N_21318,N_21048,N_20722);
xnor U21319 (N_21319,N_21002,N_20809);
and U21320 (N_21320,N_21144,N_20871);
nor U21321 (N_21321,N_21175,N_21226);
xnor U21322 (N_21322,N_20924,N_21036);
xnor U21323 (N_21323,N_20719,N_21097);
nor U21324 (N_21324,N_21042,N_21056);
nor U21325 (N_21325,N_21046,N_21080);
nand U21326 (N_21326,N_20913,N_20885);
nand U21327 (N_21327,N_20992,N_20761);
nor U21328 (N_21328,N_20769,N_20808);
xnor U21329 (N_21329,N_20978,N_20934);
nand U21330 (N_21330,N_20817,N_20957);
nor U21331 (N_21331,N_20631,N_20754);
and U21332 (N_21332,N_20766,N_21063);
nand U21333 (N_21333,N_20994,N_21225);
and U21334 (N_21334,N_21011,N_21192);
xor U21335 (N_21335,N_20673,N_20926);
xnor U21336 (N_21336,N_20954,N_20745);
xor U21337 (N_21337,N_21152,N_21227);
and U21338 (N_21338,N_21237,N_20702);
or U21339 (N_21339,N_20703,N_20647);
nor U21340 (N_21340,N_20798,N_20788);
nand U21341 (N_21341,N_21008,N_20950);
and U21342 (N_21342,N_21221,N_20995);
or U21343 (N_21343,N_20790,N_20644);
nor U21344 (N_21344,N_20880,N_20901);
and U21345 (N_21345,N_20865,N_20691);
and U21346 (N_21346,N_20812,N_20683);
nor U21347 (N_21347,N_21244,N_20767);
xnor U21348 (N_21348,N_20685,N_21086);
and U21349 (N_21349,N_20679,N_20845);
nand U21350 (N_21350,N_20660,N_21096);
or U21351 (N_21351,N_21074,N_20762);
and U21352 (N_21352,N_21209,N_21100);
nand U21353 (N_21353,N_20659,N_21053);
and U21354 (N_21354,N_20843,N_21059);
and U21355 (N_21355,N_21214,N_21190);
and U21356 (N_21356,N_21015,N_21247);
nand U21357 (N_21357,N_20723,N_21050);
xor U21358 (N_21358,N_21196,N_20864);
and U21359 (N_21359,N_21098,N_20645);
nand U21360 (N_21360,N_21241,N_21120);
nand U21361 (N_21361,N_20962,N_20856);
nor U21362 (N_21362,N_21052,N_20878);
xor U21363 (N_21363,N_21088,N_20840);
and U21364 (N_21364,N_20979,N_20772);
nor U21365 (N_21365,N_21133,N_20834);
xnor U21366 (N_21366,N_20936,N_20896);
and U21367 (N_21367,N_20872,N_20646);
nand U21368 (N_21368,N_21157,N_21041);
xor U21369 (N_21369,N_20875,N_21184);
or U21370 (N_21370,N_20893,N_20632);
nand U21371 (N_21371,N_20806,N_20847);
or U21372 (N_21372,N_21201,N_20967);
or U21373 (N_21373,N_21170,N_21171);
nand U21374 (N_21374,N_21189,N_21186);
and U21375 (N_21375,N_21076,N_20676);
xor U21376 (N_21376,N_20977,N_21105);
and U21377 (N_21377,N_20693,N_21220);
nand U21378 (N_21378,N_20814,N_20942);
xor U21379 (N_21379,N_21038,N_20751);
or U21380 (N_21380,N_20748,N_20860);
and U21381 (N_21381,N_20828,N_21067);
nand U21382 (N_21382,N_21014,N_20839);
xnor U21383 (N_21383,N_20643,N_21242);
and U21384 (N_21384,N_20727,N_21125);
xnor U21385 (N_21385,N_20833,N_21243);
xnor U21386 (N_21386,N_21239,N_20935);
or U21387 (N_21387,N_21205,N_20908);
or U21388 (N_21388,N_20876,N_21113);
nand U21389 (N_21389,N_21068,N_20958);
nand U21390 (N_21390,N_20756,N_20800);
nand U21391 (N_21391,N_21249,N_20898);
nand U21392 (N_21392,N_21108,N_21207);
or U21393 (N_21393,N_21081,N_21089);
xnor U21394 (N_21394,N_20884,N_21163);
and U21395 (N_21395,N_20768,N_21082);
nor U21396 (N_21396,N_20758,N_20862);
or U21397 (N_21397,N_21087,N_20998);
nor U21398 (N_21398,N_20746,N_21195);
nand U21399 (N_21399,N_21090,N_21182);
and U21400 (N_21400,N_20656,N_21012);
and U21401 (N_21401,N_20625,N_20662);
or U21402 (N_21402,N_20850,N_20949);
and U21403 (N_21403,N_21039,N_21058);
nand U21404 (N_21404,N_21228,N_21156);
nor U21405 (N_21405,N_21065,N_21179);
xnor U21406 (N_21406,N_20811,N_20700);
nor U21407 (N_21407,N_20914,N_20791);
nand U21408 (N_21408,N_20980,N_21215);
nor U21409 (N_21409,N_20822,N_20894);
and U21410 (N_21410,N_20779,N_21094);
and U21411 (N_21411,N_20827,N_21197);
nor U21412 (N_21412,N_20663,N_21092);
or U21413 (N_21413,N_21030,N_21017);
xnor U21414 (N_21414,N_20757,N_20922);
and U21415 (N_21415,N_21055,N_21217);
nand U21416 (N_21416,N_20710,N_21203);
or U21417 (N_21417,N_21169,N_20940);
and U21418 (N_21418,N_21099,N_20887);
and U21419 (N_21419,N_20802,N_21177);
nor U21420 (N_21420,N_20853,N_21235);
or U21421 (N_21421,N_21037,N_20639);
nand U21422 (N_21422,N_20807,N_20706);
and U21423 (N_21423,N_20717,N_20669);
nand U21424 (N_21424,N_21135,N_21150);
or U21425 (N_21425,N_20970,N_21000);
and U21426 (N_21426,N_21127,N_20912);
nor U21427 (N_21427,N_20774,N_20641);
and U21428 (N_21428,N_21238,N_20963);
xor U21429 (N_21429,N_21188,N_20972);
nor U21430 (N_21430,N_21174,N_20973);
nand U21431 (N_21431,N_21153,N_21194);
or U21432 (N_21432,N_20816,N_20670);
and U21433 (N_21433,N_20744,N_20740);
or U21434 (N_21434,N_21161,N_21062);
nand U21435 (N_21435,N_20704,N_20642);
or U21436 (N_21436,N_21114,N_20821);
nor U21437 (N_21437,N_20687,N_20959);
nor U21438 (N_21438,N_20724,N_20975);
nand U21439 (N_21439,N_20730,N_20781);
nand U21440 (N_21440,N_21180,N_21248);
xor U21441 (N_21441,N_21139,N_20951);
nor U21442 (N_21442,N_21246,N_20841);
and U21443 (N_21443,N_20866,N_21233);
xnor U21444 (N_21444,N_20735,N_20932);
xor U21445 (N_21445,N_20969,N_21040);
nand U21446 (N_21446,N_20869,N_20863);
xor U21447 (N_21447,N_21121,N_20891);
nor U21448 (N_21448,N_20799,N_21208);
nand U21449 (N_21449,N_20929,N_20755);
and U21450 (N_21450,N_20649,N_20826);
or U21451 (N_21451,N_20943,N_20630);
and U21452 (N_21452,N_20764,N_20854);
and U21453 (N_21453,N_21234,N_20844);
nand U21454 (N_21454,N_20794,N_20918);
nand U21455 (N_21455,N_20627,N_20776);
and U21456 (N_21456,N_20916,N_20681);
or U21457 (N_21457,N_21178,N_21054);
nor U21458 (N_21458,N_21023,N_20976);
nor U21459 (N_21459,N_20686,N_21151);
nand U21460 (N_21460,N_21060,N_20933);
xor U21461 (N_21461,N_20635,N_20709);
nor U21462 (N_21462,N_20797,N_20993);
or U21463 (N_21463,N_20785,N_21206);
and U21464 (N_21464,N_20778,N_21168);
or U21465 (N_21465,N_20953,N_21028);
nor U21466 (N_21466,N_20652,N_20968);
and U21467 (N_21467,N_20900,N_20640);
and U21468 (N_21468,N_20832,N_21044);
xor U21469 (N_21469,N_21004,N_20859);
xor U21470 (N_21470,N_21191,N_20657);
xnor U21471 (N_21471,N_21101,N_20895);
xnor U21472 (N_21472,N_20671,N_21025);
or U21473 (N_21473,N_21116,N_20720);
nor U21474 (N_21474,N_21181,N_20829);
xor U21475 (N_21475,N_20666,N_21079);
nor U21476 (N_21476,N_21033,N_20830);
and U21477 (N_21477,N_20892,N_20928);
nand U21478 (N_21478,N_20946,N_20930);
nand U21479 (N_21479,N_20796,N_21019);
and U21480 (N_21480,N_20801,N_20634);
xor U21481 (N_21481,N_21047,N_20674);
and U21482 (N_21482,N_21071,N_21077);
and U21483 (N_21483,N_20909,N_21240);
nor U21484 (N_21484,N_21117,N_21158);
nand U21485 (N_21485,N_21110,N_21219);
nand U21486 (N_21486,N_20825,N_20867);
xor U21487 (N_21487,N_21149,N_20780);
or U21488 (N_21488,N_20713,N_21070);
xor U21489 (N_21489,N_21223,N_21069);
nand U21490 (N_21490,N_20990,N_20711);
nand U21491 (N_21491,N_21078,N_21049);
xor U21492 (N_21492,N_21132,N_20868);
or U21493 (N_21493,N_20820,N_20725);
nand U21494 (N_21494,N_20626,N_21006);
nor U21495 (N_21495,N_20637,N_21187);
xor U21496 (N_21496,N_20986,N_20742);
or U21497 (N_21497,N_20775,N_20964);
nor U21498 (N_21498,N_21029,N_20680);
and U21499 (N_21499,N_20712,N_21083);
and U21500 (N_21500,N_21154,N_20857);
nand U21501 (N_21501,N_21051,N_20732);
nor U21502 (N_21502,N_20783,N_20694);
nor U21503 (N_21503,N_20960,N_21147);
nor U21504 (N_21504,N_20849,N_20770);
nand U21505 (N_21505,N_20721,N_21003);
or U21506 (N_21506,N_21216,N_20655);
or U21507 (N_21507,N_21111,N_20923);
nor U21508 (N_21508,N_20695,N_20733);
nand U21509 (N_21509,N_21162,N_20805);
nor U21510 (N_21510,N_20803,N_20678);
and U21511 (N_21511,N_21021,N_20701);
xor U21512 (N_21512,N_21142,N_21146);
and U21513 (N_21513,N_20810,N_20777);
and U21514 (N_21514,N_21123,N_20629);
nand U21515 (N_21515,N_20747,N_20714);
nand U21516 (N_21516,N_20658,N_20858);
or U21517 (N_21517,N_20684,N_20952);
and U21518 (N_21518,N_20987,N_21236);
or U21519 (N_21519,N_20782,N_21143);
nor U21520 (N_21520,N_21136,N_20925);
and U21521 (N_21521,N_20988,N_20835);
and U21522 (N_21522,N_20831,N_20955);
nor U21523 (N_21523,N_21137,N_20899);
nand U21524 (N_21524,N_21085,N_21222);
xnor U21525 (N_21525,N_20682,N_20708);
or U21526 (N_21526,N_20824,N_20919);
nor U21527 (N_21527,N_20819,N_20851);
nand U21528 (N_21528,N_20743,N_21164);
nor U21529 (N_21529,N_21129,N_20672);
nand U21530 (N_21530,N_21193,N_20738);
or U21531 (N_21531,N_21103,N_20636);
nand U21532 (N_21532,N_21124,N_20938);
and U21533 (N_21533,N_21005,N_21064);
and U21534 (N_21534,N_21035,N_21172);
and U21535 (N_21535,N_20773,N_20982);
and U21536 (N_21536,N_20974,N_21183);
nor U21537 (N_21537,N_20665,N_21128);
nor U21538 (N_21538,N_20689,N_20739);
or U21539 (N_21539,N_21200,N_20718);
nor U21540 (N_21540,N_21122,N_21013);
and U21541 (N_21541,N_20690,N_20996);
nand U21542 (N_21542,N_20882,N_20664);
or U21543 (N_21543,N_20716,N_20677);
or U21544 (N_21544,N_21010,N_20897);
nand U21545 (N_21545,N_21095,N_20966);
xnor U21546 (N_21546,N_20937,N_20910);
nor U21547 (N_21547,N_21245,N_21202);
nor U21548 (N_21548,N_21134,N_20961);
or U21549 (N_21549,N_21091,N_20697);
xnor U21550 (N_21550,N_21016,N_21034);
and U21551 (N_21551,N_20699,N_21230);
and U21552 (N_21552,N_20983,N_20905);
nand U21553 (N_21553,N_20920,N_21102);
nand U21554 (N_21554,N_20795,N_21118);
xnor U21555 (N_21555,N_20815,N_20760);
nand U21556 (N_21556,N_21057,N_20752);
xor U21557 (N_21557,N_21093,N_20823);
xor U21558 (N_21558,N_20888,N_20939);
xnor U21559 (N_21559,N_21104,N_21160);
and U21560 (N_21560,N_21126,N_21173);
or U21561 (N_21561,N_20879,N_20999);
or U21562 (N_21562,N_20886,N_20965);
nor U21563 (N_21563,N_21152,N_20848);
or U21564 (N_21564,N_21244,N_21177);
or U21565 (N_21565,N_20763,N_20859);
or U21566 (N_21566,N_21130,N_21143);
or U21567 (N_21567,N_21110,N_20808);
nand U21568 (N_21568,N_21205,N_21135);
xnor U21569 (N_21569,N_20944,N_20793);
and U21570 (N_21570,N_20913,N_20859);
and U21571 (N_21571,N_21048,N_20893);
and U21572 (N_21572,N_20772,N_21056);
nand U21573 (N_21573,N_21042,N_20888);
xor U21574 (N_21574,N_20670,N_21095);
nand U21575 (N_21575,N_20766,N_21218);
or U21576 (N_21576,N_21167,N_21067);
or U21577 (N_21577,N_20937,N_20789);
and U21578 (N_21578,N_20849,N_20884);
nor U21579 (N_21579,N_20689,N_20650);
nand U21580 (N_21580,N_21153,N_20831);
nor U21581 (N_21581,N_20831,N_20779);
xnor U21582 (N_21582,N_20709,N_20751);
nor U21583 (N_21583,N_20845,N_21109);
nand U21584 (N_21584,N_20694,N_21007);
xnor U21585 (N_21585,N_21039,N_21035);
xor U21586 (N_21586,N_21191,N_20679);
or U21587 (N_21587,N_20801,N_20626);
nand U21588 (N_21588,N_21049,N_20673);
nand U21589 (N_21589,N_20678,N_20750);
and U21590 (N_21590,N_21098,N_21002);
nand U21591 (N_21591,N_20861,N_20800);
or U21592 (N_21592,N_20682,N_20967);
or U21593 (N_21593,N_21038,N_20665);
or U21594 (N_21594,N_21092,N_21065);
and U21595 (N_21595,N_20974,N_21123);
xnor U21596 (N_21596,N_21162,N_21121);
nand U21597 (N_21597,N_20847,N_21208);
nand U21598 (N_21598,N_20633,N_21037);
and U21599 (N_21599,N_20857,N_20814);
or U21600 (N_21600,N_20729,N_21184);
nand U21601 (N_21601,N_20803,N_20789);
or U21602 (N_21602,N_21124,N_20982);
xor U21603 (N_21603,N_21101,N_20637);
xnor U21604 (N_21604,N_21072,N_21070);
and U21605 (N_21605,N_20837,N_21074);
and U21606 (N_21606,N_20830,N_20878);
and U21607 (N_21607,N_21239,N_21234);
nor U21608 (N_21608,N_20927,N_21036);
xnor U21609 (N_21609,N_20685,N_20763);
xnor U21610 (N_21610,N_20774,N_20824);
and U21611 (N_21611,N_20858,N_20809);
and U21612 (N_21612,N_20773,N_20660);
xnor U21613 (N_21613,N_21179,N_20797);
xor U21614 (N_21614,N_20686,N_20934);
nor U21615 (N_21615,N_20717,N_21120);
and U21616 (N_21616,N_21023,N_20907);
xnor U21617 (N_21617,N_20730,N_20926);
and U21618 (N_21618,N_20760,N_20992);
nand U21619 (N_21619,N_21024,N_20634);
and U21620 (N_21620,N_20877,N_20892);
nor U21621 (N_21621,N_21193,N_21238);
nand U21622 (N_21622,N_21063,N_20680);
nand U21623 (N_21623,N_20859,N_20981);
or U21624 (N_21624,N_21090,N_20999);
xor U21625 (N_21625,N_21155,N_20740);
nor U21626 (N_21626,N_20967,N_21101);
or U21627 (N_21627,N_20884,N_20992);
or U21628 (N_21628,N_21087,N_21181);
nand U21629 (N_21629,N_21104,N_20775);
and U21630 (N_21630,N_21040,N_21168);
nand U21631 (N_21631,N_21111,N_21050);
xor U21632 (N_21632,N_21228,N_20929);
and U21633 (N_21633,N_20908,N_20709);
and U21634 (N_21634,N_21122,N_21019);
xor U21635 (N_21635,N_20918,N_20713);
and U21636 (N_21636,N_21098,N_21182);
xor U21637 (N_21637,N_21235,N_21145);
or U21638 (N_21638,N_21045,N_21129);
nand U21639 (N_21639,N_20781,N_20740);
nor U21640 (N_21640,N_20759,N_20756);
nand U21641 (N_21641,N_20873,N_21027);
nor U21642 (N_21642,N_21006,N_20778);
and U21643 (N_21643,N_20751,N_21021);
or U21644 (N_21644,N_20737,N_20963);
or U21645 (N_21645,N_21088,N_20852);
or U21646 (N_21646,N_20944,N_21198);
xor U21647 (N_21647,N_21117,N_20912);
xnor U21648 (N_21648,N_20793,N_21077);
nand U21649 (N_21649,N_20732,N_20945);
or U21650 (N_21650,N_21057,N_20751);
and U21651 (N_21651,N_21218,N_21138);
xor U21652 (N_21652,N_21172,N_21135);
and U21653 (N_21653,N_21061,N_20979);
and U21654 (N_21654,N_21246,N_20784);
nand U21655 (N_21655,N_21017,N_20824);
nor U21656 (N_21656,N_20682,N_20917);
nand U21657 (N_21657,N_20874,N_20842);
nand U21658 (N_21658,N_20687,N_20857);
xor U21659 (N_21659,N_20689,N_20918);
xor U21660 (N_21660,N_21176,N_20854);
xor U21661 (N_21661,N_21094,N_20698);
nand U21662 (N_21662,N_20861,N_21123);
nor U21663 (N_21663,N_20795,N_20919);
nor U21664 (N_21664,N_20687,N_20751);
nor U21665 (N_21665,N_20754,N_20681);
nand U21666 (N_21666,N_20828,N_21217);
nor U21667 (N_21667,N_20953,N_20783);
nand U21668 (N_21668,N_20825,N_21083);
or U21669 (N_21669,N_20901,N_20811);
and U21670 (N_21670,N_20952,N_20773);
nor U21671 (N_21671,N_21155,N_21112);
and U21672 (N_21672,N_21119,N_21151);
nor U21673 (N_21673,N_21002,N_21069);
nor U21674 (N_21674,N_20957,N_21074);
nor U21675 (N_21675,N_20921,N_21051);
nor U21676 (N_21676,N_20929,N_20660);
xor U21677 (N_21677,N_20875,N_20775);
or U21678 (N_21678,N_20956,N_20865);
xor U21679 (N_21679,N_20875,N_20703);
nor U21680 (N_21680,N_20661,N_21218);
nor U21681 (N_21681,N_20803,N_21124);
or U21682 (N_21682,N_20667,N_20653);
nor U21683 (N_21683,N_20881,N_20777);
and U21684 (N_21684,N_20628,N_20912);
xor U21685 (N_21685,N_20909,N_21067);
nand U21686 (N_21686,N_20753,N_21084);
nand U21687 (N_21687,N_20638,N_21114);
xnor U21688 (N_21688,N_21068,N_20922);
nand U21689 (N_21689,N_20715,N_21026);
or U21690 (N_21690,N_20692,N_21220);
xor U21691 (N_21691,N_21094,N_21208);
xnor U21692 (N_21692,N_20864,N_21074);
or U21693 (N_21693,N_20805,N_21122);
nand U21694 (N_21694,N_21089,N_20739);
or U21695 (N_21695,N_21124,N_20880);
nor U21696 (N_21696,N_21005,N_21075);
and U21697 (N_21697,N_20779,N_21038);
and U21698 (N_21698,N_20800,N_20819);
and U21699 (N_21699,N_20820,N_21188);
nor U21700 (N_21700,N_21133,N_20677);
nand U21701 (N_21701,N_20687,N_20916);
xnor U21702 (N_21702,N_21062,N_21198);
nand U21703 (N_21703,N_20652,N_21102);
xor U21704 (N_21704,N_21073,N_21211);
xnor U21705 (N_21705,N_21188,N_21097);
or U21706 (N_21706,N_21045,N_20908);
or U21707 (N_21707,N_21228,N_20790);
nand U21708 (N_21708,N_21181,N_20885);
nand U21709 (N_21709,N_21128,N_20709);
nand U21710 (N_21710,N_20800,N_20823);
and U21711 (N_21711,N_21221,N_20707);
and U21712 (N_21712,N_20834,N_20690);
nor U21713 (N_21713,N_21241,N_21087);
and U21714 (N_21714,N_21177,N_21103);
and U21715 (N_21715,N_20867,N_20841);
xor U21716 (N_21716,N_21115,N_20676);
nand U21717 (N_21717,N_20833,N_21082);
nor U21718 (N_21718,N_20875,N_20867);
or U21719 (N_21719,N_20739,N_20632);
nand U21720 (N_21720,N_21148,N_20869);
or U21721 (N_21721,N_21168,N_20655);
nand U21722 (N_21722,N_20886,N_20857);
or U21723 (N_21723,N_20984,N_20932);
xnor U21724 (N_21724,N_20867,N_20805);
xnor U21725 (N_21725,N_21103,N_21116);
xor U21726 (N_21726,N_21188,N_21157);
xor U21727 (N_21727,N_20856,N_20703);
xnor U21728 (N_21728,N_20997,N_21090);
xnor U21729 (N_21729,N_20888,N_21080);
and U21730 (N_21730,N_20719,N_21196);
or U21731 (N_21731,N_21030,N_20877);
or U21732 (N_21732,N_20986,N_21072);
and U21733 (N_21733,N_20963,N_21131);
xnor U21734 (N_21734,N_20885,N_20930);
nand U21735 (N_21735,N_20926,N_20815);
or U21736 (N_21736,N_20869,N_21186);
nor U21737 (N_21737,N_21102,N_21003);
and U21738 (N_21738,N_20648,N_20909);
and U21739 (N_21739,N_21118,N_20759);
nand U21740 (N_21740,N_20734,N_20831);
xnor U21741 (N_21741,N_20771,N_20899);
xor U21742 (N_21742,N_21105,N_20694);
xor U21743 (N_21743,N_21027,N_21017);
or U21744 (N_21744,N_20945,N_20640);
and U21745 (N_21745,N_20646,N_20792);
xor U21746 (N_21746,N_21143,N_21244);
xnor U21747 (N_21747,N_20643,N_21117);
nand U21748 (N_21748,N_20727,N_20770);
xor U21749 (N_21749,N_20629,N_20856);
and U21750 (N_21750,N_20773,N_20843);
nand U21751 (N_21751,N_21235,N_21153);
or U21752 (N_21752,N_20717,N_20645);
nor U21753 (N_21753,N_20742,N_20689);
nand U21754 (N_21754,N_20718,N_20928);
nand U21755 (N_21755,N_21186,N_20804);
xor U21756 (N_21756,N_20943,N_20948);
nand U21757 (N_21757,N_21109,N_20916);
or U21758 (N_21758,N_20755,N_20657);
or U21759 (N_21759,N_21008,N_20704);
xnor U21760 (N_21760,N_20628,N_20830);
xor U21761 (N_21761,N_20714,N_21158);
xor U21762 (N_21762,N_21204,N_20754);
nand U21763 (N_21763,N_20672,N_21213);
xnor U21764 (N_21764,N_21035,N_21052);
nor U21765 (N_21765,N_20858,N_21123);
xor U21766 (N_21766,N_20974,N_21249);
or U21767 (N_21767,N_21013,N_20960);
nand U21768 (N_21768,N_20937,N_20908);
or U21769 (N_21769,N_20921,N_20817);
or U21770 (N_21770,N_20961,N_20691);
nor U21771 (N_21771,N_20889,N_21245);
and U21772 (N_21772,N_21018,N_20726);
or U21773 (N_21773,N_20830,N_20634);
and U21774 (N_21774,N_20699,N_20904);
xnor U21775 (N_21775,N_21083,N_20851);
xor U21776 (N_21776,N_21024,N_21087);
and U21777 (N_21777,N_20739,N_20793);
nand U21778 (N_21778,N_21242,N_20771);
nand U21779 (N_21779,N_21111,N_20809);
xor U21780 (N_21780,N_20874,N_20763);
nor U21781 (N_21781,N_21201,N_20818);
nand U21782 (N_21782,N_20648,N_21209);
nand U21783 (N_21783,N_20818,N_21204);
or U21784 (N_21784,N_21155,N_21023);
xor U21785 (N_21785,N_20718,N_20910);
nand U21786 (N_21786,N_20741,N_20701);
xnor U21787 (N_21787,N_20809,N_21165);
xor U21788 (N_21788,N_21037,N_21035);
or U21789 (N_21789,N_20905,N_20974);
or U21790 (N_21790,N_20743,N_20640);
xnor U21791 (N_21791,N_21198,N_21192);
xor U21792 (N_21792,N_21114,N_20922);
xor U21793 (N_21793,N_21188,N_21201);
and U21794 (N_21794,N_21226,N_20853);
and U21795 (N_21795,N_21059,N_21162);
nand U21796 (N_21796,N_20733,N_20938);
and U21797 (N_21797,N_20818,N_20977);
nand U21798 (N_21798,N_21052,N_21145);
xnor U21799 (N_21799,N_20818,N_21077);
nor U21800 (N_21800,N_20776,N_21128);
xor U21801 (N_21801,N_21146,N_20741);
nand U21802 (N_21802,N_21020,N_20690);
xnor U21803 (N_21803,N_21153,N_20695);
or U21804 (N_21804,N_21187,N_20655);
or U21805 (N_21805,N_20965,N_20756);
and U21806 (N_21806,N_20752,N_21239);
and U21807 (N_21807,N_20928,N_20846);
nor U21808 (N_21808,N_20681,N_21183);
xnor U21809 (N_21809,N_21078,N_20694);
xor U21810 (N_21810,N_20752,N_20717);
or U21811 (N_21811,N_21036,N_20786);
xor U21812 (N_21812,N_20886,N_20635);
or U21813 (N_21813,N_20813,N_21178);
nand U21814 (N_21814,N_21115,N_21219);
xnor U21815 (N_21815,N_21047,N_20877);
and U21816 (N_21816,N_20847,N_20763);
xor U21817 (N_21817,N_21155,N_21110);
nor U21818 (N_21818,N_20999,N_21103);
xor U21819 (N_21819,N_21003,N_20895);
or U21820 (N_21820,N_20953,N_20672);
or U21821 (N_21821,N_20703,N_20721);
or U21822 (N_21822,N_20972,N_21112);
nor U21823 (N_21823,N_21059,N_20719);
nand U21824 (N_21824,N_21096,N_20693);
xnor U21825 (N_21825,N_21065,N_20844);
xnor U21826 (N_21826,N_21243,N_21060);
or U21827 (N_21827,N_21012,N_21077);
xnor U21828 (N_21828,N_21013,N_21094);
xor U21829 (N_21829,N_20771,N_20927);
xnor U21830 (N_21830,N_20652,N_20676);
nand U21831 (N_21831,N_20928,N_21096);
nand U21832 (N_21832,N_21055,N_20939);
or U21833 (N_21833,N_20630,N_21188);
nor U21834 (N_21834,N_21059,N_21093);
and U21835 (N_21835,N_20644,N_20901);
and U21836 (N_21836,N_20838,N_21092);
or U21837 (N_21837,N_20969,N_21101);
xor U21838 (N_21838,N_20888,N_20886);
nor U21839 (N_21839,N_20970,N_20708);
and U21840 (N_21840,N_20656,N_21223);
nor U21841 (N_21841,N_20677,N_20703);
xnor U21842 (N_21842,N_20666,N_20927);
and U21843 (N_21843,N_20760,N_21156);
xnor U21844 (N_21844,N_20684,N_21196);
or U21845 (N_21845,N_20916,N_21247);
or U21846 (N_21846,N_20766,N_21060);
nand U21847 (N_21847,N_20881,N_21062);
xnor U21848 (N_21848,N_20991,N_21087);
and U21849 (N_21849,N_20771,N_20792);
nand U21850 (N_21850,N_20644,N_21227);
nand U21851 (N_21851,N_21194,N_21234);
xor U21852 (N_21852,N_20938,N_20799);
nor U21853 (N_21853,N_21071,N_21052);
nor U21854 (N_21854,N_21094,N_21154);
nand U21855 (N_21855,N_21015,N_21031);
xnor U21856 (N_21856,N_21156,N_21096);
and U21857 (N_21857,N_21222,N_20885);
and U21858 (N_21858,N_20716,N_20874);
or U21859 (N_21859,N_20904,N_21201);
xor U21860 (N_21860,N_21056,N_21000);
and U21861 (N_21861,N_20791,N_20626);
nor U21862 (N_21862,N_20889,N_20993);
nor U21863 (N_21863,N_21086,N_20770);
or U21864 (N_21864,N_20710,N_21220);
or U21865 (N_21865,N_20827,N_21114);
nor U21866 (N_21866,N_21141,N_20675);
nand U21867 (N_21867,N_21064,N_20925);
nor U21868 (N_21868,N_21052,N_21132);
nand U21869 (N_21869,N_20953,N_20745);
and U21870 (N_21870,N_21123,N_20863);
xor U21871 (N_21871,N_21010,N_20695);
nor U21872 (N_21872,N_21093,N_21161);
or U21873 (N_21873,N_21082,N_21167);
and U21874 (N_21874,N_20819,N_21114);
nand U21875 (N_21875,N_21659,N_21860);
nand U21876 (N_21876,N_21313,N_21324);
and U21877 (N_21877,N_21841,N_21561);
xnor U21878 (N_21878,N_21795,N_21383);
nor U21879 (N_21879,N_21868,N_21723);
nand U21880 (N_21880,N_21530,N_21271);
xor U21881 (N_21881,N_21361,N_21499);
or U21882 (N_21882,N_21785,N_21376);
and U21883 (N_21883,N_21439,N_21818);
or U21884 (N_21884,N_21745,N_21608);
or U21885 (N_21885,N_21719,N_21382);
or U21886 (N_21886,N_21472,N_21728);
or U21887 (N_21887,N_21270,N_21698);
nor U21888 (N_21888,N_21636,N_21549);
xor U21889 (N_21889,N_21465,N_21545);
and U21890 (N_21890,N_21768,N_21623);
or U21891 (N_21891,N_21337,N_21796);
xor U21892 (N_21892,N_21260,N_21718);
xor U21893 (N_21893,N_21613,N_21824);
xor U21894 (N_21894,N_21693,N_21857);
nor U21895 (N_21895,N_21327,N_21848);
nor U21896 (N_21896,N_21412,N_21488);
or U21897 (N_21897,N_21807,N_21837);
nor U21898 (N_21898,N_21655,N_21759);
nor U21899 (N_21899,N_21819,N_21476);
or U21900 (N_21900,N_21790,N_21451);
or U21901 (N_21901,N_21696,N_21832);
xor U21902 (N_21902,N_21455,N_21815);
nor U21903 (N_21903,N_21869,N_21839);
xnor U21904 (N_21904,N_21264,N_21748);
xor U21905 (N_21905,N_21304,N_21865);
nor U21906 (N_21906,N_21553,N_21385);
nor U21907 (N_21907,N_21867,N_21715);
or U21908 (N_21908,N_21544,N_21820);
and U21909 (N_21909,N_21434,N_21261);
xor U21910 (N_21910,N_21626,N_21458);
nand U21911 (N_21911,N_21285,N_21483);
or U21912 (N_21912,N_21783,N_21666);
or U21913 (N_21913,N_21317,N_21486);
and U21914 (N_21914,N_21300,N_21870);
nor U21915 (N_21915,N_21701,N_21691);
and U21916 (N_21916,N_21849,N_21532);
xnor U21917 (N_21917,N_21552,N_21631);
and U21918 (N_21918,N_21787,N_21695);
nor U21919 (N_21919,N_21834,N_21821);
or U21920 (N_21920,N_21764,N_21363);
nand U21921 (N_21921,N_21510,N_21273);
and U21922 (N_21922,N_21357,N_21755);
nand U21923 (N_21923,N_21408,N_21560);
nor U21924 (N_21924,N_21453,N_21605);
nand U21925 (N_21925,N_21296,N_21487);
nor U21926 (N_21926,N_21437,N_21491);
nand U21927 (N_21927,N_21618,N_21612);
and U21928 (N_21928,N_21781,N_21754);
xor U21929 (N_21929,N_21444,N_21752);
or U21930 (N_21930,N_21591,N_21678);
xor U21931 (N_21931,N_21812,N_21393);
or U21932 (N_21932,N_21526,N_21333);
nor U21933 (N_21933,N_21845,N_21420);
xor U21934 (N_21934,N_21474,N_21395);
and U21935 (N_21935,N_21694,N_21717);
or U21936 (N_21936,N_21684,N_21543);
and U21937 (N_21937,N_21257,N_21596);
nand U21938 (N_21938,N_21443,N_21828);
or U21939 (N_21939,N_21582,N_21550);
or U21940 (N_21940,N_21429,N_21464);
nor U21941 (N_21941,N_21531,N_21722);
nand U21942 (N_21942,N_21256,N_21725);
or U21943 (N_21943,N_21567,N_21497);
nor U21944 (N_21944,N_21388,N_21289);
xnor U21945 (N_21945,N_21836,N_21572);
and U21946 (N_21946,N_21705,N_21398);
and U21947 (N_21947,N_21417,N_21772);
or U21948 (N_21948,N_21592,N_21290);
nand U21949 (N_21949,N_21365,N_21629);
xnor U21950 (N_21950,N_21374,N_21858);
or U21951 (N_21951,N_21840,N_21616);
nor U21952 (N_21952,N_21386,N_21829);
nor U21953 (N_21953,N_21338,N_21811);
or U21954 (N_21954,N_21511,N_21320);
nor U21955 (N_21955,N_21842,N_21822);
or U21956 (N_21956,N_21419,N_21650);
nor U21957 (N_21957,N_21546,N_21354);
or U21958 (N_21958,N_21344,N_21776);
or U21959 (N_21959,N_21686,N_21283);
or U21960 (N_21960,N_21424,N_21358);
nor U21961 (N_21961,N_21527,N_21771);
xor U21962 (N_21962,N_21460,N_21797);
or U21963 (N_21963,N_21577,N_21565);
nor U21964 (N_21964,N_21287,N_21648);
or U21965 (N_21965,N_21538,N_21670);
and U21966 (N_21966,N_21607,N_21676);
and U21967 (N_21967,N_21709,N_21602);
nand U21968 (N_21968,N_21555,N_21475);
nor U21969 (N_21969,N_21319,N_21533);
or U21970 (N_21970,N_21663,N_21584);
nor U21971 (N_21971,N_21494,N_21806);
and U21972 (N_21972,N_21862,N_21833);
xnor U21973 (N_21973,N_21428,N_21665);
or U21974 (N_21974,N_21551,N_21466);
xor U21975 (N_21975,N_21254,N_21721);
or U21976 (N_21976,N_21542,N_21590);
or U21977 (N_21977,N_21432,N_21800);
nand U21978 (N_21978,N_21766,N_21547);
nand U21979 (N_21979,N_21266,N_21620);
xnor U21980 (N_21980,N_21813,N_21562);
or U21981 (N_21981,N_21353,N_21843);
xnor U21982 (N_21982,N_21816,N_21461);
xnor U21983 (N_21983,N_21263,N_21442);
nor U21984 (N_21984,N_21788,N_21568);
or U21985 (N_21985,N_21392,N_21606);
xor U21986 (N_21986,N_21431,N_21328);
and U21987 (N_21987,N_21653,N_21658);
and U21988 (N_21988,N_21803,N_21851);
nand U21989 (N_21989,N_21724,N_21765);
nor U21990 (N_21990,N_21571,N_21441);
nand U21991 (N_21991,N_21746,N_21704);
nand U21992 (N_21992,N_21447,N_21739);
nor U21993 (N_21993,N_21471,N_21651);
xnor U21994 (N_21994,N_21681,N_21307);
xnor U21995 (N_21995,N_21780,N_21347);
nand U21996 (N_21996,N_21640,N_21401);
nor U21997 (N_21997,N_21515,N_21574);
nor U21998 (N_21998,N_21864,N_21773);
xnor U21999 (N_21999,N_21610,N_21329);
nand U22000 (N_22000,N_21277,N_21762);
nand U22001 (N_22001,N_21838,N_21303);
and U22002 (N_22002,N_21258,N_21680);
xnor U22003 (N_22003,N_21378,N_21734);
nand U22004 (N_22004,N_21399,N_21570);
nor U22005 (N_22005,N_21667,N_21481);
xor U22006 (N_22006,N_21617,N_21622);
or U22007 (N_22007,N_21854,N_21334);
or U22008 (N_22008,N_21459,N_21597);
xnor U22009 (N_22009,N_21316,N_21830);
xor U22010 (N_22010,N_21331,N_21688);
and U22011 (N_22011,N_21554,N_21588);
or U22012 (N_22012,N_21402,N_21265);
xor U22013 (N_22013,N_21575,N_21438);
and U22014 (N_22014,N_21343,N_21583);
or U22015 (N_22015,N_21835,N_21740);
nor U22016 (N_22016,N_21373,N_21769);
xor U22017 (N_22017,N_21791,N_21786);
or U22018 (N_22018,N_21478,N_21528);
xnor U22019 (N_22019,N_21381,N_21844);
or U22020 (N_22020,N_21831,N_21804);
xor U22021 (N_22021,N_21578,N_21537);
xnor U22022 (N_22022,N_21673,N_21866);
nand U22023 (N_22023,N_21413,N_21517);
nor U22024 (N_22024,N_21297,N_21418);
nand U22025 (N_22025,N_21871,N_21863);
nor U22026 (N_22026,N_21782,N_21586);
or U22027 (N_22027,N_21468,N_21405);
or U22028 (N_22028,N_21284,N_21359);
nand U22029 (N_22029,N_21456,N_21262);
or U22030 (N_22030,N_21416,N_21377);
nand U22031 (N_22031,N_21855,N_21664);
nand U22032 (N_22032,N_21457,N_21332);
nor U22033 (N_22033,N_21306,N_21579);
and U22034 (N_22034,N_21825,N_21581);
xnor U22035 (N_22035,N_21339,N_21506);
nor U22036 (N_22036,N_21371,N_21730);
nand U22037 (N_22037,N_21390,N_21627);
nor U22038 (N_22038,N_21372,N_21736);
xor U22039 (N_22039,N_21817,N_21874);
or U22040 (N_22040,N_21400,N_21639);
nand U22041 (N_22041,N_21556,N_21519);
or U22042 (N_22042,N_21580,N_21326);
nand U22043 (N_22043,N_21802,N_21706);
nor U22044 (N_22044,N_21852,N_21446);
xnor U22045 (N_22045,N_21859,N_21305);
or U22046 (N_22046,N_21634,N_21774);
and U22047 (N_22047,N_21635,N_21268);
and U22048 (N_22048,N_21536,N_21861);
xnor U22049 (N_22049,N_21259,N_21793);
and U22050 (N_22050,N_21250,N_21727);
and U22051 (N_22051,N_21683,N_21741);
nand U22052 (N_22052,N_21599,N_21689);
or U22053 (N_22053,N_21614,N_21323);
or U22054 (N_22054,N_21563,N_21440);
and U22055 (N_22055,N_21710,N_21425);
or U22056 (N_22056,N_21403,N_21692);
nand U22057 (N_22057,N_21489,N_21674);
nand U22058 (N_22058,N_21362,N_21308);
and U22059 (N_22059,N_21703,N_21751);
or U22060 (N_22060,N_21348,N_21448);
xnor U22061 (N_22061,N_21801,N_21505);
nand U22062 (N_22062,N_21573,N_21540);
and U22063 (N_22063,N_21445,N_21529);
and U22064 (N_22064,N_21314,N_21702);
nor U22065 (N_22065,N_21559,N_21729);
nor U22066 (N_22066,N_21379,N_21760);
nor U22067 (N_22067,N_21593,N_21652);
or U22068 (N_22068,N_21467,N_21345);
and U22069 (N_22069,N_21604,N_21758);
nor U22070 (N_22070,N_21850,N_21414);
xor U22071 (N_22071,N_21501,N_21585);
and U22072 (N_22072,N_21375,N_21384);
or U22073 (N_22073,N_21252,N_21707);
nor U22074 (N_22074,N_21679,N_21387);
nor U22075 (N_22075,N_21473,N_21777);
xor U22076 (N_22076,N_21415,N_21669);
or U22077 (N_22077,N_21594,N_21720);
or U22078 (N_22078,N_21479,N_21394);
nor U22079 (N_22079,N_21430,N_21292);
or U22080 (N_22080,N_21856,N_21763);
or U22081 (N_22081,N_21732,N_21355);
xor U22082 (N_22082,N_21598,N_21743);
nand U22083 (N_22083,N_21294,N_21778);
and U22084 (N_22084,N_21534,N_21668);
and U22085 (N_22085,N_21566,N_21619);
or U22086 (N_22086,N_21504,N_21711);
and U22087 (N_22087,N_21496,N_21814);
or U22088 (N_22088,N_21779,N_21642);
nor U22089 (N_22089,N_21525,N_21794);
nand U22090 (N_22090,N_21310,N_21298);
nor U22091 (N_22091,N_21846,N_21675);
nand U22092 (N_22092,N_21708,N_21690);
nor U22093 (N_22093,N_21340,N_21342);
and U22094 (N_22094,N_21737,N_21823);
nand U22095 (N_22095,N_21770,N_21368);
nor U22096 (N_22096,N_21426,N_21352);
nor U22097 (N_22097,N_21280,N_21660);
nand U22098 (N_22098,N_21299,N_21495);
and U22099 (N_22099,N_21799,N_21662);
and U22100 (N_22100,N_21366,N_21433);
xnor U22101 (N_22101,N_21411,N_21253);
and U22102 (N_22102,N_21450,N_21350);
nor U22103 (N_22103,N_21436,N_21454);
and U22104 (N_22104,N_21557,N_21523);
and U22105 (N_22105,N_21435,N_21853);
or U22106 (N_22106,N_21671,N_21621);
xnor U22107 (N_22107,N_21661,N_21672);
xnor U22108 (N_22108,N_21784,N_21827);
xnor U22109 (N_22109,N_21269,N_21480);
nor U22110 (N_22110,N_21477,N_21603);
nand U22111 (N_22111,N_21847,N_21321);
nand U22112 (N_22112,N_21346,N_21498);
and U22113 (N_22113,N_21569,N_21322);
nor U22114 (N_22114,N_21315,N_21512);
and U22115 (N_22115,N_21513,N_21356);
and U22116 (N_22116,N_21389,N_21370);
or U22117 (N_22117,N_21548,N_21482);
or U22118 (N_22118,N_21600,N_21826);
xor U22119 (N_22119,N_21789,N_21539);
and U22120 (N_22120,N_21509,N_21716);
xor U22121 (N_22121,N_21463,N_21335);
and U22122 (N_22122,N_21757,N_21421);
or U22123 (N_22123,N_21756,N_21427);
and U22124 (N_22124,N_21873,N_21589);
xor U22125 (N_22125,N_21521,N_21484);
nand U22126 (N_22126,N_21485,N_21742);
nor U22127 (N_22127,N_21302,N_21470);
nand U22128 (N_22128,N_21291,N_21731);
or U22129 (N_22129,N_21391,N_21351);
and U22130 (N_22130,N_21687,N_21507);
nand U22131 (N_22131,N_21628,N_21251);
nor U22132 (N_22132,N_21514,N_21311);
and U22133 (N_22133,N_21638,N_21753);
nand U22134 (N_22134,N_21587,N_21798);
or U22135 (N_22135,N_21404,N_21792);
or U22136 (N_22136,N_21682,N_21601);
or U22137 (N_22137,N_21423,N_21407);
and U22138 (N_22138,N_21611,N_21808);
nor U22139 (N_22139,N_21276,N_21535);
or U22140 (N_22140,N_21645,N_21632);
nand U22141 (N_22141,N_21422,N_21406);
or U22142 (N_22142,N_21449,N_21685);
nand U22143 (N_22143,N_21522,N_21295);
nor U22144 (N_22144,N_21810,N_21278);
xnor U22145 (N_22145,N_21647,N_21272);
xnor U22146 (N_22146,N_21699,N_21330);
nor U22147 (N_22147,N_21309,N_21367);
nor U22148 (N_22148,N_21360,N_21749);
and U22149 (N_22149,N_21462,N_21624);
and U22150 (N_22150,N_21397,N_21646);
or U22151 (N_22151,N_21396,N_21518);
and U22152 (N_22152,N_21630,N_21644);
or U22153 (N_22153,N_21733,N_21286);
and U22154 (N_22154,N_21492,N_21767);
and U22155 (N_22155,N_21349,N_21654);
or U22156 (N_22156,N_21595,N_21369);
xnor U22157 (N_22157,N_21738,N_21452);
nand U22158 (N_22158,N_21274,N_21490);
xor U22159 (N_22159,N_21508,N_21524);
xnor U22160 (N_22160,N_21697,N_21541);
and U22161 (N_22161,N_21255,N_21712);
xnor U22162 (N_22162,N_21714,N_21641);
xor U22163 (N_22163,N_21267,N_21301);
xor U22164 (N_22164,N_21380,N_21809);
nor U22165 (N_22165,N_21469,N_21726);
or U22166 (N_22166,N_21281,N_21747);
or U22167 (N_22167,N_21677,N_21657);
nand U22168 (N_22168,N_21282,N_21516);
or U22169 (N_22169,N_21312,N_21633);
nor U22170 (N_22170,N_21750,N_21325);
and U22171 (N_22171,N_21649,N_21500);
or U22172 (N_22172,N_21503,N_21493);
nor U22173 (N_22173,N_21656,N_21615);
and U22174 (N_22174,N_21502,N_21564);
nor U22175 (N_22175,N_21744,N_21293);
and U22176 (N_22176,N_21643,N_21318);
nand U22177 (N_22177,N_21576,N_21775);
xnor U22178 (N_22178,N_21288,N_21364);
xnor U22179 (N_22179,N_21637,N_21713);
xnor U22180 (N_22180,N_21520,N_21700);
or U22181 (N_22181,N_21409,N_21625);
xor U22182 (N_22182,N_21341,N_21275);
and U22183 (N_22183,N_21558,N_21805);
nor U22184 (N_22184,N_21872,N_21761);
nor U22185 (N_22185,N_21609,N_21410);
and U22186 (N_22186,N_21279,N_21336);
or U22187 (N_22187,N_21735,N_21610);
nor U22188 (N_22188,N_21426,N_21867);
nand U22189 (N_22189,N_21367,N_21795);
and U22190 (N_22190,N_21776,N_21438);
nor U22191 (N_22191,N_21656,N_21699);
or U22192 (N_22192,N_21570,N_21845);
and U22193 (N_22193,N_21566,N_21710);
nand U22194 (N_22194,N_21500,N_21605);
and U22195 (N_22195,N_21722,N_21667);
nand U22196 (N_22196,N_21316,N_21488);
nand U22197 (N_22197,N_21601,N_21304);
nand U22198 (N_22198,N_21251,N_21256);
nand U22199 (N_22199,N_21683,N_21673);
or U22200 (N_22200,N_21845,N_21837);
and U22201 (N_22201,N_21548,N_21725);
nor U22202 (N_22202,N_21396,N_21485);
nor U22203 (N_22203,N_21608,N_21588);
nand U22204 (N_22204,N_21802,N_21682);
nand U22205 (N_22205,N_21542,N_21849);
nor U22206 (N_22206,N_21725,N_21339);
nor U22207 (N_22207,N_21374,N_21863);
or U22208 (N_22208,N_21743,N_21523);
nand U22209 (N_22209,N_21253,N_21725);
xnor U22210 (N_22210,N_21860,N_21607);
nor U22211 (N_22211,N_21711,N_21846);
nand U22212 (N_22212,N_21870,N_21770);
nand U22213 (N_22213,N_21692,N_21335);
or U22214 (N_22214,N_21671,N_21708);
and U22215 (N_22215,N_21626,N_21789);
nor U22216 (N_22216,N_21733,N_21495);
nor U22217 (N_22217,N_21730,N_21579);
xor U22218 (N_22218,N_21477,N_21673);
xor U22219 (N_22219,N_21277,N_21851);
xor U22220 (N_22220,N_21480,N_21310);
xnor U22221 (N_22221,N_21616,N_21295);
and U22222 (N_22222,N_21743,N_21720);
nand U22223 (N_22223,N_21638,N_21494);
or U22224 (N_22224,N_21592,N_21782);
nand U22225 (N_22225,N_21456,N_21714);
nand U22226 (N_22226,N_21264,N_21565);
xor U22227 (N_22227,N_21624,N_21590);
nor U22228 (N_22228,N_21735,N_21344);
or U22229 (N_22229,N_21702,N_21554);
and U22230 (N_22230,N_21720,N_21310);
xnor U22231 (N_22231,N_21706,N_21658);
nor U22232 (N_22232,N_21420,N_21422);
and U22233 (N_22233,N_21450,N_21442);
xnor U22234 (N_22234,N_21474,N_21596);
nor U22235 (N_22235,N_21367,N_21816);
nor U22236 (N_22236,N_21872,N_21821);
xor U22237 (N_22237,N_21714,N_21543);
nor U22238 (N_22238,N_21666,N_21527);
nor U22239 (N_22239,N_21342,N_21626);
nor U22240 (N_22240,N_21487,N_21404);
and U22241 (N_22241,N_21623,N_21591);
nor U22242 (N_22242,N_21758,N_21548);
and U22243 (N_22243,N_21328,N_21589);
xnor U22244 (N_22244,N_21632,N_21393);
xor U22245 (N_22245,N_21312,N_21874);
nand U22246 (N_22246,N_21588,N_21612);
nor U22247 (N_22247,N_21625,N_21696);
nand U22248 (N_22248,N_21833,N_21493);
or U22249 (N_22249,N_21566,N_21870);
nand U22250 (N_22250,N_21422,N_21568);
and U22251 (N_22251,N_21371,N_21552);
nor U22252 (N_22252,N_21602,N_21376);
and U22253 (N_22253,N_21314,N_21511);
nand U22254 (N_22254,N_21604,N_21613);
nand U22255 (N_22255,N_21322,N_21296);
or U22256 (N_22256,N_21354,N_21749);
or U22257 (N_22257,N_21286,N_21269);
nor U22258 (N_22258,N_21283,N_21757);
and U22259 (N_22259,N_21760,N_21326);
xor U22260 (N_22260,N_21502,N_21365);
xor U22261 (N_22261,N_21599,N_21343);
xnor U22262 (N_22262,N_21639,N_21408);
nand U22263 (N_22263,N_21427,N_21564);
nor U22264 (N_22264,N_21358,N_21684);
nand U22265 (N_22265,N_21629,N_21481);
and U22266 (N_22266,N_21638,N_21792);
and U22267 (N_22267,N_21633,N_21678);
xor U22268 (N_22268,N_21864,N_21406);
or U22269 (N_22269,N_21450,N_21637);
nand U22270 (N_22270,N_21440,N_21698);
and U22271 (N_22271,N_21272,N_21544);
nand U22272 (N_22272,N_21361,N_21817);
xnor U22273 (N_22273,N_21563,N_21722);
xor U22274 (N_22274,N_21725,N_21748);
and U22275 (N_22275,N_21397,N_21639);
nor U22276 (N_22276,N_21746,N_21570);
nor U22277 (N_22277,N_21845,N_21645);
nand U22278 (N_22278,N_21449,N_21334);
xor U22279 (N_22279,N_21279,N_21691);
and U22280 (N_22280,N_21719,N_21422);
and U22281 (N_22281,N_21764,N_21381);
or U22282 (N_22282,N_21780,N_21459);
nand U22283 (N_22283,N_21833,N_21457);
nor U22284 (N_22284,N_21717,N_21536);
or U22285 (N_22285,N_21837,N_21828);
xnor U22286 (N_22286,N_21793,N_21778);
nor U22287 (N_22287,N_21413,N_21612);
or U22288 (N_22288,N_21722,N_21640);
and U22289 (N_22289,N_21257,N_21594);
xnor U22290 (N_22290,N_21478,N_21653);
and U22291 (N_22291,N_21613,N_21342);
nand U22292 (N_22292,N_21651,N_21728);
nand U22293 (N_22293,N_21480,N_21821);
and U22294 (N_22294,N_21659,N_21271);
or U22295 (N_22295,N_21363,N_21361);
and U22296 (N_22296,N_21450,N_21830);
nand U22297 (N_22297,N_21728,N_21372);
and U22298 (N_22298,N_21691,N_21630);
nand U22299 (N_22299,N_21480,N_21776);
nand U22300 (N_22300,N_21324,N_21511);
or U22301 (N_22301,N_21681,N_21660);
nand U22302 (N_22302,N_21516,N_21439);
nand U22303 (N_22303,N_21368,N_21746);
nor U22304 (N_22304,N_21420,N_21301);
nand U22305 (N_22305,N_21411,N_21349);
xor U22306 (N_22306,N_21592,N_21680);
xnor U22307 (N_22307,N_21462,N_21404);
or U22308 (N_22308,N_21547,N_21480);
nor U22309 (N_22309,N_21486,N_21421);
nor U22310 (N_22310,N_21700,N_21448);
xnor U22311 (N_22311,N_21722,N_21709);
or U22312 (N_22312,N_21394,N_21771);
and U22313 (N_22313,N_21307,N_21260);
or U22314 (N_22314,N_21478,N_21572);
and U22315 (N_22315,N_21473,N_21420);
xnor U22316 (N_22316,N_21370,N_21328);
xor U22317 (N_22317,N_21502,N_21712);
nor U22318 (N_22318,N_21280,N_21695);
and U22319 (N_22319,N_21621,N_21826);
nand U22320 (N_22320,N_21259,N_21498);
or U22321 (N_22321,N_21668,N_21275);
and U22322 (N_22322,N_21316,N_21706);
nor U22323 (N_22323,N_21409,N_21716);
and U22324 (N_22324,N_21799,N_21403);
nand U22325 (N_22325,N_21539,N_21291);
xor U22326 (N_22326,N_21807,N_21808);
xor U22327 (N_22327,N_21488,N_21391);
nand U22328 (N_22328,N_21755,N_21855);
nand U22329 (N_22329,N_21836,N_21414);
or U22330 (N_22330,N_21650,N_21779);
or U22331 (N_22331,N_21464,N_21664);
nand U22332 (N_22332,N_21349,N_21475);
nor U22333 (N_22333,N_21586,N_21303);
and U22334 (N_22334,N_21568,N_21783);
and U22335 (N_22335,N_21263,N_21841);
nor U22336 (N_22336,N_21509,N_21375);
nor U22337 (N_22337,N_21867,N_21528);
nor U22338 (N_22338,N_21868,N_21526);
xnor U22339 (N_22339,N_21316,N_21384);
and U22340 (N_22340,N_21296,N_21514);
and U22341 (N_22341,N_21525,N_21353);
or U22342 (N_22342,N_21636,N_21795);
xnor U22343 (N_22343,N_21651,N_21527);
xnor U22344 (N_22344,N_21732,N_21768);
nor U22345 (N_22345,N_21668,N_21730);
and U22346 (N_22346,N_21752,N_21755);
or U22347 (N_22347,N_21416,N_21449);
nand U22348 (N_22348,N_21661,N_21793);
nor U22349 (N_22349,N_21517,N_21615);
or U22350 (N_22350,N_21871,N_21532);
and U22351 (N_22351,N_21497,N_21490);
nand U22352 (N_22352,N_21609,N_21577);
nand U22353 (N_22353,N_21579,N_21288);
nor U22354 (N_22354,N_21467,N_21312);
nand U22355 (N_22355,N_21429,N_21377);
and U22356 (N_22356,N_21614,N_21284);
nand U22357 (N_22357,N_21857,N_21785);
and U22358 (N_22358,N_21699,N_21399);
nand U22359 (N_22359,N_21655,N_21331);
nor U22360 (N_22360,N_21420,N_21308);
and U22361 (N_22361,N_21446,N_21834);
nand U22362 (N_22362,N_21570,N_21868);
or U22363 (N_22363,N_21569,N_21381);
nand U22364 (N_22364,N_21336,N_21765);
nor U22365 (N_22365,N_21607,N_21412);
nand U22366 (N_22366,N_21748,N_21652);
nor U22367 (N_22367,N_21481,N_21623);
nor U22368 (N_22368,N_21315,N_21290);
xnor U22369 (N_22369,N_21260,N_21425);
and U22370 (N_22370,N_21365,N_21772);
xor U22371 (N_22371,N_21680,N_21533);
nor U22372 (N_22372,N_21444,N_21751);
nor U22373 (N_22373,N_21457,N_21319);
nor U22374 (N_22374,N_21371,N_21535);
or U22375 (N_22375,N_21666,N_21728);
nor U22376 (N_22376,N_21377,N_21804);
or U22377 (N_22377,N_21412,N_21757);
or U22378 (N_22378,N_21421,N_21398);
nor U22379 (N_22379,N_21785,N_21679);
nor U22380 (N_22380,N_21366,N_21650);
and U22381 (N_22381,N_21253,N_21836);
and U22382 (N_22382,N_21574,N_21550);
nand U22383 (N_22383,N_21794,N_21492);
xnor U22384 (N_22384,N_21518,N_21559);
nor U22385 (N_22385,N_21551,N_21871);
or U22386 (N_22386,N_21670,N_21286);
nor U22387 (N_22387,N_21421,N_21756);
nor U22388 (N_22388,N_21344,N_21422);
nor U22389 (N_22389,N_21480,N_21315);
or U22390 (N_22390,N_21314,N_21440);
nor U22391 (N_22391,N_21481,N_21822);
xnor U22392 (N_22392,N_21558,N_21349);
and U22393 (N_22393,N_21786,N_21723);
nand U22394 (N_22394,N_21523,N_21639);
nor U22395 (N_22395,N_21618,N_21465);
nor U22396 (N_22396,N_21696,N_21500);
and U22397 (N_22397,N_21331,N_21377);
xor U22398 (N_22398,N_21750,N_21769);
and U22399 (N_22399,N_21648,N_21742);
or U22400 (N_22400,N_21578,N_21789);
and U22401 (N_22401,N_21493,N_21301);
nor U22402 (N_22402,N_21675,N_21488);
and U22403 (N_22403,N_21775,N_21550);
nor U22404 (N_22404,N_21432,N_21786);
or U22405 (N_22405,N_21673,N_21454);
nor U22406 (N_22406,N_21684,N_21393);
and U22407 (N_22407,N_21594,N_21397);
nor U22408 (N_22408,N_21406,N_21473);
and U22409 (N_22409,N_21644,N_21790);
nor U22410 (N_22410,N_21748,N_21481);
nand U22411 (N_22411,N_21590,N_21507);
nand U22412 (N_22412,N_21687,N_21590);
nand U22413 (N_22413,N_21798,N_21736);
nand U22414 (N_22414,N_21620,N_21255);
nor U22415 (N_22415,N_21350,N_21648);
nor U22416 (N_22416,N_21579,N_21538);
nand U22417 (N_22417,N_21741,N_21574);
or U22418 (N_22418,N_21315,N_21612);
nor U22419 (N_22419,N_21656,N_21722);
xnor U22420 (N_22420,N_21493,N_21671);
nor U22421 (N_22421,N_21587,N_21800);
xor U22422 (N_22422,N_21368,N_21652);
nor U22423 (N_22423,N_21844,N_21459);
and U22424 (N_22424,N_21744,N_21358);
nor U22425 (N_22425,N_21492,N_21284);
nand U22426 (N_22426,N_21501,N_21303);
nand U22427 (N_22427,N_21259,N_21803);
or U22428 (N_22428,N_21593,N_21319);
xor U22429 (N_22429,N_21811,N_21308);
nand U22430 (N_22430,N_21463,N_21360);
nand U22431 (N_22431,N_21649,N_21607);
and U22432 (N_22432,N_21737,N_21436);
and U22433 (N_22433,N_21641,N_21288);
nor U22434 (N_22434,N_21406,N_21552);
xor U22435 (N_22435,N_21594,N_21549);
nand U22436 (N_22436,N_21252,N_21581);
and U22437 (N_22437,N_21747,N_21670);
nor U22438 (N_22438,N_21292,N_21419);
xnor U22439 (N_22439,N_21472,N_21822);
and U22440 (N_22440,N_21851,N_21500);
xnor U22441 (N_22441,N_21439,N_21420);
or U22442 (N_22442,N_21539,N_21365);
xnor U22443 (N_22443,N_21702,N_21558);
nor U22444 (N_22444,N_21847,N_21530);
or U22445 (N_22445,N_21315,N_21775);
xnor U22446 (N_22446,N_21750,N_21868);
or U22447 (N_22447,N_21702,N_21736);
nand U22448 (N_22448,N_21488,N_21864);
and U22449 (N_22449,N_21868,N_21272);
xor U22450 (N_22450,N_21699,N_21796);
xnor U22451 (N_22451,N_21498,N_21287);
and U22452 (N_22452,N_21720,N_21713);
xor U22453 (N_22453,N_21438,N_21743);
or U22454 (N_22454,N_21630,N_21701);
nor U22455 (N_22455,N_21541,N_21311);
nand U22456 (N_22456,N_21478,N_21519);
or U22457 (N_22457,N_21250,N_21464);
xnor U22458 (N_22458,N_21792,N_21322);
and U22459 (N_22459,N_21603,N_21498);
nor U22460 (N_22460,N_21662,N_21599);
nand U22461 (N_22461,N_21516,N_21544);
xnor U22462 (N_22462,N_21384,N_21288);
or U22463 (N_22463,N_21575,N_21626);
and U22464 (N_22464,N_21797,N_21745);
or U22465 (N_22465,N_21605,N_21870);
nand U22466 (N_22466,N_21675,N_21278);
xor U22467 (N_22467,N_21714,N_21534);
or U22468 (N_22468,N_21761,N_21614);
xor U22469 (N_22469,N_21642,N_21409);
or U22470 (N_22470,N_21818,N_21871);
and U22471 (N_22471,N_21511,N_21315);
xnor U22472 (N_22472,N_21307,N_21794);
or U22473 (N_22473,N_21267,N_21484);
nand U22474 (N_22474,N_21806,N_21659);
nor U22475 (N_22475,N_21868,N_21250);
xnor U22476 (N_22476,N_21312,N_21409);
nor U22477 (N_22477,N_21283,N_21521);
nor U22478 (N_22478,N_21485,N_21651);
xnor U22479 (N_22479,N_21740,N_21863);
and U22480 (N_22480,N_21420,N_21286);
and U22481 (N_22481,N_21646,N_21761);
nor U22482 (N_22482,N_21375,N_21748);
nor U22483 (N_22483,N_21661,N_21546);
or U22484 (N_22484,N_21574,N_21614);
and U22485 (N_22485,N_21698,N_21612);
nand U22486 (N_22486,N_21867,N_21266);
nor U22487 (N_22487,N_21730,N_21825);
nand U22488 (N_22488,N_21339,N_21641);
or U22489 (N_22489,N_21874,N_21515);
nor U22490 (N_22490,N_21290,N_21716);
or U22491 (N_22491,N_21289,N_21628);
xor U22492 (N_22492,N_21810,N_21402);
xor U22493 (N_22493,N_21552,N_21803);
or U22494 (N_22494,N_21680,N_21590);
xnor U22495 (N_22495,N_21272,N_21368);
nor U22496 (N_22496,N_21299,N_21485);
and U22497 (N_22497,N_21448,N_21596);
nand U22498 (N_22498,N_21374,N_21588);
nand U22499 (N_22499,N_21816,N_21463);
nand U22500 (N_22500,N_22268,N_22147);
or U22501 (N_22501,N_22128,N_22409);
xnor U22502 (N_22502,N_22167,N_21907);
or U22503 (N_22503,N_22118,N_22233);
nand U22504 (N_22504,N_21910,N_21908);
or U22505 (N_22505,N_22249,N_22419);
xnor U22506 (N_22506,N_22225,N_22485);
nand U22507 (N_22507,N_22273,N_21929);
nor U22508 (N_22508,N_22113,N_22130);
nor U22509 (N_22509,N_22183,N_21946);
nor U22510 (N_22510,N_21882,N_22139);
nor U22511 (N_22511,N_22142,N_22100);
and U22512 (N_22512,N_22279,N_22383);
or U22513 (N_22513,N_22387,N_22272);
nand U22514 (N_22514,N_22017,N_22205);
and U22515 (N_22515,N_21912,N_22253);
nand U22516 (N_22516,N_22389,N_22263);
nor U22517 (N_22517,N_22022,N_22252);
xor U22518 (N_22518,N_22236,N_22226);
nand U22519 (N_22519,N_22056,N_21959);
nor U22520 (N_22520,N_22475,N_22265);
nor U22521 (N_22521,N_22498,N_22317);
or U22522 (N_22522,N_22460,N_22243);
xnor U22523 (N_22523,N_22415,N_21962);
nand U22524 (N_22524,N_22186,N_22270);
nor U22525 (N_22525,N_22166,N_21937);
xnor U22526 (N_22526,N_21881,N_22098);
nor U22527 (N_22527,N_22486,N_22020);
and U22528 (N_22528,N_22030,N_21968);
and U22529 (N_22529,N_22239,N_21961);
nor U22530 (N_22530,N_21988,N_21885);
nor U22531 (N_22531,N_22255,N_22333);
and U22532 (N_22532,N_21918,N_22032);
xor U22533 (N_22533,N_22354,N_21933);
xnor U22534 (N_22534,N_22439,N_21976);
nand U22535 (N_22535,N_21945,N_22169);
nor U22536 (N_22536,N_22002,N_21935);
or U22537 (N_22537,N_22365,N_22048);
or U22538 (N_22538,N_22384,N_22337);
nand U22539 (N_22539,N_22143,N_22036);
or U22540 (N_22540,N_22094,N_21896);
or U22541 (N_22541,N_22037,N_22442);
and U22542 (N_22542,N_22338,N_22106);
nand U22543 (N_22543,N_22040,N_22457);
nand U22544 (N_22544,N_22391,N_22479);
or U22545 (N_22545,N_22136,N_22348);
xnor U22546 (N_22546,N_22095,N_22112);
or U22547 (N_22547,N_21998,N_22119);
or U22548 (N_22548,N_22231,N_22444);
nor U22549 (N_22549,N_22286,N_21963);
or U22550 (N_22550,N_22445,N_22410);
nor U22551 (N_22551,N_22406,N_22193);
xor U22552 (N_22552,N_22257,N_21985);
and U22553 (N_22553,N_22102,N_22499);
xor U22554 (N_22554,N_21980,N_22180);
xor U22555 (N_22555,N_21971,N_22456);
nand U22556 (N_22556,N_22437,N_22114);
xnor U22557 (N_22557,N_22197,N_22206);
xnor U22558 (N_22558,N_22086,N_21887);
and U22559 (N_22559,N_22492,N_22245);
nand U22560 (N_22560,N_22079,N_22035);
xnor U22561 (N_22561,N_22140,N_22379);
xor U22562 (N_22562,N_22237,N_22052);
nand U22563 (N_22563,N_22440,N_22380);
nand U22564 (N_22564,N_22356,N_22353);
nor U22565 (N_22565,N_22378,N_22395);
nand U22566 (N_22566,N_22085,N_22244);
xnor U22567 (N_22567,N_22155,N_22224);
or U22568 (N_22568,N_21909,N_22447);
or U22569 (N_22569,N_22015,N_22152);
and U22570 (N_22570,N_22261,N_22050);
nand U22571 (N_22571,N_22133,N_22163);
and U22572 (N_22572,N_21940,N_22246);
and U22573 (N_22573,N_22123,N_22352);
xor U22574 (N_22574,N_22208,N_22459);
or U22575 (N_22575,N_22340,N_22464);
or U22576 (N_22576,N_22107,N_22179);
nand U22577 (N_22577,N_22285,N_22369);
xnor U22578 (N_22578,N_21905,N_22199);
nand U22579 (N_22579,N_21990,N_21915);
nand U22580 (N_22580,N_22271,N_21891);
and U22581 (N_22581,N_21894,N_22062);
or U22582 (N_22582,N_22221,N_22428);
nand U22583 (N_22583,N_22127,N_22481);
nand U22584 (N_22584,N_22347,N_21950);
nor U22585 (N_22585,N_21921,N_22262);
nor U22586 (N_22586,N_22463,N_21879);
and U22587 (N_22587,N_22451,N_22203);
nand U22588 (N_22588,N_21965,N_22482);
nand U22589 (N_22589,N_22138,N_22122);
nand U22590 (N_22590,N_22376,N_22018);
and U22591 (N_22591,N_21970,N_21898);
nand U22592 (N_22592,N_22311,N_22316);
and U22593 (N_22593,N_22145,N_22370);
xnor U22594 (N_22594,N_22025,N_22241);
and U22595 (N_22595,N_22397,N_22382);
or U22596 (N_22596,N_22073,N_22454);
and U22597 (N_22597,N_22364,N_22053);
and U22598 (N_22598,N_22393,N_22087);
xnor U22599 (N_22599,N_21942,N_22288);
nand U22600 (N_22600,N_21949,N_22294);
nor U22601 (N_22601,N_22297,N_22434);
xor U22602 (N_22602,N_22004,N_22493);
or U22603 (N_22603,N_22065,N_22289);
or U22604 (N_22604,N_22247,N_22054);
or U22605 (N_22605,N_21880,N_22076);
xor U22606 (N_22606,N_21982,N_21926);
or U22607 (N_22607,N_22315,N_22438);
and U22608 (N_22608,N_21927,N_21996);
xnor U22609 (N_22609,N_22398,N_22388);
nand U22610 (N_22610,N_21964,N_22309);
and U22611 (N_22611,N_22431,N_22016);
or U22612 (N_22612,N_22484,N_22371);
or U22613 (N_22613,N_22121,N_21992);
nand U22614 (N_22614,N_22325,N_22109);
nor U22615 (N_22615,N_22108,N_22495);
xnor U22616 (N_22616,N_22171,N_22013);
or U22617 (N_22617,N_22001,N_22306);
nand U22618 (N_22618,N_22471,N_22126);
xor U22619 (N_22619,N_22101,N_21947);
and U22620 (N_22620,N_22469,N_22421);
or U22621 (N_22621,N_22212,N_22024);
or U22622 (N_22622,N_22223,N_22057);
nor U22623 (N_22623,N_21958,N_22396);
nor U22624 (N_22624,N_22478,N_22060);
and U22625 (N_22625,N_22310,N_22067);
nor U22626 (N_22626,N_22425,N_22326);
xnor U22627 (N_22627,N_22343,N_21956);
nand U22628 (N_22628,N_22228,N_22468);
xnor U22629 (N_22629,N_22312,N_21906);
xor U22630 (N_22630,N_22250,N_22080);
nor U22631 (N_22631,N_22039,N_21948);
nand U22632 (N_22632,N_22227,N_22372);
and U22633 (N_22633,N_21997,N_22346);
nand U22634 (N_22634,N_22339,N_21923);
nor U22635 (N_22635,N_22209,N_22488);
xnor U22636 (N_22636,N_22099,N_22264);
or U22637 (N_22637,N_22093,N_21875);
xnor U22638 (N_22638,N_22005,N_22082);
nand U22639 (N_22639,N_22281,N_22446);
and U22640 (N_22640,N_22217,N_22220);
nand U22641 (N_22641,N_22187,N_21899);
xor U22642 (N_22642,N_22402,N_22218);
nor U22643 (N_22643,N_22427,N_22105);
nand U22644 (N_22644,N_22185,N_21886);
or U22645 (N_22645,N_22059,N_22386);
nand U22646 (N_22646,N_22313,N_21883);
xnor U22647 (N_22647,N_22474,N_22433);
nand U22648 (N_22648,N_22300,N_22328);
nor U22649 (N_22649,N_22034,N_22173);
and U22650 (N_22650,N_22117,N_22327);
nor U22651 (N_22651,N_22137,N_22473);
or U22652 (N_22652,N_22038,N_22012);
nor U22653 (N_22653,N_21930,N_22175);
and U22654 (N_22654,N_22414,N_22276);
nand U22655 (N_22655,N_22267,N_21972);
or U22656 (N_22656,N_21922,N_22307);
xor U22657 (N_22657,N_22413,N_22351);
or U22658 (N_22658,N_22051,N_21955);
xor U22659 (N_22659,N_22298,N_22091);
xnor U22660 (N_22660,N_22211,N_22222);
xnor U22661 (N_22661,N_21984,N_22003);
and U22662 (N_22662,N_22424,N_21994);
nor U22663 (N_22663,N_22071,N_22411);
or U22664 (N_22664,N_22010,N_22377);
nand U22665 (N_22665,N_22497,N_21983);
nor U22666 (N_22666,N_22070,N_22174);
nor U22667 (N_22667,N_22344,N_22305);
or U22668 (N_22668,N_22134,N_22296);
and U22669 (N_22669,N_21960,N_22321);
and U22670 (N_22670,N_22494,N_21901);
or U22671 (N_22671,N_21979,N_22234);
nand U22672 (N_22672,N_22041,N_22350);
xor U22673 (N_22673,N_22178,N_22144);
nor U22674 (N_22674,N_22329,N_22229);
nand U22675 (N_22675,N_22019,N_22066);
and U22676 (N_22676,N_22287,N_22366);
or U22677 (N_22677,N_21920,N_22238);
nand U22678 (N_22678,N_22192,N_22496);
and U22679 (N_22679,N_22213,N_22148);
xor U22680 (N_22680,N_21993,N_22284);
and U22681 (N_22681,N_21953,N_22201);
or U22682 (N_22682,N_22266,N_21884);
or U22683 (N_22683,N_22081,N_22200);
or U22684 (N_22684,N_22188,N_22031);
nand U22685 (N_22685,N_21957,N_22332);
nand U22686 (N_22686,N_22323,N_22319);
or U22687 (N_22687,N_22182,N_21913);
and U22688 (N_22688,N_22089,N_22061);
nor U22689 (N_22689,N_22042,N_22295);
nand U22690 (N_22690,N_22214,N_22450);
and U22691 (N_22691,N_22418,N_22394);
xnor U22692 (N_22692,N_22141,N_22196);
nor U22693 (N_22693,N_22189,N_22068);
and U22694 (N_22694,N_22466,N_21916);
xor U22695 (N_22695,N_21931,N_22023);
and U22696 (N_22696,N_22293,N_22170);
and U22697 (N_22697,N_21939,N_22462);
nor U22698 (N_22698,N_22280,N_22292);
or U22699 (N_22699,N_22430,N_22314);
xnor U22700 (N_22700,N_22483,N_21973);
and U22701 (N_22701,N_22453,N_22405);
nor U22702 (N_22702,N_22190,N_22006);
nor U22703 (N_22703,N_22248,N_22358);
xnor U22704 (N_22704,N_22149,N_22202);
xnor U22705 (N_22705,N_22331,N_22404);
nor U22706 (N_22706,N_21876,N_22072);
or U22707 (N_22707,N_22156,N_22111);
and U22708 (N_22708,N_22120,N_22069);
and U22709 (N_22709,N_22088,N_22172);
nor U22710 (N_22710,N_22458,N_22490);
xor U22711 (N_22711,N_22129,N_22362);
nor U22712 (N_22712,N_21975,N_22159);
nand U22713 (N_22713,N_22097,N_22355);
and U22714 (N_22714,N_22368,N_22215);
nand U22715 (N_22715,N_22063,N_21954);
and U22716 (N_22716,N_22027,N_22176);
or U22717 (N_22717,N_22043,N_21877);
or U22718 (N_22718,N_22251,N_22435);
and U22719 (N_22719,N_22291,N_22275);
or U22720 (N_22720,N_22191,N_21936);
xor U22721 (N_22721,N_22392,N_22322);
nand U22722 (N_22722,N_22318,N_22074);
nor U22723 (N_22723,N_22161,N_22058);
or U22724 (N_22724,N_21889,N_22078);
and U22725 (N_22725,N_22077,N_22461);
and U22726 (N_22726,N_22480,N_22242);
and U22727 (N_22727,N_22007,N_22124);
nor U22728 (N_22728,N_21938,N_22181);
or U22729 (N_22729,N_22282,N_22455);
and U22730 (N_22730,N_22422,N_22014);
xor U22731 (N_22731,N_22153,N_21978);
xnor U22732 (N_22732,N_22009,N_22487);
or U22733 (N_22733,N_22047,N_22049);
xnor U22734 (N_22734,N_22385,N_21925);
and U22735 (N_22735,N_22476,N_21917);
or U22736 (N_22736,N_22033,N_22416);
xnor U22737 (N_22737,N_21888,N_22408);
and U22738 (N_22738,N_22417,N_22154);
nor U22739 (N_22739,N_22367,N_22449);
and U22740 (N_22740,N_22046,N_21878);
xor U22741 (N_22741,N_22290,N_22103);
and U22742 (N_22742,N_21932,N_22302);
or U22743 (N_22743,N_21893,N_22259);
or U22744 (N_22744,N_21967,N_22096);
xor U22745 (N_22745,N_22028,N_22465);
nor U22746 (N_22746,N_22131,N_22151);
and U22747 (N_22747,N_22320,N_22345);
nand U22748 (N_22748,N_21914,N_22336);
and U22749 (N_22749,N_22055,N_22399);
nor U22750 (N_22750,N_22477,N_22083);
xor U22751 (N_22751,N_21995,N_22162);
nor U22752 (N_22752,N_22184,N_22110);
and U22753 (N_22753,N_21966,N_22165);
and U22754 (N_22754,N_22132,N_22232);
or U22755 (N_22755,N_22277,N_22135);
nand U22756 (N_22756,N_22436,N_22045);
xor U22757 (N_22757,N_21951,N_22342);
xnor U22758 (N_22758,N_22330,N_21928);
and U22759 (N_22759,N_22115,N_22403);
nand U22760 (N_22760,N_22374,N_22075);
nor U22761 (N_22761,N_21941,N_22021);
nor U22762 (N_22762,N_22168,N_22412);
nor U22763 (N_22763,N_22219,N_22084);
xnor U22764 (N_22764,N_21991,N_21999);
or U22765 (N_22765,N_22359,N_22204);
nor U22766 (N_22766,N_22278,N_22026);
nor U22767 (N_22767,N_22299,N_22283);
nand U22768 (N_22768,N_21892,N_22426);
nor U22769 (N_22769,N_22198,N_21904);
or U22770 (N_22770,N_22467,N_22341);
xor U22771 (N_22771,N_22423,N_21989);
nor U22772 (N_22772,N_22363,N_21895);
or U22773 (N_22773,N_21987,N_22432);
nor U22774 (N_22774,N_22258,N_22401);
xnor U22775 (N_22775,N_22207,N_22090);
and U22776 (N_22776,N_22308,N_22324);
nand U22777 (N_22777,N_22443,N_22452);
nor U22778 (N_22778,N_22472,N_21969);
nor U22779 (N_22779,N_22195,N_22400);
xnor U22780 (N_22780,N_22000,N_21902);
or U22781 (N_22781,N_22470,N_22240);
and U22782 (N_22782,N_22420,N_21952);
or U22783 (N_22783,N_22235,N_21981);
and U22784 (N_22784,N_22164,N_22303);
or U22785 (N_22785,N_22008,N_21934);
and U22786 (N_22786,N_21977,N_22157);
and U22787 (N_22787,N_22489,N_22146);
nand U22788 (N_22788,N_22381,N_21986);
or U22789 (N_22789,N_22375,N_21943);
nor U22790 (N_22790,N_22360,N_22104);
nand U22791 (N_22791,N_22011,N_21900);
nor U22792 (N_22792,N_22260,N_21919);
nor U22793 (N_22793,N_22254,N_22064);
nor U22794 (N_22794,N_22441,N_22158);
nand U22795 (N_22795,N_22349,N_22357);
nor U22796 (N_22796,N_22177,N_22407);
nand U22797 (N_22797,N_22269,N_22390);
nor U22798 (N_22798,N_21897,N_21924);
xnor U22799 (N_22799,N_22029,N_22373);
or U22800 (N_22800,N_22194,N_22301);
nand U22801 (N_22801,N_22116,N_21890);
nor U22802 (N_22802,N_22361,N_21944);
or U22803 (N_22803,N_22092,N_22150);
or U22804 (N_22804,N_22230,N_21974);
nand U22805 (N_22805,N_22160,N_22335);
nor U22806 (N_22806,N_22216,N_22125);
nor U22807 (N_22807,N_22256,N_22429);
nand U22808 (N_22808,N_22304,N_22210);
nor U22809 (N_22809,N_22491,N_22274);
nor U22810 (N_22810,N_21911,N_21903);
and U22811 (N_22811,N_22044,N_22448);
nand U22812 (N_22812,N_22334,N_22238);
and U22813 (N_22813,N_21997,N_22042);
or U22814 (N_22814,N_21909,N_22415);
xor U22815 (N_22815,N_22136,N_22287);
nand U22816 (N_22816,N_21943,N_22231);
xor U22817 (N_22817,N_22220,N_22131);
nand U22818 (N_22818,N_21959,N_21909);
and U22819 (N_22819,N_22047,N_22106);
nor U22820 (N_22820,N_22459,N_22409);
and U22821 (N_22821,N_21910,N_22261);
nor U22822 (N_22822,N_22340,N_22036);
nor U22823 (N_22823,N_21967,N_22074);
xor U22824 (N_22824,N_22063,N_22091);
nor U22825 (N_22825,N_22075,N_22313);
nand U22826 (N_22826,N_22327,N_22061);
nand U22827 (N_22827,N_22271,N_22030);
xor U22828 (N_22828,N_22367,N_21886);
nand U22829 (N_22829,N_21940,N_22237);
nor U22830 (N_22830,N_22043,N_22110);
or U22831 (N_22831,N_22462,N_22059);
or U22832 (N_22832,N_21999,N_22069);
and U22833 (N_22833,N_21913,N_22100);
xor U22834 (N_22834,N_21994,N_21887);
nor U22835 (N_22835,N_22311,N_22182);
and U22836 (N_22836,N_22077,N_22478);
xor U22837 (N_22837,N_21987,N_22307);
xor U22838 (N_22838,N_22101,N_22262);
nor U22839 (N_22839,N_22221,N_22258);
nor U22840 (N_22840,N_22414,N_22010);
and U22841 (N_22841,N_22232,N_21994);
and U22842 (N_22842,N_22147,N_22312);
nand U22843 (N_22843,N_22405,N_22485);
nand U22844 (N_22844,N_21888,N_22288);
or U22845 (N_22845,N_21993,N_22338);
xnor U22846 (N_22846,N_22457,N_22369);
or U22847 (N_22847,N_22415,N_22335);
and U22848 (N_22848,N_22488,N_21978);
nor U22849 (N_22849,N_22195,N_22365);
or U22850 (N_22850,N_22293,N_22234);
nor U22851 (N_22851,N_22419,N_22257);
nand U22852 (N_22852,N_22198,N_21876);
nor U22853 (N_22853,N_22145,N_22419);
or U22854 (N_22854,N_21948,N_22166);
xor U22855 (N_22855,N_21885,N_22265);
nand U22856 (N_22856,N_22008,N_22293);
or U22857 (N_22857,N_21988,N_21962);
nor U22858 (N_22858,N_22260,N_22200);
or U22859 (N_22859,N_21973,N_22148);
xnor U22860 (N_22860,N_21925,N_21946);
or U22861 (N_22861,N_22412,N_22149);
and U22862 (N_22862,N_21987,N_22237);
xor U22863 (N_22863,N_22019,N_22458);
or U22864 (N_22864,N_22109,N_22189);
or U22865 (N_22865,N_22417,N_22127);
nand U22866 (N_22866,N_22000,N_22276);
or U22867 (N_22867,N_21994,N_22281);
xor U22868 (N_22868,N_21970,N_22111);
or U22869 (N_22869,N_22433,N_22352);
and U22870 (N_22870,N_22447,N_22070);
nand U22871 (N_22871,N_22320,N_22226);
xor U22872 (N_22872,N_22446,N_22278);
nand U22873 (N_22873,N_21911,N_22247);
xor U22874 (N_22874,N_21879,N_22198);
and U22875 (N_22875,N_22396,N_21976);
nand U22876 (N_22876,N_22160,N_22071);
xnor U22877 (N_22877,N_22226,N_22382);
and U22878 (N_22878,N_22109,N_21896);
nand U22879 (N_22879,N_21951,N_22257);
nor U22880 (N_22880,N_22207,N_22105);
and U22881 (N_22881,N_22298,N_22164);
and U22882 (N_22882,N_22108,N_22368);
xor U22883 (N_22883,N_21908,N_21996);
nor U22884 (N_22884,N_22175,N_22099);
or U22885 (N_22885,N_22114,N_22207);
nor U22886 (N_22886,N_22251,N_21885);
nand U22887 (N_22887,N_22071,N_22193);
xor U22888 (N_22888,N_22186,N_22036);
xor U22889 (N_22889,N_21916,N_22196);
nor U22890 (N_22890,N_21891,N_21959);
nand U22891 (N_22891,N_22324,N_22439);
xnor U22892 (N_22892,N_22167,N_22182);
and U22893 (N_22893,N_22390,N_22210);
xor U22894 (N_22894,N_21923,N_22195);
or U22895 (N_22895,N_22007,N_21995);
or U22896 (N_22896,N_22154,N_22248);
nor U22897 (N_22897,N_22164,N_22458);
and U22898 (N_22898,N_21890,N_21905);
xnor U22899 (N_22899,N_22274,N_22392);
and U22900 (N_22900,N_22039,N_22116);
nor U22901 (N_22901,N_22397,N_21899);
and U22902 (N_22902,N_22353,N_22410);
and U22903 (N_22903,N_21992,N_22347);
or U22904 (N_22904,N_22064,N_22440);
nand U22905 (N_22905,N_22487,N_22422);
or U22906 (N_22906,N_22384,N_22205);
or U22907 (N_22907,N_21958,N_22496);
nor U22908 (N_22908,N_22315,N_22066);
nand U22909 (N_22909,N_22394,N_22496);
nor U22910 (N_22910,N_22235,N_22445);
or U22911 (N_22911,N_21883,N_21925);
xor U22912 (N_22912,N_22236,N_22482);
nand U22913 (N_22913,N_22433,N_21939);
and U22914 (N_22914,N_22345,N_22066);
or U22915 (N_22915,N_22470,N_22405);
and U22916 (N_22916,N_22051,N_21988);
and U22917 (N_22917,N_22292,N_22152);
nor U22918 (N_22918,N_22361,N_22121);
xor U22919 (N_22919,N_22180,N_22080);
nand U22920 (N_22920,N_22245,N_21912);
nand U22921 (N_22921,N_22084,N_22498);
and U22922 (N_22922,N_22195,N_22359);
xnor U22923 (N_22923,N_22388,N_22114);
and U22924 (N_22924,N_22286,N_21933);
or U22925 (N_22925,N_22167,N_22328);
and U22926 (N_22926,N_21966,N_22247);
nor U22927 (N_22927,N_22147,N_22075);
nor U22928 (N_22928,N_22289,N_22195);
xnor U22929 (N_22929,N_21915,N_21965);
and U22930 (N_22930,N_22473,N_22395);
and U22931 (N_22931,N_22459,N_22424);
nand U22932 (N_22932,N_22406,N_22362);
nor U22933 (N_22933,N_22230,N_21905);
xnor U22934 (N_22934,N_22257,N_22328);
or U22935 (N_22935,N_22078,N_21944);
nand U22936 (N_22936,N_21958,N_22348);
or U22937 (N_22937,N_22423,N_21875);
nand U22938 (N_22938,N_21946,N_22394);
nor U22939 (N_22939,N_22046,N_22070);
nor U22940 (N_22940,N_22360,N_22382);
xor U22941 (N_22941,N_22457,N_22079);
or U22942 (N_22942,N_22221,N_22324);
nor U22943 (N_22943,N_21944,N_22449);
and U22944 (N_22944,N_22051,N_21929);
xor U22945 (N_22945,N_21957,N_22288);
nor U22946 (N_22946,N_22096,N_22450);
or U22947 (N_22947,N_22380,N_22281);
xor U22948 (N_22948,N_22412,N_22300);
or U22949 (N_22949,N_21967,N_22060);
or U22950 (N_22950,N_21936,N_22188);
and U22951 (N_22951,N_22369,N_22040);
nand U22952 (N_22952,N_22158,N_22281);
nor U22953 (N_22953,N_22497,N_21974);
and U22954 (N_22954,N_22110,N_22020);
and U22955 (N_22955,N_21971,N_22335);
or U22956 (N_22956,N_22116,N_22499);
or U22957 (N_22957,N_22057,N_22306);
nand U22958 (N_22958,N_22362,N_22233);
nand U22959 (N_22959,N_22360,N_22448);
xnor U22960 (N_22960,N_22383,N_22003);
nand U22961 (N_22961,N_22444,N_22144);
nand U22962 (N_22962,N_21976,N_22441);
nor U22963 (N_22963,N_22403,N_22318);
nor U22964 (N_22964,N_22092,N_22224);
and U22965 (N_22965,N_21890,N_22429);
nor U22966 (N_22966,N_22329,N_21877);
and U22967 (N_22967,N_21934,N_22076);
or U22968 (N_22968,N_22442,N_22084);
xor U22969 (N_22969,N_22429,N_22205);
nor U22970 (N_22970,N_22453,N_22322);
and U22971 (N_22971,N_22401,N_22438);
and U22972 (N_22972,N_22027,N_22376);
nand U22973 (N_22973,N_22407,N_22365);
nor U22974 (N_22974,N_22214,N_22157);
and U22975 (N_22975,N_22003,N_22433);
or U22976 (N_22976,N_22475,N_22056);
nand U22977 (N_22977,N_22180,N_22194);
or U22978 (N_22978,N_22489,N_22437);
nand U22979 (N_22979,N_22271,N_22415);
and U22980 (N_22980,N_22057,N_22309);
nor U22981 (N_22981,N_22118,N_22499);
nor U22982 (N_22982,N_22320,N_22044);
or U22983 (N_22983,N_22273,N_21999);
or U22984 (N_22984,N_22421,N_22361);
nor U22985 (N_22985,N_22037,N_21900);
or U22986 (N_22986,N_22497,N_21967);
or U22987 (N_22987,N_22355,N_22233);
nand U22988 (N_22988,N_22065,N_22495);
nand U22989 (N_22989,N_21970,N_21884);
nor U22990 (N_22990,N_22394,N_22427);
and U22991 (N_22991,N_22190,N_21982);
nor U22992 (N_22992,N_21971,N_22471);
nand U22993 (N_22993,N_22288,N_22074);
and U22994 (N_22994,N_22063,N_22492);
nand U22995 (N_22995,N_22408,N_22358);
xnor U22996 (N_22996,N_21907,N_22143);
nand U22997 (N_22997,N_22074,N_22207);
nor U22998 (N_22998,N_22124,N_22126);
xor U22999 (N_22999,N_21913,N_22029);
nand U23000 (N_23000,N_22097,N_22222);
xnor U23001 (N_23001,N_22251,N_22227);
nor U23002 (N_23002,N_22103,N_21888);
xor U23003 (N_23003,N_21970,N_22089);
or U23004 (N_23004,N_22329,N_22287);
nand U23005 (N_23005,N_22145,N_22329);
nand U23006 (N_23006,N_22265,N_22052);
nand U23007 (N_23007,N_21890,N_21878);
or U23008 (N_23008,N_22012,N_22130);
and U23009 (N_23009,N_22090,N_22395);
and U23010 (N_23010,N_22497,N_22266);
nand U23011 (N_23011,N_22203,N_21880);
nand U23012 (N_23012,N_22215,N_22039);
xnor U23013 (N_23013,N_22398,N_21926);
nor U23014 (N_23014,N_22077,N_22322);
and U23015 (N_23015,N_22319,N_21918);
nor U23016 (N_23016,N_21886,N_22328);
nor U23017 (N_23017,N_22458,N_22244);
or U23018 (N_23018,N_21963,N_22315);
xor U23019 (N_23019,N_22299,N_22373);
xor U23020 (N_23020,N_22007,N_22426);
nor U23021 (N_23021,N_22135,N_21937);
nand U23022 (N_23022,N_22340,N_21955);
or U23023 (N_23023,N_22268,N_22409);
xnor U23024 (N_23024,N_22250,N_22311);
and U23025 (N_23025,N_22451,N_22498);
nor U23026 (N_23026,N_22104,N_22439);
nand U23027 (N_23027,N_21984,N_21889);
or U23028 (N_23028,N_22470,N_22209);
and U23029 (N_23029,N_22181,N_22066);
and U23030 (N_23030,N_22381,N_21929);
nor U23031 (N_23031,N_22439,N_22042);
and U23032 (N_23032,N_22415,N_22481);
nor U23033 (N_23033,N_21918,N_22321);
and U23034 (N_23034,N_22024,N_22333);
xor U23035 (N_23035,N_22153,N_21882);
nor U23036 (N_23036,N_22390,N_22444);
nor U23037 (N_23037,N_21877,N_22317);
xnor U23038 (N_23038,N_22027,N_22076);
and U23039 (N_23039,N_22256,N_22086);
nor U23040 (N_23040,N_21878,N_22224);
nor U23041 (N_23041,N_22218,N_22244);
and U23042 (N_23042,N_22178,N_22465);
and U23043 (N_23043,N_22478,N_22297);
nor U23044 (N_23044,N_22445,N_22406);
xor U23045 (N_23045,N_21968,N_22036);
nor U23046 (N_23046,N_21959,N_22030);
and U23047 (N_23047,N_22415,N_22209);
xor U23048 (N_23048,N_22195,N_22184);
xnor U23049 (N_23049,N_22365,N_22198);
nand U23050 (N_23050,N_22307,N_22312);
nor U23051 (N_23051,N_22001,N_21923);
and U23052 (N_23052,N_21932,N_21912);
xor U23053 (N_23053,N_21990,N_22487);
and U23054 (N_23054,N_21971,N_22418);
nand U23055 (N_23055,N_22255,N_22247);
xor U23056 (N_23056,N_22090,N_22196);
nor U23057 (N_23057,N_22434,N_22305);
xnor U23058 (N_23058,N_22112,N_22126);
or U23059 (N_23059,N_22074,N_22393);
nand U23060 (N_23060,N_22175,N_21990);
nand U23061 (N_23061,N_22347,N_22064);
or U23062 (N_23062,N_22367,N_22267);
or U23063 (N_23063,N_22158,N_22056);
or U23064 (N_23064,N_22199,N_22008);
nand U23065 (N_23065,N_21911,N_21917);
and U23066 (N_23066,N_22181,N_21964);
and U23067 (N_23067,N_22062,N_22432);
xnor U23068 (N_23068,N_22109,N_22192);
and U23069 (N_23069,N_22023,N_21892);
and U23070 (N_23070,N_22172,N_22348);
nor U23071 (N_23071,N_22481,N_21937);
nand U23072 (N_23072,N_22166,N_22329);
nor U23073 (N_23073,N_21937,N_22006);
xor U23074 (N_23074,N_22121,N_22062);
xor U23075 (N_23075,N_22475,N_22297);
and U23076 (N_23076,N_22118,N_22219);
and U23077 (N_23077,N_22358,N_21898);
or U23078 (N_23078,N_21972,N_22109);
nand U23079 (N_23079,N_21880,N_22265);
and U23080 (N_23080,N_22495,N_22481);
or U23081 (N_23081,N_22134,N_22054);
and U23082 (N_23082,N_21973,N_22323);
xor U23083 (N_23083,N_22445,N_21976);
or U23084 (N_23084,N_22383,N_22079);
nor U23085 (N_23085,N_21932,N_22172);
xnor U23086 (N_23086,N_22334,N_22104);
and U23087 (N_23087,N_21977,N_21936);
and U23088 (N_23088,N_22349,N_22334);
nor U23089 (N_23089,N_22217,N_21958);
nand U23090 (N_23090,N_22379,N_22446);
or U23091 (N_23091,N_22016,N_22354);
and U23092 (N_23092,N_22370,N_22285);
and U23093 (N_23093,N_22071,N_22163);
nand U23094 (N_23094,N_22359,N_22301);
xnor U23095 (N_23095,N_21928,N_21903);
nor U23096 (N_23096,N_22242,N_22304);
nor U23097 (N_23097,N_21912,N_22137);
or U23098 (N_23098,N_22215,N_21900);
and U23099 (N_23099,N_21898,N_22008);
xnor U23100 (N_23100,N_22191,N_22090);
xor U23101 (N_23101,N_21932,N_21939);
xnor U23102 (N_23102,N_22379,N_22035);
xnor U23103 (N_23103,N_22371,N_22473);
nand U23104 (N_23104,N_22021,N_21979);
nor U23105 (N_23105,N_22042,N_21909);
nor U23106 (N_23106,N_22153,N_21993);
and U23107 (N_23107,N_21882,N_22154);
nor U23108 (N_23108,N_22263,N_22014);
nor U23109 (N_23109,N_22259,N_22142);
nand U23110 (N_23110,N_22457,N_22055);
or U23111 (N_23111,N_21937,N_22222);
nor U23112 (N_23112,N_22178,N_22233);
and U23113 (N_23113,N_22382,N_22268);
or U23114 (N_23114,N_22328,N_22102);
nand U23115 (N_23115,N_22183,N_22055);
and U23116 (N_23116,N_22120,N_22117);
nand U23117 (N_23117,N_22152,N_21957);
xor U23118 (N_23118,N_22042,N_21947);
nand U23119 (N_23119,N_22250,N_22234);
or U23120 (N_23120,N_22264,N_22484);
xor U23121 (N_23121,N_22456,N_22122);
xor U23122 (N_23122,N_22157,N_22154);
xnor U23123 (N_23123,N_22094,N_22188);
nor U23124 (N_23124,N_22215,N_22343);
nand U23125 (N_23125,N_22764,N_22961);
or U23126 (N_23126,N_22878,N_22992);
and U23127 (N_23127,N_23111,N_22783);
xor U23128 (N_23128,N_22822,N_22780);
xnor U23129 (N_23129,N_22774,N_23005);
nand U23130 (N_23130,N_22545,N_22599);
or U23131 (N_23131,N_22862,N_23034);
nor U23132 (N_23132,N_22701,N_22768);
nor U23133 (N_23133,N_22657,N_22882);
and U23134 (N_23134,N_22567,N_22848);
nand U23135 (N_23135,N_22949,N_22631);
nor U23136 (N_23136,N_22855,N_22639);
nand U23137 (N_23137,N_22684,N_22864);
xnor U23138 (N_23138,N_22638,N_22614);
or U23139 (N_23139,N_22895,N_22813);
or U23140 (N_23140,N_22962,N_23049);
nor U23141 (N_23141,N_22620,N_22869);
nand U23142 (N_23142,N_23098,N_22951);
xnor U23143 (N_23143,N_23018,N_22630);
nor U23144 (N_23144,N_22668,N_23121);
nor U23145 (N_23145,N_22635,N_22849);
and U23146 (N_23146,N_22928,N_23031);
or U23147 (N_23147,N_22737,N_22640);
nor U23148 (N_23148,N_23024,N_22714);
nand U23149 (N_23149,N_23021,N_22659);
nor U23150 (N_23150,N_22814,N_22502);
or U23151 (N_23151,N_22979,N_22933);
and U23152 (N_23152,N_23080,N_22521);
nor U23153 (N_23153,N_22738,N_22691);
or U23154 (N_23154,N_22863,N_22528);
nor U23155 (N_23155,N_22850,N_22675);
xnor U23156 (N_23156,N_22903,N_22721);
and U23157 (N_23157,N_22572,N_22729);
nand U23158 (N_23158,N_22512,N_22840);
and U23159 (N_23159,N_22626,N_22503);
nand U23160 (N_23160,N_23051,N_22741);
or U23161 (N_23161,N_22999,N_22912);
nand U23162 (N_23162,N_22897,N_22777);
nand U23163 (N_23163,N_23085,N_22846);
xor U23164 (N_23164,N_22847,N_23017);
xnor U23165 (N_23165,N_22875,N_23022);
or U23166 (N_23166,N_22511,N_22666);
nor U23167 (N_23167,N_22637,N_22821);
nand U23168 (N_23168,N_22815,N_22947);
nor U23169 (N_23169,N_22651,N_22676);
nand U23170 (N_23170,N_22720,N_23083);
nand U23171 (N_23171,N_22942,N_22660);
xor U23172 (N_23172,N_22911,N_22574);
nor U23173 (N_23173,N_22619,N_22835);
xnor U23174 (N_23174,N_22766,N_22562);
or U23175 (N_23175,N_23073,N_22818);
and U23176 (N_23176,N_22510,N_23055);
nor U23177 (N_23177,N_22833,N_22736);
and U23178 (N_23178,N_23029,N_22885);
nand U23179 (N_23179,N_22871,N_22703);
or U23180 (N_23180,N_22646,N_22981);
nor U23181 (N_23181,N_22756,N_22532);
nand U23182 (N_23182,N_22585,N_23060);
nor U23183 (N_23183,N_22605,N_22792);
xnor U23184 (N_23184,N_23047,N_23107);
nor U23185 (N_23185,N_22834,N_22582);
and U23186 (N_23186,N_22530,N_23000);
xor U23187 (N_23187,N_22806,N_22529);
xnor U23188 (N_23188,N_22609,N_22658);
or U23189 (N_23189,N_23050,N_22986);
or U23190 (N_23190,N_22553,N_22556);
or U23191 (N_23191,N_22724,N_22971);
nand U23192 (N_23192,N_23009,N_22604);
and U23193 (N_23193,N_22851,N_23008);
or U23194 (N_23194,N_22518,N_23002);
and U23195 (N_23195,N_22622,N_22679);
nor U23196 (N_23196,N_23095,N_23099);
nor U23197 (N_23197,N_23056,N_23109);
nand U23198 (N_23198,N_23052,N_22857);
nand U23199 (N_23199,N_22688,N_22742);
or U23200 (N_23200,N_22612,N_22515);
and U23201 (N_23201,N_22994,N_23065);
and U23202 (N_23202,N_23067,N_22970);
nand U23203 (N_23203,N_22763,N_22647);
nand U23204 (N_23204,N_23001,N_23043);
or U23205 (N_23205,N_22606,N_22893);
or U23206 (N_23206,N_22925,N_22704);
and U23207 (N_23207,N_22946,N_22583);
nor U23208 (N_23208,N_22985,N_22648);
nor U23209 (N_23209,N_22727,N_22656);
and U23210 (N_23210,N_22753,N_22759);
xor U23211 (N_23211,N_22577,N_23069);
and U23212 (N_23212,N_22514,N_22811);
and U23213 (N_23213,N_23087,N_22906);
nand U23214 (N_23214,N_22953,N_22501);
xnor U23215 (N_23215,N_22749,N_22803);
xor U23216 (N_23216,N_22866,N_22570);
and U23217 (N_23217,N_22988,N_22578);
nor U23218 (N_23218,N_22709,N_22899);
or U23219 (N_23219,N_22695,N_22743);
and U23220 (N_23220,N_23011,N_22719);
and U23221 (N_23221,N_22938,N_22837);
xor U23222 (N_23222,N_22670,N_22602);
nor U23223 (N_23223,N_22819,N_22687);
and U23224 (N_23224,N_22500,N_23062);
xnor U23225 (N_23225,N_22752,N_23036);
nor U23226 (N_23226,N_22723,N_22597);
xor U23227 (N_23227,N_22625,N_22809);
or U23228 (N_23228,N_22615,N_22686);
xnor U23229 (N_23229,N_22603,N_23079);
xor U23230 (N_23230,N_22950,N_22798);
xnor U23231 (N_23231,N_22607,N_23023);
nand U23232 (N_23232,N_22836,N_22760);
and U23233 (N_23233,N_23032,N_22653);
nor U23234 (N_23234,N_22881,N_22782);
xnor U23235 (N_23235,N_22748,N_23071);
nand U23236 (N_23236,N_23072,N_22513);
nor U23237 (N_23237,N_22969,N_22544);
xnor U23238 (N_23238,N_23033,N_22824);
or U23239 (N_23239,N_22516,N_23110);
or U23240 (N_23240,N_23119,N_22931);
nor U23241 (N_23241,N_22506,N_22998);
nand U23242 (N_23242,N_22698,N_22692);
nor U23243 (N_23243,N_22874,N_22726);
or U23244 (N_23244,N_22730,N_22769);
or U23245 (N_23245,N_22802,N_22968);
nand U23246 (N_23246,N_22877,N_22735);
nand U23247 (N_23247,N_23088,N_22804);
and U23248 (N_23248,N_22523,N_22989);
nand U23249 (N_23249,N_22682,N_22601);
xnor U23250 (N_23250,N_22667,N_22873);
xor U23251 (N_23251,N_22636,N_22964);
xor U23252 (N_23252,N_23089,N_22770);
nor U23253 (N_23253,N_22681,N_22563);
xnor U23254 (N_23254,N_22936,N_22919);
and U23255 (N_23255,N_22592,N_22860);
and U23256 (N_23256,N_22901,N_22547);
nand U23257 (N_23257,N_22984,N_22879);
nand U23258 (N_23258,N_23063,N_22554);
xor U23259 (N_23259,N_23038,N_22587);
nand U23260 (N_23260,N_22654,N_22993);
nor U23261 (N_23261,N_22916,N_22926);
nand U23262 (N_23262,N_23101,N_22765);
nand U23263 (N_23263,N_22568,N_22652);
nor U23264 (N_23264,N_22894,N_22904);
nor U23265 (N_23265,N_23113,N_23010);
xor U23266 (N_23266,N_22954,N_22801);
nand U23267 (N_23267,N_22627,N_22799);
nor U23268 (N_23268,N_23124,N_22883);
or U23269 (N_23269,N_22787,N_22633);
nand U23270 (N_23270,N_22586,N_22948);
or U23271 (N_23271,N_22642,N_22543);
xor U23272 (N_23272,N_22886,N_22566);
xor U23273 (N_23273,N_23070,N_22845);
or U23274 (N_23274,N_22808,N_22584);
nor U23275 (N_23275,N_22996,N_22565);
nand U23276 (N_23276,N_23102,N_22838);
nor U23277 (N_23277,N_22579,N_22623);
xnor U23278 (N_23278,N_22941,N_23003);
nand U23279 (N_23279,N_22527,N_22778);
xor U23280 (N_23280,N_22621,N_22910);
and U23281 (N_23281,N_22940,N_22535);
xnor U23282 (N_23282,N_22674,N_23091);
nor U23283 (N_23283,N_22772,N_23082);
xnor U23284 (N_23284,N_23075,N_23120);
or U23285 (N_23285,N_23027,N_22891);
and U23286 (N_23286,N_22932,N_23118);
xor U23287 (N_23287,N_22974,N_23015);
or U23288 (N_23288,N_22796,N_22945);
or U23289 (N_23289,N_22861,N_22745);
and U23290 (N_23290,N_23092,N_22927);
nand U23291 (N_23291,N_22693,N_22569);
nand U23292 (N_23292,N_22533,N_22805);
and U23293 (N_23293,N_22575,N_23025);
nor U23294 (N_23294,N_22930,N_22816);
or U23295 (N_23295,N_23007,N_22876);
and U23296 (N_23296,N_22732,N_22618);
nor U23297 (N_23297,N_22677,N_22694);
or U23298 (N_23298,N_22747,N_22757);
nor U23299 (N_23299,N_22784,N_23046);
and U23300 (N_23300,N_22596,N_23123);
and U23301 (N_23301,N_22800,N_22924);
nand U23302 (N_23302,N_22794,N_22617);
and U23303 (N_23303,N_23028,N_22669);
nand U23304 (N_23304,N_22963,N_22884);
nand U23305 (N_23305,N_22957,N_22710);
or U23306 (N_23306,N_22826,N_23016);
and U23307 (N_23307,N_22571,N_22853);
xnor U23308 (N_23308,N_22519,N_23026);
nor U23309 (N_23309,N_22507,N_22624);
or U23310 (N_23310,N_22991,N_23053);
xor U23311 (N_23311,N_22921,N_22581);
or U23312 (N_23312,N_22972,N_22718);
nand U23313 (N_23313,N_23012,N_22744);
nand U23314 (N_23314,N_22995,N_22913);
nor U23315 (N_23315,N_22751,N_22929);
or U23316 (N_23316,N_22868,N_22634);
nor U23317 (N_23317,N_22823,N_23006);
and U23318 (N_23318,N_22702,N_23112);
nand U23319 (N_23319,N_22797,N_22920);
xnor U23320 (N_23320,N_23103,N_22917);
nand U23321 (N_23321,N_23077,N_22958);
xnor U23322 (N_23322,N_22600,N_22943);
xor U23323 (N_23323,N_22705,N_22825);
or U23324 (N_23324,N_22790,N_22548);
or U23325 (N_23325,N_22914,N_22546);
nor U23326 (N_23326,N_22965,N_22959);
nor U23327 (N_23327,N_22740,N_22611);
nor U23328 (N_23328,N_23100,N_22576);
or U23329 (N_23329,N_22696,N_22508);
or U23330 (N_23330,N_22762,N_22561);
nand U23331 (N_23331,N_23048,N_23044);
and U23332 (N_23332,N_22595,N_22700);
nor U23333 (N_23333,N_22807,N_22629);
and U23334 (N_23334,N_22645,N_23106);
xnor U23335 (N_23335,N_22831,N_22593);
nor U23336 (N_23336,N_22937,N_23004);
and U23337 (N_23337,N_22865,N_22854);
nand U23338 (N_23338,N_22504,N_22632);
xor U23339 (N_23339,N_22536,N_22649);
xnor U23340 (N_23340,N_22758,N_23066);
nand U23341 (N_23341,N_23097,N_22733);
and U23342 (N_23342,N_22786,N_22555);
nor U23343 (N_23343,N_22673,N_22839);
nor U23344 (N_23344,N_22746,N_23081);
nand U23345 (N_23345,N_22557,N_22525);
nor U23346 (N_23346,N_22842,N_22902);
or U23347 (N_23347,N_23094,N_22734);
or U23348 (N_23348,N_22793,N_23054);
or U23349 (N_23349,N_22598,N_22697);
and U23350 (N_23350,N_22767,N_23104);
and U23351 (N_23351,N_22779,N_22580);
or U23352 (N_23352,N_22559,N_22685);
and U23353 (N_23353,N_23039,N_22708);
xnor U23354 (N_23354,N_22680,N_22731);
and U23355 (N_23355,N_22956,N_22594);
xnor U23356 (N_23356,N_22689,N_23030);
or U23357 (N_23357,N_22856,N_22852);
and U23358 (N_23358,N_22655,N_22699);
or U23359 (N_23359,N_23059,N_22978);
xor U23360 (N_23360,N_22832,N_22827);
or U23361 (N_23361,N_22858,N_23045);
nand U23362 (N_23362,N_22706,N_22939);
xnor U23363 (N_23363,N_22872,N_22564);
nor U23364 (N_23364,N_22795,N_22997);
nand U23365 (N_23365,N_22717,N_22542);
nand U23366 (N_23366,N_22712,N_22841);
and U23367 (N_23367,N_23064,N_23013);
nand U23368 (N_23368,N_22890,N_22810);
nand U23369 (N_23369,N_23040,N_22952);
nor U23370 (N_23370,N_23020,N_22641);
nand U23371 (N_23371,N_22664,N_23090);
nand U23372 (N_23372,N_22983,N_22761);
or U23373 (N_23373,N_22908,N_23108);
nand U23374 (N_23374,N_22867,N_22713);
nand U23375 (N_23375,N_22540,N_22610);
or U23376 (N_23376,N_22573,N_22663);
xnor U23377 (N_23377,N_22915,N_22889);
nor U23378 (N_23378,N_22892,N_22789);
nor U23379 (N_23379,N_22905,N_22613);
xor U23380 (N_23380,N_23061,N_23057);
and U23381 (N_23381,N_22975,N_22683);
xor U23382 (N_23382,N_22907,N_22980);
nand U23383 (N_23383,N_22773,N_22589);
xnor U23384 (N_23384,N_22628,N_22534);
and U23385 (N_23385,N_22538,N_23041);
nand U23386 (N_23386,N_22520,N_23105);
and U23387 (N_23387,N_22608,N_22900);
nor U23388 (N_23388,N_22661,N_22716);
nand U23389 (N_23389,N_22918,N_23096);
nor U23390 (N_23390,N_22524,N_22967);
xnor U23391 (N_23391,N_22830,N_22844);
nor U23392 (N_23392,N_22671,N_22588);
nor U23393 (N_23393,N_22955,N_23084);
nand U23394 (N_23394,N_22537,N_23014);
or U23395 (N_23395,N_22909,N_22672);
nand U23396 (N_23396,N_22552,N_22715);
or U23397 (N_23397,N_22750,N_22880);
and U23398 (N_23398,N_22888,N_22982);
and U23399 (N_23399,N_22690,N_22616);
and U23400 (N_23400,N_23086,N_22551);
xnor U23401 (N_23401,N_23076,N_22923);
nor U23402 (N_23402,N_22560,N_22990);
nor U23403 (N_23403,N_22812,N_22973);
nand U23404 (N_23404,N_22644,N_23037);
and U23405 (N_23405,N_22591,N_22776);
nand U23406 (N_23406,N_23122,N_23042);
and U23407 (N_23407,N_22590,N_22665);
xor U23408 (N_23408,N_23035,N_22785);
and U23409 (N_23409,N_22754,N_22817);
or U23410 (N_23410,N_22887,N_23058);
xor U23411 (N_23411,N_22859,N_22539);
and U23412 (N_23412,N_22505,N_22707);
nand U23413 (N_23413,N_22722,N_22987);
nand U23414 (N_23414,N_23068,N_23093);
and U23415 (N_23415,N_22788,N_22771);
nand U23416 (N_23416,N_22531,N_22791);
nand U23417 (N_23417,N_22898,N_22558);
xnor U23418 (N_23418,N_22820,N_22829);
or U23419 (N_23419,N_23074,N_22549);
nand U23420 (N_23420,N_22739,N_22643);
and U23421 (N_23421,N_22725,N_22550);
nand U23422 (N_23422,N_22944,N_22650);
nand U23423 (N_23423,N_22711,N_23116);
xnor U23424 (N_23424,N_22960,N_22755);
xnor U23425 (N_23425,N_22522,N_22935);
nor U23426 (N_23426,N_22509,N_22728);
or U23427 (N_23427,N_22828,N_23117);
nor U23428 (N_23428,N_22870,N_23114);
nor U23429 (N_23429,N_22843,N_22966);
and U23430 (N_23430,N_23019,N_22976);
or U23431 (N_23431,N_22922,N_22526);
xor U23432 (N_23432,N_23078,N_22977);
nor U23433 (N_23433,N_22896,N_22678);
nand U23434 (N_23434,N_22662,N_22775);
nor U23435 (N_23435,N_23115,N_22517);
or U23436 (N_23436,N_22781,N_22934);
xnor U23437 (N_23437,N_22541,N_22740);
or U23438 (N_23438,N_22528,N_22993);
and U23439 (N_23439,N_22784,N_22684);
and U23440 (N_23440,N_22588,N_22557);
nor U23441 (N_23441,N_22904,N_22848);
xnor U23442 (N_23442,N_22760,N_22983);
xnor U23443 (N_23443,N_22947,N_22544);
nor U23444 (N_23444,N_22626,N_22861);
and U23445 (N_23445,N_23064,N_22729);
xnor U23446 (N_23446,N_22866,N_23079);
xnor U23447 (N_23447,N_22763,N_22532);
xnor U23448 (N_23448,N_22664,N_22792);
and U23449 (N_23449,N_22645,N_22746);
nor U23450 (N_23450,N_23017,N_23092);
nand U23451 (N_23451,N_23044,N_22630);
or U23452 (N_23452,N_22894,N_22645);
and U23453 (N_23453,N_22916,N_22594);
xor U23454 (N_23454,N_22897,N_22835);
or U23455 (N_23455,N_22865,N_22701);
and U23456 (N_23456,N_22919,N_22754);
or U23457 (N_23457,N_22970,N_23111);
nor U23458 (N_23458,N_22791,N_22981);
or U23459 (N_23459,N_22863,N_22806);
nand U23460 (N_23460,N_22543,N_22916);
and U23461 (N_23461,N_22859,N_22872);
or U23462 (N_23462,N_22660,N_23088);
nand U23463 (N_23463,N_22815,N_22638);
nor U23464 (N_23464,N_22791,N_22932);
or U23465 (N_23465,N_22979,N_22994);
or U23466 (N_23466,N_22795,N_22755);
nand U23467 (N_23467,N_22500,N_23041);
and U23468 (N_23468,N_22641,N_23006);
and U23469 (N_23469,N_22578,N_22552);
or U23470 (N_23470,N_23005,N_23027);
nand U23471 (N_23471,N_22946,N_22616);
and U23472 (N_23472,N_22702,N_22571);
nor U23473 (N_23473,N_22531,N_22755);
xor U23474 (N_23474,N_22680,N_22733);
nor U23475 (N_23475,N_23047,N_22890);
nor U23476 (N_23476,N_23014,N_22741);
nand U23477 (N_23477,N_22845,N_22895);
xor U23478 (N_23478,N_23077,N_22699);
or U23479 (N_23479,N_23082,N_22545);
or U23480 (N_23480,N_22565,N_23123);
xnor U23481 (N_23481,N_22726,N_22621);
xor U23482 (N_23482,N_22611,N_23035);
or U23483 (N_23483,N_22794,N_22896);
xor U23484 (N_23484,N_23106,N_22835);
or U23485 (N_23485,N_22509,N_22802);
nand U23486 (N_23486,N_22656,N_23089);
and U23487 (N_23487,N_22849,N_22988);
xnor U23488 (N_23488,N_22991,N_22559);
or U23489 (N_23489,N_22754,N_23052);
nand U23490 (N_23490,N_22596,N_22693);
xnor U23491 (N_23491,N_23080,N_23101);
nor U23492 (N_23492,N_22616,N_23088);
nand U23493 (N_23493,N_22611,N_22990);
or U23494 (N_23494,N_23002,N_22843);
nand U23495 (N_23495,N_23112,N_22975);
nand U23496 (N_23496,N_22808,N_23050);
and U23497 (N_23497,N_23059,N_23018);
xor U23498 (N_23498,N_22628,N_22818);
xor U23499 (N_23499,N_22613,N_22956);
nor U23500 (N_23500,N_22876,N_22610);
and U23501 (N_23501,N_22917,N_22910);
or U23502 (N_23502,N_22508,N_22882);
nor U23503 (N_23503,N_22603,N_22813);
nor U23504 (N_23504,N_22923,N_23084);
nand U23505 (N_23505,N_22573,N_22967);
and U23506 (N_23506,N_22838,N_22556);
nand U23507 (N_23507,N_22662,N_22905);
or U23508 (N_23508,N_22512,N_22893);
or U23509 (N_23509,N_22920,N_23045);
xor U23510 (N_23510,N_23091,N_22898);
or U23511 (N_23511,N_22751,N_23113);
nand U23512 (N_23512,N_22658,N_23057);
and U23513 (N_23513,N_23006,N_22836);
nand U23514 (N_23514,N_23035,N_22667);
nor U23515 (N_23515,N_22856,N_22866);
xnor U23516 (N_23516,N_23034,N_22734);
and U23517 (N_23517,N_22513,N_23115);
nor U23518 (N_23518,N_22644,N_22646);
or U23519 (N_23519,N_22520,N_22704);
and U23520 (N_23520,N_22707,N_22982);
and U23521 (N_23521,N_22626,N_22694);
or U23522 (N_23522,N_23109,N_22560);
nor U23523 (N_23523,N_22995,N_22569);
or U23524 (N_23524,N_22500,N_22958);
and U23525 (N_23525,N_22918,N_23123);
and U23526 (N_23526,N_22696,N_22668);
or U23527 (N_23527,N_22981,N_22962);
xnor U23528 (N_23528,N_22801,N_22879);
and U23529 (N_23529,N_22755,N_23051);
nand U23530 (N_23530,N_23061,N_22874);
xnor U23531 (N_23531,N_23119,N_23073);
and U23532 (N_23532,N_22878,N_23045);
or U23533 (N_23533,N_22500,N_22534);
nand U23534 (N_23534,N_22693,N_22860);
or U23535 (N_23535,N_22984,N_23085);
nand U23536 (N_23536,N_22623,N_22829);
nand U23537 (N_23537,N_22652,N_22925);
xor U23538 (N_23538,N_22720,N_22579);
xor U23539 (N_23539,N_23070,N_23000);
or U23540 (N_23540,N_22849,N_23010);
nor U23541 (N_23541,N_22657,N_22970);
nand U23542 (N_23542,N_23044,N_22528);
nand U23543 (N_23543,N_23042,N_22969);
or U23544 (N_23544,N_22892,N_22900);
or U23545 (N_23545,N_22807,N_22691);
nor U23546 (N_23546,N_22792,N_22955);
xnor U23547 (N_23547,N_22802,N_22764);
nor U23548 (N_23548,N_22678,N_22792);
nand U23549 (N_23549,N_22665,N_22879);
xnor U23550 (N_23550,N_22781,N_22618);
or U23551 (N_23551,N_22873,N_22973);
nor U23552 (N_23552,N_22879,N_23020);
and U23553 (N_23553,N_22562,N_22789);
nor U23554 (N_23554,N_22699,N_22666);
nor U23555 (N_23555,N_22534,N_22604);
nand U23556 (N_23556,N_22709,N_22919);
nor U23557 (N_23557,N_22532,N_23026);
and U23558 (N_23558,N_22749,N_22699);
nor U23559 (N_23559,N_22607,N_22646);
xnor U23560 (N_23560,N_23072,N_23091);
nor U23561 (N_23561,N_22739,N_22967);
nand U23562 (N_23562,N_22878,N_22742);
or U23563 (N_23563,N_22647,N_23062);
or U23564 (N_23564,N_22526,N_22914);
and U23565 (N_23565,N_22886,N_22739);
nor U23566 (N_23566,N_22621,N_22798);
or U23567 (N_23567,N_23070,N_22684);
or U23568 (N_23568,N_22513,N_22577);
and U23569 (N_23569,N_23121,N_22786);
nand U23570 (N_23570,N_22523,N_22546);
xor U23571 (N_23571,N_22637,N_23097);
nor U23572 (N_23572,N_23058,N_22776);
or U23573 (N_23573,N_22848,N_22623);
nand U23574 (N_23574,N_23102,N_22976);
nor U23575 (N_23575,N_23103,N_23107);
nor U23576 (N_23576,N_23109,N_23048);
and U23577 (N_23577,N_22902,N_22698);
and U23578 (N_23578,N_22947,N_22710);
nand U23579 (N_23579,N_22972,N_22884);
nor U23580 (N_23580,N_22742,N_22736);
xor U23581 (N_23581,N_22550,N_22755);
or U23582 (N_23582,N_22619,N_23086);
xnor U23583 (N_23583,N_22577,N_22742);
and U23584 (N_23584,N_22537,N_22636);
xor U23585 (N_23585,N_22693,N_22852);
or U23586 (N_23586,N_22839,N_23021);
nor U23587 (N_23587,N_22926,N_22971);
and U23588 (N_23588,N_23055,N_22545);
and U23589 (N_23589,N_22767,N_22509);
or U23590 (N_23590,N_22604,N_22879);
or U23591 (N_23591,N_22542,N_22539);
nand U23592 (N_23592,N_22830,N_22774);
xor U23593 (N_23593,N_22611,N_22594);
nor U23594 (N_23594,N_22560,N_22937);
nor U23595 (N_23595,N_23011,N_23016);
and U23596 (N_23596,N_22945,N_22754);
and U23597 (N_23597,N_22987,N_22999);
or U23598 (N_23598,N_22846,N_22981);
nand U23599 (N_23599,N_22945,N_22925);
or U23600 (N_23600,N_22867,N_23087);
or U23601 (N_23601,N_22779,N_23118);
or U23602 (N_23602,N_22881,N_23066);
nor U23603 (N_23603,N_22594,N_22917);
and U23604 (N_23604,N_22895,N_22949);
and U23605 (N_23605,N_22648,N_22922);
and U23606 (N_23606,N_23086,N_22843);
nor U23607 (N_23607,N_22646,N_22690);
nor U23608 (N_23608,N_22941,N_22730);
and U23609 (N_23609,N_23011,N_22650);
xor U23610 (N_23610,N_22814,N_22797);
nand U23611 (N_23611,N_22798,N_23102);
nor U23612 (N_23612,N_22661,N_22562);
nor U23613 (N_23613,N_22909,N_22567);
and U23614 (N_23614,N_22944,N_22792);
and U23615 (N_23615,N_22646,N_22548);
nor U23616 (N_23616,N_22860,N_22617);
nand U23617 (N_23617,N_22650,N_23076);
nor U23618 (N_23618,N_22530,N_22581);
nor U23619 (N_23619,N_22625,N_22823);
or U23620 (N_23620,N_22799,N_22596);
or U23621 (N_23621,N_22892,N_22822);
nand U23622 (N_23622,N_22954,N_22669);
nor U23623 (N_23623,N_22680,N_22967);
nand U23624 (N_23624,N_22803,N_22559);
xnor U23625 (N_23625,N_22903,N_22677);
and U23626 (N_23626,N_22580,N_22656);
nor U23627 (N_23627,N_22833,N_22733);
xor U23628 (N_23628,N_22880,N_23099);
xnor U23629 (N_23629,N_22831,N_22729);
or U23630 (N_23630,N_22562,N_22947);
or U23631 (N_23631,N_22835,N_22669);
nand U23632 (N_23632,N_22974,N_22508);
or U23633 (N_23633,N_22552,N_22605);
nand U23634 (N_23634,N_22867,N_22775);
nor U23635 (N_23635,N_22983,N_22876);
and U23636 (N_23636,N_22925,N_22764);
or U23637 (N_23637,N_22979,N_22897);
or U23638 (N_23638,N_22719,N_22942);
xnor U23639 (N_23639,N_22834,N_22948);
and U23640 (N_23640,N_22970,N_22673);
nor U23641 (N_23641,N_22658,N_22738);
nand U23642 (N_23642,N_22709,N_22906);
nor U23643 (N_23643,N_22516,N_22882);
xor U23644 (N_23644,N_22642,N_22545);
xnor U23645 (N_23645,N_22652,N_22930);
nand U23646 (N_23646,N_22608,N_22684);
or U23647 (N_23647,N_22824,N_22936);
or U23648 (N_23648,N_22808,N_22839);
nor U23649 (N_23649,N_22589,N_23076);
nor U23650 (N_23650,N_22610,N_22869);
nor U23651 (N_23651,N_22527,N_22556);
and U23652 (N_23652,N_22924,N_23103);
or U23653 (N_23653,N_23098,N_22892);
or U23654 (N_23654,N_22955,N_22908);
nand U23655 (N_23655,N_23086,N_22698);
nor U23656 (N_23656,N_22827,N_23122);
nor U23657 (N_23657,N_22924,N_22597);
xor U23658 (N_23658,N_23011,N_22620);
nor U23659 (N_23659,N_22984,N_22938);
nor U23660 (N_23660,N_22560,N_22502);
nand U23661 (N_23661,N_22592,N_23123);
xor U23662 (N_23662,N_22951,N_22858);
and U23663 (N_23663,N_23021,N_22894);
nor U23664 (N_23664,N_22864,N_22925);
nor U23665 (N_23665,N_22559,N_22642);
nand U23666 (N_23666,N_22984,N_22694);
xor U23667 (N_23667,N_22629,N_22864);
nand U23668 (N_23668,N_22623,N_23097);
nor U23669 (N_23669,N_22581,N_22903);
or U23670 (N_23670,N_23020,N_23009);
or U23671 (N_23671,N_22511,N_23059);
or U23672 (N_23672,N_22792,N_22917);
and U23673 (N_23673,N_22874,N_23014);
xor U23674 (N_23674,N_22831,N_22668);
nor U23675 (N_23675,N_23052,N_22851);
xor U23676 (N_23676,N_22778,N_22630);
nand U23677 (N_23677,N_22652,N_23018);
xnor U23678 (N_23678,N_22905,N_22515);
and U23679 (N_23679,N_22758,N_22785);
and U23680 (N_23680,N_23089,N_22585);
nor U23681 (N_23681,N_22667,N_22697);
nor U23682 (N_23682,N_22839,N_22674);
and U23683 (N_23683,N_22565,N_22741);
and U23684 (N_23684,N_23049,N_22775);
xnor U23685 (N_23685,N_22714,N_22652);
xor U23686 (N_23686,N_22724,N_22558);
or U23687 (N_23687,N_22890,N_22537);
and U23688 (N_23688,N_22839,N_22945);
or U23689 (N_23689,N_22800,N_22794);
or U23690 (N_23690,N_22657,N_22913);
nor U23691 (N_23691,N_23034,N_22894);
nor U23692 (N_23692,N_22923,N_22953);
nor U23693 (N_23693,N_22752,N_22568);
or U23694 (N_23694,N_22839,N_22890);
nand U23695 (N_23695,N_22811,N_22690);
and U23696 (N_23696,N_23047,N_23083);
nand U23697 (N_23697,N_22687,N_22501);
xor U23698 (N_23698,N_22753,N_22981);
xor U23699 (N_23699,N_22567,N_22553);
nor U23700 (N_23700,N_22778,N_22999);
or U23701 (N_23701,N_22606,N_22762);
nand U23702 (N_23702,N_22870,N_22681);
and U23703 (N_23703,N_22773,N_22643);
or U23704 (N_23704,N_22851,N_22507);
and U23705 (N_23705,N_22901,N_22623);
nand U23706 (N_23706,N_22957,N_22951);
nand U23707 (N_23707,N_22782,N_23041);
and U23708 (N_23708,N_22575,N_22726);
or U23709 (N_23709,N_22716,N_22674);
and U23710 (N_23710,N_22540,N_22644);
nand U23711 (N_23711,N_23120,N_22954);
nor U23712 (N_23712,N_22705,N_22769);
and U23713 (N_23713,N_22908,N_23025);
and U23714 (N_23714,N_22846,N_22903);
and U23715 (N_23715,N_23078,N_22817);
or U23716 (N_23716,N_23017,N_22878);
nand U23717 (N_23717,N_22936,N_22685);
or U23718 (N_23718,N_22582,N_22598);
nand U23719 (N_23719,N_23108,N_22912);
nor U23720 (N_23720,N_22977,N_22785);
xnor U23721 (N_23721,N_22794,N_22571);
nor U23722 (N_23722,N_22586,N_22963);
nor U23723 (N_23723,N_22873,N_23012);
or U23724 (N_23724,N_22781,N_22851);
nand U23725 (N_23725,N_22542,N_22787);
or U23726 (N_23726,N_22853,N_22603);
xor U23727 (N_23727,N_22880,N_22878);
or U23728 (N_23728,N_22930,N_22927);
and U23729 (N_23729,N_22786,N_22716);
xnor U23730 (N_23730,N_22984,N_22795);
nor U23731 (N_23731,N_22927,N_22835);
nor U23732 (N_23732,N_22936,N_22639);
nand U23733 (N_23733,N_22920,N_23050);
nand U23734 (N_23734,N_22970,N_23120);
nor U23735 (N_23735,N_22606,N_22860);
nor U23736 (N_23736,N_22619,N_22851);
or U23737 (N_23737,N_22556,N_22741);
nand U23738 (N_23738,N_22890,N_22745);
nor U23739 (N_23739,N_22844,N_22866);
xnor U23740 (N_23740,N_22680,N_23009);
nor U23741 (N_23741,N_22649,N_22763);
or U23742 (N_23742,N_22895,N_22953);
nor U23743 (N_23743,N_23088,N_23084);
nor U23744 (N_23744,N_22819,N_23087);
nor U23745 (N_23745,N_22991,N_22808);
nor U23746 (N_23746,N_22898,N_22835);
nor U23747 (N_23747,N_22530,N_22857);
and U23748 (N_23748,N_22691,N_22736);
or U23749 (N_23749,N_22542,N_22550);
and U23750 (N_23750,N_23331,N_23310);
nor U23751 (N_23751,N_23727,N_23293);
and U23752 (N_23752,N_23662,N_23376);
nand U23753 (N_23753,N_23301,N_23646);
or U23754 (N_23754,N_23246,N_23715);
or U23755 (N_23755,N_23157,N_23502);
or U23756 (N_23756,N_23654,N_23241);
or U23757 (N_23757,N_23744,N_23443);
or U23758 (N_23758,N_23621,N_23219);
and U23759 (N_23759,N_23426,N_23747);
and U23760 (N_23760,N_23381,N_23597);
xnor U23761 (N_23761,N_23220,N_23230);
nand U23762 (N_23762,N_23205,N_23292);
and U23763 (N_23763,N_23433,N_23337);
or U23764 (N_23764,N_23448,N_23270);
nand U23765 (N_23765,N_23445,N_23420);
nand U23766 (N_23766,N_23640,N_23555);
nor U23767 (N_23767,N_23498,N_23410);
nand U23768 (N_23768,N_23454,N_23291);
xnor U23769 (N_23769,N_23210,N_23380);
nor U23770 (N_23770,N_23284,N_23604);
and U23771 (N_23771,N_23228,N_23632);
or U23772 (N_23772,N_23685,N_23683);
or U23773 (N_23773,N_23403,N_23684);
or U23774 (N_23774,N_23608,N_23466);
nand U23775 (N_23775,N_23379,N_23355);
xnor U23776 (N_23776,N_23127,N_23728);
nor U23777 (N_23777,N_23564,N_23208);
nor U23778 (N_23778,N_23588,N_23741);
nor U23779 (N_23779,N_23706,N_23166);
nor U23780 (N_23780,N_23668,N_23492);
nand U23781 (N_23781,N_23277,N_23326);
xnor U23782 (N_23782,N_23610,N_23212);
xnor U23783 (N_23783,N_23352,N_23623);
nor U23784 (N_23784,N_23657,N_23513);
or U23785 (N_23785,N_23557,N_23427);
nand U23786 (N_23786,N_23178,N_23673);
and U23787 (N_23787,N_23351,N_23658);
nand U23788 (N_23788,N_23736,N_23384);
or U23789 (N_23789,N_23656,N_23370);
nor U23790 (N_23790,N_23360,N_23159);
xnor U23791 (N_23791,N_23451,N_23627);
xor U23792 (N_23792,N_23150,N_23132);
nand U23793 (N_23793,N_23227,N_23642);
nor U23794 (N_23794,N_23203,N_23690);
and U23795 (N_23795,N_23485,N_23174);
nor U23796 (N_23796,N_23689,N_23435);
xnor U23797 (N_23797,N_23733,N_23636);
xor U23798 (N_23798,N_23279,N_23136);
or U23799 (N_23799,N_23325,N_23573);
or U23800 (N_23800,N_23559,N_23372);
and U23801 (N_23801,N_23193,N_23211);
xor U23802 (N_23802,N_23701,N_23532);
xnor U23803 (N_23803,N_23412,N_23700);
nand U23804 (N_23804,N_23140,N_23280);
xnor U23805 (N_23805,N_23247,N_23456);
and U23806 (N_23806,N_23437,N_23734);
and U23807 (N_23807,N_23617,N_23339);
nand U23808 (N_23808,N_23192,N_23354);
nand U23809 (N_23809,N_23452,N_23184);
nand U23810 (N_23810,N_23317,N_23161);
and U23811 (N_23811,N_23664,N_23239);
xnor U23812 (N_23812,N_23424,N_23550);
or U23813 (N_23813,N_23396,N_23130);
or U23814 (N_23814,N_23674,N_23517);
xnor U23815 (N_23815,N_23399,N_23483);
xor U23816 (N_23816,N_23579,N_23204);
xor U23817 (N_23817,N_23512,N_23135);
nor U23818 (N_23818,N_23430,N_23661);
nor U23819 (N_23819,N_23669,N_23235);
and U23820 (N_23820,N_23624,N_23691);
and U23821 (N_23821,N_23322,N_23401);
or U23822 (N_23822,N_23626,N_23363);
or U23823 (N_23823,N_23476,N_23296);
or U23824 (N_23824,N_23373,N_23278);
xor U23825 (N_23825,N_23704,N_23749);
xor U23826 (N_23826,N_23538,N_23629);
and U23827 (N_23827,N_23240,N_23195);
nor U23828 (N_23828,N_23305,N_23146);
or U23829 (N_23829,N_23563,N_23288);
nor U23830 (N_23830,N_23694,N_23584);
nor U23831 (N_23831,N_23530,N_23179);
nor U23832 (N_23832,N_23329,N_23255);
xor U23833 (N_23833,N_23409,N_23631);
nand U23834 (N_23834,N_23726,N_23265);
or U23835 (N_23835,N_23745,N_23311);
xor U23836 (N_23836,N_23609,N_23251);
nor U23837 (N_23837,N_23436,N_23523);
or U23838 (N_23838,N_23333,N_23637);
or U23839 (N_23839,N_23374,N_23696);
xnor U23840 (N_23840,N_23556,N_23603);
or U23841 (N_23841,N_23599,N_23586);
and U23842 (N_23842,N_23335,N_23590);
nand U23843 (N_23843,N_23735,N_23729);
nor U23844 (N_23844,N_23461,N_23600);
nor U23845 (N_23845,N_23717,N_23431);
or U23846 (N_23846,N_23319,N_23693);
or U23847 (N_23847,N_23671,N_23306);
xnor U23848 (N_23848,N_23307,N_23666);
and U23849 (N_23849,N_23474,N_23467);
nor U23850 (N_23850,N_23562,N_23449);
nand U23851 (N_23851,N_23425,N_23257);
nor U23852 (N_23852,N_23496,N_23350);
and U23853 (N_23853,N_23183,N_23362);
nand U23854 (N_23854,N_23678,N_23197);
and U23855 (N_23855,N_23327,N_23711);
and U23856 (N_23856,N_23386,N_23371);
and U23857 (N_23857,N_23507,N_23536);
nor U23858 (N_23858,N_23236,N_23143);
and U23859 (N_23859,N_23207,N_23582);
xor U23860 (N_23860,N_23537,N_23302);
nor U23861 (N_23861,N_23273,N_23743);
xor U23862 (N_23862,N_23153,N_23432);
or U23863 (N_23863,N_23260,N_23164);
nand U23864 (N_23864,N_23406,N_23321);
nand U23865 (N_23865,N_23552,N_23149);
nor U23866 (N_23866,N_23447,N_23162);
and U23867 (N_23867,N_23639,N_23186);
nor U23868 (N_23868,N_23332,N_23414);
and U23869 (N_23869,N_23526,N_23225);
or U23870 (N_23870,N_23383,N_23402);
and U23871 (N_23871,N_23647,N_23388);
or U23872 (N_23872,N_23688,N_23269);
and U23873 (N_23873,N_23418,N_23509);
nor U23874 (N_23874,N_23580,N_23394);
nand U23875 (N_23875,N_23561,N_23546);
xor U23876 (N_23876,N_23217,N_23510);
and U23877 (N_23877,N_23377,N_23497);
nand U23878 (N_23878,N_23553,N_23385);
or U23879 (N_23879,N_23298,N_23256);
and U23880 (N_23880,N_23177,N_23272);
and U23881 (N_23881,N_23495,N_23549);
and U23882 (N_23882,N_23176,N_23679);
or U23883 (N_23883,N_23488,N_23390);
and U23884 (N_23884,N_23682,N_23316);
nor U23885 (N_23885,N_23574,N_23541);
xnor U23886 (N_23886,N_23356,N_23441);
or U23887 (N_23887,N_23165,N_23721);
xnor U23888 (N_23888,N_23528,N_23714);
nand U23889 (N_23889,N_23263,N_23576);
and U23890 (N_23890,N_23187,N_23202);
nor U23891 (N_23891,N_23725,N_23152);
and U23892 (N_23892,N_23544,N_23267);
or U23893 (N_23893,N_23473,N_23199);
xor U23894 (N_23894,N_23716,N_23172);
or U23895 (N_23895,N_23259,N_23618);
or U23896 (N_23896,N_23271,N_23665);
or U23897 (N_23897,N_23462,N_23455);
or U23898 (N_23898,N_23249,N_23397);
and U23899 (N_23899,N_23330,N_23297);
xnor U23900 (N_23900,N_23633,N_23182);
or U23901 (N_23901,N_23463,N_23547);
and U23902 (N_23902,N_23708,N_23175);
or U23903 (N_23903,N_23320,N_23232);
nor U23904 (N_23904,N_23364,N_23589);
xor U23905 (N_23905,N_23233,N_23398);
nand U23906 (N_23906,N_23194,N_23262);
nand U23907 (N_23907,N_23190,N_23648);
or U23908 (N_23908,N_23493,N_23478);
and U23909 (N_23909,N_23209,N_23196);
xor U23910 (N_23910,N_23738,N_23226);
or U23911 (N_23911,N_23534,N_23719);
nor U23912 (N_23912,N_23213,N_23421);
or U23913 (N_23913,N_23126,N_23583);
nor U23914 (N_23914,N_23154,N_23468);
xor U23915 (N_23915,N_23189,N_23341);
or U23916 (N_23916,N_23392,N_23289);
nor U23917 (N_23917,N_23514,N_23395);
and U23918 (N_23918,N_23585,N_23655);
nor U23919 (N_23919,N_23598,N_23713);
nor U23920 (N_23920,N_23254,N_23707);
or U23921 (N_23921,N_23268,N_23318);
xnor U23922 (N_23922,N_23607,N_23516);
or U23923 (N_23923,N_23419,N_23651);
and U23924 (N_23924,N_23505,N_23653);
or U23925 (N_23925,N_23264,N_23593);
and U23926 (N_23926,N_23718,N_23417);
nor U23927 (N_23927,N_23581,N_23215);
or U23928 (N_23928,N_23703,N_23334);
and U23929 (N_23929,N_23587,N_23480);
xnor U23930 (N_23930,N_23578,N_23592);
nor U23931 (N_23931,N_23628,N_23261);
and U23932 (N_23932,N_23572,N_23644);
and U23933 (N_23933,N_23676,N_23518);
and U23934 (N_23934,N_23686,N_23185);
nor U23935 (N_23935,N_23258,N_23511);
xor U23936 (N_23936,N_23635,N_23543);
or U23937 (N_23937,N_23659,N_23275);
and U23938 (N_23938,N_23560,N_23221);
nand U23939 (N_23939,N_23486,N_23542);
and U23940 (N_23940,N_23724,N_23282);
nand U23941 (N_23941,N_23338,N_23340);
xnor U23942 (N_23942,N_23141,N_23244);
or U23943 (N_23943,N_23687,N_23529);
and U23944 (N_23944,N_23612,N_23218);
nor U23945 (N_23945,N_23702,N_23229);
and U23946 (N_23946,N_23242,N_23266);
and U23947 (N_23947,N_23477,N_23133);
or U23948 (N_23948,N_23471,N_23503);
or U23949 (N_23949,N_23746,N_23324);
xor U23950 (N_23950,N_23539,N_23515);
nand U23951 (N_23951,N_23369,N_23699);
nor U23952 (N_23952,N_23641,N_23169);
or U23953 (N_23953,N_23281,N_23315);
xnor U23954 (N_23954,N_23504,N_23475);
and U23955 (N_23955,N_23416,N_23287);
and U23956 (N_23956,N_23125,N_23342);
nor U23957 (N_23957,N_23545,N_23250);
and U23958 (N_23958,N_23672,N_23611);
or U23959 (N_23959,N_23470,N_23630);
and U23960 (N_23960,N_23349,N_23167);
nor U23961 (N_23961,N_23531,N_23276);
nor U23962 (N_23962,N_23357,N_23295);
nor U23963 (N_23963,N_23314,N_23444);
nor U23964 (N_23964,N_23551,N_23575);
xnor U23965 (N_23965,N_23652,N_23252);
nand U23966 (N_23966,N_23602,N_23168);
and U23967 (N_23967,N_23299,N_23344);
or U23968 (N_23968,N_23382,N_23216);
and U23969 (N_23969,N_23308,N_23558);
nand U23970 (N_23970,N_23138,N_23439);
xnor U23971 (N_23971,N_23248,N_23411);
nor U23972 (N_23972,N_23670,N_23535);
xor U23973 (N_23973,N_23481,N_23645);
nand U23974 (N_23974,N_23160,N_23472);
and U23975 (N_23975,N_23567,N_23524);
and U23976 (N_23976,N_23519,N_23500);
or U23977 (N_23977,N_23508,N_23595);
or U23978 (N_23978,N_23730,N_23405);
xor U23979 (N_23979,N_23649,N_23290);
or U23980 (N_23980,N_23554,N_23366);
and U23981 (N_23981,N_23155,N_23732);
xnor U23982 (N_23982,N_23469,N_23156);
nand U23983 (N_23983,N_23343,N_23274);
and U23984 (N_23984,N_23137,N_23722);
and U23985 (N_23985,N_23525,N_23171);
xor U23986 (N_23986,N_23286,N_23173);
nand U23987 (N_23987,N_23442,N_23378);
xnor U23988 (N_23988,N_23365,N_23234);
nor U23989 (N_23989,N_23400,N_23566);
or U23990 (N_23990,N_23294,N_23407);
or U23991 (N_23991,N_23643,N_23742);
and U23992 (N_23992,N_23404,N_23147);
or U23993 (N_23993,N_23697,N_23491);
nor U23994 (N_23994,N_23527,N_23605);
nand U23995 (N_23995,N_23723,N_23231);
and U23996 (N_23996,N_23368,N_23303);
or U23997 (N_23997,N_23323,N_23158);
and U23998 (N_23998,N_23238,N_23328);
and U23999 (N_23999,N_23253,N_23487);
and U24000 (N_24000,N_23440,N_23345);
or U24001 (N_24001,N_23224,N_23139);
or U24002 (N_24002,N_23616,N_23348);
or U24003 (N_24003,N_23361,N_23660);
or U24004 (N_24004,N_23479,N_23438);
or U24005 (N_24005,N_23571,N_23634);
xor U24006 (N_24006,N_23460,N_23705);
xnor U24007 (N_24007,N_23522,N_23533);
nand U24008 (N_24008,N_23450,N_23606);
and U24009 (N_24009,N_23638,N_23501);
nor U24010 (N_24010,N_23300,N_23163);
or U24011 (N_24011,N_23458,N_23720);
or U24012 (N_24012,N_23170,N_23214);
and U24013 (N_24013,N_23245,N_23200);
and U24014 (N_24014,N_23748,N_23180);
or U24015 (N_24015,N_23142,N_23692);
xor U24016 (N_24016,N_23489,N_23387);
and U24017 (N_24017,N_23134,N_23465);
nor U24018 (N_24018,N_23520,N_23188);
nor U24019 (N_24019,N_23619,N_23482);
nor U24020 (N_24020,N_23413,N_23283);
and U24021 (N_24021,N_23506,N_23408);
or U24022 (N_24022,N_23680,N_23613);
nand U24023 (N_24023,N_23663,N_23347);
xor U24024 (N_24024,N_23484,N_23206);
and U24025 (N_24025,N_23548,N_23336);
xnor U24026 (N_24026,N_23237,N_23393);
nor U24027 (N_24027,N_23615,N_23144);
or U24028 (N_24028,N_23499,N_23521);
nor U24029 (N_24029,N_23565,N_23737);
nor U24030 (N_24030,N_23434,N_23540);
or U24031 (N_24031,N_23459,N_23389);
or U24032 (N_24032,N_23712,N_23191);
nor U24033 (N_24033,N_23695,N_23353);
nand U24034 (N_24034,N_23391,N_23131);
xor U24035 (N_24035,N_23569,N_23285);
nand U24036 (N_24036,N_23740,N_23698);
xor U24037 (N_24037,N_23464,N_23309);
xor U24038 (N_24038,N_23681,N_23596);
xnor U24039 (N_24039,N_23667,N_23243);
xnor U24040 (N_24040,N_23151,N_23620);
or U24041 (N_24041,N_23675,N_23198);
or U24042 (N_24042,N_23494,N_23568);
or U24043 (N_24043,N_23446,N_23145);
xor U24044 (N_24044,N_23223,N_23367);
and U24045 (N_24045,N_23614,N_23423);
nand U24046 (N_24046,N_23731,N_23359);
or U24047 (N_24047,N_23577,N_23601);
nor U24048 (N_24048,N_23201,N_23422);
and U24049 (N_24049,N_23625,N_23129);
and U24050 (N_24050,N_23415,N_23457);
xor U24051 (N_24051,N_23346,N_23181);
xor U24052 (N_24052,N_23594,N_23453);
or U24053 (N_24053,N_23222,N_23591);
and U24054 (N_24054,N_23622,N_23650);
nor U24055 (N_24055,N_23570,N_23148);
nor U24056 (N_24056,N_23709,N_23375);
and U24057 (N_24057,N_23312,N_23490);
nand U24058 (N_24058,N_23677,N_23313);
and U24059 (N_24059,N_23710,N_23428);
and U24060 (N_24060,N_23304,N_23128);
xnor U24061 (N_24061,N_23358,N_23429);
nor U24062 (N_24062,N_23739,N_23467);
and U24063 (N_24063,N_23735,N_23373);
xnor U24064 (N_24064,N_23521,N_23278);
nor U24065 (N_24065,N_23683,N_23528);
and U24066 (N_24066,N_23506,N_23137);
nand U24067 (N_24067,N_23584,N_23439);
nand U24068 (N_24068,N_23640,N_23161);
and U24069 (N_24069,N_23632,N_23247);
nand U24070 (N_24070,N_23558,N_23489);
nor U24071 (N_24071,N_23452,N_23433);
xnor U24072 (N_24072,N_23207,N_23629);
nand U24073 (N_24073,N_23586,N_23419);
nand U24074 (N_24074,N_23372,N_23260);
or U24075 (N_24075,N_23559,N_23715);
nor U24076 (N_24076,N_23158,N_23297);
nor U24077 (N_24077,N_23435,N_23714);
nand U24078 (N_24078,N_23347,N_23264);
nor U24079 (N_24079,N_23200,N_23349);
nand U24080 (N_24080,N_23612,N_23138);
nand U24081 (N_24081,N_23233,N_23747);
and U24082 (N_24082,N_23425,N_23560);
and U24083 (N_24083,N_23340,N_23197);
xnor U24084 (N_24084,N_23187,N_23266);
nand U24085 (N_24085,N_23654,N_23308);
or U24086 (N_24086,N_23498,N_23139);
nor U24087 (N_24087,N_23344,N_23545);
xor U24088 (N_24088,N_23632,N_23630);
nand U24089 (N_24089,N_23620,N_23408);
nor U24090 (N_24090,N_23742,N_23131);
xnor U24091 (N_24091,N_23278,N_23499);
and U24092 (N_24092,N_23589,N_23535);
nor U24093 (N_24093,N_23338,N_23678);
or U24094 (N_24094,N_23614,N_23575);
xor U24095 (N_24095,N_23349,N_23209);
or U24096 (N_24096,N_23166,N_23175);
nand U24097 (N_24097,N_23566,N_23287);
nor U24098 (N_24098,N_23663,N_23264);
xor U24099 (N_24099,N_23544,N_23730);
nand U24100 (N_24100,N_23150,N_23292);
xor U24101 (N_24101,N_23424,N_23738);
or U24102 (N_24102,N_23647,N_23715);
nor U24103 (N_24103,N_23411,N_23353);
xnor U24104 (N_24104,N_23604,N_23714);
nor U24105 (N_24105,N_23174,N_23137);
xor U24106 (N_24106,N_23404,N_23360);
xnor U24107 (N_24107,N_23228,N_23275);
and U24108 (N_24108,N_23563,N_23272);
xnor U24109 (N_24109,N_23218,N_23298);
or U24110 (N_24110,N_23305,N_23560);
and U24111 (N_24111,N_23460,N_23513);
and U24112 (N_24112,N_23254,N_23234);
xor U24113 (N_24113,N_23285,N_23386);
nor U24114 (N_24114,N_23300,N_23237);
nor U24115 (N_24115,N_23471,N_23259);
xnor U24116 (N_24116,N_23294,N_23194);
or U24117 (N_24117,N_23157,N_23242);
nand U24118 (N_24118,N_23641,N_23283);
and U24119 (N_24119,N_23327,N_23661);
nand U24120 (N_24120,N_23619,N_23539);
nor U24121 (N_24121,N_23642,N_23407);
nor U24122 (N_24122,N_23548,N_23745);
nor U24123 (N_24123,N_23220,N_23174);
or U24124 (N_24124,N_23258,N_23233);
nand U24125 (N_24125,N_23721,N_23264);
nand U24126 (N_24126,N_23495,N_23509);
nor U24127 (N_24127,N_23477,N_23686);
nor U24128 (N_24128,N_23255,N_23381);
and U24129 (N_24129,N_23348,N_23485);
nand U24130 (N_24130,N_23606,N_23747);
nand U24131 (N_24131,N_23347,N_23196);
and U24132 (N_24132,N_23572,N_23373);
or U24133 (N_24133,N_23486,N_23162);
nand U24134 (N_24134,N_23256,N_23188);
nor U24135 (N_24135,N_23394,N_23621);
nand U24136 (N_24136,N_23640,N_23464);
xor U24137 (N_24137,N_23585,N_23364);
and U24138 (N_24138,N_23711,N_23523);
or U24139 (N_24139,N_23386,N_23715);
or U24140 (N_24140,N_23291,N_23210);
nand U24141 (N_24141,N_23323,N_23630);
and U24142 (N_24142,N_23257,N_23154);
and U24143 (N_24143,N_23655,N_23695);
nand U24144 (N_24144,N_23628,N_23328);
nor U24145 (N_24145,N_23193,N_23392);
nor U24146 (N_24146,N_23685,N_23358);
nor U24147 (N_24147,N_23155,N_23272);
and U24148 (N_24148,N_23444,N_23178);
xor U24149 (N_24149,N_23149,N_23656);
nor U24150 (N_24150,N_23608,N_23522);
or U24151 (N_24151,N_23606,N_23595);
nand U24152 (N_24152,N_23748,N_23732);
xnor U24153 (N_24153,N_23565,N_23186);
and U24154 (N_24154,N_23745,N_23218);
or U24155 (N_24155,N_23214,N_23664);
xnor U24156 (N_24156,N_23249,N_23376);
nor U24157 (N_24157,N_23499,N_23370);
nor U24158 (N_24158,N_23337,N_23257);
or U24159 (N_24159,N_23718,N_23311);
xor U24160 (N_24160,N_23588,N_23608);
nand U24161 (N_24161,N_23678,N_23599);
and U24162 (N_24162,N_23736,N_23695);
xnor U24163 (N_24163,N_23197,N_23501);
xnor U24164 (N_24164,N_23380,N_23219);
nor U24165 (N_24165,N_23394,N_23178);
nand U24166 (N_24166,N_23651,N_23221);
and U24167 (N_24167,N_23498,N_23127);
and U24168 (N_24168,N_23133,N_23307);
and U24169 (N_24169,N_23163,N_23303);
xnor U24170 (N_24170,N_23703,N_23621);
and U24171 (N_24171,N_23169,N_23271);
or U24172 (N_24172,N_23348,N_23245);
nor U24173 (N_24173,N_23147,N_23702);
and U24174 (N_24174,N_23677,N_23341);
xor U24175 (N_24175,N_23156,N_23359);
or U24176 (N_24176,N_23392,N_23256);
and U24177 (N_24177,N_23718,N_23201);
nand U24178 (N_24178,N_23582,N_23439);
or U24179 (N_24179,N_23588,N_23647);
nor U24180 (N_24180,N_23201,N_23566);
xor U24181 (N_24181,N_23473,N_23500);
nand U24182 (N_24182,N_23413,N_23210);
xor U24183 (N_24183,N_23584,N_23488);
nand U24184 (N_24184,N_23299,N_23321);
nor U24185 (N_24185,N_23320,N_23266);
or U24186 (N_24186,N_23187,N_23397);
nor U24187 (N_24187,N_23672,N_23325);
and U24188 (N_24188,N_23235,N_23445);
nor U24189 (N_24189,N_23725,N_23567);
or U24190 (N_24190,N_23721,N_23343);
xnor U24191 (N_24191,N_23416,N_23692);
nor U24192 (N_24192,N_23626,N_23358);
xor U24193 (N_24193,N_23741,N_23460);
xnor U24194 (N_24194,N_23189,N_23541);
and U24195 (N_24195,N_23303,N_23631);
xnor U24196 (N_24196,N_23147,N_23623);
xnor U24197 (N_24197,N_23148,N_23251);
xor U24198 (N_24198,N_23240,N_23212);
nor U24199 (N_24199,N_23403,N_23183);
and U24200 (N_24200,N_23635,N_23551);
nor U24201 (N_24201,N_23428,N_23176);
xnor U24202 (N_24202,N_23273,N_23491);
xor U24203 (N_24203,N_23573,N_23249);
nor U24204 (N_24204,N_23477,N_23356);
or U24205 (N_24205,N_23127,N_23596);
nand U24206 (N_24206,N_23574,N_23146);
nor U24207 (N_24207,N_23672,N_23694);
and U24208 (N_24208,N_23643,N_23512);
xor U24209 (N_24209,N_23414,N_23657);
or U24210 (N_24210,N_23600,N_23725);
xor U24211 (N_24211,N_23590,N_23704);
and U24212 (N_24212,N_23579,N_23557);
and U24213 (N_24213,N_23681,N_23239);
nor U24214 (N_24214,N_23132,N_23240);
and U24215 (N_24215,N_23175,N_23213);
nand U24216 (N_24216,N_23443,N_23394);
nand U24217 (N_24217,N_23507,N_23185);
and U24218 (N_24218,N_23455,N_23295);
xor U24219 (N_24219,N_23669,N_23310);
xnor U24220 (N_24220,N_23433,N_23228);
and U24221 (N_24221,N_23561,N_23712);
xor U24222 (N_24222,N_23243,N_23490);
nor U24223 (N_24223,N_23695,N_23309);
nor U24224 (N_24224,N_23581,N_23367);
nor U24225 (N_24225,N_23414,N_23201);
nor U24226 (N_24226,N_23633,N_23374);
xnor U24227 (N_24227,N_23601,N_23592);
xor U24228 (N_24228,N_23239,N_23437);
or U24229 (N_24229,N_23503,N_23704);
or U24230 (N_24230,N_23469,N_23740);
nand U24231 (N_24231,N_23413,N_23479);
nor U24232 (N_24232,N_23223,N_23556);
and U24233 (N_24233,N_23347,N_23423);
nand U24234 (N_24234,N_23498,N_23373);
nor U24235 (N_24235,N_23198,N_23234);
and U24236 (N_24236,N_23748,N_23744);
and U24237 (N_24237,N_23707,N_23522);
and U24238 (N_24238,N_23141,N_23478);
or U24239 (N_24239,N_23686,N_23426);
and U24240 (N_24240,N_23704,N_23467);
and U24241 (N_24241,N_23574,N_23429);
xor U24242 (N_24242,N_23490,N_23515);
nor U24243 (N_24243,N_23469,N_23742);
and U24244 (N_24244,N_23628,N_23585);
nand U24245 (N_24245,N_23603,N_23643);
or U24246 (N_24246,N_23206,N_23397);
or U24247 (N_24247,N_23329,N_23465);
or U24248 (N_24248,N_23379,N_23572);
xor U24249 (N_24249,N_23674,N_23252);
nor U24250 (N_24250,N_23473,N_23290);
and U24251 (N_24251,N_23287,N_23519);
xnor U24252 (N_24252,N_23274,N_23339);
nor U24253 (N_24253,N_23319,N_23404);
xnor U24254 (N_24254,N_23697,N_23678);
and U24255 (N_24255,N_23132,N_23428);
and U24256 (N_24256,N_23417,N_23388);
and U24257 (N_24257,N_23555,N_23338);
nor U24258 (N_24258,N_23398,N_23700);
or U24259 (N_24259,N_23494,N_23667);
and U24260 (N_24260,N_23615,N_23559);
or U24261 (N_24261,N_23545,N_23500);
and U24262 (N_24262,N_23349,N_23590);
nor U24263 (N_24263,N_23261,N_23471);
xnor U24264 (N_24264,N_23291,N_23201);
nor U24265 (N_24265,N_23660,N_23664);
nand U24266 (N_24266,N_23433,N_23275);
or U24267 (N_24267,N_23377,N_23165);
or U24268 (N_24268,N_23530,N_23158);
or U24269 (N_24269,N_23252,N_23664);
nand U24270 (N_24270,N_23283,N_23237);
or U24271 (N_24271,N_23626,N_23147);
nor U24272 (N_24272,N_23746,N_23245);
nand U24273 (N_24273,N_23535,N_23131);
and U24274 (N_24274,N_23549,N_23697);
nand U24275 (N_24275,N_23321,N_23742);
or U24276 (N_24276,N_23690,N_23484);
xor U24277 (N_24277,N_23315,N_23251);
xnor U24278 (N_24278,N_23562,N_23258);
nor U24279 (N_24279,N_23140,N_23507);
nor U24280 (N_24280,N_23566,N_23391);
xnor U24281 (N_24281,N_23476,N_23244);
nor U24282 (N_24282,N_23521,N_23309);
nand U24283 (N_24283,N_23655,N_23565);
nor U24284 (N_24284,N_23703,N_23172);
nor U24285 (N_24285,N_23555,N_23516);
and U24286 (N_24286,N_23567,N_23385);
nor U24287 (N_24287,N_23607,N_23530);
xnor U24288 (N_24288,N_23611,N_23662);
nor U24289 (N_24289,N_23669,N_23623);
or U24290 (N_24290,N_23165,N_23502);
nor U24291 (N_24291,N_23232,N_23375);
xnor U24292 (N_24292,N_23473,N_23526);
and U24293 (N_24293,N_23418,N_23394);
nand U24294 (N_24294,N_23178,N_23143);
or U24295 (N_24295,N_23731,N_23574);
nor U24296 (N_24296,N_23480,N_23577);
xor U24297 (N_24297,N_23335,N_23691);
and U24298 (N_24298,N_23552,N_23508);
nor U24299 (N_24299,N_23240,N_23714);
and U24300 (N_24300,N_23142,N_23268);
xnor U24301 (N_24301,N_23421,N_23154);
nand U24302 (N_24302,N_23741,N_23546);
or U24303 (N_24303,N_23452,N_23171);
nand U24304 (N_24304,N_23282,N_23646);
nand U24305 (N_24305,N_23543,N_23676);
nor U24306 (N_24306,N_23579,N_23420);
or U24307 (N_24307,N_23321,N_23209);
nand U24308 (N_24308,N_23446,N_23722);
and U24309 (N_24309,N_23245,N_23664);
and U24310 (N_24310,N_23710,N_23191);
nand U24311 (N_24311,N_23225,N_23262);
xnor U24312 (N_24312,N_23535,N_23426);
and U24313 (N_24313,N_23220,N_23564);
xnor U24314 (N_24314,N_23681,N_23443);
and U24315 (N_24315,N_23188,N_23602);
or U24316 (N_24316,N_23241,N_23629);
nor U24317 (N_24317,N_23372,N_23673);
nor U24318 (N_24318,N_23305,N_23334);
or U24319 (N_24319,N_23246,N_23360);
xnor U24320 (N_24320,N_23607,N_23476);
or U24321 (N_24321,N_23283,N_23464);
or U24322 (N_24322,N_23483,N_23416);
xor U24323 (N_24323,N_23518,N_23388);
xor U24324 (N_24324,N_23192,N_23197);
nand U24325 (N_24325,N_23687,N_23254);
xnor U24326 (N_24326,N_23540,N_23431);
nor U24327 (N_24327,N_23177,N_23651);
and U24328 (N_24328,N_23518,N_23255);
or U24329 (N_24329,N_23625,N_23587);
nand U24330 (N_24330,N_23322,N_23172);
and U24331 (N_24331,N_23722,N_23318);
xor U24332 (N_24332,N_23230,N_23250);
xnor U24333 (N_24333,N_23206,N_23585);
and U24334 (N_24334,N_23162,N_23731);
nor U24335 (N_24335,N_23532,N_23748);
or U24336 (N_24336,N_23645,N_23125);
xor U24337 (N_24337,N_23614,N_23496);
xnor U24338 (N_24338,N_23590,N_23218);
or U24339 (N_24339,N_23667,N_23352);
nand U24340 (N_24340,N_23682,N_23546);
nand U24341 (N_24341,N_23706,N_23134);
nand U24342 (N_24342,N_23253,N_23620);
xnor U24343 (N_24343,N_23501,N_23431);
nor U24344 (N_24344,N_23428,N_23747);
or U24345 (N_24345,N_23263,N_23471);
or U24346 (N_24346,N_23443,N_23560);
nor U24347 (N_24347,N_23203,N_23201);
xor U24348 (N_24348,N_23618,N_23516);
or U24349 (N_24349,N_23431,N_23713);
or U24350 (N_24350,N_23338,N_23462);
nand U24351 (N_24351,N_23229,N_23648);
xnor U24352 (N_24352,N_23705,N_23683);
or U24353 (N_24353,N_23275,N_23217);
xnor U24354 (N_24354,N_23662,N_23516);
nor U24355 (N_24355,N_23459,N_23700);
or U24356 (N_24356,N_23255,N_23194);
xor U24357 (N_24357,N_23439,N_23244);
and U24358 (N_24358,N_23365,N_23722);
and U24359 (N_24359,N_23349,N_23407);
nand U24360 (N_24360,N_23256,N_23305);
and U24361 (N_24361,N_23157,N_23176);
xnor U24362 (N_24362,N_23592,N_23449);
or U24363 (N_24363,N_23673,N_23239);
nor U24364 (N_24364,N_23422,N_23196);
and U24365 (N_24365,N_23203,N_23576);
xor U24366 (N_24366,N_23312,N_23568);
nor U24367 (N_24367,N_23306,N_23507);
xor U24368 (N_24368,N_23415,N_23564);
nor U24369 (N_24369,N_23678,N_23663);
or U24370 (N_24370,N_23563,N_23494);
and U24371 (N_24371,N_23708,N_23463);
xnor U24372 (N_24372,N_23394,N_23269);
nand U24373 (N_24373,N_23538,N_23385);
xor U24374 (N_24374,N_23667,N_23612);
and U24375 (N_24375,N_24216,N_23838);
xor U24376 (N_24376,N_24018,N_24133);
or U24377 (N_24377,N_23940,N_24348);
and U24378 (N_24378,N_24286,N_24035);
or U24379 (N_24379,N_24365,N_24257);
nand U24380 (N_24380,N_24338,N_23899);
and U24381 (N_24381,N_23956,N_24290);
nor U24382 (N_24382,N_23895,N_24127);
nor U24383 (N_24383,N_24291,N_24256);
nand U24384 (N_24384,N_24011,N_24284);
xnor U24385 (N_24385,N_24179,N_24255);
xor U24386 (N_24386,N_23860,N_23997);
nor U24387 (N_24387,N_24214,N_24129);
nor U24388 (N_24388,N_24198,N_24361);
and U24389 (N_24389,N_24330,N_24200);
xnor U24390 (N_24390,N_24157,N_24050);
nand U24391 (N_24391,N_24276,N_23795);
nand U24392 (N_24392,N_24181,N_23985);
xnor U24393 (N_24393,N_24023,N_24010);
nor U24394 (N_24394,N_23821,N_24191);
and U24395 (N_24395,N_23810,N_24232);
and U24396 (N_24396,N_24340,N_24149);
or U24397 (N_24397,N_24329,N_24027);
nor U24398 (N_24398,N_24199,N_24182);
xnor U24399 (N_24399,N_23978,N_24366);
nand U24400 (N_24400,N_24034,N_24203);
nand U24401 (N_24401,N_24024,N_23909);
nand U24402 (N_24402,N_23953,N_24146);
nand U24403 (N_24403,N_24356,N_24131);
or U24404 (N_24404,N_23833,N_23786);
nand U24405 (N_24405,N_24225,N_24012);
nor U24406 (N_24406,N_23774,N_24363);
or U24407 (N_24407,N_24280,N_23801);
and U24408 (N_24408,N_24339,N_24145);
and U24409 (N_24409,N_24277,N_24115);
and U24410 (N_24410,N_23789,N_24273);
nor U24411 (N_24411,N_23906,N_23864);
or U24412 (N_24412,N_23983,N_24337);
xnor U24413 (N_24413,N_24151,N_24065);
nor U24414 (N_24414,N_24210,N_24072);
nor U24415 (N_24415,N_24292,N_23947);
and U24416 (N_24416,N_24167,N_24084);
nand U24417 (N_24417,N_24306,N_24143);
or U24418 (N_24418,N_24169,N_24021);
nand U24419 (N_24419,N_23987,N_24158);
and U24420 (N_24420,N_24208,N_24242);
nand U24421 (N_24421,N_24274,N_24042);
nor U24422 (N_24422,N_24104,N_23791);
nor U24423 (N_24423,N_23933,N_23905);
or U24424 (N_24424,N_24059,N_23792);
nand U24425 (N_24425,N_24110,N_24121);
nand U24426 (N_24426,N_24327,N_23958);
nor U24427 (N_24427,N_23826,N_24007);
and U24428 (N_24428,N_23843,N_24064);
nor U24429 (N_24429,N_23950,N_23919);
xor U24430 (N_24430,N_23959,N_23930);
nand U24431 (N_24431,N_23837,N_24196);
nor U24432 (N_24432,N_24006,N_24117);
or U24433 (N_24433,N_24358,N_23949);
and U24434 (N_24434,N_23979,N_24071);
nand U24435 (N_24435,N_24033,N_24308);
and U24436 (N_24436,N_24371,N_24185);
nand U24437 (N_24437,N_24322,N_24350);
nor U24438 (N_24438,N_23921,N_23856);
xor U24439 (N_24439,N_24248,N_23894);
nand U24440 (N_24440,N_24119,N_23824);
nand U24441 (N_24441,N_23927,N_23773);
or U24442 (N_24442,N_24353,N_24147);
or U24443 (N_24443,N_23784,N_24270);
or U24444 (N_24444,N_23819,N_24055);
nand U24445 (N_24445,N_24188,N_24295);
or U24446 (N_24446,N_23969,N_23790);
and U24447 (N_24447,N_24250,N_24036);
nor U24448 (N_24448,N_23832,N_24135);
and U24449 (N_24449,N_24300,N_24041);
xnor U24450 (N_24450,N_24152,N_24204);
nor U24451 (N_24451,N_24206,N_23858);
nor U24452 (N_24452,N_23874,N_23961);
or U24453 (N_24453,N_24192,N_24336);
nand U24454 (N_24454,N_23772,N_24357);
and U24455 (N_24455,N_24215,N_23798);
xor U24456 (N_24456,N_23952,N_24367);
nor U24457 (N_24457,N_24173,N_23765);
or U24458 (N_24458,N_24148,N_23866);
nand U24459 (N_24459,N_23929,N_24126);
nand U24460 (N_24460,N_23884,N_23771);
and U24461 (N_24461,N_24091,N_23912);
nor U24462 (N_24462,N_24175,N_24087);
nand U24463 (N_24463,N_24014,N_24243);
nand U24464 (N_24464,N_24139,N_24074);
nand U24465 (N_24465,N_24123,N_24325);
and U24466 (N_24466,N_23776,N_23751);
nor U24467 (N_24467,N_23848,N_24045);
and U24468 (N_24468,N_23989,N_24178);
or U24469 (N_24469,N_24219,N_24180);
nor U24470 (N_24470,N_24113,N_24029);
nor U24471 (N_24471,N_23924,N_24130);
xor U24472 (N_24472,N_24098,N_23913);
or U24473 (N_24473,N_23815,N_24305);
and U24474 (N_24474,N_24344,N_24230);
xor U24475 (N_24475,N_24197,N_23973);
or U24476 (N_24476,N_24205,N_23855);
nand U24477 (N_24477,N_24047,N_24092);
xor U24478 (N_24478,N_23863,N_23999);
xor U24479 (N_24479,N_23995,N_23882);
and U24480 (N_24480,N_24263,N_23910);
xnor U24481 (N_24481,N_24161,N_24106);
and U24482 (N_24482,N_23816,N_23942);
nor U24483 (N_24483,N_23840,N_24153);
xor U24484 (N_24484,N_24239,N_23917);
nand U24485 (N_24485,N_23808,N_23807);
nor U24486 (N_24486,N_23965,N_24266);
nand U24487 (N_24487,N_23971,N_24245);
nand U24488 (N_24488,N_23897,N_23875);
and U24489 (N_24489,N_24351,N_24122);
and U24490 (N_24490,N_23967,N_23862);
nand U24491 (N_24491,N_24004,N_23852);
and U24492 (N_24492,N_24299,N_24252);
and U24493 (N_24493,N_24235,N_23885);
nand U24494 (N_24494,N_24183,N_23889);
and U24495 (N_24495,N_24046,N_24307);
nor U24496 (N_24496,N_23756,N_23908);
xnor U24497 (N_24497,N_23809,N_24079);
or U24498 (N_24498,N_24083,N_24262);
nor U24499 (N_24499,N_24254,N_23900);
nor U24500 (N_24500,N_24213,N_23881);
xnor U24501 (N_24501,N_24103,N_23846);
and U24502 (N_24502,N_23793,N_24234);
or U24503 (N_24503,N_24287,N_23955);
nor U24504 (N_24504,N_24289,N_23890);
xor U24505 (N_24505,N_24170,N_23803);
nand U24506 (N_24506,N_23805,N_24053);
nand U24507 (N_24507,N_23888,N_23762);
xor U24508 (N_24508,N_23759,N_24075);
nand U24509 (N_24509,N_24224,N_24058);
nor U24510 (N_24510,N_23844,N_24026);
nor U24511 (N_24511,N_24207,N_24326);
nand U24512 (N_24512,N_24244,N_23986);
xor U24513 (N_24513,N_23813,N_23854);
and U24514 (N_24514,N_24177,N_24144);
and U24515 (N_24515,N_24323,N_24209);
nand U24516 (N_24516,N_24043,N_23828);
nor U24517 (N_24517,N_24311,N_24137);
nor U24518 (N_24518,N_24109,N_24195);
xor U24519 (N_24519,N_24189,N_23891);
or U24520 (N_24520,N_23842,N_24054);
nand U24521 (N_24521,N_24013,N_24009);
and U24522 (N_24522,N_23943,N_23932);
or U24523 (N_24523,N_23934,N_23982);
nand U24524 (N_24524,N_24260,N_24247);
and U24525 (N_24525,N_24132,N_23794);
nand U24526 (N_24526,N_23970,N_24319);
xnor U24527 (N_24527,N_23829,N_23780);
nor U24528 (N_24528,N_24194,N_23849);
and U24529 (N_24529,N_23914,N_24335);
and U24530 (N_24530,N_24304,N_23870);
or U24531 (N_24531,N_23918,N_23963);
xnor U24532 (N_24532,N_23944,N_23872);
or U24533 (N_24533,N_23850,N_23867);
or U24534 (N_24534,N_24275,N_24349);
nand U24535 (N_24535,N_23753,N_24163);
nand U24536 (N_24536,N_23814,N_24302);
and U24537 (N_24537,N_23859,N_23968);
xor U24538 (N_24538,N_24099,N_24241);
and U24539 (N_24539,N_24003,N_24328);
and U24540 (N_24540,N_23781,N_23974);
nor U24541 (N_24541,N_24202,N_23907);
and U24542 (N_24542,N_23893,N_24097);
nand U24543 (N_24543,N_24345,N_23975);
xor U24544 (N_24544,N_24221,N_24368);
nand U24545 (N_24545,N_23767,N_24112);
nand U24546 (N_24546,N_23783,N_24303);
xnor U24547 (N_24547,N_24085,N_24267);
nand U24548 (N_24548,N_23823,N_23861);
xor U24549 (N_24549,N_24310,N_23796);
and U24550 (N_24550,N_24223,N_24229);
and U24551 (N_24551,N_23936,N_23876);
xnor U24552 (N_24552,N_24222,N_23984);
and U24553 (N_24553,N_23812,N_23761);
nor U24554 (N_24554,N_24272,N_23754);
or U24555 (N_24555,N_24271,N_24114);
xnor U24556 (N_24556,N_24116,N_24237);
nand U24557 (N_24557,N_24076,N_23851);
nor U24558 (N_24558,N_24360,N_23951);
or U24559 (N_24559,N_23752,N_23758);
nor U24560 (N_24560,N_24283,N_23886);
nor U24561 (N_24561,N_23988,N_23766);
nand U24562 (N_24562,N_23916,N_24096);
nor U24563 (N_24563,N_23865,N_24355);
or U24564 (N_24564,N_24296,N_24373);
nand U24565 (N_24565,N_24128,N_23937);
nor U24566 (N_24566,N_23948,N_24077);
and U24567 (N_24567,N_24193,N_24251);
xor U24568 (N_24568,N_24293,N_23991);
or U24569 (N_24569,N_24278,N_23777);
nand U24570 (N_24570,N_24136,N_24155);
or U24571 (N_24571,N_23841,N_24238);
xor U24572 (N_24572,N_23868,N_23779);
or U24573 (N_24573,N_24141,N_23818);
nand U24574 (N_24574,N_24067,N_24312);
and U24575 (N_24575,N_24282,N_23898);
xnor U24576 (N_24576,N_23788,N_24333);
nor U24577 (N_24577,N_23928,N_24259);
nor U24578 (N_24578,N_23763,N_24342);
nor U24579 (N_24579,N_24020,N_24002);
and U24580 (N_24580,N_24314,N_23847);
nand U24581 (N_24581,N_24264,N_24346);
nand U24582 (N_24582,N_24028,N_24080);
xor U24583 (N_24583,N_24364,N_24168);
nand U24584 (N_24584,N_24000,N_24125);
xor U24585 (N_24585,N_24037,N_24253);
or U24586 (N_24586,N_24031,N_24268);
xor U24587 (N_24587,N_24017,N_24298);
nor U24588 (N_24588,N_24332,N_24334);
xnor U24589 (N_24589,N_24231,N_23992);
or U24590 (N_24590,N_24347,N_24052);
nor U24591 (N_24591,N_23901,N_23834);
and U24592 (N_24592,N_24082,N_24019);
nand U24593 (N_24593,N_23804,N_23993);
nor U24594 (N_24594,N_23811,N_23925);
and U24595 (N_24595,N_24162,N_24176);
or U24596 (N_24596,N_24309,N_24240);
or U24597 (N_24597,N_24318,N_24258);
nor U24598 (N_24598,N_23931,N_23782);
and U24599 (N_24599,N_24374,N_24369);
xor U24600 (N_24600,N_23915,N_23760);
and U24601 (N_24601,N_24166,N_23896);
nand U24602 (N_24602,N_23990,N_23757);
xor U24603 (N_24603,N_24081,N_24088);
and U24604 (N_24604,N_23962,N_24105);
nor U24605 (N_24605,N_23887,N_24317);
and U24606 (N_24606,N_24134,N_24341);
xnor U24607 (N_24607,N_23857,N_23903);
xnor U24608 (N_24608,N_24201,N_23960);
nand U24609 (N_24609,N_24359,N_24093);
nand U24610 (N_24610,N_24070,N_24165);
or U24611 (N_24611,N_24281,N_24186);
xnor U24612 (N_24612,N_24279,N_23799);
nand U24613 (N_24613,N_23764,N_24016);
nor U24614 (N_24614,N_24269,N_23957);
xnor U24615 (N_24615,N_24044,N_24086);
nor U24616 (N_24616,N_24142,N_23922);
nand U24617 (N_24617,N_24184,N_24032);
and U24618 (N_24618,N_23994,N_23770);
nor U24619 (N_24619,N_24138,N_23904);
and U24620 (N_24620,N_23769,N_23981);
nand U24621 (N_24621,N_24040,N_24217);
nor U24622 (N_24622,N_23750,N_23946);
xor U24623 (N_24623,N_24001,N_24352);
nor U24624 (N_24624,N_24078,N_24294);
nor U24625 (N_24625,N_23825,N_23802);
xnor U24626 (N_24626,N_23883,N_23873);
nor U24627 (N_24627,N_24066,N_23945);
and U24628 (N_24628,N_24372,N_24073);
or U24629 (N_24629,N_23830,N_24324);
and U24630 (N_24630,N_24102,N_24297);
and U24631 (N_24631,N_23920,N_24261);
nand U24632 (N_24632,N_23902,N_24288);
nor U24633 (N_24633,N_23938,N_24107);
nor U24634 (N_24634,N_23954,N_24190);
nor U24635 (N_24635,N_24187,N_23879);
nand U24636 (N_24636,N_23836,N_24301);
and U24637 (N_24637,N_24062,N_24095);
nand U24638 (N_24638,N_24025,N_23911);
nor U24639 (N_24639,N_24150,N_23935);
and U24640 (N_24640,N_23892,N_24038);
xor U24641 (N_24641,N_24089,N_24218);
nor U24642 (N_24642,N_24265,N_23775);
nand U24643 (N_24643,N_24100,N_23941);
nand U24644 (N_24644,N_24090,N_23877);
or U24645 (N_24645,N_23806,N_24063);
or U24646 (N_24646,N_24068,N_24108);
nor U24647 (N_24647,N_24159,N_23755);
or U24648 (N_24648,N_24228,N_24069);
or U24649 (N_24649,N_23835,N_23827);
or U24650 (N_24650,N_24160,N_23768);
xnor U24651 (N_24651,N_23878,N_24154);
or U24652 (N_24652,N_24048,N_23785);
nand U24653 (N_24653,N_23778,N_24171);
nor U24654 (N_24654,N_23869,N_24211);
and U24655 (N_24655,N_24118,N_23839);
nor U24656 (N_24656,N_24236,N_24156);
xor U24657 (N_24657,N_24343,N_23964);
nor U24658 (N_24658,N_24313,N_23880);
xnor U24659 (N_24659,N_24030,N_24320);
xnor U24660 (N_24660,N_23797,N_23831);
nand U24661 (N_24661,N_24049,N_24022);
and U24662 (N_24662,N_24056,N_24039);
nand U24663 (N_24663,N_24124,N_24370);
or U24664 (N_24664,N_23972,N_24164);
nor U24665 (N_24665,N_23977,N_23923);
nor U24666 (N_24666,N_23976,N_24101);
nand U24667 (N_24667,N_23996,N_24331);
and U24668 (N_24668,N_24094,N_24174);
or U24669 (N_24669,N_24249,N_24362);
and U24670 (N_24670,N_24354,N_24220);
xor U24671 (N_24671,N_23998,N_24285);
nor U24672 (N_24672,N_24061,N_24051);
nand U24673 (N_24673,N_23800,N_24227);
or U24674 (N_24674,N_24315,N_23787);
xor U24675 (N_24675,N_23853,N_23817);
nand U24676 (N_24676,N_24057,N_23980);
nor U24677 (N_24677,N_24233,N_24111);
nand U24678 (N_24678,N_24008,N_23939);
or U24679 (N_24679,N_24316,N_24005);
and U24680 (N_24680,N_23820,N_24120);
or U24681 (N_24681,N_23845,N_24172);
and U24682 (N_24682,N_24246,N_24226);
xnor U24683 (N_24683,N_23871,N_24140);
nor U24684 (N_24684,N_23966,N_24015);
nand U24685 (N_24685,N_24321,N_24212);
xor U24686 (N_24686,N_23822,N_24060);
nand U24687 (N_24687,N_23926,N_23964);
xor U24688 (N_24688,N_23763,N_24113);
nor U24689 (N_24689,N_24137,N_23845);
nand U24690 (N_24690,N_23964,N_23854);
nand U24691 (N_24691,N_24089,N_23984);
nand U24692 (N_24692,N_24305,N_23963);
or U24693 (N_24693,N_23763,N_24209);
nand U24694 (N_24694,N_23902,N_24141);
nor U24695 (N_24695,N_23997,N_23898);
or U24696 (N_24696,N_24021,N_24336);
xnor U24697 (N_24697,N_24268,N_24187);
xor U24698 (N_24698,N_24190,N_24372);
nor U24699 (N_24699,N_23904,N_24157);
xnor U24700 (N_24700,N_24243,N_23769);
nand U24701 (N_24701,N_24341,N_23772);
nor U24702 (N_24702,N_24133,N_24070);
or U24703 (N_24703,N_24255,N_24137);
xor U24704 (N_24704,N_24374,N_23764);
nor U24705 (N_24705,N_24126,N_24337);
nor U24706 (N_24706,N_23910,N_23943);
and U24707 (N_24707,N_24006,N_24207);
nor U24708 (N_24708,N_24074,N_24174);
nand U24709 (N_24709,N_24098,N_23861);
and U24710 (N_24710,N_24347,N_23950);
and U24711 (N_24711,N_23876,N_24196);
or U24712 (N_24712,N_23829,N_24103);
nor U24713 (N_24713,N_24042,N_24324);
and U24714 (N_24714,N_24185,N_24159);
nand U24715 (N_24715,N_23774,N_24272);
nand U24716 (N_24716,N_24250,N_23899);
nand U24717 (N_24717,N_24285,N_24086);
or U24718 (N_24718,N_23986,N_24298);
nor U24719 (N_24719,N_24251,N_24145);
or U24720 (N_24720,N_24356,N_24329);
or U24721 (N_24721,N_24107,N_24077);
xnor U24722 (N_24722,N_23765,N_23948);
nor U24723 (N_24723,N_24254,N_24218);
xnor U24724 (N_24724,N_24101,N_24371);
and U24725 (N_24725,N_23792,N_24223);
nor U24726 (N_24726,N_24106,N_24138);
or U24727 (N_24727,N_24346,N_24120);
nor U24728 (N_24728,N_24030,N_24315);
and U24729 (N_24729,N_24021,N_23928);
xor U24730 (N_24730,N_24102,N_23913);
and U24731 (N_24731,N_24288,N_24345);
nand U24732 (N_24732,N_23845,N_24029);
nand U24733 (N_24733,N_24282,N_24143);
or U24734 (N_24734,N_24045,N_23797);
nor U24735 (N_24735,N_24136,N_24042);
and U24736 (N_24736,N_24251,N_23957);
or U24737 (N_24737,N_24185,N_23942);
or U24738 (N_24738,N_24361,N_24257);
nor U24739 (N_24739,N_23788,N_24260);
and U24740 (N_24740,N_24148,N_23996);
nand U24741 (N_24741,N_23865,N_23758);
and U24742 (N_24742,N_24240,N_24340);
or U24743 (N_24743,N_24132,N_23844);
or U24744 (N_24744,N_24165,N_24035);
nand U24745 (N_24745,N_23855,N_24230);
nor U24746 (N_24746,N_23750,N_23867);
xnor U24747 (N_24747,N_24188,N_24001);
nor U24748 (N_24748,N_24042,N_24296);
and U24749 (N_24749,N_24230,N_23875);
xnor U24750 (N_24750,N_24276,N_24300);
xnor U24751 (N_24751,N_24300,N_24181);
nor U24752 (N_24752,N_24157,N_23903);
xor U24753 (N_24753,N_24269,N_24371);
xor U24754 (N_24754,N_23769,N_24030);
and U24755 (N_24755,N_24059,N_23905);
or U24756 (N_24756,N_23808,N_24370);
or U24757 (N_24757,N_24362,N_24157);
nand U24758 (N_24758,N_24266,N_23873);
nor U24759 (N_24759,N_24191,N_23988);
nor U24760 (N_24760,N_23956,N_24099);
nand U24761 (N_24761,N_24093,N_23868);
xor U24762 (N_24762,N_24277,N_23900);
or U24763 (N_24763,N_23966,N_23882);
xnor U24764 (N_24764,N_23895,N_23915);
or U24765 (N_24765,N_24069,N_23797);
xor U24766 (N_24766,N_23995,N_24137);
or U24767 (N_24767,N_23768,N_24245);
or U24768 (N_24768,N_24364,N_24169);
and U24769 (N_24769,N_24134,N_23902);
nand U24770 (N_24770,N_23896,N_24273);
nor U24771 (N_24771,N_24247,N_24334);
nand U24772 (N_24772,N_23891,N_24198);
nor U24773 (N_24773,N_24154,N_24073);
nand U24774 (N_24774,N_24220,N_24221);
or U24775 (N_24775,N_23872,N_23764);
or U24776 (N_24776,N_23947,N_24312);
nor U24777 (N_24777,N_24062,N_24367);
xor U24778 (N_24778,N_23957,N_24188);
nand U24779 (N_24779,N_24246,N_24236);
nor U24780 (N_24780,N_23969,N_24178);
nand U24781 (N_24781,N_23888,N_24295);
or U24782 (N_24782,N_24335,N_23935);
nand U24783 (N_24783,N_24169,N_23978);
nand U24784 (N_24784,N_24282,N_24314);
nor U24785 (N_24785,N_24112,N_23831);
nand U24786 (N_24786,N_24087,N_24110);
xnor U24787 (N_24787,N_24013,N_24278);
nand U24788 (N_24788,N_24081,N_23849);
nand U24789 (N_24789,N_23859,N_23770);
and U24790 (N_24790,N_24347,N_24315);
and U24791 (N_24791,N_24115,N_24082);
nand U24792 (N_24792,N_24200,N_24176);
and U24793 (N_24793,N_24103,N_23965);
nand U24794 (N_24794,N_24171,N_24283);
and U24795 (N_24795,N_24145,N_24144);
and U24796 (N_24796,N_24361,N_23979);
xor U24797 (N_24797,N_24253,N_24144);
nand U24798 (N_24798,N_23895,N_24237);
and U24799 (N_24799,N_24117,N_24177);
or U24800 (N_24800,N_23869,N_24205);
nor U24801 (N_24801,N_24263,N_24126);
xnor U24802 (N_24802,N_23817,N_23807);
or U24803 (N_24803,N_23973,N_23850);
and U24804 (N_24804,N_24040,N_23750);
nor U24805 (N_24805,N_23933,N_23984);
nand U24806 (N_24806,N_23886,N_24321);
nand U24807 (N_24807,N_24270,N_23786);
and U24808 (N_24808,N_23836,N_24256);
xor U24809 (N_24809,N_24249,N_24013);
nand U24810 (N_24810,N_24122,N_24260);
nand U24811 (N_24811,N_23919,N_24315);
or U24812 (N_24812,N_23939,N_24199);
nor U24813 (N_24813,N_24155,N_24008);
and U24814 (N_24814,N_24088,N_24163);
xnor U24815 (N_24815,N_24037,N_24054);
and U24816 (N_24816,N_23779,N_24016);
or U24817 (N_24817,N_24287,N_23908);
xor U24818 (N_24818,N_23892,N_24145);
xor U24819 (N_24819,N_24303,N_24358);
or U24820 (N_24820,N_23965,N_24097);
and U24821 (N_24821,N_23913,N_24056);
xnor U24822 (N_24822,N_24320,N_24342);
nand U24823 (N_24823,N_24022,N_23941);
or U24824 (N_24824,N_23874,N_23793);
xor U24825 (N_24825,N_24148,N_24309);
nand U24826 (N_24826,N_24350,N_24282);
and U24827 (N_24827,N_24330,N_24096);
or U24828 (N_24828,N_24091,N_24028);
nand U24829 (N_24829,N_24236,N_23779);
and U24830 (N_24830,N_24257,N_24053);
and U24831 (N_24831,N_23822,N_24199);
or U24832 (N_24832,N_23760,N_24205);
and U24833 (N_24833,N_23776,N_24200);
nor U24834 (N_24834,N_23961,N_24107);
or U24835 (N_24835,N_24219,N_24159);
xnor U24836 (N_24836,N_24128,N_24201);
nand U24837 (N_24837,N_24332,N_23857);
nor U24838 (N_24838,N_23866,N_24309);
xnor U24839 (N_24839,N_23876,N_23963);
xor U24840 (N_24840,N_23890,N_24089);
nor U24841 (N_24841,N_24367,N_24211);
nand U24842 (N_24842,N_23945,N_24295);
and U24843 (N_24843,N_23826,N_23983);
nor U24844 (N_24844,N_24028,N_23851);
nor U24845 (N_24845,N_24106,N_24329);
or U24846 (N_24846,N_23843,N_24363);
nor U24847 (N_24847,N_24033,N_23762);
nand U24848 (N_24848,N_23914,N_23970);
or U24849 (N_24849,N_24135,N_24307);
or U24850 (N_24850,N_24051,N_24004);
nand U24851 (N_24851,N_24109,N_24363);
and U24852 (N_24852,N_23980,N_24275);
and U24853 (N_24853,N_24182,N_23976);
nand U24854 (N_24854,N_23751,N_23967);
xor U24855 (N_24855,N_24171,N_23773);
and U24856 (N_24856,N_23969,N_24102);
or U24857 (N_24857,N_24206,N_23789);
xnor U24858 (N_24858,N_23831,N_24054);
nand U24859 (N_24859,N_23960,N_24257);
or U24860 (N_24860,N_24297,N_24274);
xnor U24861 (N_24861,N_23864,N_24108);
xor U24862 (N_24862,N_24175,N_24217);
xor U24863 (N_24863,N_23954,N_23892);
nand U24864 (N_24864,N_24082,N_23855);
nand U24865 (N_24865,N_24202,N_23965);
and U24866 (N_24866,N_23947,N_23954);
nand U24867 (N_24867,N_24068,N_23816);
nor U24868 (N_24868,N_23900,N_24065);
nor U24869 (N_24869,N_23878,N_23943);
xnor U24870 (N_24870,N_23905,N_24118);
nor U24871 (N_24871,N_24246,N_23963);
xor U24872 (N_24872,N_23981,N_23805);
nor U24873 (N_24873,N_24010,N_24299);
and U24874 (N_24874,N_23842,N_24244);
and U24875 (N_24875,N_23816,N_23764);
nand U24876 (N_24876,N_24077,N_24126);
xor U24877 (N_24877,N_23808,N_23855);
xnor U24878 (N_24878,N_24347,N_24104);
xor U24879 (N_24879,N_24278,N_24083);
nand U24880 (N_24880,N_24073,N_23882);
or U24881 (N_24881,N_23844,N_24096);
nand U24882 (N_24882,N_24136,N_24079);
and U24883 (N_24883,N_23907,N_24295);
xor U24884 (N_24884,N_23813,N_24255);
xnor U24885 (N_24885,N_24102,N_24132);
or U24886 (N_24886,N_24134,N_23791);
xor U24887 (N_24887,N_24329,N_23845);
xnor U24888 (N_24888,N_23825,N_24208);
or U24889 (N_24889,N_24199,N_24251);
and U24890 (N_24890,N_24012,N_24189);
xnor U24891 (N_24891,N_24263,N_23833);
or U24892 (N_24892,N_23808,N_24365);
nor U24893 (N_24893,N_23849,N_24252);
or U24894 (N_24894,N_24124,N_23847);
xnor U24895 (N_24895,N_23834,N_24311);
or U24896 (N_24896,N_24014,N_23972);
or U24897 (N_24897,N_23896,N_24159);
and U24898 (N_24898,N_24362,N_23960);
or U24899 (N_24899,N_23943,N_23924);
or U24900 (N_24900,N_23767,N_23930);
xnor U24901 (N_24901,N_23985,N_23899);
and U24902 (N_24902,N_23840,N_24354);
nand U24903 (N_24903,N_24345,N_23818);
or U24904 (N_24904,N_24202,N_23758);
and U24905 (N_24905,N_23923,N_23840);
or U24906 (N_24906,N_23797,N_24244);
and U24907 (N_24907,N_23805,N_24149);
xor U24908 (N_24908,N_24374,N_24144);
or U24909 (N_24909,N_24047,N_23816);
or U24910 (N_24910,N_23911,N_24306);
or U24911 (N_24911,N_23761,N_24307);
and U24912 (N_24912,N_24120,N_24227);
and U24913 (N_24913,N_23875,N_24309);
or U24914 (N_24914,N_24271,N_23788);
nor U24915 (N_24915,N_24066,N_24166);
nor U24916 (N_24916,N_23824,N_23912);
and U24917 (N_24917,N_24366,N_24093);
nand U24918 (N_24918,N_24037,N_23956);
nor U24919 (N_24919,N_24347,N_23988);
and U24920 (N_24920,N_23846,N_23997);
xnor U24921 (N_24921,N_24186,N_23849);
nand U24922 (N_24922,N_23760,N_23889);
and U24923 (N_24923,N_24314,N_24179);
nand U24924 (N_24924,N_23843,N_24077);
or U24925 (N_24925,N_24143,N_23899);
or U24926 (N_24926,N_24164,N_23976);
and U24927 (N_24927,N_24211,N_24327);
nand U24928 (N_24928,N_23837,N_23995);
nand U24929 (N_24929,N_24091,N_23911);
xnor U24930 (N_24930,N_24110,N_23792);
or U24931 (N_24931,N_23887,N_24087);
nor U24932 (N_24932,N_24158,N_24264);
nor U24933 (N_24933,N_23751,N_24286);
nand U24934 (N_24934,N_23785,N_24031);
nand U24935 (N_24935,N_24146,N_24072);
nor U24936 (N_24936,N_23980,N_24308);
or U24937 (N_24937,N_23788,N_24089);
nor U24938 (N_24938,N_23773,N_24353);
xor U24939 (N_24939,N_24270,N_24059);
nor U24940 (N_24940,N_24268,N_23757);
xnor U24941 (N_24941,N_24255,N_24357);
xor U24942 (N_24942,N_24289,N_24004);
nand U24943 (N_24943,N_24108,N_23750);
or U24944 (N_24944,N_24079,N_24127);
and U24945 (N_24945,N_24190,N_24044);
xnor U24946 (N_24946,N_23988,N_24013);
nor U24947 (N_24947,N_24325,N_24354);
xnor U24948 (N_24948,N_23815,N_23939);
nand U24949 (N_24949,N_24260,N_24031);
and U24950 (N_24950,N_23779,N_24271);
and U24951 (N_24951,N_24321,N_24301);
nor U24952 (N_24952,N_23841,N_23953);
and U24953 (N_24953,N_24355,N_24322);
nand U24954 (N_24954,N_23958,N_24316);
and U24955 (N_24955,N_24070,N_24250);
nor U24956 (N_24956,N_24313,N_23825);
nor U24957 (N_24957,N_23950,N_23854);
xor U24958 (N_24958,N_24203,N_24025);
or U24959 (N_24959,N_24128,N_23992);
nor U24960 (N_24960,N_24239,N_24175);
xor U24961 (N_24961,N_23751,N_24094);
xor U24962 (N_24962,N_23946,N_23932);
nor U24963 (N_24963,N_23859,N_24066);
nor U24964 (N_24964,N_24126,N_24334);
or U24965 (N_24965,N_24351,N_24115);
nand U24966 (N_24966,N_24131,N_23881);
xor U24967 (N_24967,N_23785,N_24065);
and U24968 (N_24968,N_23782,N_23933);
nor U24969 (N_24969,N_24151,N_24361);
nand U24970 (N_24970,N_23838,N_24016);
or U24971 (N_24971,N_23829,N_24148);
nor U24972 (N_24972,N_24118,N_24080);
nand U24973 (N_24973,N_24252,N_24187);
xor U24974 (N_24974,N_23815,N_24004);
nand U24975 (N_24975,N_24288,N_23796);
and U24976 (N_24976,N_24160,N_23979);
and U24977 (N_24977,N_24260,N_24201);
or U24978 (N_24978,N_23803,N_23850);
xnor U24979 (N_24979,N_24247,N_24204);
and U24980 (N_24980,N_24317,N_23757);
xnor U24981 (N_24981,N_24372,N_24307);
nand U24982 (N_24982,N_24239,N_24154);
and U24983 (N_24983,N_24258,N_23902);
or U24984 (N_24984,N_23918,N_24309);
xnor U24985 (N_24985,N_24329,N_24344);
and U24986 (N_24986,N_24328,N_24165);
or U24987 (N_24987,N_23902,N_24298);
and U24988 (N_24988,N_23854,N_23895);
or U24989 (N_24989,N_24295,N_24292);
nand U24990 (N_24990,N_24292,N_24311);
nand U24991 (N_24991,N_24185,N_24309);
xor U24992 (N_24992,N_23895,N_23896);
nand U24993 (N_24993,N_24126,N_24246);
nand U24994 (N_24994,N_24173,N_24100);
xor U24995 (N_24995,N_23905,N_23865);
nor U24996 (N_24996,N_24258,N_24211);
nor U24997 (N_24997,N_24316,N_24356);
and U24998 (N_24998,N_24322,N_24036);
xnor U24999 (N_24999,N_23944,N_23952);
nor UO_0 (O_0,N_24644,N_24971);
or UO_1 (O_1,N_24915,N_24758);
xnor UO_2 (O_2,N_24428,N_24496);
nand UO_3 (O_3,N_24567,N_24499);
xnor UO_4 (O_4,N_24625,N_24489);
and UO_5 (O_5,N_24526,N_24498);
or UO_6 (O_6,N_24539,N_24637);
nor UO_7 (O_7,N_24694,N_24586);
nor UO_8 (O_8,N_24587,N_24550);
nor UO_9 (O_9,N_24707,N_24668);
and UO_10 (O_10,N_24522,N_24782);
nand UO_11 (O_11,N_24438,N_24899);
xor UO_12 (O_12,N_24389,N_24440);
nand UO_13 (O_13,N_24685,N_24749);
nand UO_14 (O_14,N_24659,N_24859);
and UO_15 (O_15,N_24677,N_24926);
nand UO_16 (O_16,N_24503,N_24381);
nand UO_17 (O_17,N_24549,N_24741);
nor UO_18 (O_18,N_24444,N_24736);
or UO_19 (O_19,N_24601,N_24999);
and UO_20 (O_20,N_24593,N_24865);
and UO_21 (O_21,N_24477,N_24472);
xnor UO_22 (O_22,N_24730,N_24589);
and UO_23 (O_23,N_24632,N_24913);
and UO_24 (O_24,N_24907,N_24604);
or UO_25 (O_25,N_24555,N_24824);
and UO_26 (O_26,N_24717,N_24921);
xnor UO_27 (O_27,N_24518,N_24946);
nand UO_28 (O_28,N_24618,N_24402);
nand UO_29 (O_29,N_24948,N_24822);
or UO_30 (O_30,N_24556,N_24666);
nor UO_31 (O_31,N_24862,N_24885);
or UO_32 (O_32,N_24757,N_24655);
and UO_33 (O_33,N_24533,N_24953);
and UO_34 (O_34,N_24712,N_24765);
and UO_35 (O_35,N_24379,N_24722);
xnor UO_36 (O_36,N_24799,N_24917);
and UO_37 (O_37,N_24537,N_24821);
and UO_38 (O_38,N_24572,N_24720);
nor UO_39 (O_39,N_24935,N_24390);
xnor UO_40 (O_40,N_24497,N_24959);
xor UO_41 (O_41,N_24861,N_24848);
or UO_42 (O_42,N_24798,N_24780);
and UO_43 (O_43,N_24789,N_24453);
or UO_44 (O_44,N_24967,N_24403);
and UO_45 (O_45,N_24462,N_24635);
nor UO_46 (O_46,N_24648,N_24690);
and UO_47 (O_47,N_24998,N_24426);
nand UO_48 (O_48,N_24711,N_24647);
or UO_49 (O_49,N_24564,N_24981);
nor UO_50 (O_50,N_24442,N_24542);
nand UO_51 (O_51,N_24450,N_24591);
or UO_52 (O_52,N_24396,N_24698);
nand UO_53 (O_53,N_24531,N_24830);
nand UO_54 (O_54,N_24613,N_24762);
and UO_55 (O_55,N_24929,N_24705);
nand UO_56 (O_56,N_24775,N_24986);
nand UO_57 (O_57,N_24943,N_24742);
nor UO_58 (O_58,N_24923,N_24582);
and UO_59 (O_59,N_24561,N_24552);
nor UO_60 (O_60,N_24599,N_24812);
nand UO_61 (O_61,N_24558,N_24755);
and UO_62 (O_62,N_24973,N_24502);
nand UO_63 (O_63,N_24393,N_24597);
and UO_64 (O_64,N_24709,N_24810);
and UO_65 (O_65,N_24422,N_24731);
and UO_66 (O_66,N_24874,N_24557);
or UO_67 (O_67,N_24454,N_24884);
nand UO_68 (O_68,N_24793,N_24787);
xor UO_69 (O_69,N_24804,N_24876);
xor UO_70 (O_70,N_24476,N_24528);
and UO_71 (O_71,N_24983,N_24576);
or UO_72 (O_72,N_24776,N_24455);
and UO_73 (O_73,N_24541,N_24735);
xnor UO_74 (O_74,N_24691,N_24554);
and UO_75 (O_75,N_24585,N_24763);
and UO_76 (O_76,N_24387,N_24507);
nand UO_77 (O_77,N_24553,N_24424);
nand UO_78 (O_78,N_24517,N_24430);
nor UO_79 (O_79,N_24609,N_24485);
nand UO_80 (O_80,N_24759,N_24845);
xor UO_81 (O_81,N_24512,N_24473);
xnor UO_82 (O_82,N_24504,N_24431);
and UO_83 (O_83,N_24910,N_24847);
or UO_84 (O_84,N_24409,N_24680);
nand UO_85 (O_85,N_24594,N_24652);
or UO_86 (O_86,N_24596,N_24624);
and UO_87 (O_87,N_24616,N_24629);
and UO_88 (O_88,N_24617,N_24975);
nand UO_89 (O_89,N_24933,N_24457);
nand UO_90 (O_90,N_24844,N_24883);
xor UO_91 (O_91,N_24997,N_24737);
or UO_92 (O_92,N_24702,N_24559);
or UO_93 (O_93,N_24952,N_24856);
and UO_94 (O_94,N_24945,N_24785);
xnor UO_95 (O_95,N_24828,N_24397);
xor UO_96 (O_96,N_24871,N_24744);
xor UO_97 (O_97,N_24683,N_24902);
xnor UO_98 (O_98,N_24827,N_24951);
xnor UO_99 (O_99,N_24535,N_24928);
xnor UO_100 (O_100,N_24980,N_24638);
and UO_101 (O_101,N_24656,N_24375);
xnor UO_102 (O_102,N_24615,N_24949);
and UO_103 (O_103,N_24919,N_24942);
and UO_104 (O_104,N_24460,N_24429);
xnor UO_105 (O_105,N_24819,N_24574);
or UO_106 (O_106,N_24376,N_24699);
and UO_107 (O_107,N_24463,N_24905);
xor UO_108 (O_108,N_24739,N_24486);
and UO_109 (O_109,N_24488,N_24954);
xor UO_110 (O_110,N_24813,N_24480);
or UO_111 (O_111,N_24872,N_24882);
and UO_112 (O_112,N_24962,N_24937);
nand UO_113 (O_113,N_24740,N_24456);
nand UO_114 (O_114,N_24725,N_24818);
or UO_115 (O_115,N_24815,N_24808);
nand UO_116 (O_116,N_24748,N_24723);
nand UO_117 (O_117,N_24569,N_24727);
and UO_118 (O_118,N_24568,N_24714);
xnor UO_119 (O_119,N_24448,N_24688);
xnor UO_120 (O_120,N_24612,N_24888);
or UO_121 (O_121,N_24417,N_24832);
nor UO_122 (O_122,N_24420,N_24781);
xor UO_123 (O_123,N_24639,N_24588);
or UO_124 (O_124,N_24605,N_24619);
and UO_125 (O_125,N_24546,N_24383);
nand UO_126 (O_126,N_24511,N_24443);
xnor UO_127 (O_127,N_24916,N_24726);
nor UO_128 (O_128,N_24501,N_24492);
or UO_129 (O_129,N_24825,N_24678);
nor UO_130 (O_130,N_24852,N_24996);
nand UO_131 (O_131,N_24769,N_24406);
and UO_132 (O_132,N_24932,N_24738);
nor UO_133 (O_133,N_24670,N_24817);
nand UO_134 (O_134,N_24895,N_24858);
nand UO_135 (O_135,N_24446,N_24548);
nor UO_136 (O_136,N_24607,N_24689);
and UO_137 (O_137,N_24718,N_24598);
xnor UO_138 (O_138,N_24530,N_24675);
nor UO_139 (O_139,N_24764,N_24743);
nand UO_140 (O_140,N_24491,N_24835);
and UO_141 (O_141,N_24408,N_24879);
nor UO_142 (O_142,N_24665,N_24660);
and UO_143 (O_143,N_24425,N_24977);
xor UO_144 (O_144,N_24966,N_24704);
and UO_145 (O_145,N_24990,N_24944);
nand UO_146 (O_146,N_24445,N_24754);
nor UO_147 (O_147,N_24965,N_24918);
or UO_148 (O_148,N_24797,N_24377);
xor UO_149 (O_149,N_24860,N_24437);
or UO_150 (O_150,N_24771,N_24469);
or UO_151 (O_151,N_24398,N_24912);
or UO_152 (O_152,N_24796,N_24385);
and UO_153 (O_153,N_24686,N_24706);
nand UO_154 (O_154,N_24681,N_24490);
or UO_155 (O_155,N_24989,N_24672);
or UO_156 (O_156,N_24386,N_24620);
xor UO_157 (O_157,N_24449,N_24663);
and UO_158 (O_158,N_24521,N_24838);
or UO_159 (O_159,N_24479,N_24878);
nand UO_160 (O_160,N_24992,N_24696);
nor UO_161 (O_161,N_24724,N_24651);
nand UO_162 (O_162,N_24674,N_24684);
or UO_163 (O_163,N_24809,N_24747);
or UO_164 (O_164,N_24642,N_24693);
and UO_165 (O_165,N_24745,N_24534);
xnor UO_166 (O_166,N_24662,N_24514);
nor UO_167 (O_167,N_24843,N_24471);
nand UO_168 (O_168,N_24692,N_24968);
nor UO_169 (O_169,N_24566,N_24461);
xor UO_170 (O_170,N_24695,N_24520);
nor UO_171 (O_171,N_24500,N_24767);
xnor UO_172 (O_172,N_24846,N_24993);
nand UO_173 (O_173,N_24939,N_24657);
or UO_174 (O_174,N_24893,N_24467);
nand UO_175 (O_175,N_24654,N_24777);
nand UO_176 (O_176,N_24433,N_24719);
nor UO_177 (O_177,N_24525,N_24877);
nor UO_178 (O_178,N_24415,N_24760);
or UO_179 (O_179,N_24887,N_24608);
and UO_180 (O_180,N_24658,N_24536);
nor UO_181 (O_181,N_24510,N_24784);
nand UO_182 (O_182,N_24853,N_24487);
xnor UO_183 (O_183,N_24421,N_24701);
and UO_184 (O_184,N_24898,N_24728);
nand UO_185 (O_185,N_24636,N_24661);
and UO_186 (O_186,N_24404,N_24697);
or UO_187 (O_187,N_24631,N_24603);
or UO_188 (O_188,N_24419,N_24938);
and UO_189 (O_189,N_24543,N_24988);
nand UO_190 (O_190,N_24894,N_24994);
or UO_191 (O_191,N_24896,N_24423);
xnor UO_192 (O_192,N_24900,N_24547);
nor UO_193 (O_193,N_24653,N_24405);
nor UO_194 (O_194,N_24577,N_24873);
nor UO_195 (O_195,N_24523,N_24590);
nor UO_196 (O_196,N_24509,N_24447);
xnor UO_197 (O_197,N_24930,N_24710);
and UO_198 (O_198,N_24700,N_24484);
and UO_199 (O_199,N_24881,N_24578);
or UO_200 (O_200,N_24880,N_24413);
nand UO_201 (O_201,N_24671,N_24914);
xnor UO_202 (O_202,N_24972,N_24482);
or UO_203 (O_203,N_24669,N_24791);
nand UO_204 (O_204,N_24388,N_24527);
and UO_205 (O_205,N_24579,N_24478);
nor UO_206 (O_206,N_24934,N_24909);
xnor UO_207 (O_207,N_24435,N_24468);
nand UO_208 (O_208,N_24753,N_24532);
or UO_209 (O_209,N_24451,N_24384);
or UO_210 (O_210,N_24545,N_24628);
nand UO_211 (O_211,N_24783,N_24750);
or UO_212 (O_212,N_24958,N_24600);
xnor UO_213 (O_213,N_24924,N_24950);
and UO_214 (O_214,N_24459,N_24427);
xor UO_215 (O_215,N_24602,N_24964);
nor UO_216 (O_216,N_24575,N_24940);
nor UO_217 (O_217,N_24544,N_24378);
nand UO_218 (O_218,N_24849,N_24801);
and UO_219 (O_219,N_24626,N_24540);
and UO_220 (O_220,N_24399,N_24716);
nand UO_221 (O_221,N_24855,N_24925);
or UO_222 (O_222,N_24866,N_24904);
nor UO_223 (O_223,N_24703,N_24562);
and UO_224 (O_224,N_24790,N_24400);
xnor UO_225 (O_225,N_24766,N_24868);
nor UO_226 (O_226,N_24464,N_24851);
and UO_227 (O_227,N_24770,N_24792);
and UO_228 (O_228,N_24831,N_24957);
nor UO_229 (O_229,N_24412,N_24524);
and UO_230 (O_230,N_24826,N_24622);
and UO_231 (O_231,N_24401,N_24850);
or UO_232 (O_232,N_24779,N_24867);
or UO_233 (O_233,N_24611,N_24643);
nor UO_234 (O_234,N_24955,N_24519);
xor UO_235 (O_235,N_24708,N_24960);
nor UO_236 (O_236,N_24573,N_24839);
nand UO_237 (O_237,N_24411,N_24956);
and UO_238 (O_238,N_24800,N_24465);
and UO_239 (O_239,N_24920,N_24645);
nor UO_240 (O_240,N_24565,N_24976);
nand UO_241 (O_241,N_24650,N_24664);
nand UO_242 (O_242,N_24614,N_24441);
nand UO_243 (O_243,N_24458,N_24995);
nor UO_244 (O_244,N_24987,N_24772);
or UO_245 (O_245,N_24515,N_24969);
and UO_246 (O_246,N_24392,N_24833);
and UO_247 (O_247,N_24595,N_24991);
xor UO_248 (O_248,N_24729,N_24908);
nand UO_249 (O_249,N_24814,N_24778);
or UO_250 (O_250,N_24394,N_24516);
nor UO_251 (O_251,N_24982,N_24970);
nor UO_252 (O_252,N_24495,N_24687);
xnor UO_253 (O_253,N_24841,N_24840);
nor UO_254 (O_254,N_24816,N_24836);
xor UO_255 (O_255,N_24560,N_24416);
nor UO_256 (O_256,N_24870,N_24834);
and UO_257 (O_257,N_24434,N_24439);
or UO_258 (O_258,N_24806,N_24947);
xor UO_259 (O_259,N_24890,N_24829);
xnor UO_260 (O_260,N_24649,N_24505);
xnor UO_261 (O_261,N_24584,N_24768);
xnor UO_262 (O_262,N_24786,N_24961);
and UO_263 (O_263,N_24864,N_24922);
nor UO_264 (O_264,N_24470,N_24820);
nor UO_265 (O_265,N_24580,N_24641);
xor UO_266 (O_266,N_24436,N_24713);
xnor UO_267 (O_267,N_24979,N_24673);
nand UO_268 (O_268,N_24571,N_24506);
and UO_269 (O_269,N_24911,N_24756);
nand UO_270 (O_270,N_24391,N_24733);
xor UO_271 (O_271,N_24774,N_24802);
nor UO_272 (O_272,N_24623,N_24432);
xor UO_273 (O_273,N_24889,N_24903);
or UO_274 (O_274,N_24985,N_24752);
xnor UO_275 (O_275,N_24746,N_24529);
and UO_276 (O_276,N_24795,N_24513);
xor UO_277 (O_277,N_24494,N_24875);
xor UO_278 (O_278,N_24773,N_24538);
and UO_279 (O_279,N_24869,N_24667);
nand UO_280 (O_280,N_24842,N_24592);
nor UO_281 (O_281,N_24886,N_24418);
nor UO_282 (O_282,N_24805,N_24721);
or UO_283 (O_283,N_24640,N_24936);
or UO_284 (O_284,N_24854,N_24563);
and UO_285 (O_285,N_24508,N_24380);
nor UO_286 (O_286,N_24901,N_24676);
nor UO_287 (O_287,N_24978,N_24941);
and UO_288 (O_288,N_24984,N_24621);
or UO_289 (O_289,N_24634,N_24803);
or UO_290 (O_290,N_24857,N_24583);
or UO_291 (O_291,N_24837,N_24627);
or UO_292 (O_292,N_24475,N_24963);
nand UO_293 (O_293,N_24823,N_24481);
nor UO_294 (O_294,N_24551,N_24732);
xnor UO_295 (O_295,N_24474,N_24382);
and UO_296 (O_296,N_24794,N_24682);
or UO_297 (O_297,N_24931,N_24891);
xor UO_298 (O_298,N_24395,N_24974);
and UO_299 (O_299,N_24761,N_24452);
xor UO_300 (O_300,N_24633,N_24715);
xnor UO_301 (O_301,N_24751,N_24897);
nand UO_302 (O_302,N_24788,N_24466);
or UO_303 (O_303,N_24630,N_24414);
xnor UO_304 (O_304,N_24679,N_24734);
nand UO_305 (O_305,N_24807,N_24811);
or UO_306 (O_306,N_24646,N_24407);
xor UO_307 (O_307,N_24606,N_24570);
nor UO_308 (O_308,N_24927,N_24410);
nor UO_309 (O_309,N_24892,N_24863);
xor UO_310 (O_310,N_24493,N_24581);
nand UO_311 (O_311,N_24610,N_24483);
xor UO_312 (O_312,N_24906,N_24688);
nor UO_313 (O_313,N_24435,N_24594);
nand UO_314 (O_314,N_24983,N_24783);
and UO_315 (O_315,N_24680,N_24582);
and UO_316 (O_316,N_24522,N_24850);
and UO_317 (O_317,N_24487,N_24845);
xnor UO_318 (O_318,N_24458,N_24746);
and UO_319 (O_319,N_24399,N_24683);
and UO_320 (O_320,N_24618,N_24780);
nand UO_321 (O_321,N_24707,N_24498);
xor UO_322 (O_322,N_24600,N_24825);
and UO_323 (O_323,N_24381,N_24845);
and UO_324 (O_324,N_24419,N_24932);
xnor UO_325 (O_325,N_24688,N_24459);
nand UO_326 (O_326,N_24849,N_24664);
xor UO_327 (O_327,N_24975,N_24824);
or UO_328 (O_328,N_24566,N_24539);
xnor UO_329 (O_329,N_24967,N_24634);
nor UO_330 (O_330,N_24556,N_24639);
or UO_331 (O_331,N_24554,N_24616);
or UO_332 (O_332,N_24988,N_24451);
xnor UO_333 (O_333,N_24474,N_24548);
nand UO_334 (O_334,N_24707,N_24648);
xnor UO_335 (O_335,N_24577,N_24505);
and UO_336 (O_336,N_24444,N_24620);
nand UO_337 (O_337,N_24645,N_24462);
nand UO_338 (O_338,N_24834,N_24406);
xnor UO_339 (O_339,N_24902,N_24592);
nand UO_340 (O_340,N_24995,N_24892);
or UO_341 (O_341,N_24666,N_24956);
and UO_342 (O_342,N_24671,N_24570);
and UO_343 (O_343,N_24810,N_24917);
xnor UO_344 (O_344,N_24814,N_24458);
and UO_345 (O_345,N_24911,N_24561);
and UO_346 (O_346,N_24557,N_24798);
nand UO_347 (O_347,N_24589,N_24590);
nand UO_348 (O_348,N_24539,N_24645);
and UO_349 (O_349,N_24745,N_24439);
nor UO_350 (O_350,N_24726,N_24889);
xor UO_351 (O_351,N_24736,N_24525);
and UO_352 (O_352,N_24425,N_24593);
nor UO_353 (O_353,N_24762,N_24501);
nor UO_354 (O_354,N_24572,N_24539);
nor UO_355 (O_355,N_24712,N_24836);
nand UO_356 (O_356,N_24426,N_24700);
or UO_357 (O_357,N_24806,N_24697);
xnor UO_358 (O_358,N_24660,N_24440);
xor UO_359 (O_359,N_24517,N_24394);
xor UO_360 (O_360,N_24959,N_24915);
nor UO_361 (O_361,N_24601,N_24389);
nand UO_362 (O_362,N_24521,N_24505);
or UO_363 (O_363,N_24559,N_24707);
nand UO_364 (O_364,N_24651,N_24772);
xnor UO_365 (O_365,N_24937,N_24822);
nand UO_366 (O_366,N_24526,N_24616);
xnor UO_367 (O_367,N_24744,N_24845);
and UO_368 (O_368,N_24564,N_24835);
xnor UO_369 (O_369,N_24418,N_24994);
or UO_370 (O_370,N_24585,N_24451);
xor UO_371 (O_371,N_24415,N_24542);
nor UO_372 (O_372,N_24810,N_24495);
xor UO_373 (O_373,N_24874,N_24664);
xnor UO_374 (O_374,N_24601,N_24576);
nand UO_375 (O_375,N_24796,N_24756);
or UO_376 (O_376,N_24695,N_24565);
nand UO_377 (O_377,N_24671,N_24589);
nand UO_378 (O_378,N_24397,N_24990);
or UO_379 (O_379,N_24482,N_24556);
xor UO_380 (O_380,N_24423,N_24683);
xnor UO_381 (O_381,N_24596,N_24810);
nor UO_382 (O_382,N_24559,N_24912);
or UO_383 (O_383,N_24429,N_24951);
nor UO_384 (O_384,N_24757,N_24946);
or UO_385 (O_385,N_24600,N_24420);
and UO_386 (O_386,N_24813,N_24797);
and UO_387 (O_387,N_24502,N_24675);
xnor UO_388 (O_388,N_24409,N_24463);
nor UO_389 (O_389,N_24932,N_24580);
and UO_390 (O_390,N_24631,N_24480);
nor UO_391 (O_391,N_24801,N_24668);
nor UO_392 (O_392,N_24583,N_24889);
nor UO_393 (O_393,N_24914,N_24770);
or UO_394 (O_394,N_24649,N_24703);
or UO_395 (O_395,N_24669,N_24519);
or UO_396 (O_396,N_24977,N_24899);
and UO_397 (O_397,N_24753,N_24544);
nor UO_398 (O_398,N_24618,N_24772);
xor UO_399 (O_399,N_24874,N_24498);
and UO_400 (O_400,N_24826,N_24856);
or UO_401 (O_401,N_24568,N_24790);
nand UO_402 (O_402,N_24624,N_24694);
and UO_403 (O_403,N_24636,N_24986);
xnor UO_404 (O_404,N_24450,N_24801);
and UO_405 (O_405,N_24376,N_24583);
nor UO_406 (O_406,N_24834,N_24728);
and UO_407 (O_407,N_24464,N_24961);
or UO_408 (O_408,N_24653,N_24756);
or UO_409 (O_409,N_24544,N_24868);
or UO_410 (O_410,N_24483,N_24950);
nor UO_411 (O_411,N_24847,N_24633);
or UO_412 (O_412,N_24710,N_24979);
xor UO_413 (O_413,N_24892,N_24964);
xnor UO_414 (O_414,N_24781,N_24840);
xor UO_415 (O_415,N_24464,N_24962);
xnor UO_416 (O_416,N_24699,N_24530);
xor UO_417 (O_417,N_24469,N_24944);
nor UO_418 (O_418,N_24773,N_24532);
nand UO_419 (O_419,N_24683,N_24811);
nand UO_420 (O_420,N_24801,N_24598);
or UO_421 (O_421,N_24833,N_24561);
xnor UO_422 (O_422,N_24454,N_24550);
nor UO_423 (O_423,N_24584,N_24994);
nand UO_424 (O_424,N_24741,N_24660);
nand UO_425 (O_425,N_24571,N_24836);
xor UO_426 (O_426,N_24876,N_24954);
and UO_427 (O_427,N_24628,N_24956);
nor UO_428 (O_428,N_24621,N_24565);
nand UO_429 (O_429,N_24391,N_24534);
nor UO_430 (O_430,N_24962,N_24599);
nor UO_431 (O_431,N_24606,N_24949);
nor UO_432 (O_432,N_24657,N_24828);
xnor UO_433 (O_433,N_24562,N_24945);
nor UO_434 (O_434,N_24613,N_24381);
nand UO_435 (O_435,N_24454,N_24938);
or UO_436 (O_436,N_24663,N_24730);
and UO_437 (O_437,N_24643,N_24748);
and UO_438 (O_438,N_24491,N_24886);
or UO_439 (O_439,N_24604,N_24485);
xnor UO_440 (O_440,N_24458,N_24612);
or UO_441 (O_441,N_24771,N_24647);
nor UO_442 (O_442,N_24808,N_24556);
nor UO_443 (O_443,N_24956,N_24427);
nor UO_444 (O_444,N_24537,N_24382);
and UO_445 (O_445,N_24997,N_24796);
and UO_446 (O_446,N_24896,N_24899);
xor UO_447 (O_447,N_24718,N_24681);
xnor UO_448 (O_448,N_24378,N_24718);
and UO_449 (O_449,N_24753,N_24857);
or UO_450 (O_450,N_24779,N_24586);
xor UO_451 (O_451,N_24625,N_24804);
nor UO_452 (O_452,N_24984,N_24899);
xor UO_453 (O_453,N_24387,N_24426);
xnor UO_454 (O_454,N_24398,N_24907);
and UO_455 (O_455,N_24956,N_24931);
nor UO_456 (O_456,N_24589,N_24857);
and UO_457 (O_457,N_24676,N_24906);
xor UO_458 (O_458,N_24825,N_24398);
or UO_459 (O_459,N_24426,N_24617);
nand UO_460 (O_460,N_24487,N_24624);
or UO_461 (O_461,N_24932,N_24786);
or UO_462 (O_462,N_24763,N_24792);
nand UO_463 (O_463,N_24836,N_24808);
nor UO_464 (O_464,N_24550,N_24999);
nand UO_465 (O_465,N_24532,N_24530);
nand UO_466 (O_466,N_24930,N_24908);
nor UO_467 (O_467,N_24605,N_24680);
and UO_468 (O_468,N_24885,N_24790);
and UO_469 (O_469,N_24584,N_24716);
or UO_470 (O_470,N_24501,N_24551);
nand UO_471 (O_471,N_24800,N_24925);
nor UO_472 (O_472,N_24620,N_24827);
nand UO_473 (O_473,N_24542,N_24763);
and UO_474 (O_474,N_24922,N_24963);
xnor UO_475 (O_475,N_24900,N_24769);
or UO_476 (O_476,N_24705,N_24887);
nor UO_477 (O_477,N_24609,N_24782);
or UO_478 (O_478,N_24769,N_24766);
nand UO_479 (O_479,N_24684,N_24770);
or UO_480 (O_480,N_24873,N_24866);
nor UO_481 (O_481,N_24806,N_24499);
and UO_482 (O_482,N_24580,N_24651);
nand UO_483 (O_483,N_24710,N_24464);
nor UO_484 (O_484,N_24489,N_24700);
and UO_485 (O_485,N_24660,N_24714);
and UO_486 (O_486,N_24816,N_24743);
nor UO_487 (O_487,N_24424,N_24926);
and UO_488 (O_488,N_24485,N_24800);
nand UO_489 (O_489,N_24612,N_24923);
or UO_490 (O_490,N_24794,N_24507);
nor UO_491 (O_491,N_24998,N_24569);
or UO_492 (O_492,N_24953,N_24688);
nand UO_493 (O_493,N_24838,N_24439);
nand UO_494 (O_494,N_24612,N_24853);
nor UO_495 (O_495,N_24476,N_24990);
nand UO_496 (O_496,N_24775,N_24806);
and UO_497 (O_497,N_24384,N_24718);
nor UO_498 (O_498,N_24438,N_24799);
nand UO_499 (O_499,N_24832,N_24951);
nor UO_500 (O_500,N_24700,N_24385);
or UO_501 (O_501,N_24680,N_24913);
nor UO_502 (O_502,N_24503,N_24758);
nand UO_503 (O_503,N_24412,N_24638);
and UO_504 (O_504,N_24986,N_24893);
xnor UO_505 (O_505,N_24672,N_24819);
xor UO_506 (O_506,N_24850,N_24671);
or UO_507 (O_507,N_24607,N_24477);
or UO_508 (O_508,N_24569,N_24677);
and UO_509 (O_509,N_24527,N_24412);
nand UO_510 (O_510,N_24777,N_24992);
or UO_511 (O_511,N_24720,N_24578);
nor UO_512 (O_512,N_24488,N_24447);
or UO_513 (O_513,N_24759,N_24705);
xor UO_514 (O_514,N_24925,N_24526);
nor UO_515 (O_515,N_24986,N_24732);
nand UO_516 (O_516,N_24879,N_24933);
nand UO_517 (O_517,N_24488,N_24923);
xor UO_518 (O_518,N_24834,N_24913);
nor UO_519 (O_519,N_24797,N_24535);
or UO_520 (O_520,N_24706,N_24578);
and UO_521 (O_521,N_24421,N_24697);
nand UO_522 (O_522,N_24705,N_24725);
xor UO_523 (O_523,N_24684,N_24756);
xor UO_524 (O_524,N_24477,N_24869);
nand UO_525 (O_525,N_24947,N_24935);
nand UO_526 (O_526,N_24999,N_24791);
xor UO_527 (O_527,N_24713,N_24490);
xor UO_528 (O_528,N_24433,N_24857);
or UO_529 (O_529,N_24905,N_24727);
or UO_530 (O_530,N_24584,N_24539);
and UO_531 (O_531,N_24447,N_24461);
xor UO_532 (O_532,N_24722,N_24614);
or UO_533 (O_533,N_24715,N_24643);
or UO_534 (O_534,N_24636,N_24895);
nand UO_535 (O_535,N_24887,N_24818);
nand UO_536 (O_536,N_24990,N_24927);
nand UO_537 (O_537,N_24628,N_24754);
and UO_538 (O_538,N_24975,N_24900);
nor UO_539 (O_539,N_24977,N_24570);
and UO_540 (O_540,N_24621,N_24748);
and UO_541 (O_541,N_24766,N_24689);
or UO_542 (O_542,N_24603,N_24868);
xor UO_543 (O_543,N_24520,N_24540);
xnor UO_544 (O_544,N_24561,N_24389);
nand UO_545 (O_545,N_24483,N_24513);
xor UO_546 (O_546,N_24550,N_24599);
xor UO_547 (O_547,N_24847,N_24873);
nand UO_548 (O_548,N_24448,N_24612);
nand UO_549 (O_549,N_24937,N_24603);
xor UO_550 (O_550,N_24927,N_24807);
or UO_551 (O_551,N_24428,N_24442);
xor UO_552 (O_552,N_24619,N_24487);
nor UO_553 (O_553,N_24451,N_24763);
xor UO_554 (O_554,N_24811,N_24698);
nor UO_555 (O_555,N_24752,N_24525);
and UO_556 (O_556,N_24546,N_24748);
xor UO_557 (O_557,N_24944,N_24834);
or UO_558 (O_558,N_24932,N_24629);
and UO_559 (O_559,N_24715,N_24818);
xor UO_560 (O_560,N_24531,N_24780);
and UO_561 (O_561,N_24879,N_24723);
xnor UO_562 (O_562,N_24726,N_24658);
nor UO_563 (O_563,N_24464,N_24926);
nor UO_564 (O_564,N_24420,N_24775);
xnor UO_565 (O_565,N_24781,N_24415);
nor UO_566 (O_566,N_24642,N_24747);
xnor UO_567 (O_567,N_24722,N_24602);
nor UO_568 (O_568,N_24478,N_24794);
and UO_569 (O_569,N_24446,N_24733);
or UO_570 (O_570,N_24531,N_24397);
nand UO_571 (O_571,N_24579,N_24778);
and UO_572 (O_572,N_24796,N_24421);
xnor UO_573 (O_573,N_24775,N_24929);
or UO_574 (O_574,N_24673,N_24545);
nor UO_575 (O_575,N_24530,N_24823);
or UO_576 (O_576,N_24939,N_24641);
or UO_577 (O_577,N_24613,N_24670);
nor UO_578 (O_578,N_24808,N_24771);
or UO_579 (O_579,N_24563,N_24866);
nor UO_580 (O_580,N_24438,N_24762);
nand UO_581 (O_581,N_24865,N_24514);
or UO_582 (O_582,N_24702,N_24869);
and UO_583 (O_583,N_24509,N_24952);
xnor UO_584 (O_584,N_24859,N_24381);
xnor UO_585 (O_585,N_24951,N_24834);
and UO_586 (O_586,N_24546,N_24737);
xor UO_587 (O_587,N_24819,N_24527);
nand UO_588 (O_588,N_24814,N_24475);
xor UO_589 (O_589,N_24927,N_24842);
nor UO_590 (O_590,N_24948,N_24429);
nor UO_591 (O_591,N_24903,N_24665);
or UO_592 (O_592,N_24914,N_24691);
nand UO_593 (O_593,N_24450,N_24688);
xnor UO_594 (O_594,N_24804,N_24637);
nand UO_595 (O_595,N_24719,N_24603);
nor UO_596 (O_596,N_24903,N_24721);
xnor UO_597 (O_597,N_24507,N_24397);
and UO_598 (O_598,N_24392,N_24696);
nor UO_599 (O_599,N_24834,N_24765);
or UO_600 (O_600,N_24839,N_24638);
nand UO_601 (O_601,N_24465,N_24633);
xnor UO_602 (O_602,N_24548,N_24939);
nor UO_603 (O_603,N_24654,N_24566);
xnor UO_604 (O_604,N_24946,N_24554);
and UO_605 (O_605,N_24513,N_24416);
nand UO_606 (O_606,N_24464,N_24542);
xor UO_607 (O_607,N_24599,N_24921);
and UO_608 (O_608,N_24407,N_24616);
nand UO_609 (O_609,N_24427,N_24786);
and UO_610 (O_610,N_24735,N_24480);
or UO_611 (O_611,N_24979,N_24945);
and UO_612 (O_612,N_24428,N_24437);
xor UO_613 (O_613,N_24536,N_24879);
or UO_614 (O_614,N_24755,N_24519);
xor UO_615 (O_615,N_24428,N_24869);
or UO_616 (O_616,N_24498,N_24770);
nor UO_617 (O_617,N_24988,N_24502);
nand UO_618 (O_618,N_24737,N_24485);
and UO_619 (O_619,N_24972,N_24401);
or UO_620 (O_620,N_24435,N_24838);
and UO_621 (O_621,N_24707,N_24808);
and UO_622 (O_622,N_24816,N_24911);
xor UO_623 (O_623,N_24830,N_24734);
or UO_624 (O_624,N_24619,N_24477);
xor UO_625 (O_625,N_24603,N_24397);
nor UO_626 (O_626,N_24584,N_24881);
nor UO_627 (O_627,N_24836,N_24917);
xnor UO_628 (O_628,N_24622,N_24795);
nand UO_629 (O_629,N_24790,N_24979);
xnor UO_630 (O_630,N_24617,N_24608);
or UO_631 (O_631,N_24425,N_24684);
nand UO_632 (O_632,N_24669,N_24504);
and UO_633 (O_633,N_24970,N_24679);
nand UO_634 (O_634,N_24823,N_24719);
or UO_635 (O_635,N_24391,N_24877);
or UO_636 (O_636,N_24862,N_24395);
xor UO_637 (O_637,N_24992,N_24855);
nor UO_638 (O_638,N_24768,N_24989);
or UO_639 (O_639,N_24917,N_24419);
and UO_640 (O_640,N_24964,N_24659);
xor UO_641 (O_641,N_24978,N_24533);
nand UO_642 (O_642,N_24581,N_24651);
nand UO_643 (O_643,N_24674,N_24930);
nand UO_644 (O_644,N_24739,N_24619);
nand UO_645 (O_645,N_24593,N_24676);
and UO_646 (O_646,N_24404,N_24559);
nand UO_647 (O_647,N_24654,N_24406);
nor UO_648 (O_648,N_24787,N_24385);
or UO_649 (O_649,N_24511,N_24838);
or UO_650 (O_650,N_24921,N_24895);
and UO_651 (O_651,N_24449,N_24632);
xnor UO_652 (O_652,N_24513,N_24893);
nand UO_653 (O_653,N_24676,N_24660);
nand UO_654 (O_654,N_24394,N_24434);
xnor UO_655 (O_655,N_24800,N_24893);
nand UO_656 (O_656,N_24478,N_24731);
and UO_657 (O_657,N_24783,N_24646);
and UO_658 (O_658,N_24963,N_24869);
and UO_659 (O_659,N_24560,N_24665);
or UO_660 (O_660,N_24954,N_24711);
nor UO_661 (O_661,N_24920,N_24651);
and UO_662 (O_662,N_24906,N_24978);
nor UO_663 (O_663,N_24515,N_24796);
and UO_664 (O_664,N_24881,N_24382);
or UO_665 (O_665,N_24417,N_24623);
nand UO_666 (O_666,N_24527,N_24695);
xnor UO_667 (O_667,N_24879,N_24680);
or UO_668 (O_668,N_24813,N_24650);
and UO_669 (O_669,N_24663,N_24638);
xor UO_670 (O_670,N_24861,N_24414);
nor UO_671 (O_671,N_24722,N_24535);
nor UO_672 (O_672,N_24707,N_24891);
and UO_673 (O_673,N_24933,N_24673);
and UO_674 (O_674,N_24849,N_24537);
and UO_675 (O_675,N_24658,N_24381);
nand UO_676 (O_676,N_24742,N_24557);
nor UO_677 (O_677,N_24817,N_24823);
and UO_678 (O_678,N_24849,N_24559);
and UO_679 (O_679,N_24749,N_24648);
nand UO_680 (O_680,N_24706,N_24428);
xnor UO_681 (O_681,N_24393,N_24586);
xor UO_682 (O_682,N_24595,N_24412);
or UO_683 (O_683,N_24653,N_24616);
xnor UO_684 (O_684,N_24927,N_24558);
nand UO_685 (O_685,N_24693,N_24377);
nand UO_686 (O_686,N_24385,N_24408);
nor UO_687 (O_687,N_24850,N_24943);
and UO_688 (O_688,N_24700,N_24634);
or UO_689 (O_689,N_24967,N_24666);
nor UO_690 (O_690,N_24810,N_24974);
xnor UO_691 (O_691,N_24693,N_24835);
nor UO_692 (O_692,N_24954,N_24655);
xnor UO_693 (O_693,N_24858,N_24585);
or UO_694 (O_694,N_24658,N_24920);
and UO_695 (O_695,N_24574,N_24640);
and UO_696 (O_696,N_24579,N_24477);
and UO_697 (O_697,N_24814,N_24421);
xnor UO_698 (O_698,N_24624,N_24437);
or UO_699 (O_699,N_24847,N_24986);
nand UO_700 (O_700,N_24991,N_24598);
nand UO_701 (O_701,N_24887,N_24630);
nor UO_702 (O_702,N_24792,N_24380);
nor UO_703 (O_703,N_24812,N_24419);
nand UO_704 (O_704,N_24386,N_24524);
nor UO_705 (O_705,N_24602,N_24756);
xnor UO_706 (O_706,N_24735,N_24935);
nand UO_707 (O_707,N_24881,N_24722);
nor UO_708 (O_708,N_24942,N_24681);
and UO_709 (O_709,N_24603,N_24614);
nor UO_710 (O_710,N_24576,N_24669);
or UO_711 (O_711,N_24412,N_24569);
or UO_712 (O_712,N_24816,N_24871);
or UO_713 (O_713,N_24413,N_24611);
or UO_714 (O_714,N_24655,N_24493);
or UO_715 (O_715,N_24529,N_24976);
or UO_716 (O_716,N_24910,N_24709);
nor UO_717 (O_717,N_24455,N_24382);
xor UO_718 (O_718,N_24763,N_24700);
and UO_719 (O_719,N_24838,N_24908);
nor UO_720 (O_720,N_24533,N_24868);
nor UO_721 (O_721,N_24973,N_24489);
xor UO_722 (O_722,N_24568,N_24472);
xnor UO_723 (O_723,N_24484,N_24377);
and UO_724 (O_724,N_24379,N_24551);
xor UO_725 (O_725,N_24894,N_24996);
or UO_726 (O_726,N_24446,N_24903);
xor UO_727 (O_727,N_24527,N_24499);
nor UO_728 (O_728,N_24375,N_24820);
and UO_729 (O_729,N_24725,N_24762);
xnor UO_730 (O_730,N_24499,N_24530);
and UO_731 (O_731,N_24991,N_24850);
or UO_732 (O_732,N_24890,N_24786);
or UO_733 (O_733,N_24958,N_24876);
xnor UO_734 (O_734,N_24995,N_24495);
xor UO_735 (O_735,N_24416,N_24861);
or UO_736 (O_736,N_24826,N_24714);
nand UO_737 (O_737,N_24864,N_24466);
or UO_738 (O_738,N_24582,N_24689);
xor UO_739 (O_739,N_24952,N_24569);
or UO_740 (O_740,N_24431,N_24591);
nor UO_741 (O_741,N_24730,N_24512);
and UO_742 (O_742,N_24670,N_24665);
nor UO_743 (O_743,N_24540,N_24648);
nor UO_744 (O_744,N_24907,N_24658);
nand UO_745 (O_745,N_24607,N_24716);
nand UO_746 (O_746,N_24531,N_24846);
xnor UO_747 (O_747,N_24386,N_24911);
nand UO_748 (O_748,N_24886,N_24500);
nand UO_749 (O_749,N_24627,N_24930);
or UO_750 (O_750,N_24515,N_24727);
nor UO_751 (O_751,N_24903,N_24984);
and UO_752 (O_752,N_24605,N_24867);
nor UO_753 (O_753,N_24511,N_24891);
and UO_754 (O_754,N_24735,N_24966);
nor UO_755 (O_755,N_24581,N_24850);
nand UO_756 (O_756,N_24756,N_24835);
or UO_757 (O_757,N_24573,N_24445);
and UO_758 (O_758,N_24605,N_24572);
or UO_759 (O_759,N_24739,N_24861);
or UO_760 (O_760,N_24494,N_24668);
xor UO_761 (O_761,N_24855,N_24763);
xor UO_762 (O_762,N_24644,N_24611);
xnor UO_763 (O_763,N_24972,N_24592);
and UO_764 (O_764,N_24453,N_24897);
or UO_765 (O_765,N_24775,N_24750);
nand UO_766 (O_766,N_24672,N_24487);
nor UO_767 (O_767,N_24684,N_24602);
nand UO_768 (O_768,N_24469,N_24791);
nor UO_769 (O_769,N_24655,N_24931);
nand UO_770 (O_770,N_24767,N_24494);
or UO_771 (O_771,N_24970,N_24460);
or UO_772 (O_772,N_24769,N_24930);
xor UO_773 (O_773,N_24910,N_24762);
nand UO_774 (O_774,N_24832,N_24698);
xor UO_775 (O_775,N_24396,N_24630);
xor UO_776 (O_776,N_24833,N_24431);
and UO_777 (O_777,N_24557,N_24788);
and UO_778 (O_778,N_24469,N_24806);
nand UO_779 (O_779,N_24382,N_24884);
xor UO_780 (O_780,N_24397,N_24972);
nor UO_781 (O_781,N_24733,N_24638);
and UO_782 (O_782,N_24397,N_24439);
and UO_783 (O_783,N_24893,N_24714);
or UO_784 (O_784,N_24997,N_24560);
xor UO_785 (O_785,N_24590,N_24418);
nand UO_786 (O_786,N_24720,N_24952);
and UO_787 (O_787,N_24569,N_24558);
xnor UO_788 (O_788,N_24859,N_24921);
nor UO_789 (O_789,N_24590,N_24584);
xnor UO_790 (O_790,N_24911,N_24453);
or UO_791 (O_791,N_24390,N_24998);
nand UO_792 (O_792,N_24443,N_24915);
xnor UO_793 (O_793,N_24492,N_24429);
nand UO_794 (O_794,N_24910,N_24905);
nand UO_795 (O_795,N_24884,N_24503);
xor UO_796 (O_796,N_24893,N_24950);
or UO_797 (O_797,N_24642,N_24769);
or UO_798 (O_798,N_24725,N_24720);
and UO_799 (O_799,N_24842,N_24883);
nand UO_800 (O_800,N_24998,N_24444);
xnor UO_801 (O_801,N_24487,N_24486);
nand UO_802 (O_802,N_24644,N_24630);
xor UO_803 (O_803,N_24964,N_24995);
and UO_804 (O_804,N_24394,N_24677);
or UO_805 (O_805,N_24844,N_24706);
nor UO_806 (O_806,N_24637,N_24659);
or UO_807 (O_807,N_24840,N_24725);
and UO_808 (O_808,N_24456,N_24707);
nand UO_809 (O_809,N_24424,N_24563);
xnor UO_810 (O_810,N_24476,N_24526);
or UO_811 (O_811,N_24414,N_24797);
nor UO_812 (O_812,N_24996,N_24913);
nor UO_813 (O_813,N_24902,N_24652);
or UO_814 (O_814,N_24669,N_24724);
or UO_815 (O_815,N_24805,N_24587);
or UO_816 (O_816,N_24783,N_24375);
nor UO_817 (O_817,N_24401,N_24495);
xor UO_818 (O_818,N_24777,N_24983);
xor UO_819 (O_819,N_24756,N_24988);
or UO_820 (O_820,N_24400,N_24377);
nand UO_821 (O_821,N_24379,N_24386);
or UO_822 (O_822,N_24912,N_24505);
xnor UO_823 (O_823,N_24475,N_24798);
xor UO_824 (O_824,N_24626,N_24902);
nor UO_825 (O_825,N_24678,N_24598);
nand UO_826 (O_826,N_24401,N_24934);
or UO_827 (O_827,N_24807,N_24614);
nand UO_828 (O_828,N_24758,N_24401);
or UO_829 (O_829,N_24869,N_24405);
or UO_830 (O_830,N_24657,N_24863);
xnor UO_831 (O_831,N_24786,N_24698);
nor UO_832 (O_832,N_24948,N_24749);
and UO_833 (O_833,N_24650,N_24756);
and UO_834 (O_834,N_24406,N_24640);
xor UO_835 (O_835,N_24536,N_24680);
or UO_836 (O_836,N_24670,N_24772);
and UO_837 (O_837,N_24475,N_24480);
nor UO_838 (O_838,N_24512,N_24376);
xnor UO_839 (O_839,N_24488,N_24696);
nand UO_840 (O_840,N_24593,N_24843);
nor UO_841 (O_841,N_24803,N_24893);
xnor UO_842 (O_842,N_24685,N_24674);
and UO_843 (O_843,N_24962,N_24719);
and UO_844 (O_844,N_24544,N_24611);
nor UO_845 (O_845,N_24676,N_24945);
xnor UO_846 (O_846,N_24392,N_24827);
or UO_847 (O_847,N_24867,N_24489);
or UO_848 (O_848,N_24861,N_24749);
nor UO_849 (O_849,N_24546,N_24629);
xnor UO_850 (O_850,N_24824,N_24598);
xor UO_851 (O_851,N_24661,N_24475);
or UO_852 (O_852,N_24406,N_24651);
nand UO_853 (O_853,N_24564,N_24488);
nand UO_854 (O_854,N_24839,N_24836);
and UO_855 (O_855,N_24409,N_24712);
or UO_856 (O_856,N_24517,N_24835);
nor UO_857 (O_857,N_24916,N_24684);
nor UO_858 (O_858,N_24694,N_24534);
xnor UO_859 (O_859,N_24576,N_24525);
xor UO_860 (O_860,N_24964,N_24739);
or UO_861 (O_861,N_24378,N_24517);
or UO_862 (O_862,N_24901,N_24756);
xnor UO_863 (O_863,N_24411,N_24817);
nand UO_864 (O_864,N_24774,N_24886);
xnor UO_865 (O_865,N_24769,N_24552);
or UO_866 (O_866,N_24433,N_24727);
or UO_867 (O_867,N_24538,N_24662);
and UO_868 (O_868,N_24647,N_24899);
or UO_869 (O_869,N_24769,N_24595);
xnor UO_870 (O_870,N_24570,N_24489);
and UO_871 (O_871,N_24597,N_24516);
and UO_872 (O_872,N_24778,N_24604);
nand UO_873 (O_873,N_24586,N_24502);
xnor UO_874 (O_874,N_24601,N_24771);
nor UO_875 (O_875,N_24914,N_24684);
or UO_876 (O_876,N_24702,N_24835);
and UO_877 (O_877,N_24667,N_24908);
nand UO_878 (O_878,N_24617,N_24553);
and UO_879 (O_879,N_24526,N_24883);
nor UO_880 (O_880,N_24747,N_24683);
nor UO_881 (O_881,N_24947,N_24758);
nand UO_882 (O_882,N_24638,N_24563);
and UO_883 (O_883,N_24852,N_24620);
xor UO_884 (O_884,N_24667,N_24944);
xor UO_885 (O_885,N_24614,N_24693);
nor UO_886 (O_886,N_24777,N_24755);
nand UO_887 (O_887,N_24930,N_24875);
and UO_888 (O_888,N_24962,N_24821);
nor UO_889 (O_889,N_24568,N_24728);
nor UO_890 (O_890,N_24402,N_24892);
or UO_891 (O_891,N_24978,N_24546);
nor UO_892 (O_892,N_24624,N_24645);
nand UO_893 (O_893,N_24610,N_24468);
or UO_894 (O_894,N_24680,N_24421);
or UO_895 (O_895,N_24494,N_24568);
xnor UO_896 (O_896,N_24625,N_24544);
xor UO_897 (O_897,N_24556,N_24408);
and UO_898 (O_898,N_24445,N_24998);
xor UO_899 (O_899,N_24987,N_24465);
or UO_900 (O_900,N_24754,N_24707);
nor UO_901 (O_901,N_24804,N_24990);
or UO_902 (O_902,N_24879,N_24926);
nor UO_903 (O_903,N_24816,N_24937);
nand UO_904 (O_904,N_24982,N_24460);
nor UO_905 (O_905,N_24544,N_24703);
or UO_906 (O_906,N_24707,N_24533);
nand UO_907 (O_907,N_24474,N_24556);
and UO_908 (O_908,N_24852,N_24710);
or UO_909 (O_909,N_24781,N_24959);
nand UO_910 (O_910,N_24997,N_24486);
nand UO_911 (O_911,N_24499,N_24579);
nor UO_912 (O_912,N_24555,N_24738);
nor UO_913 (O_913,N_24974,N_24510);
xnor UO_914 (O_914,N_24780,N_24755);
or UO_915 (O_915,N_24783,N_24622);
nor UO_916 (O_916,N_24431,N_24902);
and UO_917 (O_917,N_24588,N_24813);
nor UO_918 (O_918,N_24791,N_24445);
or UO_919 (O_919,N_24508,N_24916);
or UO_920 (O_920,N_24710,N_24600);
xor UO_921 (O_921,N_24502,N_24643);
xor UO_922 (O_922,N_24582,N_24439);
nor UO_923 (O_923,N_24955,N_24550);
nor UO_924 (O_924,N_24663,N_24744);
or UO_925 (O_925,N_24422,N_24728);
and UO_926 (O_926,N_24456,N_24379);
nand UO_927 (O_927,N_24620,N_24937);
xnor UO_928 (O_928,N_24818,N_24428);
and UO_929 (O_929,N_24480,N_24658);
and UO_930 (O_930,N_24608,N_24388);
nor UO_931 (O_931,N_24844,N_24986);
xor UO_932 (O_932,N_24747,N_24625);
or UO_933 (O_933,N_24976,N_24980);
xnor UO_934 (O_934,N_24921,N_24647);
and UO_935 (O_935,N_24457,N_24577);
and UO_936 (O_936,N_24554,N_24466);
xnor UO_937 (O_937,N_24765,N_24684);
and UO_938 (O_938,N_24525,N_24886);
or UO_939 (O_939,N_24644,N_24712);
or UO_940 (O_940,N_24739,N_24390);
xor UO_941 (O_941,N_24923,N_24731);
or UO_942 (O_942,N_24881,N_24473);
xor UO_943 (O_943,N_24999,N_24377);
and UO_944 (O_944,N_24753,N_24812);
nor UO_945 (O_945,N_24727,N_24414);
and UO_946 (O_946,N_24942,N_24522);
and UO_947 (O_947,N_24420,N_24440);
nand UO_948 (O_948,N_24576,N_24455);
nor UO_949 (O_949,N_24783,N_24572);
nor UO_950 (O_950,N_24554,N_24644);
nand UO_951 (O_951,N_24631,N_24486);
nand UO_952 (O_952,N_24864,N_24846);
nor UO_953 (O_953,N_24725,N_24566);
nand UO_954 (O_954,N_24799,N_24386);
and UO_955 (O_955,N_24576,N_24550);
and UO_956 (O_956,N_24841,N_24843);
nand UO_957 (O_957,N_24734,N_24512);
nor UO_958 (O_958,N_24394,N_24755);
nand UO_959 (O_959,N_24846,N_24376);
nor UO_960 (O_960,N_24713,N_24639);
nor UO_961 (O_961,N_24906,N_24540);
nor UO_962 (O_962,N_24741,N_24663);
xor UO_963 (O_963,N_24457,N_24589);
or UO_964 (O_964,N_24470,N_24951);
nor UO_965 (O_965,N_24503,N_24511);
and UO_966 (O_966,N_24912,N_24711);
nand UO_967 (O_967,N_24888,N_24872);
xnor UO_968 (O_968,N_24959,N_24605);
xnor UO_969 (O_969,N_24578,N_24648);
nor UO_970 (O_970,N_24808,N_24716);
and UO_971 (O_971,N_24382,N_24704);
and UO_972 (O_972,N_24903,N_24583);
xor UO_973 (O_973,N_24461,N_24781);
xor UO_974 (O_974,N_24546,N_24711);
and UO_975 (O_975,N_24435,N_24451);
nand UO_976 (O_976,N_24419,N_24867);
and UO_977 (O_977,N_24918,N_24582);
nor UO_978 (O_978,N_24776,N_24416);
or UO_979 (O_979,N_24968,N_24719);
and UO_980 (O_980,N_24811,N_24907);
or UO_981 (O_981,N_24492,N_24780);
or UO_982 (O_982,N_24507,N_24968);
or UO_983 (O_983,N_24921,N_24958);
and UO_984 (O_984,N_24720,N_24624);
nor UO_985 (O_985,N_24838,N_24550);
and UO_986 (O_986,N_24470,N_24691);
and UO_987 (O_987,N_24476,N_24792);
or UO_988 (O_988,N_24516,N_24985);
and UO_989 (O_989,N_24835,N_24820);
nand UO_990 (O_990,N_24874,N_24876);
and UO_991 (O_991,N_24751,N_24831);
nand UO_992 (O_992,N_24852,N_24756);
and UO_993 (O_993,N_24561,N_24774);
nand UO_994 (O_994,N_24609,N_24827);
and UO_995 (O_995,N_24692,N_24703);
or UO_996 (O_996,N_24932,N_24842);
xnor UO_997 (O_997,N_24615,N_24545);
xnor UO_998 (O_998,N_24924,N_24814);
and UO_999 (O_999,N_24395,N_24416);
nor UO_1000 (O_1000,N_24407,N_24557);
and UO_1001 (O_1001,N_24420,N_24924);
or UO_1002 (O_1002,N_24947,N_24729);
or UO_1003 (O_1003,N_24502,N_24791);
nor UO_1004 (O_1004,N_24795,N_24738);
or UO_1005 (O_1005,N_24562,N_24608);
xor UO_1006 (O_1006,N_24990,N_24492);
xnor UO_1007 (O_1007,N_24394,N_24944);
nand UO_1008 (O_1008,N_24515,N_24842);
and UO_1009 (O_1009,N_24898,N_24968);
and UO_1010 (O_1010,N_24843,N_24417);
nor UO_1011 (O_1011,N_24507,N_24833);
xnor UO_1012 (O_1012,N_24848,N_24741);
or UO_1013 (O_1013,N_24956,N_24839);
nand UO_1014 (O_1014,N_24502,N_24854);
nor UO_1015 (O_1015,N_24902,N_24549);
nor UO_1016 (O_1016,N_24947,N_24897);
and UO_1017 (O_1017,N_24676,N_24540);
xor UO_1018 (O_1018,N_24954,N_24391);
nand UO_1019 (O_1019,N_24615,N_24661);
xor UO_1020 (O_1020,N_24434,N_24592);
nand UO_1021 (O_1021,N_24513,N_24889);
xor UO_1022 (O_1022,N_24628,N_24467);
or UO_1023 (O_1023,N_24724,N_24389);
nand UO_1024 (O_1024,N_24605,N_24676);
nor UO_1025 (O_1025,N_24710,N_24681);
nand UO_1026 (O_1026,N_24867,N_24955);
nor UO_1027 (O_1027,N_24605,N_24571);
nor UO_1028 (O_1028,N_24998,N_24423);
and UO_1029 (O_1029,N_24804,N_24875);
xnor UO_1030 (O_1030,N_24781,N_24595);
and UO_1031 (O_1031,N_24651,N_24865);
nand UO_1032 (O_1032,N_24646,N_24812);
nand UO_1033 (O_1033,N_24551,N_24559);
nor UO_1034 (O_1034,N_24631,N_24468);
or UO_1035 (O_1035,N_24496,N_24594);
xnor UO_1036 (O_1036,N_24850,N_24493);
nor UO_1037 (O_1037,N_24532,N_24868);
nand UO_1038 (O_1038,N_24834,N_24499);
nand UO_1039 (O_1039,N_24463,N_24415);
nor UO_1040 (O_1040,N_24904,N_24938);
nand UO_1041 (O_1041,N_24689,N_24473);
and UO_1042 (O_1042,N_24523,N_24560);
and UO_1043 (O_1043,N_24465,N_24892);
nand UO_1044 (O_1044,N_24667,N_24658);
or UO_1045 (O_1045,N_24599,N_24530);
xnor UO_1046 (O_1046,N_24722,N_24771);
nand UO_1047 (O_1047,N_24450,N_24605);
xnor UO_1048 (O_1048,N_24413,N_24617);
or UO_1049 (O_1049,N_24884,N_24560);
or UO_1050 (O_1050,N_24868,N_24466);
or UO_1051 (O_1051,N_24540,N_24432);
or UO_1052 (O_1052,N_24773,N_24832);
and UO_1053 (O_1053,N_24619,N_24551);
and UO_1054 (O_1054,N_24545,N_24956);
or UO_1055 (O_1055,N_24617,N_24959);
xor UO_1056 (O_1056,N_24655,N_24637);
nor UO_1057 (O_1057,N_24557,N_24966);
and UO_1058 (O_1058,N_24560,N_24955);
xor UO_1059 (O_1059,N_24541,N_24658);
nand UO_1060 (O_1060,N_24387,N_24747);
and UO_1061 (O_1061,N_24668,N_24392);
or UO_1062 (O_1062,N_24845,N_24978);
xnor UO_1063 (O_1063,N_24480,N_24561);
or UO_1064 (O_1064,N_24673,N_24489);
and UO_1065 (O_1065,N_24668,N_24640);
and UO_1066 (O_1066,N_24997,N_24464);
and UO_1067 (O_1067,N_24861,N_24799);
and UO_1068 (O_1068,N_24872,N_24399);
nor UO_1069 (O_1069,N_24595,N_24929);
and UO_1070 (O_1070,N_24993,N_24524);
and UO_1071 (O_1071,N_24983,N_24864);
and UO_1072 (O_1072,N_24694,N_24568);
nor UO_1073 (O_1073,N_24675,N_24536);
nand UO_1074 (O_1074,N_24997,N_24387);
nand UO_1075 (O_1075,N_24679,N_24776);
or UO_1076 (O_1076,N_24524,N_24745);
nand UO_1077 (O_1077,N_24811,N_24832);
nand UO_1078 (O_1078,N_24750,N_24967);
nand UO_1079 (O_1079,N_24702,N_24843);
nand UO_1080 (O_1080,N_24486,N_24882);
xor UO_1081 (O_1081,N_24965,N_24937);
and UO_1082 (O_1082,N_24440,N_24603);
or UO_1083 (O_1083,N_24732,N_24799);
nor UO_1084 (O_1084,N_24604,N_24696);
nor UO_1085 (O_1085,N_24553,N_24392);
or UO_1086 (O_1086,N_24987,N_24719);
and UO_1087 (O_1087,N_24614,N_24905);
nor UO_1088 (O_1088,N_24892,N_24602);
nor UO_1089 (O_1089,N_24726,N_24780);
xor UO_1090 (O_1090,N_24982,N_24783);
and UO_1091 (O_1091,N_24935,N_24671);
nand UO_1092 (O_1092,N_24442,N_24580);
nor UO_1093 (O_1093,N_24691,N_24737);
or UO_1094 (O_1094,N_24618,N_24627);
nand UO_1095 (O_1095,N_24540,N_24896);
nor UO_1096 (O_1096,N_24993,N_24994);
and UO_1097 (O_1097,N_24873,N_24832);
and UO_1098 (O_1098,N_24908,N_24767);
nand UO_1099 (O_1099,N_24579,N_24892);
or UO_1100 (O_1100,N_24737,N_24738);
or UO_1101 (O_1101,N_24435,N_24913);
or UO_1102 (O_1102,N_24913,N_24535);
xor UO_1103 (O_1103,N_24932,N_24566);
and UO_1104 (O_1104,N_24392,N_24425);
nand UO_1105 (O_1105,N_24394,N_24774);
and UO_1106 (O_1106,N_24629,N_24648);
nand UO_1107 (O_1107,N_24845,N_24957);
nor UO_1108 (O_1108,N_24984,N_24945);
or UO_1109 (O_1109,N_24867,N_24993);
nor UO_1110 (O_1110,N_24769,N_24688);
nor UO_1111 (O_1111,N_24723,N_24535);
nand UO_1112 (O_1112,N_24496,N_24980);
and UO_1113 (O_1113,N_24668,N_24404);
nand UO_1114 (O_1114,N_24998,N_24720);
xor UO_1115 (O_1115,N_24921,N_24798);
and UO_1116 (O_1116,N_24504,N_24560);
xor UO_1117 (O_1117,N_24648,N_24647);
nand UO_1118 (O_1118,N_24472,N_24821);
xnor UO_1119 (O_1119,N_24445,N_24463);
nor UO_1120 (O_1120,N_24471,N_24605);
nand UO_1121 (O_1121,N_24945,N_24792);
nand UO_1122 (O_1122,N_24380,N_24554);
and UO_1123 (O_1123,N_24648,N_24953);
or UO_1124 (O_1124,N_24878,N_24615);
and UO_1125 (O_1125,N_24988,N_24625);
or UO_1126 (O_1126,N_24549,N_24672);
nand UO_1127 (O_1127,N_24457,N_24533);
nor UO_1128 (O_1128,N_24382,N_24821);
nand UO_1129 (O_1129,N_24782,N_24733);
xnor UO_1130 (O_1130,N_24473,N_24574);
nand UO_1131 (O_1131,N_24691,N_24478);
and UO_1132 (O_1132,N_24434,N_24803);
or UO_1133 (O_1133,N_24377,N_24637);
or UO_1134 (O_1134,N_24837,N_24497);
and UO_1135 (O_1135,N_24982,N_24829);
xnor UO_1136 (O_1136,N_24741,N_24472);
nand UO_1137 (O_1137,N_24889,N_24594);
nand UO_1138 (O_1138,N_24942,N_24503);
and UO_1139 (O_1139,N_24955,N_24449);
xor UO_1140 (O_1140,N_24690,N_24591);
nor UO_1141 (O_1141,N_24960,N_24909);
nor UO_1142 (O_1142,N_24481,N_24667);
xnor UO_1143 (O_1143,N_24970,N_24855);
nand UO_1144 (O_1144,N_24392,N_24530);
nor UO_1145 (O_1145,N_24524,N_24474);
and UO_1146 (O_1146,N_24824,N_24557);
and UO_1147 (O_1147,N_24652,N_24702);
or UO_1148 (O_1148,N_24440,N_24954);
nand UO_1149 (O_1149,N_24959,N_24380);
nor UO_1150 (O_1150,N_24402,N_24769);
xnor UO_1151 (O_1151,N_24864,N_24860);
nor UO_1152 (O_1152,N_24905,N_24885);
and UO_1153 (O_1153,N_24402,N_24635);
or UO_1154 (O_1154,N_24550,N_24469);
xor UO_1155 (O_1155,N_24660,N_24782);
or UO_1156 (O_1156,N_24988,N_24699);
or UO_1157 (O_1157,N_24788,N_24919);
or UO_1158 (O_1158,N_24923,N_24433);
xnor UO_1159 (O_1159,N_24378,N_24646);
xor UO_1160 (O_1160,N_24691,N_24454);
or UO_1161 (O_1161,N_24798,N_24391);
xnor UO_1162 (O_1162,N_24926,N_24383);
xor UO_1163 (O_1163,N_24510,N_24461);
xnor UO_1164 (O_1164,N_24827,N_24954);
and UO_1165 (O_1165,N_24604,N_24825);
xor UO_1166 (O_1166,N_24580,N_24432);
nor UO_1167 (O_1167,N_24420,N_24586);
xnor UO_1168 (O_1168,N_24677,N_24920);
and UO_1169 (O_1169,N_24568,N_24724);
or UO_1170 (O_1170,N_24495,N_24655);
xnor UO_1171 (O_1171,N_24552,N_24793);
nand UO_1172 (O_1172,N_24957,N_24883);
nand UO_1173 (O_1173,N_24457,N_24834);
nor UO_1174 (O_1174,N_24717,N_24749);
and UO_1175 (O_1175,N_24726,N_24580);
or UO_1176 (O_1176,N_24454,N_24877);
nand UO_1177 (O_1177,N_24960,N_24575);
xor UO_1178 (O_1178,N_24565,N_24718);
xnor UO_1179 (O_1179,N_24800,N_24633);
nand UO_1180 (O_1180,N_24937,N_24602);
or UO_1181 (O_1181,N_24426,N_24499);
and UO_1182 (O_1182,N_24442,N_24985);
nor UO_1183 (O_1183,N_24705,N_24563);
xor UO_1184 (O_1184,N_24989,N_24963);
or UO_1185 (O_1185,N_24496,N_24696);
and UO_1186 (O_1186,N_24558,N_24378);
nor UO_1187 (O_1187,N_24804,N_24691);
or UO_1188 (O_1188,N_24747,N_24974);
or UO_1189 (O_1189,N_24600,N_24931);
and UO_1190 (O_1190,N_24491,N_24824);
nand UO_1191 (O_1191,N_24993,N_24961);
nor UO_1192 (O_1192,N_24636,N_24876);
xnor UO_1193 (O_1193,N_24497,N_24867);
or UO_1194 (O_1194,N_24401,N_24670);
xor UO_1195 (O_1195,N_24815,N_24388);
nand UO_1196 (O_1196,N_24408,N_24934);
nor UO_1197 (O_1197,N_24850,N_24712);
or UO_1198 (O_1198,N_24872,N_24936);
nor UO_1199 (O_1199,N_24532,N_24845);
and UO_1200 (O_1200,N_24736,N_24726);
nor UO_1201 (O_1201,N_24409,N_24580);
or UO_1202 (O_1202,N_24550,N_24530);
xor UO_1203 (O_1203,N_24466,N_24616);
and UO_1204 (O_1204,N_24686,N_24472);
xor UO_1205 (O_1205,N_24860,N_24668);
nor UO_1206 (O_1206,N_24552,N_24628);
nand UO_1207 (O_1207,N_24619,N_24707);
nor UO_1208 (O_1208,N_24728,N_24748);
xor UO_1209 (O_1209,N_24649,N_24658);
or UO_1210 (O_1210,N_24637,N_24664);
and UO_1211 (O_1211,N_24655,N_24895);
nand UO_1212 (O_1212,N_24507,N_24566);
or UO_1213 (O_1213,N_24830,N_24792);
and UO_1214 (O_1214,N_24450,N_24944);
nor UO_1215 (O_1215,N_24972,N_24551);
nand UO_1216 (O_1216,N_24974,N_24896);
xnor UO_1217 (O_1217,N_24863,N_24747);
xnor UO_1218 (O_1218,N_24903,N_24470);
and UO_1219 (O_1219,N_24763,N_24567);
xor UO_1220 (O_1220,N_24757,N_24564);
xor UO_1221 (O_1221,N_24399,N_24484);
nor UO_1222 (O_1222,N_24751,N_24655);
and UO_1223 (O_1223,N_24802,N_24502);
nor UO_1224 (O_1224,N_24779,N_24761);
nand UO_1225 (O_1225,N_24440,N_24788);
and UO_1226 (O_1226,N_24784,N_24439);
nor UO_1227 (O_1227,N_24957,N_24669);
nand UO_1228 (O_1228,N_24426,N_24487);
nand UO_1229 (O_1229,N_24690,N_24872);
nor UO_1230 (O_1230,N_24617,N_24960);
and UO_1231 (O_1231,N_24858,N_24496);
xor UO_1232 (O_1232,N_24436,N_24766);
nor UO_1233 (O_1233,N_24895,N_24766);
nor UO_1234 (O_1234,N_24826,N_24487);
and UO_1235 (O_1235,N_24938,N_24759);
xor UO_1236 (O_1236,N_24610,N_24572);
and UO_1237 (O_1237,N_24872,N_24569);
and UO_1238 (O_1238,N_24898,N_24819);
nand UO_1239 (O_1239,N_24844,N_24390);
xor UO_1240 (O_1240,N_24655,N_24382);
and UO_1241 (O_1241,N_24424,N_24698);
and UO_1242 (O_1242,N_24705,N_24668);
or UO_1243 (O_1243,N_24389,N_24413);
xor UO_1244 (O_1244,N_24734,N_24528);
nand UO_1245 (O_1245,N_24514,N_24771);
xor UO_1246 (O_1246,N_24675,N_24841);
xor UO_1247 (O_1247,N_24656,N_24668);
xor UO_1248 (O_1248,N_24791,N_24891);
or UO_1249 (O_1249,N_24996,N_24671);
or UO_1250 (O_1250,N_24711,N_24861);
or UO_1251 (O_1251,N_24495,N_24585);
nor UO_1252 (O_1252,N_24701,N_24449);
nand UO_1253 (O_1253,N_24459,N_24385);
nand UO_1254 (O_1254,N_24861,N_24766);
nand UO_1255 (O_1255,N_24716,N_24599);
nor UO_1256 (O_1256,N_24499,N_24756);
xor UO_1257 (O_1257,N_24505,N_24426);
nand UO_1258 (O_1258,N_24820,N_24846);
nand UO_1259 (O_1259,N_24557,N_24642);
or UO_1260 (O_1260,N_24813,N_24642);
nor UO_1261 (O_1261,N_24813,N_24682);
nor UO_1262 (O_1262,N_24558,N_24867);
or UO_1263 (O_1263,N_24415,N_24518);
or UO_1264 (O_1264,N_24505,N_24922);
nor UO_1265 (O_1265,N_24914,N_24594);
or UO_1266 (O_1266,N_24623,N_24692);
nand UO_1267 (O_1267,N_24765,N_24539);
or UO_1268 (O_1268,N_24942,N_24581);
nand UO_1269 (O_1269,N_24734,N_24707);
nor UO_1270 (O_1270,N_24414,N_24931);
and UO_1271 (O_1271,N_24753,N_24383);
xor UO_1272 (O_1272,N_24969,N_24878);
nand UO_1273 (O_1273,N_24386,N_24808);
nand UO_1274 (O_1274,N_24644,N_24845);
nor UO_1275 (O_1275,N_24555,N_24457);
and UO_1276 (O_1276,N_24491,N_24969);
xnor UO_1277 (O_1277,N_24901,N_24438);
xnor UO_1278 (O_1278,N_24641,N_24619);
xor UO_1279 (O_1279,N_24868,N_24837);
and UO_1280 (O_1280,N_24649,N_24811);
nor UO_1281 (O_1281,N_24702,N_24813);
nor UO_1282 (O_1282,N_24428,N_24523);
nand UO_1283 (O_1283,N_24401,N_24651);
or UO_1284 (O_1284,N_24421,N_24912);
xor UO_1285 (O_1285,N_24697,N_24701);
nand UO_1286 (O_1286,N_24803,N_24400);
nor UO_1287 (O_1287,N_24952,N_24986);
or UO_1288 (O_1288,N_24458,N_24530);
nand UO_1289 (O_1289,N_24510,N_24485);
nor UO_1290 (O_1290,N_24647,N_24450);
nand UO_1291 (O_1291,N_24614,N_24426);
nor UO_1292 (O_1292,N_24773,N_24957);
or UO_1293 (O_1293,N_24733,N_24686);
nand UO_1294 (O_1294,N_24601,N_24714);
nand UO_1295 (O_1295,N_24512,N_24964);
nor UO_1296 (O_1296,N_24378,N_24968);
nand UO_1297 (O_1297,N_24436,N_24917);
or UO_1298 (O_1298,N_24767,N_24710);
nand UO_1299 (O_1299,N_24763,N_24922);
xnor UO_1300 (O_1300,N_24533,N_24687);
nand UO_1301 (O_1301,N_24680,N_24638);
nand UO_1302 (O_1302,N_24853,N_24950);
or UO_1303 (O_1303,N_24607,N_24445);
or UO_1304 (O_1304,N_24761,N_24758);
nor UO_1305 (O_1305,N_24447,N_24756);
nor UO_1306 (O_1306,N_24837,N_24987);
xor UO_1307 (O_1307,N_24906,N_24466);
nand UO_1308 (O_1308,N_24591,N_24803);
xnor UO_1309 (O_1309,N_24449,N_24734);
xor UO_1310 (O_1310,N_24824,N_24514);
and UO_1311 (O_1311,N_24498,N_24517);
nor UO_1312 (O_1312,N_24859,N_24710);
nand UO_1313 (O_1313,N_24610,N_24451);
and UO_1314 (O_1314,N_24604,N_24930);
xnor UO_1315 (O_1315,N_24713,N_24894);
nor UO_1316 (O_1316,N_24706,N_24535);
xor UO_1317 (O_1317,N_24813,N_24995);
and UO_1318 (O_1318,N_24900,N_24949);
xnor UO_1319 (O_1319,N_24836,N_24441);
xor UO_1320 (O_1320,N_24584,N_24510);
xor UO_1321 (O_1321,N_24633,N_24985);
xor UO_1322 (O_1322,N_24892,N_24881);
and UO_1323 (O_1323,N_24926,N_24423);
or UO_1324 (O_1324,N_24946,N_24906);
nor UO_1325 (O_1325,N_24890,N_24539);
or UO_1326 (O_1326,N_24470,N_24532);
and UO_1327 (O_1327,N_24657,N_24631);
xnor UO_1328 (O_1328,N_24943,N_24825);
or UO_1329 (O_1329,N_24900,N_24625);
nand UO_1330 (O_1330,N_24741,N_24945);
nand UO_1331 (O_1331,N_24544,N_24733);
or UO_1332 (O_1332,N_24606,N_24463);
and UO_1333 (O_1333,N_24681,N_24810);
and UO_1334 (O_1334,N_24637,N_24580);
or UO_1335 (O_1335,N_24675,N_24925);
or UO_1336 (O_1336,N_24696,N_24806);
and UO_1337 (O_1337,N_24665,N_24914);
or UO_1338 (O_1338,N_24626,N_24938);
nor UO_1339 (O_1339,N_24909,N_24832);
xor UO_1340 (O_1340,N_24552,N_24563);
nor UO_1341 (O_1341,N_24730,N_24661);
nor UO_1342 (O_1342,N_24488,N_24432);
nor UO_1343 (O_1343,N_24704,N_24526);
and UO_1344 (O_1344,N_24774,N_24573);
and UO_1345 (O_1345,N_24400,N_24575);
nand UO_1346 (O_1346,N_24556,N_24413);
nand UO_1347 (O_1347,N_24995,N_24568);
xor UO_1348 (O_1348,N_24573,N_24756);
xnor UO_1349 (O_1349,N_24641,N_24676);
and UO_1350 (O_1350,N_24724,N_24782);
xor UO_1351 (O_1351,N_24642,N_24487);
nand UO_1352 (O_1352,N_24418,N_24774);
nor UO_1353 (O_1353,N_24570,N_24864);
and UO_1354 (O_1354,N_24584,N_24862);
xor UO_1355 (O_1355,N_24996,N_24692);
nand UO_1356 (O_1356,N_24565,N_24484);
xnor UO_1357 (O_1357,N_24618,N_24934);
or UO_1358 (O_1358,N_24926,N_24394);
nor UO_1359 (O_1359,N_24430,N_24523);
and UO_1360 (O_1360,N_24610,N_24427);
or UO_1361 (O_1361,N_24988,N_24899);
nand UO_1362 (O_1362,N_24680,N_24469);
nor UO_1363 (O_1363,N_24973,N_24388);
xnor UO_1364 (O_1364,N_24654,N_24762);
xnor UO_1365 (O_1365,N_24618,N_24859);
and UO_1366 (O_1366,N_24394,N_24930);
and UO_1367 (O_1367,N_24662,N_24467);
or UO_1368 (O_1368,N_24798,N_24969);
nor UO_1369 (O_1369,N_24773,N_24750);
and UO_1370 (O_1370,N_24778,N_24649);
nor UO_1371 (O_1371,N_24527,N_24641);
xor UO_1372 (O_1372,N_24433,N_24519);
xnor UO_1373 (O_1373,N_24618,N_24865);
and UO_1374 (O_1374,N_24867,N_24666);
and UO_1375 (O_1375,N_24421,N_24991);
nor UO_1376 (O_1376,N_24725,N_24518);
xnor UO_1377 (O_1377,N_24783,N_24556);
and UO_1378 (O_1378,N_24541,N_24805);
or UO_1379 (O_1379,N_24816,N_24979);
nand UO_1380 (O_1380,N_24947,N_24996);
xnor UO_1381 (O_1381,N_24576,N_24944);
nand UO_1382 (O_1382,N_24465,N_24445);
or UO_1383 (O_1383,N_24766,N_24515);
xnor UO_1384 (O_1384,N_24387,N_24951);
nand UO_1385 (O_1385,N_24807,N_24802);
nor UO_1386 (O_1386,N_24403,N_24409);
and UO_1387 (O_1387,N_24911,N_24704);
nor UO_1388 (O_1388,N_24773,N_24414);
xnor UO_1389 (O_1389,N_24956,N_24870);
nor UO_1390 (O_1390,N_24993,N_24939);
xnor UO_1391 (O_1391,N_24852,N_24475);
or UO_1392 (O_1392,N_24851,N_24566);
and UO_1393 (O_1393,N_24660,N_24680);
and UO_1394 (O_1394,N_24775,N_24996);
nor UO_1395 (O_1395,N_24527,N_24567);
xnor UO_1396 (O_1396,N_24761,N_24579);
and UO_1397 (O_1397,N_24880,N_24714);
and UO_1398 (O_1398,N_24797,N_24568);
nand UO_1399 (O_1399,N_24495,N_24831);
nor UO_1400 (O_1400,N_24605,N_24936);
xor UO_1401 (O_1401,N_24440,N_24988);
and UO_1402 (O_1402,N_24484,N_24793);
and UO_1403 (O_1403,N_24516,N_24859);
or UO_1404 (O_1404,N_24670,N_24815);
and UO_1405 (O_1405,N_24810,N_24507);
and UO_1406 (O_1406,N_24941,N_24767);
nand UO_1407 (O_1407,N_24934,N_24971);
and UO_1408 (O_1408,N_24717,N_24920);
nand UO_1409 (O_1409,N_24873,N_24446);
nor UO_1410 (O_1410,N_24460,N_24418);
or UO_1411 (O_1411,N_24469,N_24784);
and UO_1412 (O_1412,N_24570,N_24967);
nor UO_1413 (O_1413,N_24413,N_24659);
and UO_1414 (O_1414,N_24568,N_24539);
and UO_1415 (O_1415,N_24763,N_24802);
and UO_1416 (O_1416,N_24582,N_24735);
and UO_1417 (O_1417,N_24523,N_24414);
nand UO_1418 (O_1418,N_24744,N_24561);
xor UO_1419 (O_1419,N_24756,N_24857);
nor UO_1420 (O_1420,N_24766,N_24422);
xnor UO_1421 (O_1421,N_24414,N_24777);
xnor UO_1422 (O_1422,N_24938,N_24477);
nand UO_1423 (O_1423,N_24385,N_24660);
or UO_1424 (O_1424,N_24809,N_24577);
or UO_1425 (O_1425,N_24833,N_24699);
xnor UO_1426 (O_1426,N_24873,N_24800);
xor UO_1427 (O_1427,N_24487,N_24574);
and UO_1428 (O_1428,N_24441,N_24822);
nor UO_1429 (O_1429,N_24464,N_24380);
nand UO_1430 (O_1430,N_24416,N_24825);
and UO_1431 (O_1431,N_24763,N_24898);
nand UO_1432 (O_1432,N_24665,N_24754);
and UO_1433 (O_1433,N_24938,N_24786);
xor UO_1434 (O_1434,N_24496,N_24973);
nand UO_1435 (O_1435,N_24424,N_24834);
nor UO_1436 (O_1436,N_24810,N_24627);
or UO_1437 (O_1437,N_24547,N_24969);
and UO_1438 (O_1438,N_24748,N_24813);
nor UO_1439 (O_1439,N_24717,N_24459);
nand UO_1440 (O_1440,N_24485,N_24384);
nand UO_1441 (O_1441,N_24702,N_24990);
and UO_1442 (O_1442,N_24486,N_24465);
nor UO_1443 (O_1443,N_24871,N_24942);
or UO_1444 (O_1444,N_24550,N_24452);
and UO_1445 (O_1445,N_24813,N_24975);
and UO_1446 (O_1446,N_24663,N_24418);
and UO_1447 (O_1447,N_24432,N_24692);
xnor UO_1448 (O_1448,N_24832,N_24627);
nand UO_1449 (O_1449,N_24628,N_24471);
and UO_1450 (O_1450,N_24685,N_24486);
xor UO_1451 (O_1451,N_24497,N_24953);
or UO_1452 (O_1452,N_24902,N_24767);
and UO_1453 (O_1453,N_24749,N_24744);
nand UO_1454 (O_1454,N_24967,N_24580);
nor UO_1455 (O_1455,N_24568,N_24466);
xor UO_1456 (O_1456,N_24563,N_24380);
nand UO_1457 (O_1457,N_24853,N_24869);
xnor UO_1458 (O_1458,N_24485,N_24590);
nand UO_1459 (O_1459,N_24876,N_24786);
xnor UO_1460 (O_1460,N_24470,N_24593);
or UO_1461 (O_1461,N_24897,N_24809);
nand UO_1462 (O_1462,N_24541,N_24513);
nor UO_1463 (O_1463,N_24547,N_24828);
nor UO_1464 (O_1464,N_24543,N_24646);
nand UO_1465 (O_1465,N_24949,N_24928);
nor UO_1466 (O_1466,N_24701,N_24874);
and UO_1467 (O_1467,N_24459,N_24680);
nand UO_1468 (O_1468,N_24767,N_24762);
or UO_1469 (O_1469,N_24966,N_24620);
or UO_1470 (O_1470,N_24623,N_24907);
xor UO_1471 (O_1471,N_24991,N_24787);
nand UO_1472 (O_1472,N_24501,N_24748);
nand UO_1473 (O_1473,N_24878,N_24794);
nor UO_1474 (O_1474,N_24648,N_24877);
or UO_1475 (O_1475,N_24720,N_24736);
and UO_1476 (O_1476,N_24614,N_24455);
nor UO_1477 (O_1477,N_24749,N_24797);
nand UO_1478 (O_1478,N_24472,N_24907);
or UO_1479 (O_1479,N_24534,N_24435);
nand UO_1480 (O_1480,N_24583,N_24538);
and UO_1481 (O_1481,N_24777,N_24609);
or UO_1482 (O_1482,N_24537,N_24767);
or UO_1483 (O_1483,N_24487,N_24421);
or UO_1484 (O_1484,N_24852,N_24628);
or UO_1485 (O_1485,N_24585,N_24553);
xnor UO_1486 (O_1486,N_24469,N_24789);
or UO_1487 (O_1487,N_24762,N_24536);
xor UO_1488 (O_1488,N_24543,N_24792);
or UO_1489 (O_1489,N_24903,N_24572);
xnor UO_1490 (O_1490,N_24740,N_24869);
nand UO_1491 (O_1491,N_24974,N_24450);
or UO_1492 (O_1492,N_24413,N_24791);
xnor UO_1493 (O_1493,N_24823,N_24407);
xnor UO_1494 (O_1494,N_24620,N_24748);
nand UO_1495 (O_1495,N_24928,N_24501);
and UO_1496 (O_1496,N_24854,N_24519);
nor UO_1497 (O_1497,N_24656,N_24526);
or UO_1498 (O_1498,N_24388,N_24796);
and UO_1499 (O_1499,N_24898,N_24952);
and UO_1500 (O_1500,N_24629,N_24813);
xor UO_1501 (O_1501,N_24808,N_24839);
nand UO_1502 (O_1502,N_24680,N_24964);
xor UO_1503 (O_1503,N_24501,N_24674);
and UO_1504 (O_1504,N_24989,N_24830);
nand UO_1505 (O_1505,N_24947,N_24802);
nor UO_1506 (O_1506,N_24894,N_24673);
nor UO_1507 (O_1507,N_24467,N_24777);
nand UO_1508 (O_1508,N_24662,N_24731);
and UO_1509 (O_1509,N_24608,N_24475);
nand UO_1510 (O_1510,N_24391,N_24757);
or UO_1511 (O_1511,N_24544,N_24464);
or UO_1512 (O_1512,N_24746,N_24539);
and UO_1513 (O_1513,N_24932,N_24892);
or UO_1514 (O_1514,N_24588,N_24917);
nand UO_1515 (O_1515,N_24722,N_24470);
and UO_1516 (O_1516,N_24776,N_24580);
nor UO_1517 (O_1517,N_24578,N_24859);
nor UO_1518 (O_1518,N_24578,N_24709);
nand UO_1519 (O_1519,N_24695,N_24413);
xor UO_1520 (O_1520,N_24651,N_24949);
xnor UO_1521 (O_1521,N_24974,N_24855);
or UO_1522 (O_1522,N_24819,N_24944);
nor UO_1523 (O_1523,N_24840,N_24457);
or UO_1524 (O_1524,N_24433,N_24504);
nor UO_1525 (O_1525,N_24569,N_24416);
or UO_1526 (O_1526,N_24743,N_24890);
or UO_1527 (O_1527,N_24446,N_24772);
or UO_1528 (O_1528,N_24868,N_24459);
nor UO_1529 (O_1529,N_24913,N_24484);
and UO_1530 (O_1530,N_24498,N_24676);
nand UO_1531 (O_1531,N_24702,N_24598);
and UO_1532 (O_1532,N_24923,N_24806);
or UO_1533 (O_1533,N_24703,N_24384);
nor UO_1534 (O_1534,N_24962,N_24918);
and UO_1535 (O_1535,N_24792,N_24932);
nand UO_1536 (O_1536,N_24626,N_24932);
and UO_1537 (O_1537,N_24708,N_24840);
xnor UO_1538 (O_1538,N_24728,N_24517);
or UO_1539 (O_1539,N_24984,N_24986);
and UO_1540 (O_1540,N_24663,N_24666);
or UO_1541 (O_1541,N_24730,N_24945);
and UO_1542 (O_1542,N_24965,N_24926);
nand UO_1543 (O_1543,N_24729,N_24834);
nand UO_1544 (O_1544,N_24649,N_24422);
nand UO_1545 (O_1545,N_24875,N_24823);
nor UO_1546 (O_1546,N_24770,N_24671);
xor UO_1547 (O_1547,N_24388,N_24825);
xor UO_1548 (O_1548,N_24891,N_24781);
nand UO_1549 (O_1549,N_24755,N_24812);
or UO_1550 (O_1550,N_24965,N_24586);
nor UO_1551 (O_1551,N_24847,N_24723);
and UO_1552 (O_1552,N_24480,N_24662);
nor UO_1553 (O_1553,N_24688,N_24793);
nand UO_1554 (O_1554,N_24417,N_24917);
xor UO_1555 (O_1555,N_24593,N_24760);
or UO_1556 (O_1556,N_24507,N_24760);
nor UO_1557 (O_1557,N_24419,N_24631);
and UO_1558 (O_1558,N_24415,N_24991);
and UO_1559 (O_1559,N_24969,N_24770);
nand UO_1560 (O_1560,N_24927,N_24453);
xor UO_1561 (O_1561,N_24819,N_24867);
and UO_1562 (O_1562,N_24866,N_24968);
or UO_1563 (O_1563,N_24378,N_24549);
and UO_1564 (O_1564,N_24611,N_24480);
or UO_1565 (O_1565,N_24685,N_24553);
xnor UO_1566 (O_1566,N_24852,N_24414);
and UO_1567 (O_1567,N_24574,N_24867);
nand UO_1568 (O_1568,N_24844,N_24442);
or UO_1569 (O_1569,N_24747,N_24418);
or UO_1570 (O_1570,N_24916,N_24822);
nand UO_1571 (O_1571,N_24695,N_24766);
and UO_1572 (O_1572,N_24950,N_24472);
nand UO_1573 (O_1573,N_24952,N_24771);
or UO_1574 (O_1574,N_24632,N_24945);
nand UO_1575 (O_1575,N_24648,N_24730);
nor UO_1576 (O_1576,N_24792,N_24677);
xnor UO_1577 (O_1577,N_24584,N_24502);
xor UO_1578 (O_1578,N_24975,N_24530);
or UO_1579 (O_1579,N_24375,N_24928);
or UO_1580 (O_1580,N_24782,N_24625);
or UO_1581 (O_1581,N_24923,N_24427);
nor UO_1582 (O_1582,N_24545,N_24785);
nor UO_1583 (O_1583,N_24500,N_24435);
nor UO_1584 (O_1584,N_24538,N_24771);
nand UO_1585 (O_1585,N_24521,N_24520);
nor UO_1586 (O_1586,N_24886,N_24771);
xor UO_1587 (O_1587,N_24469,N_24851);
xnor UO_1588 (O_1588,N_24983,N_24776);
nand UO_1589 (O_1589,N_24757,N_24797);
nor UO_1590 (O_1590,N_24465,N_24382);
and UO_1591 (O_1591,N_24759,N_24553);
and UO_1592 (O_1592,N_24784,N_24899);
xor UO_1593 (O_1593,N_24792,N_24393);
nor UO_1594 (O_1594,N_24397,N_24899);
or UO_1595 (O_1595,N_24412,N_24692);
or UO_1596 (O_1596,N_24565,N_24435);
nand UO_1597 (O_1597,N_24863,N_24575);
or UO_1598 (O_1598,N_24497,N_24754);
nor UO_1599 (O_1599,N_24994,N_24548);
or UO_1600 (O_1600,N_24433,N_24730);
nand UO_1601 (O_1601,N_24662,N_24880);
or UO_1602 (O_1602,N_24643,N_24674);
xor UO_1603 (O_1603,N_24924,N_24547);
nor UO_1604 (O_1604,N_24793,N_24985);
or UO_1605 (O_1605,N_24431,N_24393);
nand UO_1606 (O_1606,N_24406,N_24683);
xor UO_1607 (O_1607,N_24998,N_24903);
and UO_1608 (O_1608,N_24472,N_24639);
nor UO_1609 (O_1609,N_24528,N_24564);
or UO_1610 (O_1610,N_24671,N_24618);
nand UO_1611 (O_1611,N_24867,N_24588);
or UO_1612 (O_1612,N_24475,N_24618);
nor UO_1613 (O_1613,N_24690,N_24458);
or UO_1614 (O_1614,N_24422,N_24569);
xor UO_1615 (O_1615,N_24556,N_24481);
nor UO_1616 (O_1616,N_24897,N_24535);
nor UO_1617 (O_1617,N_24998,N_24573);
nand UO_1618 (O_1618,N_24967,N_24759);
and UO_1619 (O_1619,N_24475,N_24772);
and UO_1620 (O_1620,N_24556,N_24421);
nand UO_1621 (O_1621,N_24905,N_24863);
or UO_1622 (O_1622,N_24438,N_24408);
nor UO_1623 (O_1623,N_24497,N_24399);
and UO_1624 (O_1624,N_24982,N_24686);
and UO_1625 (O_1625,N_24730,N_24520);
and UO_1626 (O_1626,N_24743,N_24783);
xor UO_1627 (O_1627,N_24834,N_24544);
nand UO_1628 (O_1628,N_24921,N_24660);
or UO_1629 (O_1629,N_24562,N_24550);
nand UO_1630 (O_1630,N_24960,N_24952);
and UO_1631 (O_1631,N_24728,N_24777);
nor UO_1632 (O_1632,N_24488,N_24780);
and UO_1633 (O_1633,N_24850,N_24550);
or UO_1634 (O_1634,N_24637,N_24915);
or UO_1635 (O_1635,N_24599,N_24787);
nand UO_1636 (O_1636,N_24610,N_24533);
nand UO_1637 (O_1637,N_24375,N_24705);
nor UO_1638 (O_1638,N_24541,N_24891);
nor UO_1639 (O_1639,N_24584,N_24486);
nand UO_1640 (O_1640,N_24579,N_24395);
and UO_1641 (O_1641,N_24720,N_24627);
xnor UO_1642 (O_1642,N_24975,N_24957);
or UO_1643 (O_1643,N_24438,N_24999);
or UO_1644 (O_1644,N_24866,N_24483);
and UO_1645 (O_1645,N_24774,N_24528);
nand UO_1646 (O_1646,N_24568,N_24627);
and UO_1647 (O_1647,N_24649,N_24835);
nor UO_1648 (O_1648,N_24424,N_24874);
nand UO_1649 (O_1649,N_24780,N_24522);
nor UO_1650 (O_1650,N_24450,N_24618);
or UO_1651 (O_1651,N_24902,N_24385);
nand UO_1652 (O_1652,N_24637,N_24879);
and UO_1653 (O_1653,N_24699,N_24746);
nor UO_1654 (O_1654,N_24929,N_24408);
nand UO_1655 (O_1655,N_24922,N_24982);
nand UO_1656 (O_1656,N_24810,N_24640);
nor UO_1657 (O_1657,N_24565,N_24397);
or UO_1658 (O_1658,N_24668,N_24745);
xnor UO_1659 (O_1659,N_24970,N_24713);
and UO_1660 (O_1660,N_24673,N_24420);
xnor UO_1661 (O_1661,N_24850,N_24870);
nor UO_1662 (O_1662,N_24445,N_24472);
and UO_1663 (O_1663,N_24816,N_24457);
xnor UO_1664 (O_1664,N_24992,N_24472);
and UO_1665 (O_1665,N_24712,N_24773);
and UO_1666 (O_1666,N_24723,N_24933);
or UO_1667 (O_1667,N_24831,N_24790);
and UO_1668 (O_1668,N_24994,N_24881);
nor UO_1669 (O_1669,N_24453,N_24945);
xor UO_1670 (O_1670,N_24719,N_24648);
or UO_1671 (O_1671,N_24877,N_24910);
nand UO_1672 (O_1672,N_24620,N_24658);
nor UO_1673 (O_1673,N_24762,N_24653);
nor UO_1674 (O_1674,N_24684,N_24585);
or UO_1675 (O_1675,N_24648,N_24594);
nand UO_1676 (O_1676,N_24586,N_24958);
and UO_1677 (O_1677,N_24842,N_24494);
or UO_1678 (O_1678,N_24872,N_24741);
nor UO_1679 (O_1679,N_24619,N_24749);
xor UO_1680 (O_1680,N_24673,N_24418);
xor UO_1681 (O_1681,N_24868,N_24434);
and UO_1682 (O_1682,N_24854,N_24527);
nor UO_1683 (O_1683,N_24725,N_24388);
nand UO_1684 (O_1684,N_24682,N_24768);
nand UO_1685 (O_1685,N_24636,N_24556);
nor UO_1686 (O_1686,N_24921,N_24954);
or UO_1687 (O_1687,N_24513,N_24778);
or UO_1688 (O_1688,N_24952,N_24706);
or UO_1689 (O_1689,N_24868,N_24680);
and UO_1690 (O_1690,N_24749,N_24987);
and UO_1691 (O_1691,N_24489,N_24546);
and UO_1692 (O_1692,N_24612,N_24878);
or UO_1693 (O_1693,N_24463,N_24508);
or UO_1694 (O_1694,N_24674,N_24688);
or UO_1695 (O_1695,N_24591,N_24717);
nor UO_1696 (O_1696,N_24599,N_24741);
nor UO_1697 (O_1697,N_24688,N_24858);
nor UO_1698 (O_1698,N_24423,N_24710);
xnor UO_1699 (O_1699,N_24622,N_24391);
xnor UO_1700 (O_1700,N_24618,N_24777);
or UO_1701 (O_1701,N_24666,N_24653);
or UO_1702 (O_1702,N_24450,N_24957);
and UO_1703 (O_1703,N_24383,N_24624);
or UO_1704 (O_1704,N_24800,N_24562);
nand UO_1705 (O_1705,N_24791,N_24670);
or UO_1706 (O_1706,N_24786,N_24905);
and UO_1707 (O_1707,N_24694,N_24393);
nand UO_1708 (O_1708,N_24806,N_24509);
nand UO_1709 (O_1709,N_24387,N_24525);
or UO_1710 (O_1710,N_24433,N_24908);
nand UO_1711 (O_1711,N_24445,N_24609);
and UO_1712 (O_1712,N_24466,N_24681);
and UO_1713 (O_1713,N_24927,N_24392);
and UO_1714 (O_1714,N_24926,N_24977);
xnor UO_1715 (O_1715,N_24800,N_24639);
or UO_1716 (O_1716,N_24489,N_24941);
nand UO_1717 (O_1717,N_24608,N_24471);
xor UO_1718 (O_1718,N_24794,N_24625);
xor UO_1719 (O_1719,N_24690,N_24532);
nor UO_1720 (O_1720,N_24484,N_24633);
or UO_1721 (O_1721,N_24673,N_24448);
or UO_1722 (O_1722,N_24696,N_24579);
nand UO_1723 (O_1723,N_24416,N_24598);
nor UO_1724 (O_1724,N_24661,N_24727);
nand UO_1725 (O_1725,N_24844,N_24448);
nand UO_1726 (O_1726,N_24892,N_24454);
nand UO_1727 (O_1727,N_24637,N_24903);
and UO_1728 (O_1728,N_24540,N_24598);
nor UO_1729 (O_1729,N_24815,N_24555);
nand UO_1730 (O_1730,N_24567,N_24834);
nand UO_1731 (O_1731,N_24579,N_24529);
and UO_1732 (O_1732,N_24832,N_24508);
nand UO_1733 (O_1733,N_24715,N_24505);
nand UO_1734 (O_1734,N_24901,N_24971);
xor UO_1735 (O_1735,N_24585,N_24754);
nor UO_1736 (O_1736,N_24891,N_24534);
xor UO_1737 (O_1737,N_24614,N_24563);
or UO_1738 (O_1738,N_24411,N_24445);
or UO_1739 (O_1739,N_24897,N_24963);
nand UO_1740 (O_1740,N_24420,N_24991);
nor UO_1741 (O_1741,N_24774,N_24906);
xor UO_1742 (O_1742,N_24790,N_24395);
or UO_1743 (O_1743,N_24947,N_24592);
nor UO_1744 (O_1744,N_24723,N_24631);
nand UO_1745 (O_1745,N_24883,N_24948);
and UO_1746 (O_1746,N_24968,N_24585);
or UO_1747 (O_1747,N_24473,N_24662);
nand UO_1748 (O_1748,N_24742,N_24779);
nand UO_1749 (O_1749,N_24667,N_24465);
nor UO_1750 (O_1750,N_24917,N_24454);
or UO_1751 (O_1751,N_24846,N_24796);
nand UO_1752 (O_1752,N_24432,N_24978);
and UO_1753 (O_1753,N_24465,N_24478);
nor UO_1754 (O_1754,N_24708,N_24496);
nor UO_1755 (O_1755,N_24848,N_24694);
and UO_1756 (O_1756,N_24898,N_24824);
and UO_1757 (O_1757,N_24518,N_24734);
xor UO_1758 (O_1758,N_24857,N_24680);
nor UO_1759 (O_1759,N_24863,N_24959);
xor UO_1760 (O_1760,N_24382,N_24507);
xnor UO_1761 (O_1761,N_24625,N_24884);
xor UO_1762 (O_1762,N_24738,N_24428);
xnor UO_1763 (O_1763,N_24485,N_24392);
and UO_1764 (O_1764,N_24537,N_24967);
xor UO_1765 (O_1765,N_24862,N_24711);
and UO_1766 (O_1766,N_24801,N_24524);
xor UO_1767 (O_1767,N_24803,N_24563);
nor UO_1768 (O_1768,N_24833,N_24660);
xnor UO_1769 (O_1769,N_24515,N_24711);
nand UO_1770 (O_1770,N_24960,N_24959);
and UO_1771 (O_1771,N_24469,N_24657);
and UO_1772 (O_1772,N_24537,N_24792);
nor UO_1773 (O_1773,N_24513,N_24425);
nand UO_1774 (O_1774,N_24424,N_24870);
xor UO_1775 (O_1775,N_24409,N_24749);
xor UO_1776 (O_1776,N_24494,N_24794);
nor UO_1777 (O_1777,N_24638,N_24411);
xnor UO_1778 (O_1778,N_24420,N_24649);
xor UO_1779 (O_1779,N_24788,N_24760);
or UO_1780 (O_1780,N_24900,N_24668);
or UO_1781 (O_1781,N_24964,N_24595);
and UO_1782 (O_1782,N_24720,N_24845);
nand UO_1783 (O_1783,N_24865,N_24624);
nand UO_1784 (O_1784,N_24615,N_24947);
xnor UO_1785 (O_1785,N_24825,N_24531);
nor UO_1786 (O_1786,N_24378,N_24586);
or UO_1787 (O_1787,N_24630,N_24669);
xor UO_1788 (O_1788,N_24801,N_24777);
xnor UO_1789 (O_1789,N_24904,N_24775);
nor UO_1790 (O_1790,N_24782,N_24501);
nand UO_1791 (O_1791,N_24461,N_24992);
xor UO_1792 (O_1792,N_24657,N_24981);
and UO_1793 (O_1793,N_24922,N_24844);
or UO_1794 (O_1794,N_24978,N_24427);
or UO_1795 (O_1795,N_24408,N_24566);
xnor UO_1796 (O_1796,N_24531,N_24907);
nand UO_1797 (O_1797,N_24435,N_24711);
xnor UO_1798 (O_1798,N_24723,N_24801);
xor UO_1799 (O_1799,N_24520,N_24578);
or UO_1800 (O_1800,N_24581,N_24767);
and UO_1801 (O_1801,N_24463,N_24885);
xor UO_1802 (O_1802,N_24914,N_24470);
and UO_1803 (O_1803,N_24493,N_24726);
xnor UO_1804 (O_1804,N_24500,N_24402);
nor UO_1805 (O_1805,N_24952,N_24520);
nand UO_1806 (O_1806,N_24900,N_24956);
nand UO_1807 (O_1807,N_24739,N_24679);
nor UO_1808 (O_1808,N_24860,N_24475);
and UO_1809 (O_1809,N_24663,N_24749);
nor UO_1810 (O_1810,N_24508,N_24629);
or UO_1811 (O_1811,N_24885,N_24893);
and UO_1812 (O_1812,N_24544,N_24744);
xnor UO_1813 (O_1813,N_24811,N_24728);
xnor UO_1814 (O_1814,N_24960,N_24779);
xnor UO_1815 (O_1815,N_24542,N_24378);
nor UO_1816 (O_1816,N_24529,N_24626);
nor UO_1817 (O_1817,N_24561,N_24995);
nor UO_1818 (O_1818,N_24495,N_24774);
and UO_1819 (O_1819,N_24714,N_24662);
nand UO_1820 (O_1820,N_24679,N_24571);
nor UO_1821 (O_1821,N_24447,N_24716);
nor UO_1822 (O_1822,N_24841,N_24980);
or UO_1823 (O_1823,N_24916,N_24387);
or UO_1824 (O_1824,N_24392,N_24785);
xnor UO_1825 (O_1825,N_24830,N_24529);
nand UO_1826 (O_1826,N_24428,N_24583);
or UO_1827 (O_1827,N_24528,N_24601);
and UO_1828 (O_1828,N_24718,N_24379);
or UO_1829 (O_1829,N_24748,N_24497);
or UO_1830 (O_1830,N_24544,N_24721);
nand UO_1831 (O_1831,N_24402,N_24617);
and UO_1832 (O_1832,N_24398,N_24385);
nor UO_1833 (O_1833,N_24551,N_24861);
and UO_1834 (O_1834,N_24904,N_24777);
nand UO_1835 (O_1835,N_24790,N_24619);
nor UO_1836 (O_1836,N_24752,N_24402);
nand UO_1837 (O_1837,N_24385,N_24774);
nor UO_1838 (O_1838,N_24744,N_24689);
or UO_1839 (O_1839,N_24890,N_24960);
nor UO_1840 (O_1840,N_24640,N_24875);
nand UO_1841 (O_1841,N_24514,N_24742);
nand UO_1842 (O_1842,N_24418,N_24782);
and UO_1843 (O_1843,N_24436,N_24516);
xnor UO_1844 (O_1844,N_24718,N_24513);
xnor UO_1845 (O_1845,N_24400,N_24672);
nand UO_1846 (O_1846,N_24385,N_24921);
xor UO_1847 (O_1847,N_24525,N_24475);
or UO_1848 (O_1848,N_24614,N_24593);
nand UO_1849 (O_1849,N_24640,N_24681);
xor UO_1850 (O_1850,N_24757,N_24382);
xnor UO_1851 (O_1851,N_24802,N_24404);
nand UO_1852 (O_1852,N_24988,N_24979);
nand UO_1853 (O_1853,N_24827,N_24458);
xnor UO_1854 (O_1854,N_24897,N_24875);
or UO_1855 (O_1855,N_24631,N_24886);
nand UO_1856 (O_1856,N_24702,N_24996);
and UO_1857 (O_1857,N_24632,N_24390);
nand UO_1858 (O_1858,N_24430,N_24713);
xnor UO_1859 (O_1859,N_24812,N_24402);
xnor UO_1860 (O_1860,N_24647,N_24403);
nand UO_1861 (O_1861,N_24826,N_24530);
or UO_1862 (O_1862,N_24501,N_24974);
and UO_1863 (O_1863,N_24662,N_24736);
nor UO_1864 (O_1864,N_24981,N_24879);
nand UO_1865 (O_1865,N_24470,N_24882);
or UO_1866 (O_1866,N_24883,N_24755);
or UO_1867 (O_1867,N_24832,N_24572);
and UO_1868 (O_1868,N_24874,N_24564);
nor UO_1869 (O_1869,N_24962,N_24900);
xor UO_1870 (O_1870,N_24755,N_24743);
xnor UO_1871 (O_1871,N_24707,N_24709);
nand UO_1872 (O_1872,N_24508,N_24461);
nor UO_1873 (O_1873,N_24440,N_24763);
and UO_1874 (O_1874,N_24691,N_24376);
and UO_1875 (O_1875,N_24427,N_24501);
nand UO_1876 (O_1876,N_24894,N_24808);
or UO_1877 (O_1877,N_24740,N_24951);
xor UO_1878 (O_1878,N_24919,N_24907);
or UO_1879 (O_1879,N_24430,N_24486);
or UO_1880 (O_1880,N_24480,N_24424);
and UO_1881 (O_1881,N_24671,N_24688);
nand UO_1882 (O_1882,N_24792,N_24414);
xor UO_1883 (O_1883,N_24460,N_24591);
nand UO_1884 (O_1884,N_24949,N_24527);
xnor UO_1885 (O_1885,N_24685,N_24573);
xnor UO_1886 (O_1886,N_24994,N_24962);
nand UO_1887 (O_1887,N_24818,N_24492);
or UO_1888 (O_1888,N_24869,N_24921);
and UO_1889 (O_1889,N_24861,N_24916);
nor UO_1890 (O_1890,N_24393,N_24630);
nand UO_1891 (O_1891,N_24472,N_24998);
or UO_1892 (O_1892,N_24827,N_24552);
or UO_1893 (O_1893,N_24566,N_24590);
nand UO_1894 (O_1894,N_24544,N_24858);
nor UO_1895 (O_1895,N_24420,N_24482);
nor UO_1896 (O_1896,N_24721,N_24706);
and UO_1897 (O_1897,N_24824,N_24660);
xor UO_1898 (O_1898,N_24808,N_24647);
nor UO_1899 (O_1899,N_24406,N_24397);
nor UO_1900 (O_1900,N_24457,N_24522);
nand UO_1901 (O_1901,N_24400,N_24629);
nand UO_1902 (O_1902,N_24406,N_24635);
xor UO_1903 (O_1903,N_24383,N_24423);
or UO_1904 (O_1904,N_24394,N_24429);
xnor UO_1905 (O_1905,N_24630,N_24994);
or UO_1906 (O_1906,N_24523,N_24902);
xnor UO_1907 (O_1907,N_24679,N_24845);
nand UO_1908 (O_1908,N_24641,N_24523);
nor UO_1909 (O_1909,N_24381,N_24460);
xnor UO_1910 (O_1910,N_24902,N_24502);
xnor UO_1911 (O_1911,N_24528,N_24674);
or UO_1912 (O_1912,N_24387,N_24412);
and UO_1913 (O_1913,N_24592,N_24994);
or UO_1914 (O_1914,N_24873,N_24571);
or UO_1915 (O_1915,N_24571,N_24907);
xor UO_1916 (O_1916,N_24883,N_24774);
xnor UO_1917 (O_1917,N_24811,N_24837);
nor UO_1918 (O_1918,N_24922,N_24809);
nor UO_1919 (O_1919,N_24930,N_24636);
nand UO_1920 (O_1920,N_24614,N_24561);
xnor UO_1921 (O_1921,N_24935,N_24456);
xnor UO_1922 (O_1922,N_24812,N_24911);
and UO_1923 (O_1923,N_24902,N_24720);
nor UO_1924 (O_1924,N_24393,N_24623);
xnor UO_1925 (O_1925,N_24739,N_24433);
or UO_1926 (O_1926,N_24519,N_24997);
nand UO_1927 (O_1927,N_24844,N_24504);
and UO_1928 (O_1928,N_24507,N_24999);
xor UO_1929 (O_1929,N_24914,N_24907);
or UO_1930 (O_1930,N_24930,N_24485);
or UO_1931 (O_1931,N_24638,N_24747);
or UO_1932 (O_1932,N_24641,N_24882);
xnor UO_1933 (O_1933,N_24568,N_24430);
and UO_1934 (O_1934,N_24678,N_24756);
or UO_1935 (O_1935,N_24633,N_24659);
nor UO_1936 (O_1936,N_24492,N_24567);
or UO_1937 (O_1937,N_24528,N_24603);
nand UO_1938 (O_1938,N_24603,N_24800);
nand UO_1939 (O_1939,N_24411,N_24787);
xor UO_1940 (O_1940,N_24456,N_24598);
and UO_1941 (O_1941,N_24725,N_24478);
nand UO_1942 (O_1942,N_24743,N_24770);
nor UO_1943 (O_1943,N_24714,N_24862);
xor UO_1944 (O_1944,N_24704,N_24422);
or UO_1945 (O_1945,N_24442,N_24464);
and UO_1946 (O_1946,N_24975,N_24933);
or UO_1947 (O_1947,N_24609,N_24412);
nand UO_1948 (O_1948,N_24436,N_24954);
xor UO_1949 (O_1949,N_24505,N_24651);
nand UO_1950 (O_1950,N_24436,N_24502);
nand UO_1951 (O_1951,N_24576,N_24922);
nor UO_1952 (O_1952,N_24782,N_24534);
nand UO_1953 (O_1953,N_24481,N_24559);
and UO_1954 (O_1954,N_24764,N_24827);
nand UO_1955 (O_1955,N_24628,N_24594);
xnor UO_1956 (O_1956,N_24648,N_24945);
xnor UO_1957 (O_1957,N_24433,N_24486);
nor UO_1958 (O_1958,N_24799,N_24746);
xnor UO_1959 (O_1959,N_24641,N_24615);
nand UO_1960 (O_1960,N_24812,N_24851);
or UO_1961 (O_1961,N_24708,N_24963);
and UO_1962 (O_1962,N_24968,N_24853);
nor UO_1963 (O_1963,N_24964,N_24960);
xnor UO_1964 (O_1964,N_24956,N_24635);
nand UO_1965 (O_1965,N_24728,N_24493);
nand UO_1966 (O_1966,N_24470,N_24625);
nor UO_1967 (O_1967,N_24541,N_24980);
or UO_1968 (O_1968,N_24518,N_24645);
or UO_1969 (O_1969,N_24636,N_24520);
nor UO_1970 (O_1970,N_24729,N_24993);
xnor UO_1971 (O_1971,N_24712,N_24973);
xnor UO_1972 (O_1972,N_24410,N_24550);
and UO_1973 (O_1973,N_24628,N_24444);
nand UO_1974 (O_1974,N_24965,N_24777);
or UO_1975 (O_1975,N_24918,N_24628);
nand UO_1976 (O_1976,N_24701,N_24870);
xor UO_1977 (O_1977,N_24803,N_24821);
nor UO_1978 (O_1978,N_24504,N_24978);
or UO_1979 (O_1979,N_24943,N_24721);
nor UO_1980 (O_1980,N_24433,N_24631);
or UO_1981 (O_1981,N_24803,N_24402);
or UO_1982 (O_1982,N_24460,N_24714);
nor UO_1983 (O_1983,N_24912,N_24928);
and UO_1984 (O_1984,N_24933,N_24891);
or UO_1985 (O_1985,N_24438,N_24381);
xnor UO_1986 (O_1986,N_24401,N_24827);
xor UO_1987 (O_1987,N_24476,N_24844);
xnor UO_1988 (O_1988,N_24935,N_24433);
and UO_1989 (O_1989,N_24798,N_24544);
and UO_1990 (O_1990,N_24486,N_24440);
and UO_1991 (O_1991,N_24914,N_24784);
xor UO_1992 (O_1992,N_24869,N_24975);
nand UO_1993 (O_1993,N_24378,N_24529);
and UO_1994 (O_1994,N_24436,N_24473);
nand UO_1995 (O_1995,N_24469,N_24646);
xnor UO_1996 (O_1996,N_24741,N_24988);
nand UO_1997 (O_1997,N_24840,N_24869);
or UO_1998 (O_1998,N_24823,N_24899);
or UO_1999 (O_1999,N_24479,N_24868);
nand UO_2000 (O_2000,N_24835,N_24923);
nor UO_2001 (O_2001,N_24603,N_24968);
nor UO_2002 (O_2002,N_24903,N_24803);
nor UO_2003 (O_2003,N_24505,N_24485);
or UO_2004 (O_2004,N_24667,N_24597);
or UO_2005 (O_2005,N_24622,N_24848);
xnor UO_2006 (O_2006,N_24528,N_24556);
and UO_2007 (O_2007,N_24508,N_24599);
nand UO_2008 (O_2008,N_24786,N_24904);
nor UO_2009 (O_2009,N_24421,N_24507);
nor UO_2010 (O_2010,N_24936,N_24783);
and UO_2011 (O_2011,N_24516,N_24688);
xnor UO_2012 (O_2012,N_24801,N_24669);
and UO_2013 (O_2013,N_24663,N_24805);
or UO_2014 (O_2014,N_24902,N_24785);
and UO_2015 (O_2015,N_24418,N_24564);
xor UO_2016 (O_2016,N_24797,N_24522);
or UO_2017 (O_2017,N_24621,N_24521);
or UO_2018 (O_2018,N_24801,N_24545);
xnor UO_2019 (O_2019,N_24846,N_24931);
or UO_2020 (O_2020,N_24913,N_24932);
and UO_2021 (O_2021,N_24740,N_24781);
nand UO_2022 (O_2022,N_24813,N_24376);
and UO_2023 (O_2023,N_24732,N_24745);
and UO_2024 (O_2024,N_24880,N_24781);
or UO_2025 (O_2025,N_24954,N_24779);
or UO_2026 (O_2026,N_24617,N_24955);
nor UO_2027 (O_2027,N_24981,N_24540);
nand UO_2028 (O_2028,N_24521,N_24923);
nor UO_2029 (O_2029,N_24903,N_24740);
and UO_2030 (O_2030,N_24636,N_24526);
or UO_2031 (O_2031,N_24644,N_24786);
and UO_2032 (O_2032,N_24545,N_24776);
or UO_2033 (O_2033,N_24742,N_24919);
and UO_2034 (O_2034,N_24795,N_24925);
nor UO_2035 (O_2035,N_24771,N_24499);
xnor UO_2036 (O_2036,N_24419,N_24870);
xnor UO_2037 (O_2037,N_24393,N_24951);
nand UO_2038 (O_2038,N_24489,N_24601);
and UO_2039 (O_2039,N_24775,N_24454);
xnor UO_2040 (O_2040,N_24806,N_24660);
and UO_2041 (O_2041,N_24380,N_24987);
and UO_2042 (O_2042,N_24809,N_24965);
nor UO_2043 (O_2043,N_24642,N_24930);
nor UO_2044 (O_2044,N_24749,N_24407);
and UO_2045 (O_2045,N_24939,N_24780);
or UO_2046 (O_2046,N_24857,N_24859);
xor UO_2047 (O_2047,N_24542,N_24887);
nor UO_2048 (O_2048,N_24721,N_24428);
nor UO_2049 (O_2049,N_24628,N_24650);
nor UO_2050 (O_2050,N_24468,N_24816);
and UO_2051 (O_2051,N_24496,N_24882);
or UO_2052 (O_2052,N_24934,N_24557);
nand UO_2053 (O_2053,N_24792,N_24616);
nor UO_2054 (O_2054,N_24926,N_24573);
nand UO_2055 (O_2055,N_24430,N_24583);
or UO_2056 (O_2056,N_24923,N_24468);
nand UO_2057 (O_2057,N_24705,N_24409);
nor UO_2058 (O_2058,N_24469,N_24790);
or UO_2059 (O_2059,N_24684,N_24562);
and UO_2060 (O_2060,N_24467,N_24980);
xor UO_2061 (O_2061,N_24941,N_24716);
nand UO_2062 (O_2062,N_24394,N_24503);
xor UO_2063 (O_2063,N_24391,N_24581);
or UO_2064 (O_2064,N_24714,N_24804);
nand UO_2065 (O_2065,N_24628,N_24776);
xor UO_2066 (O_2066,N_24908,N_24779);
xor UO_2067 (O_2067,N_24639,N_24453);
xnor UO_2068 (O_2068,N_24894,N_24893);
xnor UO_2069 (O_2069,N_24694,N_24757);
nand UO_2070 (O_2070,N_24498,N_24731);
nor UO_2071 (O_2071,N_24809,N_24993);
nand UO_2072 (O_2072,N_24998,N_24977);
and UO_2073 (O_2073,N_24383,N_24840);
and UO_2074 (O_2074,N_24534,N_24569);
nor UO_2075 (O_2075,N_24908,N_24653);
and UO_2076 (O_2076,N_24643,N_24645);
or UO_2077 (O_2077,N_24476,N_24965);
and UO_2078 (O_2078,N_24806,N_24968);
and UO_2079 (O_2079,N_24436,N_24476);
and UO_2080 (O_2080,N_24889,N_24489);
xor UO_2081 (O_2081,N_24376,N_24419);
and UO_2082 (O_2082,N_24663,N_24645);
xor UO_2083 (O_2083,N_24715,N_24458);
or UO_2084 (O_2084,N_24393,N_24722);
or UO_2085 (O_2085,N_24857,N_24925);
or UO_2086 (O_2086,N_24783,N_24889);
nor UO_2087 (O_2087,N_24636,N_24726);
nand UO_2088 (O_2088,N_24695,N_24631);
nand UO_2089 (O_2089,N_24961,N_24536);
xor UO_2090 (O_2090,N_24602,N_24795);
or UO_2091 (O_2091,N_24375,N_24377);
nor UO_2092 (O_2092,N_24536,N_24765);
and UO_2093 (O_2093,N_24735,N_24514);
xnor UO_2094 (O_2094,N_24537,N_24459);
nor UO_2095 (O_2095,N_24887,N_24538);
nor UO_2096 (O_2096,N_24727,N_24772);
nor UO_2097 (O_2097,N_24645,N_24780);
and UO_2098 (O_2098,N_24875,N_24942);
nand UO_2099 (O_2099,N_24869,N_24948);
and UO_2100 (O_2100,N_24535,N_24388);
xor UO_2101 (O_2101,N_24721,N_24789);
nand UO_2102 (O_2102,N_24779,N_24561);
and UO_2103 (O_2103,N_24620,N_24727);
xor UO_2104 (O_2104,N_24996,N_24508);
xor UO_2105 (O_2105,N_24952,N_24593);
nor UO_2106 (O_2106,N_24541,N_24378);
nor UO_2107 (O_2107,N_24553,N_24771);
nand UO_2108 (O_2108,N_24645,N_24862);
xnor UO_2109 (O_2109,N_24986,N_24431);
xor UO_2110 (O_2110,N_24838,N_24544);
nor UO_2111 (O_2111,N_24855,N_24733);
and UO_2112 (O_2112,N_24945,N_24579);
and UO_2113 (O_2113,N_24735,N_24556);
nand UO_2114 (O_2114,N_24690,N_24788);
nor UO_2115 (O_2115,N_24839,N_24457);
nand UO_2116 (O_2116,N_24764,N_24535);
or UO_2117 (O_2117,N_24822,N_24998);
nand UO_2118 (O_2118,N_24791,N_24996);
or UO_2119 (O_2119,N_24779,N_24570);
nor UO_2120 (O_2120,N_24831,N_24935);
nor UO_2121 (O_2121,N_24422,N_24972);
nor UO_2122 (O_2122,N_24772,N_24943);
xor UO_2123 (O_2123,N_24597,N_24542);
and UO_2124 (O_2124,N_24860,N_24899);
xor UO_2125 (O_2125,N_24534,N_24886);
xor UO_2126 (O_2126,N_24915,N_24494);
nor UO_2127 (O_2127,N_24871,N_24552);
xor UO_2128 (O_2128,N_24712,N_24786);
and UO_2129 (O_2129,N_24385,N_24653);
or UO_2130 (O_2130,N_24420,N_24539);
and UO_2131 (O_2131,N_24899,N_24869);
nor UO_2132 (O_2132,N_24818,N_24801);
and UO_2133 (O_2133,N_24835,N_24993);
or UO_2134 (O_2134,N_24720,N_24464);
xnor UO_2135 (O_2135,N_24390,N_24910);
or UO_2136 (O_2136,N_24749,N_24736);
and UO_2137 (O_2137,N_24643,N_24450);
or UO_2138 (O_2138,N_24963,N_24675);
and UO_2139 (O_2139,N_24949,N_24605);
xnor UO_2140 (O_2140,N_24431,N_24497);
xor UO_2141 (O_2141,N_24496,N_24917);
nor UO_2142 (O_2142,N_24709,N_24929);
nor UO_2143 (O_2143,N_24710,N_24630);
or UO_2144 (O_2144,N_24841,N_24457);
or UO_2145 (O_2145,N_24562,N_24709);
nand UO_2146 (O_2146,N_24645,N_24579);
nand UO_2147 (O_2147,N_24462,N_24441);
nor UO_2148 (O_2148,N_24983,N_24686);
xnor UO_2149 (O_2149,N_24613,N_24630);
nor UO_2150 (O_2150,N_24451,N_24683);
and UO_2151 (O_2151,N_24444,N_24424);
nor UO_2152 (O_2152,N_24447,N_24597);
or UO_2153 (O_2153,N_24894,N_24390);
nor UO_2154 (O_2154,N_24815,N_24668);
nor UO_2155 (O_2155,N_24475,N_24810);
or UO_2156 (O_2156,N_24701,N_24842);
xor UO_2157 (O_2157,N_24790,N_24518);
or UO_2158 (O_2158,N_24896,N_24814);
nor UO_2159 (O_2159,N_24535,N_24990);
and UO_2160 (O_2160,N_24530,N_24833);
or UO_2161 (O_2161,N_24470,N_24941);
xnor UO_2162 (O_2162,N_24544,N_24896);
and UO_2163 (O_2163,N_24471,N_24655);
nor UO_2164 (O_2164,N_24583,N_24860);
xnor UO_2165 (O_2165,N_24796,N_24847);
xnor UO_2166 (O_2166,N_24700,N_24994);
and UO_2167 (O_2167,N_24454,N_24744);
nand UO_2168 (O_2168,N_24859,N_24505);
xnor UO_2169 (O_2169,N_24426,N_24960);
or UO_2170 (O_2170,N_24427,N_24471);
xor UO_2171 (O_2171,N_24657,N_24739);
nand UO_2172 (O_2172,N_24722,N_24861);
nor UO_2173 (O_2173,N_24708,N_24380);
or UO_2174 (O_2174,N_24650,N_24419);
xor UO_2175 (O_2175,N_24466,N_24964);
nor UO_2176 (O_2176,N_24894,N_24969);
or UO_2177 (O_2177,N_24867,N_24942);
nand UO_2178 (O_2178,N_24796,N_24592);
or UO_2179 (O_2179,N_24524,N_24407);
nand UO_2180 (O_2180,N_24613,N_24911);
nand UO_2181 (O_2181,N_24764,N_24664);
nor UO_2182 (O_2182,N_24541,N_24859);
and UO_2183 (O_2183,N_24832,N_24509);
xor UO_2184 (O_2184,N_24659,N_24398);
or UO_2185 (O_2185,N_24889,N_24718);
or UO_2186 (O_2186,N_24382,N_24875);
xor UO_2187 (O_2187,N_24726,N_24878);
or UO_2188 (O_2188,N_24935,N_24933);
nand UO_2189 (O_2189,N_24666,N_24669);
or UO_2190 (O_2190,N_24725,N_24798);
nand UO_2191 (O_2191,N_24475,N_24794);
and UO_2192 (O_2192,N_24649,N_24479);
xor UO_2193 (O_2193,N_24622,N_24605);
xnor UO_2194 (O_2194,N_24793,N_24915);
xnor UO_2195 (O_2195,N_24966,N_24518);
nand UO_2196 (O_2196,N_24699,N_24489);
nor UO_2197 (O_2197,N_24984,N_24843);
and UO_2198 (O_2198,N_24579,N_24860);
xor UO_2199 (O_2199,N_24858,N_24958);
or UO_2200 (O_2200,N_24682,N_24638);
or UO_2201 (O_2201,N_24649,N_24812);
nand UO_2202 (O_2202,N_24981,N_24634);
and UO_2203 (O_2203,N_24384,N_24854);
xor UO_2204 (O_2204,N_24797,N_24392);
nand UO_2205 (O_2205,N_24570,N_24491);
and UO_2206 (O_2206,N_24829,N_24558);
and UO_2207 (O_2207,N_24630,N_24502);
nor UO_2208 (O_2208,N_24882,N_24472);
or UO_2209 (O_2209,N_24864,N_24895);
nor UO_2210 (O_2210,N_24487,N_24948);
xor UO_2211 (O_2211,N_24825,N_24456);
and UO_2212 (O_2212,N_24702,N_24399);
or UO_2213 (O_2213,N_24441,N_24770);
nor UO_2214 (O_2214,N_24460,N_24786);
and UO_2215 (O_2215,N_24378,N_24563);
and UO_2216 (O_2216,N_24769,N_24486);
nor UO_2217 (O_2217,N_24700,N_24537);
nand UO_2218 (O_2218,N_24420,N_24964);
nand UO_2219 (O_2219,N_24425,N_24729);
xnor UO_2220 (O_2220,N_24704,N_24604);
nor UO_2221 (O_2221,N_24533,N_24979);
nand UO_2222 (O_2222,N_24590,N_24697);
or UO_2223 (O_2223,N_24569,N_24730);
and UO_2224 (O_2224,N_24534,N_24999);
nor UO_2225 (O_2225,N_24877,N_24749);
nand UO_2226 (O_2226,N_24413,N_24534);
or UO_2227 (O_2227,N_24900,N_24471);
and UO_2228 (O_2228,N_24464,N_24805);
xor UO_2229 (O_2229,N_24591,N_24722);
or UO_2230 (O_2230,N_24557,N_24990);
nor UO_2231 (O_2231,N_24821,N_24833);
nand UO_2232 (O_2232,N_24472,N_24632);
nand UO_2233 (O_2233,N_24590,N_24751);
or UO_2234 (O_2234,N_24453,N_24841);
xor UO_2235 (O_2235,N_24912,N_24772);
nor UO_2236 (O_2236,N_24675,N_24884);
xnor UO_2237 (O_2237,N_24663,N_24750);
and UO_2238 (O_2238,N_24942,N_24864);
xor UO_2239 (O_2239,N_24500,N_24810);
nor UO_2240 (O_2240,N_24583,N_24447);
nand UO_2241 (O_2241,N_24733,N_24752);
or UO_2242 (O_2242,N_24950,N_24585);
and UO_2243 (O_2243,N_24716,N_24486);
or UO_2244 (O_2244,N_24639,N_24875);
xor UO_2245 (O_2245,N_24465,N_24882);
and UO_2246 (O_2246,N_24547,N_24496);
or UO_2247 (O_2247,N_24765,N_24622);
xnor UO_2248 (O_2248,N_24996,N_24747);
and UO_2249 (O_2249,N_24775,N_24923);
nor UO_2250 (O_2250,N_24850,N_24795);
nand UO_2251 (O_2251,N_24795,N_24990);
xnor UO_2252 (O_2252,N_24548,N_24776);
and UO_2253 (O_2253,N_24484,N_24642);
nor UO_2254 (O_2254,N_24461,N_24463);
xnor UO_2255 (O_2255,N_24490,N_24676);
nand UO_2256 (O_2256,N_24836,N_24949);
xnor UO_2257 (O_2257,N_24773,N_24949);
nand UO_2258 (O_2258,N_24498,N_24906);
nor UO_2259 (O_2259,N_24937,N_24931);
nor UO_2260 (O_2260,N_24383,N_24812);
nand UO_2261 (O_2261,N_24899,N_24832);
nand UO_2262 (O_2262,N_24919,N_24951);
xor UO_2263 (O_2263,N_24810,N_24832);
or UO_2264 (O_2264,N_24699,N_24425);
or UO_2265 (O_2265,N_24705,N_24561);
and UO_2266 (O_2266,N_24745,N_24902);
nor UO_2267 (O_2267,N_24746,N_24443);
and UO_2268 (O_2268,N_24953,N_24835);
or UO_2269 (O_2269,N_24584,N_24582);
or UO_2270 (O_2270,N_24808,N_24914);
nor UO_2271 (O_2271,N_24874,N_24853);
and UO_2272 (O_2272,N_24999,N_24702);
xnor UO_2273 (O_2273,N_24480,N_24601);
nand UO_2274 (O_2274,N_24710,N_24640);
and UO_2275 (O_2275,N_24766,N_24401);
and UO_2276 (O_2276,N_24820,N_24893);
nand UO_2277 (O_2277,N_24418,N_24772);
nor UO_2278 (O_2278,N_24864,N_24448);
nor UO_2279 (O_2279,N_24377,N_24387);
and UO_2280 (O_2280,N_24467,N_24785);
or UO_2281 (O_2281,N_24894,N_24638);
xor UO_2282 (O_2282,N_24469,N_24887);
xor UO_2283 (O_2283,N_24645,N_24791);
or UO_2284 (O_2284,N_24928,N_24468);
xor UO_2285 (O_2285,N_24385,N_24581);
nand UO_2286 (O_2286,N_24772,N_24665);
and UO_2287 (O_2287,N_24955,N_24979);
xor UO_2288 (O_2288,N_24840,N_24402);
and UO_2289 (O_2289,N_24982,N_24823);
nand UO_2290 (O_2290,N_24647,N_24994);
and UO_2291 (O_2291,N_24712,N_24556);
and UO_2292 (O_2292,N_24711,N_24437);
nor UO_2293 (O_2293,N_24439,N_24809);
or UO_2294 (O_2294,N_24967,N_24604);
or UO_2295 (O_2295,N_24850,N_24378);
or UO_2296 (O_2296,N_24413,N_24792);
nand UO_2297 (O_2297,N_24665,N_24994);
or UO_2298 (O_2298,N_24803,N_24993);
nor UO_2299 (O_2299,N_24854,N_24970);
or UO_2300 (O_2300,N_24532,N_24730);
or UO_2301 (O_2301,N_24713,N_24384);
nor UO_2302 (O_2302,N_24673,N_24720);
nor UO_2303 (O_2303,N_24653,N_24878);
nor UO_2304 (O_2304,N_24967,N_24508);
xnor UO_2305 (O_2305,N_24853,N_24419);
xor UO_2306 (O_2306,N_24950,N_24724);
xnor UO_2307 (O_2307,N_24709,N_24583);
nand UO_2308 (O_2308,N_24682,N_24966);
or UO_2309 (O_2309,N_24436,N_24868);
nor UO_2310 (O_2310,N_24666,N_24686);
nor UO_2311 (O_2311,N_24404,N_24868);
nor UO_2312 (O_2312,N_24400,N_24495);
nor UO_2313 (O_2313,N_24609,N_24793);
or UO_2314 (O_2314,N_24386,N_24883);
nor UO_2315 (O_2315,N_24603,N_24775);
or UO_2316 (O_2316,N_24625,N_24954);
xnor UO_2317 (O_2317,N_24746,N_24541);
nor UO_2318 (O_2318,N_24831,N_24919);
xnor UO_2319 (O_2319,N_24591,N_24709);
nor UO_2320 (O_2320,N_24522,N_24837);
nand UO_2321 (O_2321,N_24751,N_24714);
and UO_2322 (O_2322,N_24441,N_24699);
nor UO_2323 (O_2323,N_24390,N_24436);
nor UO_2324 (O_2324,N_24808,N_24889);
or UO_2325 (O_2325,N_24691,N_24918);
nor UO_2326 (O_2326,N_24733,N_24622);
nor UO_2327 (O_2327,N_24710,N_24731);
and UO_2328 (O_2328,N_24475,N_24824);
and UO_2329 (O_2329,N_24601,N_24704);
xnor UO_2330 (O_2330,N_24451,N_24537);
nor UO_2331 (O_2331,N_24521,N_24813);
and UO_2332 (O_2332,N_24559,N_24407);
xnor UO_2333 (O_2333,N_24408,N_24698);
and UO_2334 (O_2334,N_24977,N_24594);
nor UO_2335 (O_2335,N_24866,N_24787);
and UO_2336 (O_2336,N_24487,N_24780);
nor UO_2337 (O_2337,N_24863,N_24578);
nor UO_2338 (O_2338,N_24898,N_24788);
or UO_2339 (O_2339,N_24604,N_24614);
or UO_2340 (O_2340,N_24721,N_24672);
nand UO_2341 (O_2341,N_24571,N_24376);
or UO_2342 (O_2342,N_24398,N_24679);
and UO_2343 (O_2343,N_24382,N_24812);
nor UO_2344 (O_2344,N_24524,N_24659);
or UO_2345 (O_2345,N_24596,N_24557);
or UO_2346 (O_2346,N_24623,N_24485);
xor UO_2347 (O_2347,N_24533,N_24684);
and UO_2348 (O_2348,N_24824,N_24988);
or UO_2349 (O_2349,N_24838,N_24791);
xnor UO_2350 (O_2350,N_24750,N_24561);
and UO_2351 (O_2351,N_24740,N_24876);
and UO_2352 (O_2352,N_24449,N_24833);
xnor UO_2353 (O_2353,N_24760,N_24483);
or UO_2354 (O_2354,N_24607,N_24936);
or UO_2355 (O_2355,N_24641,N_24796);
nor UO_2356 (O_2356,N_24417,N_24413);
nand UO_2357 (O_2357,N_24508,N_24542);
or UO_2358 (O_2358,N_24683,N_24972);
nor UO_2359 (O_2359,N_24580,N_24839);
and UO_2360 (O_2360,N_24755,N_24560);
and UO_2361 (O_2361,N_24770,N_24477);
and UO_2362 (O_2362,N_24573,N_24595);
xor UO_2363 (O_2363,N_24657,N_24481);
or UO_2364 (O_2364,N_24865,N_24842);
xnor UO_2365 (O_2365,N_24789,N_24585);
xnor UO_2366 (O_2366,N_24984,N_24649);
and UO_2367 (O_2367,N_24440,N_24896);
or UO_2368 (O_2368,N_24547,N_24541);
xor UO_2369 (O_2369,N_24556,N_24426);
nor UO_2370 (O_2370,N_24702,N_24690);
xor UO_2371 (O_2371,N_24497,N_24516);
or UO_2372 (O_2372,N_24499,N_24517);
nand UO_2373 (O_2373,N_24544,N_24529);
nand UO_2374 (O_2374,N_24963,N_24881);
nor UO_2375 (O_2375,N_24514,N_24913);
nand UO_2376 (O_2376,N_24862,N_24993);
xor UO_2377 (O_2377,N_24419,N_24503);
nor UO_2378 (O_2378,N_24396,N_24398);
xor UO_2379 (O_2379,N_24977,N_24909);
nand UO_2380 (O_2380,N_24522,N_24421);
xor UO_2381 (O_2381,N_24756,N_24444);
nand UO_2382 (O_2382,N_24405,N_24944);
nor UO_2383 (O_2383,N_24677,N_24624);
nand UO_2384 (O_2384,N_24612,N_24421);
and UO_2385 (O_2385,N_24586,N_24517);
nor UO_2386 (O_2386,N_24644,N_24919);
or UO_2387 (O_2387,N_24825,N_24533);
nand UO_2388 (O_2388,N_24950,N_24613);
nor UO_2389 (O_2389,N_24510,N_24971);
nand UO_2390 (O_2390,N_24414,N_24736);
xor UO_2391 (O_2391,N_24972,N_24874);
and UO_2392 (O_2392,N_24767,N_24488);
nor UO_2393 (O_2393,N_24629,N_24573);
xnor UO_2394 (O_2394,N_24720,N_24863);
nor UO_2395 (O_2395,N_24784,N_24945);
xnor UO_2396 (O_2396,N_24452,N_24467);
nor UO_2397 (O_2397,N_24399,N_24434);
nor UO_2398 (O_2398,N_24547,N_24993);
nor UO_2399 (O_2399,N_24817,N_24770);
nand UO_2400 (O_2400,N_24836,N_24845);
nand UO_2401 (O_2401,N_24955,N_24680);
and UO_2402 (O_2402,N_24523,N_24861);
nor UO_2403 (O_2403,N_24550,N_24704);
nand UO_2404 (O_2404,N_24865,N_24517);
nor UO_2405 (O_2405,N_24491,N_24452);
nand UO_2406 (O_2406,N_24661,N_24836);
or UO_2407 (O_2407,N_24506,N_24986);
nand UO_2408 (O_2408,N_24589,N_24984);
nand UO_2409 (O_2409,N_24858,N_24871);
or UO_2410 (O_2410,N_24727,N_24898);
and UO_2411 (O_2411,N_24592,N_24976);
and UO_2412 (O_2412,N_24898,N_24553);
and UO_2413 (O_2413,N_24977,N_24836);
nor UO_2414 (O_2414,N_24379,N_24830);
xnor UO_2415 (O_2415,N_24576,N_24431);
xor UO_2416 (O_2416,N_24394,N_24560);
nor UO_2417 (O_2417,N_24630,N_24962);
nor UO_2418 (O_2418,N_24634,N_24726);
or UO_2419 (O_2419,N_24982,N_24707);
xor UO_2420 (O_2420,N_24836,N_24999);
nand UO_2421 (O_2421,N_24732,N_24716);
or UO_2422 (O_2422,N_24618,N_24481);
and UO_2423 (O_2423,N_24905,N_24690);
xor UO_2424 (O_2424,N_24646,N_24387);
or UO_2425 (O_2425,N_24551,N_24854);
or UO_2426 (O_2426,N_24504,N_24375);
nand UO_2427 (O_2427,N_24410,N_24781);
nand UO_2428 (O_2428,N_24421,N_24751);
or UO_2429 (O_2429,N_24921,N_24740);
or UO_2430 (O_2430,N_24996,N_24469);
nor UO_2431 (O_2431,N_24708,N_24887);
nand UO_2432 (O_2432,N_24625,N_24574);
nand UO_2433 (O_2433,N_24978,N_24893);
xnor UO_2434 (O_2434,N_24849,N_24478);
nand UO_2435 (O_2435,N_24896,N_24846);
or UO_2436 (O_2436,N_24859,N_24957);
nor UO_2437 (O_2437,N_24922,N_24425);
xnor UO_2438 (O_2438,N_24774,N_24733);
or UO_2439 (O_2439,N_24747,N_24621);
or UO_2440 (O_2440,N_24811,N_24872);
nand UO_2441 (O_2441,N_24876,N_24573);
xnor UO_2442 (O_2442,N_24445,N_24978);
or UO_2443 (O_2443,N_24565,N_24769);
xnor UO_2444 (O_2444,N_24415,N_24875);
and UO_2445 (O_2445,N_24386,N_24843);
and UO_2446 (O_2446,N_24715,N_24470);
nand UO_2447 (O_2447,N_24509,N_24391);
or UO_2448 (O_2448,N_24762,N_24512);
nand UO_2449 (O_2449,N_24889,N_24545);
nand UO_2450 (O_2450,N_24692,N_24966);
or UO_2451 (O_2451,N_24684,N_24514);
xnor UO_2452 (O_2452,N_24727,N_24857);
and UO_2453 (O_2453,N_24956,N_24872);
nor UO_2454 (O_2454,N_24666,N_24634);
and UO_2455 (O_2455,N_24732,N_24840);
nand UO_2456 (O_2456,N_24890,N_24612);
and UO_2457 (O_2457,N_24708,N_24964);
nand UO_2458 (O_2458,N_24673,N_24934);
or UO_2459 (O_2459,N_24924,N_24700);
xnor UO_2460 (O_2460,N_24534,N_24839);
and UO_2461 (O_2461,N_24620,N_24681);
or UO_2462 (O_2462,N_24383,N_24490);
nor UO_2463 (O_2463,N_24689,N_24460);
xnor UO_2464 (O_2464,N_24390,N_24843);
xor UO_2465 (O_2465,N_24592,N_24811);
nand UO_2466 (O_2466,N_24583,N_24641);
nor UO_2467 (O_2467,N_24861,N_24846);
xnor UO_2468 (O_2468,N_24510,N_24698);
or UO_2469 (O_2469,N_24815,N_24747);
or UO_2470 (O_2470,N_24880,N_24980);
xor UO_2471 (O_2471,N_24728,N_24819);
or UO_2472 (O_2472,N_24821,N_24817);
nor UO_2473 (O_2473,N_24379,N_24859);
xnor UO_2474 (O_2474,N_24672,N_24903);
xor UO_2475 (O_2475,N_24491,N_24692);
nand UO_2476 (O_2476,N_24641,N_24762);
nand UO_2477 (O_2477,N_24913,N_24541);
nor UO_2478 (O_2478,N_24596,N_24463);
nand UO_2479 (O_2479,N_24674,N_24690);
nand UO_2480 (O_2480,N_24580,N_24544);
or UO_2481 (O_2481,N_24900,N_24648);
and UO_2482 (O_2482,N_24827,N_24770);
nand UO_2483 (O_2483,N_24388,N_24404);
and UO_2484 (O_2484,N_24562,N_24931);
nor UO_2485 (O_2485,N_24445,N_24990);
nand UO_2486 (O_2486,N_24461,N_24583);
nand UO_2487 (O_2487,N_24865,N_24827);
nand UO_2488 (O_2488,N_24499,N_24449);
xnor UO_2489 (O_2489,N_24607,N_24533);
nor UO_2490 (O_2490,N_24943,N_24939);
xnor UO_2491 (O_2491,N_24685,N_24851);
or UO_2492 (O_2492,N_24911,N_24414);
and UO_2493 (O_2493,N_24620,N_24611);
and UO_2494 (O_2494,N_24393,N_24747);
and UO_2495 (O_2495,N_24493,N_24731);
and UO_2496 (O_2496,N_24702,N_24957);
xor UO_2497 (O_2497,N_24783,N_24929);
nor UO_2498 (O_2498,N_24982,N_24436);
or UO_2499 (O_2499,N_24547,N_24699);
nor UO_2500 (O_2500,N_24484,N_24890);
nand UO_2501 (O_2501,N_24581,N_24749);
and UO_2502 (O_2502,N_24945,N_24928);
and UO_2503 (O_2503,N_24933,N_24762);
nor UO_2504 (O_2504,N_24898,N_24535);
and UO_2505 (O_2505,N_24548,N_24473);
nor UO_2506 (O_2506,N_24737,N_24455);
xnor UO_2507 (O_2507,N_24888,N_24974);
and UO_2508 (O_2508,N_24429,N_24800);
nor UO_2509 (O_2509,N_24822,N_24619);
nand UO_2510 (O_2510,N_24748,N_24952);
nor UO_2511 (O_2511,N_24786,N_24559);
and UO_2512 (O_2512,N_24979,N_24502);
xor UO_2513 (O_2513,N_24972,N_24971);
nor UO_2514 (O_2514,N_24826,N_24793);
nand UO_2515 (O_2515,N_24907,N_24584);
and UO_2516 (O_2516,N_24997,N_24615);
nor UO_2517 (O_2517,N_24704,N_24846);
xor UO_2518 (O_2518,N_24571,N_24490);
or UO_2519 (O_2519,N_24578,N_24593);
and UO_2520 (O_2520,N_24861,N_24569);
nand UO_2521 (O_2521,N_24487,N_24885);
xnor UO_2522 (O_2522,N_24743,N_24635);
nand UO_2523 (O_2523,N_24821,N_24661);
nor UO_2524 (O_2524,N_24880,N_24440);
nand UO_2525 (O_2525,N_24472,N_24990);
nand UO_2526 (O_2526,N_24960,N_24666);
nand UO_2527 (O_2527,N_24956,N_24564);
nand UO_2528 (O_2528,N_24984,N_24390);
and UO_2529 (O_2529,N_24965,N_24837);
and UO_2530 (O_2530,N_24793,N_24964);
xnor UO_2531 (O_2531,N_24802,N_24534);
xor UO_2532 (O_2532,N_24867,N_24918);
nor UO_2533 (O_2533,N_24995,N_24636);
xor UO_2534 (O_2534,N_24390,N_24854);
nand UO_2535 (O_2535,N_24646,N_24382);
nand UO_2536 (O_2536,N_24456,N_24415);
nand UO_2537 (O_2537,N_24817,N_24981);
nand UO_2538 (O_2538,N_24709,N_24798);
or UO_2539 (O_2539,N_24923,N_24616);
nand UO_2540 (O_2540,N_24810,N_24610);
xor UO_2541 (O_2541,N_24980,N_24808);
xor UO_2542 (O_2542,N_24844,N_24907);
xnor UO_2543 (O_2543,N_24502,N_24759);
nor UO_2544 (O_2544,N_24625,N_24721);
xor UO_2545 (O_2545,N_24544,N_24705);
nor UO_2546 (O_2546,N_24475,N_24803);
or UO_2547 (O_2547,N_24931,N_24568);
nor UO_2548 (O_2548,N_24485,N_24693);
xnor UO_2549 (O_2549,N_24981,N_24594);
nand UO_2550 (O_2550,N_24804,N_24915);
or UO_2551 (O_2551,N_24972,N_24700);
and UO_2552 (O_2552,N_24949,N_24707);
or UO_2553 (O_2553,N_24809,N_24595);
or UO_2554 (O_2554,N_24834,N_24602);
nand UO_2555 (O_2555,N_24661,N_24903);
xnor UO_2556 (O_2556,N_24944,N_24573);
and UO_2557 (O_2557,N_24920,N_24899);
or UO_2558 (O_2558,N_24926,N_24758);
xnor UO_2559 (O_2559,N_24486,N_24583);
xnor UO_2560 (O_2560,N_24540,N_24376);
xor UO_2561 (O_2561,N_24912,N_24803);
nand UO_2562 (O_2562,N_24499,N_24955);
or UO_2563 (O_2563,N_24868,N_24584);
xor UO_2564 (O_2564,N_24822,N_24517);
nand UO_2565 (O_2565,N_24516,N_24875);
nand UO_2566 (O_2566,N_24634,N_24952);
xnor UO_2567 (O_2567,N_24441,N_24784);
nand UO_2568 (O_2568,N_24743,N_24750);
or UO_2569 (O_2569,N_24794,N_24976);
nor UO_2570 (O_2570,N_24614,N_24820);
or UO_2571 (O_2571,N_24695,N_24772);
nand UO_2572 (O_2572,N_24868,N_24982);
nand UO_2573 (O_2573,N_24828,N_24948);
xor UO_2574 (O_2574,N_24937,N_24760);
and UO_2575 (O_2575,N_24959,N_24792);
xor UO_2576 (O_2576,N_24794,N_24400);
or UO_2577 (O_2577,N_24781,N_24970);
xor UO_2578 (O_2578,N_24729,N_24498);
and UO_2579 (O_2579,N_24825,N_24524);
nand UO_2580 (O_2580,N_24890,N_24686);
xnor UO_2581 (O_2581,N_24397,N_24872);
nor UO_2582 (O_2582,N_24876,N_24406);
nand UO_2583 (O_2583,N_24560,N_24741);
and UO_2584 (O_2584,N_24740,N_24580);
xnor UO_2585 (O_2585,N_24888,N_24620);
nand UO_2586 (O_2586,N_24562,N_24782);
xnor UO_2587 (O_2587,N_24976,N_24639);
and UO_2588 (O_2588,N_24514,N_24745);
and UO_2589 (O_2589,N_24779,N_24935);
nor UO_2590 (O_2590,N_24584,N_24770);
xor UO_2591 (O_2591,N_24574,N_24631);
nor UO_2592 (O_2592,N_24651,N_24955);
and UO_2593 (O_2593,N_24688,N_24924);
nor UO_2594 (O_2594,N_24598,N_24473);
nand UO_2595 (O_2595,N_24539,N_24996);
xnor UO_2596 (O_2596,N_24590,N_24909);
nand UO_2597 (O_2597,N_24727,N_24498);
nor UO_2598 (O_2598,N_24499,N_24629);
nor UO_2599 (O_2599,N_24690,N_24937);
xor UO_2600 (O_2600,N_24790,N_24843);
nor UO_2601 (O_2601,N_24737,N_24925);
xnor UO_2602 (O_2602,N_24445,N_24545);
nor UO_2603 (O_2603,N_24979,N_24792);
xor UO_2604 (O_2604,N_24750,N_24412);
and UO_2605 (O_2605,N_24460,N_24481);
xnor UO_2606 (O_2606,N_24810,N_24588);
or UO_2607 (O_2607,N_24504,N_24819);
or UO_2608 (O_2608,N_24540,N_24946);
nand UO_2609 (O_2609,N_24388,N_24855);
nand UO_2610 (O_2610,N_24692,N_24755);
nand UO_2611 (O_2611,N_24595,N_24377);
xor UO_2612 (O_2612,N_24979,N_24774);
or UO_2613 (O_2613,N_24995,N_24616);
and UO_2614 (O_2614,N_24491,N_24821);
nor UO_2615 (O_2615,N_24893,N_24532);
xnor UO_2616 (O_2616,N_24568,N_24898);
or UO_2617 (O_2617,N_24992,N_24418);
nor UO_2618 (O_2618,N_24903,N_24961);
xnor UO_2619 (O_2619,N_24967,N_24777);
nor UO_2620 (O_2620,N_24712,N_24451);
or UO_2621 (O_2621,N_24510,N_24722);
and UO_2622 (O_2622,N_24441,N_24725);
nor UO_2623 (O_2623,N_24830,N_24731);
nor UO_2624 (O_2624,N_24691,N_24621);
and UO_2625 (O_2625,N_24832,N_24386);
or UO_2626 (O_2626,N_24409,N_24480);
xor UO_2627 (O_2627,N_24687,N_24457);
or UO_2628 (O_2628,N_24603,N_24597);
nand UO_2629 (O_2629,N_24979,N_24415);
and UO_2630 (O_2630,N_24948,N_24912);
or UO_2631 (O_2631,N_24380,N_24796);
nor UO_2632 (O_2632,N_24639,N_24751);
nand UO_2633 (O_2633,N_24980,N_24717);
and UO_2634 (O_2634,N_24579,N_24614);
nor UO_2635 (O_2635,N_24729,N_24720);
nand UO_2636 (O_2636,N_24721,N_24558);
nand UO_2637 (O_2637,N_24806,N_24582);
nand UO_2638 (O_2638,N_24944,N_24500);
xnor UO_2639 (O_2639,N_24899,N_24493);
or UO_2640 (O_2640,N_24650,N_24456);
nor UO_2641 (O_2641,N_24969,N_24982);
or UO_2642 (O_2642,N_24821,N_24546);
xor UO_2643 (O_2643,N_24659,N_24938);
nand UO_2644 (O_2644,N_24934,N_24891);
xor UO_2645 (O_2645,N_24876,N_24632);
nor UO_2646 (O_2646,N_24626,N_24797);
xor UO_2647 (O_2647,N_24596,N_24465);
or UO_2648 (O_2648,N_24891,N_24376);
and UO_2649 (O_2649,N_24705,N_24920);
or UO_2650 (O_2650,N_24989,N_24542);
or UO_2651 (O_2651,N_24624,N_24702);
nor UO_2652 (O_2652,N_24677,N_24764);
or UO_2653 (O_2653,N_24403,N_24676);
or UO_2654 (O_2654,N_24634,N_24641);
and UO_2655 (O_2655,N_24477,N_24597);
or UO_2656 (O_2656,N_24820,N_24499);
or UO_2657 (O_2657,N_24865,N_24877);
nand UO_2658 (O_2658,N_24616,N_24408);
or UO_2659 (O_2659,N_24622,N_24802);
and UO_2660 (O_2660,N_24781,N_24768);
or UO_2661 (O_2661,N_24410,N_24761);
xnor UO_2662 (O_2662,N_24843,N_24855);
xnor UO_2663 (O_2663,N_24519,N_24505);
or UO_2664 (O_2664,N_24879,N_24848);
and UO_2665 (O_2665,N_24402,N_24417);
or UO_2666 (O_2666,N_24425,N_24702);
and UO_2667 (O_2667,N_24783,N_24651);
or UO_2668 (O_2668,N_24624,N_24781);
or UO_2669 (O_2669,N_24378,N_24990);
and UO_2670 (O_2670,N_24551,N_24544);
nand UO_2671 (O_2671,N_24878,N_24916);
nor UO_2672 (O_2672,N_24554,N_24674);
or UO_2673 (O_2673,N_24813,N_24538);
nor UO_2674 (O_2674,N_24858,N_24651);
or UO_2675 (O_2675,N_24636,N_24795);
nand UO_2676 (O_2676,N_24407,N_24975);
nor UO_2677 (O_2677,N_24606,N_24617);
or UO_2678 (O_2678,N_24376,N_24386);
xor UO_2679 (O_2679,N_24666,N_24592);
nand UO_2680 (O_2680,N_24652,N_24779);
or UO_2681 (O_2681,N_24835,N_24753);
nor UO_2682 (O_2682,N_24985,N_24911);
or UO_2683 (O_2683,N_24821,N_24999);
nand UO_2684 (O_2684,N_24558,N_24582);
nand UO_2685 (O_2685,N_24940,N_24787);
or UO_2686 (O_2686,N_24439,N_24885);
xor UO_2687 (O_2687,N_24628,N_24969);
and UO_2688 (O_2688,N_24475,N_24921);
nor UO_2689 (O_2689,N_24699,N_24645);
nand UO_2690 (O_2690,N_24915,N_24549);
xor UO_2691 (O_2691,N_24772,N_24776);
nor UO_2692 (O_2692,N_24561,N_24467);
nor UO_2693 (O_2693,N_24499,N_24544);
or UO_2694 (O_2694,N_24771,N_24835);
xnor UO_2695 (O_2695,N_24436,N_24380);
nor UO_2696 (O_2696,N_24466,N_24817);
nor UO_2697 (O_2697,N_24667,N_24854);
xnor UO_2698 (O_2698,N_24395,N_24854);
or UO_2699 (O_2699,N_24472,N_24523);
or UO_2700 (O_2700,N_24658,N_24934);
and UO_2701 (O_2701,N_24944,N_24504);
and UO_2702 (O_2702,N_24766,N_24882);
nand UO_2703 (O_2703,N_24908,N_24501);
nor UO_2704 (O_2704,N_24410,N_24997);
nor UO_2705 (O_2705,N_24886,N_24748);
and UO_2706 (O_2706,N_24971,N_24640);
or UO_2707 (O_2707,N_24712,N_24903);
nor UO_2708 (O_2708,N_24671,N_24894);
nand UO_2709 (O_2709,N_24433,N_24402);
nor UO_2710 (O_2710,N_24651,N_24462);
or UO_2711 (O_2711,N_24890,N_24709);
and UO_2712 (O_2712,N_24494,N_24696);
nor UO_2713 (O_2713,N_24860,N_24800);
or UO_2714 (O_2714,N_24387,N_24418);
and UO_2715 (O_2715,N_24399,N_24932);
xnor UO_2716 (O_2716,N_24598,N_24448);
or UO_2717 (O_2717,N_24909,N_24783);
or UO_2718 (O_2718,N_24884,N_24651);
xnor UO_2719 (O_2719,N_24580,N_24887);
or UO_2720 (O_2720,N_24584,N_24799);
or UO_2721 (O_2721,N_24791,N_24655);
and UO_2722 (O_2722,N_24976,N_24468);
xnor UO_2723 (O_2723,N_24974,N_24839);
and UO_2724 (O_2724,N_24735,N_24435);
and UO_2725 (O_2725,N_24956,N_24523);
nand UO_2726 (O_2726,N_24914,N_24905);
xor UO_2727 (O_2727,N_24427,N_24514);
or UO_2728 (O_2728,N_24592,N_24638);
or UO_2729 (O_2729,N_24898,N_24825);
nand UO_2730 (O_2730,N_24477,N_24854);
nor UO_2731 (O_2731,N_24604,N_24787);
and UO_2732 (O_2732,N_24866,N_24804);
and UO_2733 (O_2733,N_24609,N_24791);
and UO_2734 (O_2734,N_24841,N_24694);
and UO_2735 (O_2735,N_24542,N_24701);
and UO_2736 (O_2736,N_24754,N_24746);
and UO_2737 (O_2737,N_24434,N_24509);
nand UO_2738 (O_2738,N_24505,N_24883);
nor UO_2739 (O_2739,N_24915,N_24952);
nand UO_2740 (O_2740,N_24842,N_24562);
nor UO_2741 (O_2741,N_24594,N_24608);
xor UO_2742 (O_2742,N_24966,N_24536);
or UO_2743 (O_2743,N_24601,N_24891);
or UO_2744 (O_2744,N_24436,N_24964);
xnor UO_2745 (O_2745,N_24786,N_24852);
and UO_2746 (O_2746,N_24492,N_24568);
and UO_2747 (O_2747,N_24854,N_24443);
and UO_2748 (O_2748,N_24721,N_24933);
xor UO_2749 (O_2749,N_24780,N_24592);
nand UO_2750 (O_2750,N_24541,N_24503);
nand UO_2751 (O_2751,N_24921,N_24832);
nand UO_2752 (O_2752,N_24462,N_24959);
nor UO_2753 (O_2753,N_24505,N_24406);
and UO_2754 (O_2754,N_24377,N_24621);
nand UO_2755 (O_2755,N_24653,N_24394);
or UO_2756 (O_2756,N_24471,N_24815);
nand UO_2757 (O_2757,N_24991,N_24463);
nand UO_2758 (O_2758,N_24557,N_24988);
nand UO_2759 (O_2759,N_24870,N_24881);
or UO_2760 (O_2760,N_24897,N_24969);
xnor UO_2761 (O_2761,N_24808,N_24502);
nor UO_2762 (O_2762,N_24837,N_24886);
nor UO_2763 (O_2763,N_24449,N_24630);
or UO_2764 (O_2764,N_24471,N_24890);
and UO_2765 (O_2765,N_24601,N_24724);
nor UO_2766 (O_2766,N_24607,N_24879);
or UO_2767 (O_2767,N_24805,N_24392);
or UO_2768 (O_2768,N_24607,N_24669);
nor UO_2769 (O_2769,N_24659,N_24601);
nand UO_2770 (O_2770,N_24656,N_24913);
nand UO_2771 (O_2771,N_24513,N_24890);
nand UO_2772 (O_2772,N_24436,N_24899);
nand UO_2773 (O_2773,N_24430,N_24923);
or UO_2774 (O_2774,N_24938,N_24660);
and UO_2775 (O_2775,N_24616,N_24499);
or UO_2776 (O_2776,N_24708,N_24483);
xor UO_2777 (O_2777,N_24883,N_24446);
nor UO_2778 (O_2778,N_24426,N_24596);
xor UO_2779 (O_2779,N_24510,N_24804);
and UO_2780 (O_2780,N_24548,N_24851);
or UO_2781 (O_2781,N_24750,N_24642);
nor UO_2782 (O_2782,N_24557,N_24648);
xnor UO_2783 (O_2783,N_24600,N_24486);
nor UO_2784 (O_2784,N_24453,N_24895);
xnor UO_2785 (O_2785,N_24396,N_24400);
nand UO_2786 (O_2786,N_24783,N_24999);
nand UO_2787 (O_2787,N_24459,N_24451);
nor UO_2788 (O_2788,N_24942,N_24396);
or UO_2789 (O_2789,N_24957,N_24607);
xor UO_2790 (O_2790,N_24775,N_24670);
xor UO_2791 (O_2791,N_24674,N_24780);
and UO_2792 (O_2792,N_24521,N_24397);
nor UO_2793 (O_2793,N_24584,N_24659);
nand UO_2794 (O_2794,N_24537,N_24787);
and UO_2795 (O_2795,N_24795,N_24408);
or UO_2796 (O_2796,N_24630,N_24703);
xor UO_2797 (O_2797,N_24562,N_24914);
and UO_2798 (O_2798,N_24994,N_24536);
nand UO_2799 (O_2799,N_24968,N_24879);
xnor UO_2800 (O_2800,N_24594,N_24716);
and UO_2801 (O_2801,N_24541,N_24608);
or UO_2802 (O_2802,N_24657,N_24655);
xnor UO_2803 (O_2803,N_24775,N_24749);
nand UO_2804 (O_2804,N_24623,N_24721);
xnor UO_2805 (O_2805,N_24950,N_24944);
nand UO_2806 (O_2806,N_24588,N_24485);
nor UO_2807 (O_2807,N_24671,N_24432);
or UO_2808 (O_2808,N_24841,N_24635);
nand UO_2809 (O_2809,N_24824,N_24501);
nand UO_2810 (O_2810,N_24429,N_24574);
or UO_2811 (O_2811,N_24424,N_24733);
or UO_2812 (O_2812,N_24838,N_24861);
nand UO_2813 (O_2813,N_24711,N_24397);
xor UO_2814 (O_2814,N_24491,N_24424);
and UO_2815 (O_2815,N_24645,N_24837);
xnor UO_2816 (O_2816,N_24662,N_24819);
nor UO_2817 (O_2817,N_24727,N_24493);
xor UO_2818 (O_2818,N_24565,N_24846);
xnor UO_2819 (O_2819,N_24872,N_24990);
or UO_2820 (O_2820,N_24402,N_24962);
and UO_2821 (O_2821,N_24547,N_24955);
nand UO_2822 (O_2822,N_24566,N_24587);
nand UO_2823 (O_2823,N_24873,N_24478);
xor UO_2824 (O_2824,N_24540,N_24616);
nor UO_2825 (O_2825,N_24884,N_24670);
and UO_2826 (O_2826,N_24376,N_24944);
nand UO_2827 (O_2827,N_24406,N_24825);
nor UO_2828 (O_2828,N_24665,N_24643);
or UO_2829 (O_2829,N_24778,N_24577);
xnor UO_2830 (O_2830,N_24688,N_24563);
xnor UO_2831 (O_2831,N_24890,N_24606);
xor UO_2832 (O_2832,N_24902,N_24750);
nor UO_2833 (O_2833,N_24889,N_24407);
nand UO_2834 (O_2834,N_24852,N_24972);
nor UO_2835 (O_2835,N_24407,N_24718);
xor UO_2836 (O_2836,N_24445,N_24696);
and UO_2837 (O_2837,N_24728,N_24441);
xnor UO_2838 (O_2838,N_24518,N_24540);
nor UO_2839 (O_2839,N_24871,N_24791);
nor UO_2840 (O_2840,N_24897,N_24504);
and UO_2841 (O_2841,N_24482,N_24919);
nor UO_2842 (O_2842,N_24889,N_24452);
nor UO_2843 (O_2843,N_24882,N_24712);
or UO_2844 (O_2844,N_24991,N_24539);
xor UO_2845 (O_2845,N_24665,N_24773);
xor UO_2846 (O_2846,N_24714,N_24534);
and UO_2847 (O_2847,N_24901,N_24844);
nand UO_2848 (O_2848,N_24450,N_24928);
nor UO_2849 (O_2849,N_24757,N_24965);
xnor UO_2850 (O_2850,N_24691,N_24770);
nor UO_2851 (O_2851,N_24483,N_24379);
xor UO_2852 (O_2852,N_24702,N_24533);
xor UO_2853 (O_2853,N_24488,N_24388);
or UO_2854 (O_2854,N_24629,N_24608);
xor UO_2855 (O_2855,N_24450,N_24932);
or UO_2856 (O_2856,N_24865,N_24609);
and UO_2857 (O_2857,N_24575,N_24571);
or UO_2858 (O_2858,N_24831,N_24724);
nand UO_2859 (O_2859,N_24770,N_24960);
and UO_2860 (O_2860,N_24682,N_24993);
or UO_2861 (O_2861,N_24807,N_24390);
nor UO_2862 (O_2862,N_24870,N_24561);
nand UO_2863 (O_2863,N_24391,N_24834);
or UO_2864 (O_2864,N_24534,N_24661);
and UO_2865 (O_2865,N_24720,N_24632);
or UO_2866 (O_2866,N_24610,N_24874);
or UO_2867 (O_2867,N_24778,N_24523);
nor UO_2868 (O_2868,N_24497,N_24797);
nand UO_2869 (O_2869,N_24590,N_24814);
xnor UO_2870 (O_2870,N_24558,N_24430);
nand UO_2871 (O_2871,N_24806,N_24815);
xor UO_2872 (O_2872,N_24720,N_24840);
nor UO_2873 (O_2873,N_24669,N_24755);
or UO_2874 (O_2874,N_24476,N_24570);
nand UO_2875 (O_2875,N_24661,N_24403);
nand UO_2876 (O_2876,N_24739,N_24755);
nand UO_2877 (O_2877,N_24438,N_24852);
or UO_2878 (O_2878,N_24460,N_24798);
or UO_2879 (O_2879,N_24725,N_24611);
xor UO_2880 (O_2880,N_24792,N_24624);
nand UO_2881 (O_2881,N_24564,N_24434);
xnor UO_2882 (O_2882,N_24772,N_24500);
or UO_2883 (O_2883,N_24649,N_24831);
or UO_2884 (O_2884,N_24448,N_24997);
nand UO_2885 (O_2885,N_24424,N_24728);
xnor UO_2886 (O_2886,N_24791,N_24884);
or UO_2887 (O_2887,N_24528,N_24492);
or UO_2888 (O_2888,N_24785,N_24654);
xor UO_2889 (O_2889,N_24753,N_24656);
xnor UO_2890 (O_2890,N_24490,N_24940);
nor UO_2891 (O_2891,N_24758,N_24412);
xnor UO_2892 (O_2892,N_24867,N_24719);
nand UO_2893 (O_2893,N_24541,N_24858);
or UO_2894 (O_2894,N_24563,N_24706);
nand UO_2895 (O_2895,N_24619,N_24716);
and UO_2896 (O_2896,N_24448,N_24660);
xnor UO_2897 (O_2897,N_24557,N_24606);
nand UO_2898 (O_2898,N_24502,N_24920);
nor UO_2899 (O_2899,N_24774,N_24705);
and UO_2900 (O_2900,N_24996,N_24401);
xor UO_2901 (O_2901,N_24653,N_24969);
nand UO_2902 (O_2902,N_24774,N_24922);
nand UO_2903 (O_2903,N_24915,N_24656);
nand UO_2904 (O_2904,N_24621,N_24882);
or UO_2905 (O_2905,N_24680,N_24585);
xor UO_2906 (O_2906,N_24999,N_24751);
nand UO_2907 (O_2907,N_24652,N_24667);
nor UO_2908 (O_2908,N_24781,N_24952);
xnor UO_2909 (O_2909,N_24657,N_24421);
xnor UO_2910 (O_2910,N_24687,N_24531);
nor UO_2911 (O_2911,N_24849,N_24515);
and UO_2912 (O_2912,N_24766,N_24991);
or UO_2913 (O_2913,N_24515,N_24415);
or UO_2914 (O_2914,N_24658,N_24626);
xor UO_2915 (O_2915,N_24679,N_24750);
and UO_2916 (O_2916,N_24701,N_24755);
and UO_2917 (O_2917,N_24680,N_24801);
xor UO_2918 (O_2918,N_24438,N_24955);
nand UO_2919 (O_2919,N_24590,N_24416);
nor UO_2920 (O_2920,N_24498,N_24788);
and UO_2921 (O_2921,N_24743,N_24659);
nand UO_2922 (O_2922,N_24975,N_24854);
and UO_2923 (O_2923,N_24542,N_24678);
or UO_2924 (O_2924,N_24537,N_24919);
nand UO_2925 (O_2925,N_24879,N_24630);
or UO_2926 (O_2926,N_24797,N_24603);
nand UO_2927 (O_2927,N_24663,N_24734);
nand UO_2928 (O_2928,N_24775,N_24404);
nand UO_2929 (O_2929,N_24596,N_24852);
and UO_2930 (O_2930,N_24842,N_24678);
nand UO_2931 (O_2931,N_24819,N_24676);
and UO_2932 (O_2932,N_24540,N_24770);
nand UO_2933 (O_2933,N_24617,N_24568);
or UO_2934 (O_2934,N_24563,N_24968);
or UO_2935 (O_2935,N_24815,N_24842);
nand UO_2936 (O_2936,N_24656,N_24606);
or UO_2937 (O_2937,N_24408,N_24593);
and UO_2938 (O_2938,N_24527,N_24953);
nand UO_2939 (O_2939,N_24772,N_24716);
nor UO_2940 (O_2940,N_24755,N_24909);
nor UO_2941 (O_2941,N_24686,N_24867);
xor UO_2942 (O_2942,N_24704,N_24505);
nor UO_2943 (O_2943,N_24800,N_24406);
or UO_2944 (O_2944,N_24828,N_24999);
or UO_2945 (O_2945,N_24864,N_24518);
xor UO_2946 (O_2946,N_24423,N_24572);
or UO_2947 (O_2947,N_24719,N_24510);
and UO_2948 (O_2948,N_24386,N_24851);
or UO_2949 (O_2949,N_24732,N_24901);
nand UO_2950 (O_2950,N_24732,N_24823);
nor UO_2951 (O_2951,N_24805,N_24914);
nand UO_2952 (O_2952,N_24876,N_24813);
or UO_2953 (O_2953,N_24736,N_24670);
and UO_2954 (O_2954,N_24432,N_24401);
xor UO_2955 (O_2955,N_24901,N_24787);
nor UO_2956 (O_2956,N_24540,N_24759);
or UO_2957 (O_2957,N_24606,N_24509);
or UO_2958 (O_2958,N_24663,N_24654);
and UO_2959 (O_2959,N_24462,N_24916);
and UO_2960 (O_2960,N_24528,N_24467);
nand UO_2961 (O_2961,N_24405,N_24790);
or UO_2962 (O_2962,N_24890,N_24457);
nor UO_2963 (O_2963,N_24827,N_24868);
nor UO_2964 (O_2964,N_24912,N_24572);
and UO_2965 (O_2965,N_24812,N_24982);
xnor UO_2966 (O_2966,N_24753,N_24818);
or UO_2967 (O_2967,N_24878,N_24542);
nand UO_2968 (O_2968,N_24440,N_24800);
and UO_2969 (O_2969,N_24430,N_24903);
or UO_2970 (O_2970,N_24921,N_24662);
nor UO_2971 (O_2971,N_24657,N_24744);
xnor UO_2972 (O_2972,N_24694,N_24977);
or UO_2973 (O_2973,N_24388,N_24723);
nand UO_2974 (O_2974,N_24526,N_24912);
or UO_2975 (O_2975,N_24409,N_24450);
or UO_2976 (O_2976,N_24418,N_24793);
xnor UO_2977 (O_2977,N_24897,N_24566);
nor UO_2978 (O_2978,N_24449,N_24496);
and UO_2979 (O_2979,N_24518,N_24998);
nand UO_2980 (O_2980,N_24882,N_24841);
and UO_2981 (O_2981,N_24422,N_24452);
and UO_2982 (O_2982,N_24739,N_24741);
and UO_2983 (O_2983,N_24390,N_24686);
xnor UO_2984 (O_2984,N_24758,N_24840);
or UO_2985 (O_2985,N_24755,N_24420);
xnor UO_2986 (O_2986,N_24805,N_24680);
or UO_2987 (O_2987,N_24425,N_24738);
xor UO_2988 (O_2988,N_24635,N_24932);
and UO_2989 (O_2989,N_24504,N_24474);
and UO_2990 (O_2990,N_24765,N_24681);
and UO_2991 (O_2991,N_24552,N_24577);
and UO_2992 (O_2992,N_24756,N_24972);
nand UO_2993 (O_2993,N_24573,N_24574);
nand UO_2994 (O_2994,N_24745,N_24483);
nand UO_2995 (O_2995,N_24758,N_24644);
or UO_2996 (O_2996,N_24599,N_24467);
nand UO_2997 (O_2997,N_24753,N_24435);
nand UO_2998 (O_2998,N_24776,N_24928);
or UO_2999 (O_2999,N_24927,N_24645);
endmodule