module basic_1000_10000_1500_2_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5005,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5018,N_5019,N_5020,N_5021,N_5022,N_5024,N_5028,N_5030,N_5031,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5046,N_5047,N_5048,N_5049,N_5052,N_5054,N_5055,N_5056,N_5057,N_5058,N_5060,N_5062,N_5064,N_5067,N_5068,N_5070,N_5074,N_5078,N_5080,N_5081,N_5083,N_5084,N_5087,N_5088,N_5090,N_5093,N_5094,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5105,N_5109,N_5110,N_5111,N_5112,N_5114,N_5115,N_5116,N_5118,N_5119,N_5120,N_5121,N_5123,N_5125,N_5126,N_5127,N_5128,N_5129,N_5134,N_5135,N_5136,N_5138,N_5139,N_5141,N_5142,N_5143,N_5144,N_5146,N_5147,N_5150,N_5151,N_5153,N_5155,N_5158,N_5159,N_5160,N_5161,N_5163,N_5165,N_5167,N_5168,N_5169,N_5170,N_5172,N_5173,N_5177,N_5178,N_5180,N_5181,N_5183,N_5185,N_5186,N_5188,N_5189,N_5190,N_5192,N_5194,N_5196,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5207,N_5208,N_5209,N_5213,N_5214,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5231,N_5233,N_5234,N_5238,N_5239,N_5242,N_5245,N_5247,N_5248,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5263,N_5264,N_5265,N_5266,N_5267,N_5269,N_5270,N_5271,N_5273,N_5274,N_5275,N_5276,N_5277,N_5280,N_5281,N_5283,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5294,N_5297,N_5298,N_5299,N_5301,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5311,N_5313,N_5317,N_5318,N_5321,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5332,N_5333,N_5334,N_5335,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5348,N_5351,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5360,N_5361,N_5362,N_5363,N_5366,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5375,N_5377,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5391,N_5398,N_5400,N_5401,N_5403,N_5406,N_5407,N_5408,N_5413,N_5415,N_5418,N_5419,N_5421,N_5425,N_5426,N_5427,N_5428,N_5430,N_5432,N_5433,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5443,N_5445,N_5446,N_5450,N_5452,N_5456,N_5458,N_5460,N_5461,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5476,N_5478,N_5480,N_5481,N_5482,N_5486,N_5487,N_5488,N_5492,N_5493,N_5497,N_5500,N_5501,N_5503,N_5505,N_5506,N_5507,N_5508,N_5509,N_5511,N_5512,N_5513,N_5514,N_5517,N_5518,N_5519,N_5521,N_5522,N_5523,N_5524,N_5526,N_5527,N_5531,N_5532,N_5533,N_5536,N_5538,N_5539,N_5540,N_5541,N_5544,N_5545,N_5548,N_5551,N_5554,N_5560,N_5563,N_5564,N_5567,N_5568,N_5571,N_5572,N_5573,N_5576,N_5577,N_5579,N_5582,N_5583,N_5587,N_5588,N_5589,N_5591,N_5594,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5603,N_5604,N_5606,N_5607,N_5608,N_5609,N_5610,N_5616,N_5619,N_5620,N_5621,N_5622,N_5625,N_5626,N_5627,N_5628,N_5630,N_5631,N_5632,N_5634,N_5637,N_5639,N_5640,N_5644,N_5645,N_5646,N_5651,N_5652,N_5653,N_5654,N_5655,N_5658,N_5659,N_5660,N_5661,N_5662,N_5664,N_5665,N_5666,N_5668,N_5671,N_5672,N_5673,N_5677,N_5680,N_5681,N_5683,N_5685,N_5686,N_5688,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5701,N_5705,N_5707,N_5708,N_5709,N_5711,N_5713,N_5714,N_5715,N_5717,N_5718,N_5722,N_5723,N_5725,N_5726,N_5728,N_5730,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5741,N_5742,N_5743,N_5746,N_5748,N_5749,N_5751,N_5756,N_5757,N_5758,N_5759,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5769,N_5770,N_5771,N_5772,N_5774,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5786,N_5791,N_5793,N_5795,N_5796,N_5797,N_5800,N_5801,N_5802,N_5804,N_5806,N_5807,N_5810,N_5811,N_5813,N_5814,N_5816,N_5820,N_5821,N_5822,N_5823,N_5824,N_5826,N_5828,N_5829,N_5830,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5842,N_5844,N_5845,N_5846,N_5847,N_5848,N_5851,N_5852,N_5858,N_5859,N_5862,N_5863,N_5864,N_5865,N_5866,N_5868,N_5869,N_5870,N_5873,N_5874,N_5876,N_5877,N_5878,N_5879,N_5881,N_5883,N_5885,N_5886,N_5888,N_5891,N_5892,N_5895,N_5897,N_5899,N_5900,N_5902,N_5905,N_5908,N_5910,N_5912,N_5915,N_5916,N_5917,N_5918,N_5920,N_5921,N_5924,N_5925,N_5927,N_5930,N_5932,N_5933,N_5935,N_5936,N_5938,N_5939,N_5941,N_5942,N_5943,N_5944,N_5946,N_5947,N_5949,N_5951,N_5952,N_5954,N_5955,N_5956,N_5958,N_5959,N_5960,N_5962,N_5964,N_5965,N_5967,N_5968,N_5970,N_5971,N_5972,N_5975,N_5976,N_5977,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5989,N_5992,N_5993,N_5994,N_5996,N_5997,N_5998,N_6000,N_6001,N_6002,N_6003,N_6005,N_6007,N_6008,N_6010,N_6017,N_6019,N_6023,N_6024,N_6025,N_6026,N_6028,N_6030,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6044,N_6047,N_6049,N_6053,N_6056,N_6057,N_6060,N_6061,N_6063,N_6069,N_6071,N_6073,N_6075,N_6076,N_6078,N_6079,N_6080,N_6081,N_6082,N_6088,N_6092,N_6093,N_6094,N_6095,N_6097,N_6098,N_6099,N_6100,N_6103,N_6104,N_6106,N_6107,N_6109,N_6110,N_6111,N_6112,N_6115,N_6116,N_6117,N_6120,N_6121,N_6122,N_6125,N_6126,N_6127,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6139,N_6140,N_6142,N_6143,N_6146,N_6147,N_6151,N_6153,N_6155,N_6156,N_6157,N_6160,N_6161,N_6163,N_6164,N_6166,N_6167,N_6168,N_6171,N_6172,N_6176,N_6177,N_6180,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6192,N_6193,N_6195,N_6196,N_6197,N_6198,N_6202,N_6205,N_6209,N_6210,N_6211,N_6212,N_6213,N_6217,N_6218,N_6219,N_6220,N_6222,N_6223,N_6224,N_6225,N_6228,N_6229,N_6232,N_6235,N_6237,N_6238,N_6239,N_6241,N_6242,N_6243,N_6245,N_6249,N_6250,N_6254,N_6255,N_6256,N_6259,N_6260,N_6263,N_6264,N_6267,N_6268,N_6269,N_6270,N_6271,N_6273,N_6275,N_6279,N_6281,N_6284,N_6288,N_6289,N_6292,N_6293,N_6295,N_6296,N_6297,N_6298,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6318,N_6320,N_6321,N_6322,N_6325,N_6327,N_6328,N_6330,N_6331,N_6332,N_6334,N_6335,N_6336,N_6338,N_6339,N_6340,N_6344,N_6345,N_6346,N_6347,N_6351,N_6353,N_6354,N_6356,N_6357,N_6361,N_6362,N_6363,N_6369,N_6371,N_6372,N_6373,N_6378,N_6379,N_6381,N_6384,N_6385,N_6386,N_6387,N_6390,N_6391,N_6393,N_6394,N_6395,N_6398,N_6400,N_6401,N_6403,N_6405,N_6406,N_6408,N_6409,N_6411,N_6413,N_6414,N_6415,N_6417,N_6418,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6428,N_6429,N_6431,N_6433,N_6436,N_6440,N_6441,N_6443,N_6445,N_6447,N_6448,N_6451,N_6453,N_6455,N_6456,N_6458,N_6459,N_6463,N_6464,N_6465,N_6467,N_6468,N_6469,N_6470,N_6473,N_6474,N_6475,N_6477,N_6481,N_6484,N_6485,N_6488,N_6490,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6501,N_6502,N_6503,N_6504,N_6505,N_6508,N_6510,N_6512,N_6515,N_6516,N_6517,N_6518,N_6520,N_6521,N_6522,N_6523,N_6525,N_6526,N_6527,N_6528,N_6530,N_6532,N_6533,N_6534,N_6536,N_6539,N_6540,N_6541,N_6542,N_6547,N_6549,N_6557,N_6558,N_6559,N_6560,N_6561,N_6563,N_6564,N_6565,N_6566,N_6568,N_6569,N_6572,N_6573,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6583,N_6584,N_6587,N_6592,N_6595,N_6596,N_6598,N_6599,N_6601,N_6602,N_6607,N_6608,N_6609,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6619,N_6620,N_6621,N_6622,N_6624,N_6626,N_6629,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6640,N_6641,N_6643,N_6645,N_6647,N_6650,N_6651,N_6653,N_6655,N_6656,N_6658,N_6659,N_6660,N_6661,N_6663,N_6665,N_6667,N_6668,N_6672,N_6674,N_6675,N_6676,N_6677,N_6678,N_6680,N_6681,N_6682,N_6683,N_6687,N_6690,N_6692,N_6694,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6705,N_6707,N_6708,N_6709,N_6710,N_6711,N_6713,N_6714,N_6715,N_6716,N_6717,N_6719,N_6720,N_6723,N_6725,N_6727,N_6729,N_6732,N_6734,N_6735,N_6736,N_6737,N_6738,N_6740,N_6742,N_6745,N_6749,N_6750,N_6752,N_6755,N_6757,N_6760,N_6761,N_6764,N_6765,N_6766,N_6767,N_6768,N_6770,N_6771,N_6773,N_6774,N_6776,N_6777,N_6779,N_6780,N_6781,N_6782,N_6783,N_6786,N_6787,N_6789,N_6791,N_6793,N_6794,N_6795,N_6796,N_6798,N_6799,N_6801,N_6802,N_6804,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6823,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6833,N_6834,N_6835,N_6837,N_6838,N_6840,N_6846,N_6848,N_6852,N_6853,N_6854,N_6855,N_6857,N_6858,N_6859,N_6860,N_6863,N_6864,N_6865,N_6866,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6875,N_6877,N_6878,N_6880,N_6883,N_6884,N_6885,N_6887,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6899,N_6900,N_6901,N_6903,N_6905,N_6906,N_6908,N_6912,N_6913,N_6914,N_6918,N_6919,N_6922,N_6923,N_6927,N_6930,N_6935,N_6937,N_6939,N_6941,N_6942,N_6943,N_6944,N_6948,N_6949,N_6951,N_6954,N_6955,N_6956,N_6959,N_6960,N_6961,N_6962,N_6963,N_6965,N_6967,N_6968,N_6969,N_6971,N_6972,N_6973,N_6975,N_6976,N_6981,N_6982,N_6984,N_6987,N_6988,N_6989,N_6990,N_6994,N_6995,N_6996,N_6998,N_7000,N_7002,N_7003,N_7004,N_7005,N_7006,N_7008,N_7009,N_7010,N_7013,N_7014,N_7015,N_7018,N_7019,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7028,N_7029,N_7032,N_7033,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7043,N_7044,N_7045,N_7046,N_7048,N_7049,N_7051,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7061,N_7062,N_7065,N_7066,N_7067,N_7068,N_7069,N_7071,N_7072,N_7074,N_7075,N_7077,N_7079,N_7080,N_7082,N_7083,N_7084,N_7085,N_7090,N_7091,N_7092,N_7094,N_7095,N_7096,N_7097,N_7099,N_7101,N_7102,N_7104,N_7105,N_7106,N_7109,N_7111,N_7112,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7124,N_7128,N_7131,N_7132,N_7133,N_7137,N_7139,N_7142,N_7144,N_7146,N_7148,N_7149,N_7152,N_7154,N_7155,N_7156,N_7162,N_7163,N_7168,N_7169,N_7170,N_7173,N_7174,N_7175,N_7176,N_7179,N_7180,N_7182,N_7184,N_7185,N_7186,N_7188,N_7189,N_7191,N_7194,N_7195,N_7196,N_7198,N_7200,N_7202,N_7203,N_7204,N_7205,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7217,N_7220,N_7221,N_7222,N_7224,N_7225,N_7226,N_7229,N_7233,N_7235,N_7236,N_7237,N_7240,N_7242,N_7243,N_7246,N_7248,N_7249,N_7250,N_7252,N_7253,N_7257,N_7261,N_7262,N_7263,N_7265,N_7266,N_7269,N_7270,N_7272,N_7273,N_7275,N_7276,N_7277,N_7279,N_7280,N_7282,N_7283,N_7285,N_7288,N_7289,N_7290,N_7292,N_7293,N_7295,N_7296,N_7297,N_7298,N_7302,N_7303,N_7305,N_7306,N_7307,N_7310,N_7313,N_7317,N_7318,N_7320,N_7325,N_7327,N_7328,N_7330,N_7332,N_7336,N_7338,N_7341,N_7342,N_7343,N_7344,N_7347,N_7348,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7360,N_7361,N_7362,N_7366,N_7367,N_7369,N_7370,N_7371,N_7372,N_7373,N_7375,N_7378,N_7380,N_7383,N_7384,N_7388,N_7391,N_7393,N_7396,N_7397,N_7400,N_7401,N_7402,N_7403,N_7405,N_7409,N_7413,N_7414,N_7416,N_7417,N_7420,N_7421,N_7424,N_7425,N_7427,N_7428,N_7431,N_7432,N_7433,N_7434,N_7436,N_7438,N_7439,N_7440,N_7442,N_7444,N_7450,N_7451,N_7454,N_7455,N_7457,N_7458,N_7460,N_7461,N_7463,N_7464,N_7466,N_7468,N_7470,N_7471,N_7475,N_7476,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7488,N_7490,N_7492,N_7493,N_7494,N_7495,N_7497,N_7498,N_7500,N_7501,N_7502,N_7503,N_7506,N_7508,N_7509,N_7510,N_7511,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7522,N_7523,N_7524,N_7525,N_7526,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7536,N_7537,N_7539,N_7542,N_7544,N_7545,N_7547,N_7548,N_7549,N_7550,N_7552,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7569,N_7570,N_7573,N_7574,N_7578,N_7579,N_7580,N_7582,N_7583,N_7586,N_7587,N_7588,N_7590,N_7591,N_7595,N_7596,N_7597,N_7598,N_7600,N_7602,N_7603,N_7604,N_7606,N_7607,N_7609,N_7610,N_7611,N_7614,N_7617,N_7618,N_7620,N_7623,N_7624,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7634,N_7636,N_7637,N_7638,N_7639,N_7641,N_7643,N_7647,N_7650,N_7651,N_7652,N_7653,N_7655,N_7657,N_7658,N_7659,N_7662,N_7663,N_7665,N_7668,N_7670,N_7672,N_7673,N_7675,N_7677,N_7678,N_7679,N_7681,N_7682,N_7683,N_7685,N_7686,N_7688,N_7689,N_7690,N_7692,N_7693,N_7695,N_7697,N_7698,N_7704,N_7705,N_7706,N_7708,N_7709,N_7710,N_7711,N_7712,N_7714,N_7716,N_7717,N_7718,N_7720,N_7725,N_7726,N_7727,N_7728,N_7731,N_7732,N_7733,N_7735,N_7736,N_7739,N_7740,N_7741,N_7742,N_7745,N_7746,N_7747,N_7749,N_7752,N_7753,N_7754,N_7755,N_7757,N_7758,N_7760,N_7761,N_7764,N_7765,N_7767,N_7770,N_7772,N_7773,N_7778,N_7779,N_7781,N_7783,N_7785,N_7787,N_7790,N_7793,N_7794,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7805,N_7806,N_7808,N_7809,N_7812,N_7813,N_7815,N_7816,N_7818,N_7819,N_7820,N_7823,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7836,N_7838,N_7839,N_7840,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7853,N_7855,N_7856,N_7857,N_7859,N_7861,N_7862,N_7865,N_7866,N_7869,N_7870,N_7871,N_7873,N_7874,N_7879,N_7880,N_7882,N_7883,N_7886,N_7887,N_7889,N_7892,N_7893,N_7895,N_7896,N_7898,N_7900,N_7902,N_7903,N_7906,N_7907,N_7908,N_7910,N_7911,N_7912,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7923,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7943,N_7945,N_7947,N_7948,N_7949,N_7952,N_7955,N_7957,N_7958,N_7960,N_7961,N_7962,N_7964,N_7966,N_7967,N_7968,N_7969,N_7971,N_7974,N_7976,N_7978,N_7979,N_7981,N_7983,N_7984,N_7985,N_7987,N_7988,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7999,N_8001,N_8002,N_8003,N_8005,N_8014,N_8015,N_8016,N_8017,N_8019,N_8020,N_8022,N_8024,N_8027,N_8028,N_8030,N_8031,N_8032,N_8034,N_8036,N_8037,N_8039,N_8043,N_8045,N_8046,N_8048,N_8050,N_8051,N_8052,N_8053,N_8054,N_8056,N_8058,N_8059,N_8061,N_8062,N_8064,N_8065,N_8066,N_8067,N_8070,N_8071,N_8073,N_8074,N_8075,N_8076,N_8078,N_8079,N_8081,N_8086,N_8087,N_8088,N_8089,N_8090,N_8094,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8114,N_8115,N_8117,N_8118,N_8119,N_8124,N_8125,N_8126,N_8127,N_8128,N_8130,N_8131,N_8132,N_8134,N_8136,N_8137,N_8138,N_8143,N_8144,N_8145,N_8146,N_8147,N_8149,N_8150,N_8155,N_8156,N_8160,N_8162,N_8164,N_8165,N_8166,N_8168,N_8171,N_8176,N_8180,N_8183,N_8184,N_8186,N_8187,N_8188,N_8191,N_8193,N_8194,N_8196,N_8200,N_8201,N_8202,N_8203,N_8204,N_8206,N_8210,N_8212,N_8213,N_8214,N_8215,N_8219,N_8220,N_8223,N_8226,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8240,N_8241,N_8245,N_8246,N_8247,N_8250,N_8253,N_8254,N_8256,N_8257,N_8260,N_8261,N_8262,N_8265,N_8266,N_8268,N_8271,N_8272,N_8273,N_8276,N_8278,N_8279,N_8280,N_8281,N_8282,N_8285,N_8288,N_8290,N_8292,N_8293,N_8294,N_8295,N_8296,N_8299,N_8300,N_8303,N_8305,N_8306,N_8308,N_8309,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8322,N_8323,N_8325,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8334,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8343,N_8344,N_8345,N_8346,N_8348,N_8349,N_8350,N_8352,N_8354,N_8355,N_8356,N_8357,N_8359,N_8360,N_8361,N_8362,N_8363,N_8366,N_8368,N_8374,N_8375,N_8376,N_8378,N_8380,N_8381,N_8382,N_8385,N_8386,N_8387,N_8389,N_8390,N_8391,N_8392,N_8394,N_8395,N_8397,N_8398,N_8400,N_8401,N_8404,N_8405,N_8406,N_8407,N_8408,N_8410,N_8411,N_8412,N_8413,N_8414,N_8419,N_8420,N_8422,N_8423,N_8424,N_8425,N_8427,N_8429,N_8430,N_8431,N_8434,N_8437,N_8444,N_8446,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8457,N_8460,N_8461,N_8466,N_8469,N_8471,N_8475,N_8477,N_8478,N_8480,N_8481,N_8482,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8494,N_8495,N_8496,N_8497,N_8498,N_8500,N_8501,N_8502,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8513,N_8515,N_8516,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8530,N_8531,N_8532,N_8534,N_8535,N_8537,N_8538,N_8539,N_8540,N_8543,N_8544,N_8545,N_8547,N_8548,N_8549,N_8550,N_8551,N_8553,N_8554,N_8556,N_8559,N_8560,N_8561,N_8562,N_8564,N_8565,N_8566,N_8568,N_8569,N_8570,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8582,N_8583,N_8584,N_8586,N_8587,N_8589,N_8591,N_8592,N_8597,N_8598,N_8599,N_8602,N_8603,N_8604,N_8605,N_8606,N_8608,N_8610,N_8612,N_8614,N_8616,N_8617,N_8618,N_8619,N_8620,N_8622,N_8624,N_8626,N_8627,N_8628,N_8631,N_8632,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8641,N_8643,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8652,N_8653,N_8655,N_8657,N_8659,N_8660,N_8662,N_8665,N_8667,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8676,N_8677,N_8680,N_8681,N_8683,N_8684,N_8686,N_8688,N_8689,N_8690,N_8691,N_8693,N_8694,N_8696,N_8697,N_8698,N_8699,N_8701,N_8702,N_8703,N_8704,N_8705,N_8707,N_8712,N_8713,N_8714,N_8715,N_8718,N_8720,N_8722,N_8728,N_8730,N_8731,N_8732,N_8734,N_8735,N_8736,N_8737,N_8739,N_8740,N_8742,N_8743,N_8749,N_8752,N_8753,N_8754,N_8755,N_8757,N_8758,N_8759,N_8761,N_8763,N_8764,N_8766,N_8768,N_8770,N_8772,N_8773,N_8775,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8787,N_8788,N_8790,N_8793,N_8794,N_8796,N_8797,N_8800,N_8804,N_8806,N_8808,N_8809,N_8815,N_8816,N_8819,N_8820,N_8821,N_8822,N_8823,N_8826,N_8827,N_8829,N_8830,N_8831,N_8833,N_8836,N_8837,N_8838,N_8840,N_8843,N_8844,N_8847,N_8850,N_8852,N_8853,N_8854,N_8857,N_8858,N_8862,N_8865,N_8868,N_8870,N_8871,N_8872,N_8873,N_8875,N_8876,N_8880,N_8881,N_8884,N_8885,N_8887,N_8889,N_8890,N_8891,N_8892,N_8896,N_8898,N_8899,N_8900,N_8902,N_8903,N_8904,N_8906,N_8908,N_8909,N_8910,N_8914,N_8916,N_8922,N_8923,N_8924,N_8926,N_8929,N_8930,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8940,N_8941,N_8942,N_8943,N_8948,N_8949,N_8950,N_8952,N_8954,N_8956,N_8957,N_8959,N_8960,N_8961,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8971,N_8972,N_8975,N_8976,N_8977,N_8979,N_8980,N_8981,N_8982,N_8984,N_8985,N_8986,N_8987,N_8988,N_8990,N_8991,N_8994,N_8995,N_8996,N_9000,N_9003,N_9004,N_9005,N_9006,N_9008,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9018,N_9019,N_9021,N_9022,N_9023,N_9024,N_9026,N_9027,N_9028,N_9029,N_9030,N_9032,N_9035,N_9040,N_9041,N_9042,N_9043,N_9045,N_9046,N_9048,N_9050,N_9051,N_9054,N_9056,N_9058,N_9059,N_9060,N_9064,N_9066,N_9067,N_9070,N_9073,N_9074,N_9076,N_9078,N_9079,N_9080,N_9087,N_9089,N_9090,N_9091,N_9092,N_9093,N_9095,N_9097,N_9098,N_9099,N_9100,N_9103,N_9104,N_9105,N_9107,N_9111,N_9113,N_9116,N_9118,N_9119,N_9121,N_9122,N_9126,N_9128,N_9130,N_9131,N_9133,N_9135,N_9136,N_9138,N_9139,N_9141,N_9142,N_9143,N_9144,N_9146,N_9147,N_9151,N_9154,N_9156,N_9157,N_9159,N_9160,N_9161,N_9166,N_9167,N_9168,N_9169,N_9172,N_9173,N_9177,N_9181,N_9184,N_9186,N_9187,N_9188,N_9189,N_9190,N_9192,N_9194,N_9195,N_9196,N_9197,N_9200,N_9202,N_9205,N_9206,N_9207,N_9208,N_9210,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9222,N_9224,N_9225,N_9226,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9238,N_9239,N_9241,N_9243,N_9244,N_9245,N_9246,N_9250,N_9251,N_9252,N_9253,N_9257,N_9258,N_9263,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9275,N_9276,N_9277,N_9278,N_9280,N_9282,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9297,N_9298,N_9299,N_9302,N_9306,N_9307,N_9308,N_9312,N_9315,N_9316,N_9317,N_9318,N_9320,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9337,N_9338,N_9339,N_9340,N_9341,N_9343,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9353,N_9355,N_9357,N_9358,N_9360,N_9363,N_9367,N_9369,N_9371,N_9372,N_9374,N_9377,N_9379,N_9380,N_9381,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9390,N_9397,N_9398,N_9400,N_9401,N_9402,N_9404,N_9406,N_9412,N_9413,N_9415,N_9418,N_9422,N_9424,N_9425,N_9426,N_9427,N_9430,N_9431,N_9432,N_9433,N_9435,N_9436,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9448,N_9449,N_9451,N_9453,N_9454,N_9455,N_9457,N_9458,N_9459,N_9460,N_9461,N_9465,N_9466,N_9467,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9477,N_9478,N_9480,N_9481,N_9482,N_9483,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9496,N_9497,N_9498,N_9501,N_9503,N_9505,N_9507,N_9509,N_9510,N_9513,N_9514,N_9516,N_9518,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9527,N_9528,N_9530,N_9532,N_9533,N_9534,N_9536,N_9537,N_9544,N_9545,N_9546,N_9549,N_9550,N_9556,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9567,N_9569,N_9570,N_9573,N_9574,N_9575,N_9578,N_9580,N_9581,N_9582,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9595,N_9597,N_9598,N_9599,N_9600,N_9601,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9611,N_9612,N_9613,N_9614,N_9618,N_9619,N_9621,N_9623,N_9624,N_9625,N_9626,N_9629,N_9631,N_9632,N_9633,N_9635,N_9638,N_9639,N_9641,N_9642,N_9643,N_9644,N_9646,N_9649,N_9650,N_9651,N_9652,N_9655,N_9659,N_9661,N_9662,N_9665,N_9666,N_9669,N_9670,N_9672,N_9673,N_9675,N_9676,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9686,N_9688,N_9689,N_9690,N_9692,N_9694,N_9695,N_9697,N_9698,N_9699,N_9700,N_9702,N_9703,N_9704,N_9705,N_9706,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9719,N_9722,N_9724,N_9725,N_9726,N_9727,N_9729,N_9730,N_9731,N_9735,N_9737,N_9738,N_9740,N_9741,N_9742,N_9744,N_9745,N_9747,N_9748,N_9749,N_9751,N_9755,N_9756,N_9757,N_9758,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9770,N_9771,N_9772,N_9774,N_9775,N_9776,N_9778,N_9780,N_9781,N_9783,N_9784,N_9785,N_9786,N_9789,N_9790,N_9791,N_9792,N_9794,N_9795,N_9796,N_9799,N_9801,N_9802,N_9805,N_9806,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9817,N_9818,N_9820,N_9822,N_9824,N_9825,N_9827,N_9828,N_9830,N_9832,N_9833,N_9835,N_9837,N_9838,N_9840,N_9841,N_9842,N_9845,N_9846,N_9850,N_9851,N_9852,N_9856,N_9858,N_9860,N_9861,N_9862,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9872,N_9873,N_9875,N_9876,N_9878,N_9879,N_9880,N_9882,N_9883,N_9885,N_9888,N_9889,N_9891,N_9893,N_9894,N_9897,N_9899,N_9900,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9911,N_9912,N_9913,N_9915,N_9918,N_9919,N_9920,N_9922,N_9923,N_9924,N_9925,N_9926,N_9929,N_9935,N_9936,N_9937,N_9938,N_9940,N_9941,N_9942,N_9944,N_9947,N_9950,N_9951,N_9953,N_9954,N_9956,N_9958,N_9959,N_9962,N_9963,N_9968,N_9970,N_9971,N_9972,N_9974,N_9975,N_9976,N_9979,N_9980,N_9982,N_9985,N_9986,N_9987,N_9990,N_9992,N_9995,N_9996,N_9998,N_9999;
nand U0 (N_0,In_172,In_826);
xnor U1 (N_1,In_47,In_565);
nor U2 (N_2,In_898,In_653);
and U3 (N_3,In_243,In_261);
nand U4 (N_4,In_500,In_603);
and U5 (N_5,In_964,In_840);
nor U6 (N_6,In_893,In_525);
or U7 (N_7,In_389,In_360);
nor U8 (N_8,In_775,In_599);
nand U9 (N_9,In_288,In_585);
and U10 (N_10,In_274,In_221);
or U11 (N_11,In_999,In_395);
nand U12 (N_12,In_43,In_91);
or U13 (N_13,In_861,In_841);
nor U14 (N_14,In_75,In_535);
nor U15 (N_15,In_687,In_33);
and U16 (N_16,In_204,In_141);
nor U17 (N_17,In_988,In_2);
nor U18 (N_18,In_680,In_758);
nand U19 (N_19,In_304,In_386);
or U20 (N_20,In_921,In_245);
and U21 (N_21,In_991,In_662);
nand U22 (N_22,In_798,In_875);
nand U23 (N_23,In_786,In_588);
or U24 (N_24,In_96,In_617);
or U25 (N_25,In_441,In_517);
or U26 (N_26,In_495,In_300);
nand U27 (N_27,In_628,In_374);
and U28 (N_28,In_199,In_170);
nor U29 (N_29,In_709,In_895);
nor U30 (N_30,In_416,In_472);
or U31 (N_31,In_747,In_338);
nor U32 (N_32,In_460,In_498);
nor U33 (N_33,In_524,In_166);
and U34 (N_34,In_636,In_11);
nor U35 (N_35,In_244,In_275);
and U36 (N_36,In_570,In_787);
and U37 (N_37,In_18,In_104);
nand U38 (N_38,In_185,In_849);
and U39 (N_39,In_228,In_337);
nand U40 (N_40,In_986,In_555);
nor U41 (N_41,In_331,In_522);
or U42 (N_42,In_82,In_449);
or U43 (N_43,In_865,In_324);
nor U44 (N_44,In_349,In_982);
and U45 (N_45,In_286,In_150);
and U46 (N_46,In_812,In_891);
nor U47 (N_47,In_962,In_76);
and U48 (N_48,In_423,In_39);
nand U49 (N_49,In_216,In_607);
and U50 (N_50,In_147,In_435);
and U51 (N_51,In_790,In_480);
nand U52 (N_52,In_897,In_259);
nor U53 (N_53,In_579,In_698);
or U54 (N_54,In_487,In_720);
nor U55 (N_55,In_795,In_377);
nand U56 (N_56,In_192,In_551);
and U57 (N_57,In_239,In_542);
or U58 (N_58,In_410,In_268);
and U59 (N_59,In_92,In_685);
nor U60 (N_60,In_129,In_618);
nand U61 (N_61,In_792,In_208);
or U62 (N_62,In_568,In_142);
and U63 (N_63,In_538,In_572);
nor U64 (N_64,In_691,In_532);
nand U65 (N_65,In_944,In_526);
xnor U66 (N_66,In_753,In_871);
nor U67 (N_67,In_120,In_347);
or U68 (N_68,In_706,In_272);
or U69 (N_69,In_462,In_649);
nor U70 (N_70,In_146,In_137);
and U71 (N_71,In_844,In_143);
nor U72 (N_72,In_475,In_598);
and U73 (N_73,In_519,In_317);
nand U74 (N_74,In_101,In_877);
nand U75 (N_75,In_868,In_589);
or U76 (N_76,In_132,In_866);
nand U77 (N_77,In_486,In_333);
and U78 (N_78,In_631,In_520);
nor U79 (N_79,In_556,In_455);
and U80 (N_80,In_447,In_413);
and U81 (N_81,In_906,In_408);
or U82 (N_82,In_515,In_796);
nor U83 (N_83,In_94,In_181);
nand U84 (N_84,In_914,In_443);
nor U85 (N_85,In_332,In_38);
or U86 (N_86,In_434,In_432);
and U87 (N_87,In_516,In_828);
nor U88 (N_88,In_483,In_390);
and U89 (N_89,In_7,In_123);
nor U90 (N_90,In_417,In_64);
or U91 (N_91,In_811,In_270);
xor U92 (N_92,In_450,In_543);
nor U93 (N_93,In_567,In_174);
and U94 (N_94,In_552,In_260);
and U95 (N_95,In_289,In_399);
or U96 (N_96,In_477,In_665);
nor U97 (N_97,In_754,In_683);
nor U98 (N_98,In_514,In_308);
nand U99 (N_99,In_630,In_148);
and U100 (N_100,In_739,In_712);
nand U101 (N_101,In_819,In_452);
and U102 (N_102,In_501,In_666);
xnor U103 (N_103,In_87,In_160);
nor U104 (N_104,In_122,In_98);
and U105 (N_105,In_79,In_801);
nand U106 (N_106,In_206,In_207);
nand U107 (N_107,In_745,In_909);
nor U108 (N_108,In_257,In_523);
nor U109 (N_109,In_505,In_521);
nor U110 (N_110,In_113,In_127);
or U111 (N_111,In_643,In_211);
nor U112 (N_112,In_121,In_886);
and U113 (N_113,In_365,In_664);
and U114 (N_114,In_156,In_608);
nand U115 (N_115,In_717,In_729);
or U116 (N_116,In_346,In_913);
or U117 (N_117,In_470,In_320);
or U118 (N_118,In_985,In_917);
nor U119 (N_119,In_702,In_529);
and U120 (N_120,In_103,In_230);
nand U121 (N_121,In_345,In_135);
nand U122 (N_122,In_357,In_380);
and U123 (N_123,In_836,In_864);
or U124 (N_124,In_961,In_249);
nand U125 (N_125,In_610,In_157);
or U126 (N_126,In_454,In_387);
and U127 (N_127,In_298,In_492);
nand U128 (N_128,In_488,In_158);
nand U129 (N_129,In_634,In_889);
nor U130 (N_130,In_838,In_496);
nand U131 (N_131,In_9,In_553);
and U132 (N_132,In_167,In_918);
or U133 (N_133,In_959,In_409);
and U134 (N_134,In_303,In_214);
nor U135 (N_135,In_932,In_301);
and U136 (N_136,In_433,In_892);
and U137 (N_137,In_266,In_925);
nor U138 (N_138,In_419,In_837);
or U139 (N_139,In_90,In_253);
nand U140 (N_140,In_48,In_859);
and U141 (N_141,In_30,In_537);
and U142 (N_142,In_15,In_931);
or U143 (N_143,In_130,In_993);
xnor U144 (N_144,In_863,In_491);
and U145 (N_145,In_686,In_88);
nand U146 (N_146,In_267,In_651);
and U147 (N_147,In_363,In_471);
and U148 (N_148,In_581,In_466);
or U149 (N_149,In_707,In_963);
or U150 (N_150,In_518,In_392);
nand U151 (N_151,In_912,In_592);
or U152 (N_152,In_883,In_933);
nor U153 (N_153,In_546,In_670);
and U154 (N_154,In_711,In_995);
nand U155 (N_155,In_590,In_955);
or U156 (N_156,In_847,In_42);
or U157 (N_157,In_809,In_149);
nor U158 (N_158,In_557,In_330);
or U159 (N_159,In_671,In_764);
or U160 (N_160,In_641,In_766);
nand U161 (N_161,In_839,In_922);
nor U162 (N_162,In_726,In_852);
and U163 (N_163,In_222,In_705);
nor U164 (N_164,In_58,In_759);
or U165 (N_165,In_371,In_278);
nor U166 (N_166,In_956,In_545);
or U167 (N_167,In_252,In_818);
or U168 (N_168,In_297,In_139);
nand U169 (N_169,In_689,In_153);
and U170 (N_170,In_508,In_507);
nand U171 (N_171,In_782,In_623);
nand U172 (N_172,In_165,In_5);
or U173 (N_173,In_669,In_894);
nor U174 (N_174,In_478,In_601);
or U175 (N_175,In_700,In_315);
nand U176 (N_176,In_305,In_737);
xnor U177 (N_177,In_824,In_247);
or U178 (N_178,In_973,In_456);
and U179 (N_179,In_976,In_559);
or U180 (N_180,In_348,In_370);
nand U181 (N_181,In_611,In_202);
nand U182 (N_182,In_731,In_406);
and U183 (N_183,In_95,In_437);
and U184 (N_184,In_888,In_342);
nand U185 (N_185,In_168,In_781);
or U186 (N_186,In_509,In_162);
and U187 (N_187,In_882,In_548);
or U188 (N_188,In_860,In_924);
and U189 (N_189,In_69,In_242);
and U190 (N_190,In_372,In_210);
and U191 (N_191,In_177,In_996);
or U192 (N_192,In_646,In_562);
nor U193 (N_193,In_458,In_41);
and U194 (N_194,In_476,In_779);
or U195 (N_195,In_527,In_264);
nand U196 (N_196,In_53,In_533);
or U197 (N_197,In_436,In_547);
and U198 (N_198,In_85,In_269);
or U199 (N_199,In_904,In_960);
and U200 (N_200,In_953,In_391);
or U201 (N_201,In_12,In_594);
nand U202 (N_202,In_979,In_424);
and U203 (N_203,In_738,In_970);
and U204 (N_204,In_614,In_334);
and U205 (N_205,In_639,In_299);
or U206 (N_206,In_273,In_195);
nor U207 (N_207,In_684,In_474);
nor U208 (N_208,In_901,In_655);
and U209 (N_209,In_439,In_171);
nand U210 (N_210,In_13,In_81);
nand U211 (N_211,In_695,In_540);
nor U212 (N_212,In_549,In_55);
nor U213 (N_213,In_226,In_874);
or U214 (N_214,In_727,In_715);
and U215 (N_215,In_341,In_907);
nand U216 (N_216,In_791,In_678);
nand U217 (N_217,In_23,In_378);
or U218 (N_218,In_743,In_881);
or U219 (N_219,In_654,In_279);
nor U220 (N_220,In_635,In_93);
and U221 (N_221,In_28,In_934);
nand U222 (N_222,In_760,In_251);
nand U223 (N_223,In_822,In_708);
nor U224 (N_224,In_459,In_644);
nand U225 (N_225,In_701,In_312);
and U226 (N_226,In_780,In_319);
or U227 (N_227,In_994,In_998);
nor U228 (N_228,In_848,In_750);
nand U229 (N_229,In_144,In_867);
or U230 (N_230,In_975,In_248);
and U231 (N_231,In_350,In_952);
or U232 (N_232,In_612,In_600);
nand U233 (N_233,In_935,In_554);
or U234 (N_234,In_770,In_367);
and U235 (N_235,In_361,In_619);
xnor U236 (N_236,In_971,In_467);
nand U237 (N_237,In_605,In_677);
and U238 (N_238,In_663,In_650);
or U239 (N_239,In_930,In_566);
and U240 (N_240,In_421,In_311);
or U241 (N_241,In_783,In_464);
and U242 (N_242,In_400,In_37);
or U243 (N_243,In_942,In_70);
and U244 (N_244,In_788,In_673);
nor U245 (N_245,In_203,In_768);
nand U246 (N_246,In_173,In_744);
nand U247 (N_247,In_870,In_723);
nor U248 (N_248,In_806,In_52);
nor U249 (N_249,In_675,In_394);
or U250 (N_250,In_880,In_558);
nor U251 (N_251,In_494,In_564);
nand U252 (N_252,In_544,In_989);
nor U253 (N_253,In_68,In_481);
and U254 (N_254,In_746,In_100);
and U255 (N_255,In_929,In_180);
nor U256 (N_256,In_418,In_777);
or U257 (N_257,In_896,In_984);
nor U258 (N_258,In_794,In_957);
or U259 (N_259,In_280,In_80);
and U260 (N_260,In_941,In_969);
and U261 (N_261,In_159,In_78);
nor U262 (N_262,In_306,In_106);
or U263 (N_263,In_232,In_722);
or U264 (N_264,In_164,In_107);
nand U265 (N_265,In_696,In_108);
and U266 (N_266,In_429,In_110);
nor U267 (N_267,In_10,In_17);
or U268 (N_268,In_490,In_352);
nor U269 (N_269,In_182,In_679);
or U270 (N_270,In_974,In_937);
nor U271 (N_271,In_749,In_31);
nand U272 (N_272,In_1,In_858);
and U273 (N_273,In_613,In_947);
nor U274 (N_274,In_234,In_927);
or U275 (N_275,In_431,In_940);
or U276 (N_276,In_810,In_294);
and U277 (N_277,In_152,In_807);
and U278 (N_278,In_595,In_569);
or U279 (N_279,In_189,In_624);
or U280 (N_280,In_813,In_936);
xor U281 (N_281,In_329,In_710);
and U282 (N_282,In_339,In_19);
and U283 (N_283,In_682,In_425);
or U284 (N_284,In_946,In_577);
and U285 (N_285,In_161,In_29);
and U286 (N_286,In_111,In_402);
nor U287 (N_287,In_560,In_125);
and U288 (N_288,In_676,In_427);
nand U289 (N_289,In_51,In_405);
or U290 (N_290,In_49,In_422);
or U291 (N_291,In_194,In_283);
nand U292 (N_292,In_178,In_183);
nand U293 (N_293,In_902,In_850);
nand U294 (N_294,In_923,In_154);
nor U295 (N_295,In_528,In_815);
or U296 (N_296,In_659,In_797);
nand U297 (N_297,In_733,In_384);
and U298 (N_298,In_116,In_948);
or U299 (N_299,In_295,In_151);
or U300 (N_300,In_622,In_531);
or U301 (N_301,In_714,In_713);
or U302 (N_302,In_6,In_784);
nand U303 (N_303,In_401,In_224);
nand U304 (N_304,In_276,In_939);
nor U305 (N_305,In_366,In_382);
nor U306 (N_306,In_716,In_851);
nor U307 (N_307,In_503,In_642);
or U308 (N_308,In_905,In_328);
or U309 (N_309,In_415,In_582);
nor U310 (N_310,In_128,In_992);
and U311 (N_311,In_778,In_314);
nand U312 (N_312,In_751,In_351);
nor U313 (N_313,In_291,In_219);
and U314 (N_314,In_246,In_225);
nand U315 (N_315,In_661,In_561);
nor U316 (N_316,In_853,In_184);
nor U317 (N_317,In_626,In_587);
and U318 (N_318,In_950,In_536);
or U319 (N_319,In_463,In_752);
nand U320 (N_320,In_385,In_198);
or U321 (N_321,In_854,In_430);
xor U322 (N_322,In_40,In_951);
nand U323 (N_323,In_97,In_802);
nand U324 (N_324,In_602,In_823);
and U325 (N_325,In_117,In_24);
and U326 (N_326,In_857,In_187);
or U327 (N_327,In_292,In_61);
nand U328 (N_328,In_282,In_681);
nand U329 (N_329,In_445,In_223);
and U330 (N_330,In_911,In_502);
nand U331 (N_331,In_672,In_571);
xnor U332 (N_332,In_379,In_878);
nand U333 (N_333,In_205,In_145);
and U334 (N_334,In_284,In_647);
nor U335 (N_335,In_648,In_965);
nor U336 (N_336,In_265,In_3);
and U337 (N_337,In_489,In_943);
or U338 (N_338,In_240,In_772);
nor U339 (N_339,In_736,In_426);
nand U340 (N_340,In_8,In_972);
and U341 (N_341,In_534,In_668);
and U342 (N_342,In_115,In_469);
and U343 (N_343,In_725,In_584);
and U344 (N_344,In_591,In_14);
nor U345 (N_345,In_296,In_359);
or U346 (N_346,In_468,In_461);
and U347 (N_347,In_163,In_50);
and U348 (N_348,In_321,In_322);
or U349 (N_349,In_46,In_393);
nor U350 (N_350,In_465,In_484);
nor U351 (N_351,In_215,In_704);
and U352 (N_352,In_511,In_218);
and U353 (N_353,In_541,In_313);
nor U354 (N_354,In_945,In_621);
and U355 (N_355,In_916,In_769);
nand U356 (N_356,In_74,In_735);
or U357 (N_357,In_302,In_285);
nor U358 (N_358,In_938,In_829);
and U359 (N_359,In_212,In_949);
nand U360 (N_360,In_381,In_86);
and U361 (N_361,In_827,In_420);
and U362 (N_362,In_660,In_620);
nor U363 (N_363,In_200,In_99);
or U364 (N_364,In_869,In_638);
nor U365 (N_365,In_411,In_834);
nor U366 (N_366,In_134,In_136);
nand U367 (N_367,In_550,In_616);
nor U368 (N_368,In_287,In_112);
nand U369 (N_369,In_699,In_118);
nor U370 (N_370,In_697,In_318);
and U371 (N_371,In_473,In_830);
and U372 (N_372,In_343,In_263);
nor U373 (N_373,In_658,In_803);
nor U374 (N_374,In_293,In_977);
xnor U375 (N_375,In_27,In_504);
nor U376 (N_376,In_748,In_444);
nor U377 (N_377,In_271,In_606);
nor U378 (N_378,In_499,In_482);
or U379 (N_379,In_133,In_241);
nor U380 (N_380,In_138,In_887);
and U381 (N_381,In_583,In_220);
or U382 (N_382,In_71,In_404);
nor U383 (N_383,In_236,In_250);
or U384 (N_384,In_765,In_997);
and U385 (N_385,In_336,In_44);
nor U386 (N_386,In_67,In_958);
xor U387 (N_387,In_625,In_21);
nand U388 (N_388,In_693,In_89);
nand U389 (N_389,In_899,In_862);
nand U390 (N_390,In_0,In_35);
or U391 (N_391,In_910,In_821);
and U392 (N_392,In_176,In_926);
nor U393 (N_393,In_510,In_186);
or U394 (N_394,In_325,In_609);
nand U395 (N_395,In_373,In_175);
nor U396 (N_396,In_190,In_479);
nor U397 (N_397,In_109,In_364);
or U398 (N_398,In_83,In_873);
and U399 (N_399,In_513,In_774);
nand U400 (N_400,In_831,In_84);
or U401 (N_401,In_277,In_309);
and U402 (N_402,In_354,In_846);
nand U403 (N_403,In_451,In_805);
nor U404 (N_404,In_179,In_843);
or U405 (N_405,In_217,In_485);
and U406 (N_406,In_383,In_580);
nand U407 (N_407,In_820,In_640);
or U408 (N_408,In_124,In_966);
nor U409 (N_409,In_398,In_563);
xor U410 (N_410,In_356,In_637);
and U411 (N_411,In_690,In_310);
nand U412 (N_412,In_632,In_20);
nand U413 (N_413,In_539,In_344);
xnor U414 (N_414,In_928,In_692);
and U415 (N_415,In_119,In_721);
nor U416 (N_416,In_493,In_808);
xor U417 (N_417,In_512,In_335);
and U418 (N_418,In_340,In_231);
and U419 (N_419,In_789,In_573);
and U420 (N_420,In_978,In_229);
nor U421 (N_421,In_730,In_732);
and U422 (N_422,In_316,In_281);
or U423 (N_423,In_442,In_457);
and U424 (N_424,In_890,In_63);
nand U425 (N_425,In_734,In_412);
nand U426 (N_426,In_593,In_793);
or U427 (N_427,In_233,In_771);
and U428 (N_428,In_799,In_105);
nand U429 (N_429,In_440,In_724);
nor U430 (N_430,In_987,In_196);
or U431 (N_431,In_576,In_66);
nand U432 (N_432,In_741,In_54);
nand U433 (N_433,In_855,In_968);
nor U434 (N_434,In_397,In_327);
nor U435 (N_435,In_355,In_742);
nor U436 (N_436,In_256,In_627);
nand U437 (N_437,In_140,In_376);
nor U438 (N_438,In_65,In_845);
or U439 (N_439,In_258,In_396);
nand U440 (N_440,In_703,In_816);
nor U441 (N_441,In_72,In_983);
nor U442 (N_442,In_169,In_767);
nor U443 (N_443,In_967,In_756);
or U444 (N_444,In_633,In_428);
nor U445 (N_445,In_497,In_57);
nor U446 (N_446,In_448,In_761);
nor U447 (N_447,In_667,In_407);
nand U448 (N_448,In_825,In_353);
nor U449 (N_449,In_990,In_255);
or U450 (N_450,In_102,In_688);
and U451 (N_451,In_323,In_59);
or U452 (N_452,In_718,In_842);
or U453 (N_453,In_506,In_586);
nor U454 (N_454,In_209,In_757);
nor U455 (N_455,In_530,In_574);
nor U456 (N_456,In_656,In_155);
or U457 (N_457,In_438,In_4);
or U458 (N_458,In_657,In_615);
nand U459 (N_459,In_307,In_77);
and U460 (N_460,In_25,In_22);
xnor U461 (N_461,In_446,In_645);
or U462 (N_462,In_32,In_254);
or U463 (N_463,In_197,In_915);
or U464 (N_464,In_876,In_73);
or U465 (N_465,In_981,In_227);
nor U466 (N_466,In_919,In_326);
and U467 (N_467,In_694,In_900);
nor U468 (N_468,In_763,In_740);
nand U469 (N_469,In_833,In_36);
or U470 (N_470,In_879,In_578);
and U471 (N_471,In_16,In_835);
and U472 (N_472,In_604,In_804);
nor U473 (N_473,In_776,In_56);
nor U474 (N_474,In_856,In_188);
xor U475 (N_475,In_596,In_62);
or U476 (N_476,In_262,In_60);
and U477 (N_477,In_728,In_980);
or U478 (N_478,In_45,In_885);
or U479 (N_479,In_652,In_238);
nand U480 (N_480,In_800,In_597);
and U481 (N_481,In_785,In_201);
and U482 (N_482,In_369,In_388);
and U483 (N_483,In_954,In_237);
nor U484 (N_484,In_358,In_773);
nor U485 (N_485,In_920,In_817);
nand U486 (N_486,In_903,In_126);
or U487 (N_487,In_453,In_34);
and U488 (N_488,In_719,In_629);
and U489 (N_489,In_832,In_235);
nor U490 (N_490,In_872,In_403);
nor U491 (N_491,In_362,In_26);
nand U492 (N_492,In_755,In_193);
and U493 (N_493,In_213,In_191);
xor U494 (N_494,In_674,In_884);
xor U495 (N_495,In_814,In_131);
nor U496 (N_496,In_375,In_908);
nand U497 (N_497,In_114,In_575);
nand U498 (N_498,In_290,In_414);
nand U499 (N_499,In_762,In_368);
nand U500 (N_500,In_172,In_22);
nand U501 (N_501,In_587,In_797);
and U502 (N_502,In_151,In_95);
nand U503 (N_503,In_865,In_2);
nand U504 (N_504,In_503,In_582);
or U505 (N_505,In_278,In_615);
and U506 (N_506,In_752,In_426);
and U507 (N_507,In_347,In_854);
nor U508 (N_508,In_205,In_990);
and U509 (N_509,In_706,In_749);
or U510 (N_510,In_803,In_471);
or U511 (N_511,In_760,In_304);
nor U512 (N_512,In_178,In_459);
nand U513 (N_513,In_971,In_90);
and U514 (N_514,In_104,In_405);
or U515 (N_515,In_878,In_121);
or U516 (N_516,In_170,In_400);
and U517 (N_517,In_735,In_310);
nor U518 (N_518,In_694,In_212);
nor U519 (N_519,In_633,In_617);
nand U520 (N_520,In_199,In_978);
nand U521 (N_521,In_588,In_828);
nor U522 (N_522,In_927,In_911);
and U523 (N_523,In_15,In_452);
or U524 (N_524,In_306,In_970);
xnor U525 (N_525,In_4,In_700);
or U526 (N_526,In_151,In_419);
and U527 (N_527,In_357,In_794);
nand U528 (N_528,In_251,In_430);
or U529 (N_529,In_616,In_758);
or U530 (N_530,In_812,In_395);
and U531 (N_531,In_248,In_934);
and U532 (N_532,In_890,In_522);
nand U533 (N_533,In_887,In_110);
nand U534 (N_534,In_892,In_882);
nand U535 (N_535,In_680,In_420);
and U536 (N_536,In_836,In_38);
nand U537 (N_537,In_762,In_264);
or U538 (N_538,In_93,In_184);
nand U539 (N_539,In_274,In_255);
and U540 (N_540,In_939,In_858);
or U541 (N_541,In_934,In_753);
or U542 (N_542,In_311,In_920);
nand U543 (N_543,In_878,In_796);
and U544 (N_544,In_488,In_700);
and U545 (N_545,In_533,In_426);
or U546 (N_546,In_771,In_788);
nor U547 (N_547,In_246,In_140);
and U548 (N_548,In_68,In_945);
nand U549 (N_549,In_237,In_185);
nor U550 (N_550,In_767,In_256);
nand U551 (N_551,In_388,In_655);
xor U552 (N_552,In_483,In_237);
nor U553 (N_553,In_202,In_97);
or U554 (N_554,In_68,In_792);
nand U555 (N_555,In_122,In_958);
nand U556 (N_556,In_636,In_879);
and U557 (N_557,In_595,In_86);
or U558 (N_558,In_269,In_570);
or U559 (N_559,In_881,In_175);
and U560 (N_560,In_257,In_903);
or U561 (N_561,In_377,In_492);
nor U562 (N_562,In_921,In_496);
or U563 (N_563,In_974,In_334);
nor U564 (N_564,In_664,In_372);
nor U565 (N_565,In_34,In_397);
nand U566 (N_566,In_321,In_591);
nand U567 (N_567,In_497,In_567);
nor U568 (N_568,In_392,In_615);
nand U569 (N_569,In_969,In_415);
or U570 (N_570,In_384,In_532);
nor U571 (N_571,In_972,In_260);
nand U572 (N_572,In_188,In_24);
and U573 (N_573,In_700,In_633);
and U574 (N_574,In_874,In_927);
or U575 (N_575,In_939,In_777);
nand U576 (N_576,In_373,In_278);
and U577 (N_577,In_642,In_938);
nand U578 (N_578,In_909,In_377);
nand U579 (N_579,In_166,In_670);
nand U580 (N_580,In_234,In_648);
and U581 (N_581,In_509,In_631);
and U582 (N_582,In_235,In_282);
and U583 (N_583,In_240,In_231);
and U584 (N_584,In_32,In_749);
or U585 (N_585,In_154,In_786);
and U586 (N_586,In_590,In_440);
nand U587 (N_587,In_908,In_373);
nor U588 (N_588,In_702,In_37);
xor U589 (N_589,In_974,In_383);
or U590 (N_590,In_110,In_439);
nor U591 (N_591,In_554,In_701);
and U592 (N_592,In_832,In_312);
nor U593 (N_593,In_247,In_972);
and U594 (N_594,In_6,In_706);
nor U595 (N_595,In_559,In_788);
and U596 (N_596,In_32,In_922);
and U597 (N_597,In_514,In_324);
nand U598 (N_598,In_178,In_731);
nor U599 (N_599,In_11,In_439);
nand U600 (N_600,In_101,In_439);
nand U601 (N_601,In_390,In_505);
and U602 (N_602,In_481,In_59);
and U603 (N_603,In_52,In_717);
nand U604 (N_604,In_613,In_807);
nor U605 (N_605,In_87,In_414);
nor U606 (N_606,In_80,In_991);
or U607 (N_607,In_468,In_973);
and U608 (N_608,In_495,In_915);
and U609 (N_609,In_442,In_408);
nor U610 (N_610,In_812,In_532);
nor U611 (N_611,In_606,In_999);
and U612 (N_612,In_64,In_462);
or U613 (N_613,In_855,In_304);
nor U614 (N_614,In_230,In_362);
or U615 (N_615,In_653,In_69);
nand U616 (N_616,In_719,In_855);
xnor U617 (N_617,In_6,In_844);
or U618 (N_618,In_504,In_657);
and U619 (N_619,In_315,In_470);
nand U620 (N_620,In_530,In_453);
nand U621 (N_621,In_102,In_793);
or U622 (N_622,In_103,In_911);
or U623 (N_623,In_535,In_732);
nand U624 (N_624,In_658,In_334);
and U625 (N_625,In_812,In_874);
or U626 (N_626,In_28,In_127);
or U627 (N_627,In_974,In_992);
and U628 (N_628,In_591,In_99);
or U629 (N_629,In_258,In_826);
and U630 (N_630,In_772,In_663);
and U631 (N_631,In_550,In_685);
nand U632 (N_632,In_35,In_301);
or U633 (N_633,In_767,In_140);
xnor U634 (N_634,In_280,In_987);
or U635 (N_635,In_570,In_207);
nor U636 (N_636,In_112,In_467);
and U637 (N_637,In_798,In_778);
nand U638 (N_638,In_6,In_66);
or U639 (N_639,In_778,In_11);
or U640 (N_640,In_182,In_665);
or U641 (N_641,In_871,In_38);
and U642 (N_642,In_454,In_901);
nand U643 (N_643,In_851,In_453);
xor U644 (N_644,In_818,In_354);
nand U645 (N_645,In_952,In_795);
nor U646 (N_646,In_670,In_694);
nand U647 (N_647,In_608,In_453);
and U648 (N_648,In_724,In_558);
nand U649 (N_649,In_558,In_691);
nor U650 (N_650,In_829,In_199);
and U651 (N_651,In_8,In_821);
or U652 (N_652,In_773,In_64);
nand U653 (N_653,In_746,In_809);
xnor U654 (N_654,In_904,In_26);
and U655 (N_655,In_331,In_194);
and U656 (N_656,In_258,In_370);
and U657 (N_657,In_641,In_727);
nand U658 (N_658,In_320,In_397);
nor U659 (N_659,In_2,In_639);
and U660 (N_660,In_108,In_292);
or U661 (N_661,In_786,In_369);
nand U662 (N_662,In_243,In_358);
nand U663 (N_663,In_950,In_841);
nor U664 (N_664,In_339,In_294);
or U665 (N_665,In_105,In_838);
and U666 (N_666,In_886,In_956);
and U667 (N_667,In_156,In_470);
xor U668 (N_668,In_685,In_455);
nor U669 (N_669,In_376,In_879);
or U670 (N_670,In_293,In_16);
and U671 (N_671,In_91,In_517);
nand U672 (N_672,In_509,In_246);
nand U673 (N_673,In_665,In_341);
xnor U674 (N_674,In_176,In_436);
or U675 (N_675,In_872,In_816);
nand U676 (N_676,In_639,In_315);
and U677 (N_677,In_736,In_540);
or U678 (N_678,In_894,In_330);
nor U679 (N_679,In_99,In_124);
or U680 (N_680,In_192,In_167);
nor U681 (N_681,In_351,In_299);
nor U682 (N_682,In_884,In_29);
or U683 (N_683,In_387,In_704);
nor U684 (N_684,In_586,In_91);
or U685 (N_685,In_120,In_436);
nor U686 (N_686,In_756,In_907);
nand U687 (N_687,In_862,In_452);
and U688 (N_688,In_91,In_873);
and U689 (N_689,In_347,In_161);
nor U690 (N_690,In_12,In_91);
and U691 (N_691,In_467,In_829);
nand U692 (N_692,In_797,In_25);
nand U693 (N_693,In_971,In_435);
nand U694 (N_694,In_407,In_19);
nand U695 (N_695,In_128,In_68);
and U696 (N_696,In_758,In_175);
xnor U697 (N_697,In_210,In_788);
nand U698 (N_698,In_194,In_791);
and U699 (N_699,In_781,In_218);
and U700 (N_700,In_262,In_392);
nand U701 (N_701,In_197,In_358);
xor U702 (N_702,In_847,In_716);
and U703 (N_703,In_14,In_65);
nand U704 (N_704,In_336,In_301);
nand U705 (N_705,In_30,In_73);
or U706 (N_706,In_377,In_791);
or U707 (N_707,In_530,In_746);
and U708 (N_708,In_919,In_974);
nor U709 (N_709,In_409,In_996);
nand U710 (N_710,In_524,In_958);
nor U711 (N_711,In_876,In_421);
or U712 (N_712,In_519,In_136);
nand U713 (N_713,In_490,In_541);
and U714 (N_714,In_521,In_800);
nand U715 (N_715,In_737,In_678);
and U716 (N_716,In_861,In_378);
or U717 (N_717,In_265,In_302);
nor U718 (N_718,In_863,In_278);
nand U719 (N_719,In_691,In_136);
nand U720 (N_720,In_666,In_536);
nor U721 (N_721,In_871,In_538);
or U722 (N_722,In_710,In_346);
or U723 (N_723,In_39,In_866);
nand U724 (N_724,In_999,In_684);
and U725 (N_725,In_138,In_677);
and U726 (N_726,In_569,In_964);
or U727 (N_727,In_798,In_301);
nor U728 (N_728,In_607,In_806);
or U729 (N_729,In_962,In_84);
nor U730 (N_730,In_486,In_638);
nand U731 (N_731,In_730,In_550);
xor U732 (N_732,In_371,In_304);
or U733 (N_733,In_57,In_954);
nor U734 (N_734,In_599,In_473);
nor U735 (N_735,In_629,In_93);
nand U736 (N_736,In_254,In_870);
nand U737 (N_737,In_564,In_577);
or U738 (N_738,In_196,In_986);
and U739 (N_739,In_167,In_204);
and U740 (N_740,In_797,In_871);
nor U741 (N_741,In_188,In_257);
and U742 (N_742,In_838,In_611);
nor U743 (N_743,In_337,In_398);
or U744 (N_744,In_821,In_11);
nand U745 (N_745,In_476,In_315);
nor U746 (N_746,In_188,In_539);
nand U747 (N_747,In_382,In_314);
and U748 (N_748,In_872,In_93);
xor U749 (N_749,In_420,In_24);
nand U750 (N_750,In_158,In_327);
and U751 (N_751,In_708,In_457);
and U752 (N_752,In_409,In_590);
and U753 (N_753,In_697,In_621);
nor U754 (N_754,In_440,In_492);
and U755 (N_755,In_514,In_228);
nor U756 (N_756,In_77,In_346);
nand U757 (N_757,In_982,In_210);
nand U758 (N_758,In_276,In_133);
nand U759 (N_759,In_193,In_664);
nand U760 (N_760,In_749,In_74);
or U761 (N_761,In_939,In_448);
xnor U762 (N_762,In_407,In_160);
or U763 (N_763,In_351,In_993);
nand U764 (N_764,In_979,In_76);
nor U765 (N_765,In_213,In_867);
nand U766 (N_766,In_370,In_937);
nor U767 (N_767,In_901,In_130);
nor U768 (N_768,In_75,In_154);
xnor U769 (N_769,In_561,In_920);
or U770 (N_770,In_163,In_796);
nor U771 (N_771,In_595,In_577);
or U772 (N_772,In_723,In_228);
nand U773 (N_773,In_914,In_384);
nor U774 (N_774,In_447,In_878);
or U775 (N_775,In_931,In_989);
and U776 (N_776,In_461,In_694);
nor U777 (N_777,In_61,In_886);
or U778 (N_778,In_674,In_871);
nand U779 (N_779,In_270,In_509);
nor U780 (N_780,In_461,In_449);
or U781 (N_781,In_605,In_24);
nor U782 (N_782,In_889,In_277);
nor U783 (N_783,In_952,In_417);
xor U784 (N_784,In_334,In_355);
nand U785 (N_785,In_640,In_769);
or U786 (N_786,In_76,In_769);
nor U787 (N_787,In_155,In_57);
or U788 (N_788,In_428,In_527);
and U789 (N_789,In_929,In_396);
nand U790 (N_790,In_500,In_324);
xor U791 (N_791,In_340,In_422);
nand U792 (N_792,In_174,In_199);
or U793 (N_793,In_102,In_38);
and U794 (N_794,In_946,In_594);
nand U795 (N_795,In_978,In_315);
nand U796 (N_796,In_196,In_869);
and U797 (N_797,In_703,In_149);
nand U798 (N_798,In_90,In_977);
nand U799 (N_799,In_771,In_590);
or U800 (N_800,In_336,In_901);
nand U801 (N_801,In_646,In_787);
nor U802 (N_802,In_32,In_769);
and U803 (N_803,In_320,In_596);
xor U804 (N_804,In_288,In_550);
nor U805 (N_805,In_335,In_816);
and U806 (N_806,In_864,In_318);
nand U807 (N_807,In_291,In_861);
nand U808 (N_808,In_150,In_408);
nor U809 (N_809,In_164,In_536);
nor U810 (N_810,In_784,In_536);
or U811 (N_811,In_882,In_14);
and U812 (N_812,In_106,In_988);
nor U813 (N_813,In_471,In_59);
nor U814 (N_814,In_958,In_780);
or U815 (N_815,In_685,In_672);
nor U816 (N_816,In_163,In_966);
or U817 (N_817,In_608,In_468);
and U818 (N_818,In_422,In_844);
or U819 (N_819,In_485,In_338);
nor U820 (N_820,In_209,In_591);
or U821 (N_821,In_452,In_600);
and U822 (N_822,In_930,In_158);
nand U823 (N_823,In_888,In_996);
or U824 (N_824,In_86,In_645);
and U825 (N_825,In_807,In_627);
nand U826 (N_826,In_975,In_689);
or U827 (N_827,In_897,In_951);
and U828 (N_828,In_989,In_635);
and U829 (N_829,In_226,In_374);
and U830 (N_830,In_111,In_981);
nand U831 (N_831,In_682,In_969);
or U832 (N_832,In_587,In_230);
and U833 (N_833,In_389,In_290);
xnor U834 (N_834,In_381,In_254);
or U835 (N_835,In_622,In_281);
nor U836 (N_836,In_899,In_185);
nand U837 (N_837,In_632,In_127);
nand U838 (N_838,In_908,In_369);
nor U839 (N_839,In_202,In_810);
nand U840 (N_840,In_679,In_454);
nand U841 (N_841,In_709,In_924);
and U842 (N_842,In_82,In_269);
and U843 (N_843,In_355,In_33);
nand U844 (N_844,In_635,In_187);
or U845 (N_845,In_132,In_544);
nor U846 (N_846,In_74,In_656);
and U847 (N_847,In_844,In_463);
nor U848 (N_848,In_87,In_53);
nor U849 (N_849,In_824,In_437);
nand U850 (N_850,In_847,In_915);
nor U851 (N_851,In_218,In_346);
nor U852 (N_852,In_621,In_485);
and U853 (N_853,In_139,In_189);
and U854 (N_854,In_664,In_568);
or U855 (N_855,In_279,In_697);
nor U856 (N_856,In_910,In_998);
or U857 (N_857,In_218,In_420);
and U858 (N_858,In_311,In_965);
and U859 (N_859,In_778,In_181);
nand U860 (N_860,In_544,In_654);
nand U861 (N_861,In_817,In_380);
nor U862 (N_862,In_959,In_89);
nand U863 (N_863,In_3,In_79);
nor U864 (N_864,In_473,In_370);
and U865 (N_865,In_663,In_911);
or U866 (N_866,In_815,In_473);
and U867 (N_867,In_837,In_166);
and U868 (N_868,In_3,In_8);
and U869 (N_869,In_921,In_321);
or U870 (N_870,In_609,In_118);
or U871 (N_871,In_47,In_470);
or U872 (N_872,In_477,In_192);
or U873 (N_873,In_60,In_504);
xnor U874 (N_874,In_190,In_791);
nor U875 (N_875,In_782,In_167);
nand U876 (N_876,In_371,In_997);
or U877 (N_877,In_793,In_497);
nand U878 (N_878,In_59,In_922);
nor U879 (N_879,In_595,In_908);
nand U880 (N_880,In_215,In_933);
or U881 (N_881,In_14,In_316);
nand U882 (N_882,In_93,In_559);
or U883 (N_883,In_791,In_429);
nor U884 (N_884,In_424,In_133);
or U885 (N_885,In_918,In_234);
nand U886 (N_886,In_215,In_332);
nor U887 (N_887,In_160,In_451);
nor U888 (N_888,In_702,In_548);
and U889 (N_889,In_266,In_559);
nor U890 (N_890,In_898,In_918);
nor U891 (N_891,In_782,In_96);
nand U892 (N_892,In_514,In_480);
nand U893 (N_893,In_34,In_719);
and U894 (N_894,In_88,In_192);
xor U895 (N_895,In_142,In_463);
nor U896 (N_896,In_11,In_518);
nor U897 (N_897,In_620,In_729);
nor U898 (N_898,In_949,In_642);
or U899 (N_899,In_524,In_673);
and U900 (N_900,In_194,In_766);
and U901 (N_901,In_410,In_832);
and U902 (N_902,In_675,In_533);
nand U903 (N_903,In_773,In_261);
and U904 (N_904,In_876,In_911);
or U905 (N_905,In_473,In_986);
or U906 (N_906,In_761,In_141);
nand U907 (N_907,In_762,In_51);
nand U908 (N_908,In_662,In_870);
nand U909 (N_909,In_139,In_78);
and U910 (N_910,In_205,In_794);
or U911 (N_911,In_213,In_793);
nor U912 (N_912,In_479,In_594);
and U913 (N_913,In_12,In_307);
and U914 (N_914,In_442,In_486);
or U915 (N_915,In_859,In_696);
and U916 (N_916,In_397,In_774);
or U917 (N_917,In_43,In_637);
or U918 (N_918,In_279,In_787);
nand U919 (N_919,In_697,In_476);
nand U920 (N_920,In_498,In_12);
nand U921 (N_921,In_517,In_926);
or U922 (N_922,In_320,In_571);
and U923 (N_923,In_821,In_336);
and U924 (N_924,In_728,In_273);
nor U925 (N_925,In_855,In_956);
and U926 (N_926,In_779,In_196);
xnor U927 (N_927,In_565,In_840);
nor U928 (N_928,In_198,In_97);
and U929 (N_929,In_752,In_112);
nor U930 (N_930,In_744,In_419);
nand U931 (N_931,In_794,In_598);
nand U932 (N_932,In_847,In_586);
or U933 (N_933,In_470,In_449);
or U934 (N_934,In_189,In_826);
nand U935 (N_935,In_615,In_488);
nand U936 (N_936,In_867,In_927);
or U937 (N_937,In_528,In_785);
or U938 (N_938,In_650,In_721);
nor U939 (N_939,In_734,In_828);
xnor U940 (N_940,In_904,In_70);
or U941 (N_941,In_232,In_475);
nand U942 (N_942,In_331,In_339);
nand U943 (N_943,In_285,In_197);
and U944 (N_944,In_225,In_268);
nand U945 (N_945,In_223,In_476);
or U946 (N_946,In_769,In_482);
nand U947 (N_947,In_884,In_59);
and U948 (N_948,In_959,In_768);
or U949 (N_949,In_831,In_524);
nand U950 (N_950,In_287,In_235);
or U951 (N_951,In_824,In_578);
nor U952 (N_952,In_697,In_494);
nand U953 (N_953,In_196,In_160);
and U954 (N_954,In_577,In_919);
and U955 (N_955,In_923,In_171);
nand U956 (N_956,In_151,In_332);
or U957 (N_957,In_372,In_311);
or U958 (N_958,In_115,In_459);
and U959 (N_959,In_551,In_105);
and U960 (N_960,In_832,In_284);
or U961 (N_961,In_735,In_53);
nor U962 (N_962,In_149,In_753);
nor U963 (N_963,In_72,In_919);
and U964 (N_964,In_299,In_748);
nand U965 (N_965,In_337,In_681);
or U966 (N_966,In_493,In_755);
or U967 (N_967,In_855,In_331);
or U968 (N_968,In_543,In_190);
nor U969 (N_969,In_841,In_883);
or U970 (N_970,In_475,In_374);
or U971 (N_971,In_346,In_371);
and U972 (N_972,In_560,In_438);
nand U973 (N_973,In_439,In_988);
xor U974 (N_974,In_675,In_588);
and U975 (N_975,In_762,In_71);
nand U976 (N_976,In_344,In_999);
nand U977 (N_977,In_889,In_408);
or U978 (N_978,In_496,In_292);
or U979 (N_979,In_503,In_686);
and U980 (N_980,In_703,In_182);
and U981 (N_981,In_765,In_273);
and U982 (N_982,In_264,In_121);
nand U983 (N_983,In_743,In_550);
or U984 (N_984,In_8,In_191);
or U985 (N_985,In_541,In_223);
nor U986 (N_986,In_366,In_898);
and U987 (N_987,In_394,In_847);
or U988 (N_988,In_370,In_271);
nor U989 (N_989,In_386,In_460);
nand U990 (N_990,In_468,In_935);
and U991 (N_991,In_620,In_569);
or U992 (N_992,In_540,In_977);
nor U993 (N_993,In_111,In_848);
and U994 (N_994,In_529,In_869);
or U995 (N_995,In_605,In_483);
or U996 (N_996,In_528,In_568);
nor U997 (N_997,In_542,In_960);
and U998 (N_998,In_736,In_134);
nand U999 (N_999,In_163,In_749);
or U1000 (N_1000,In_650,In_354);
nand U1001 (N_1001,In_260,In_490);
and U1002 (N_1002,In_304,In_245);
nand U1003 (N_1003,In_909,In_397);
nand U1004 (N_1004,In_522,In_66);
or U1005 (N_1005,In_541,In_150);
or U1006 (N_1006,In_106,In_155);
nand U1007 (N_1007,In_995,In_869);
nand U1008 (N_1008,In_532,In_466);
nand U1009 (N_1009,In_505,In_446);
nor U1010 (N_1010,In_365,In_988);
nor U1011 (N_1011,In_21,In_385);
and U1012 (N_1012,In_564,In_512);
nor U1013 (N_1013,In_940,In_983);
and U1014 (N_1014,In_234,In_803);
nand U1015 (N_1015,In_512,In_381);
nor U1016 (N_1016,In_812,In_346);
nand U1017 (N_1017,In_507,In_736);
nor U1018 (N_1018,In_422,In_752);
and U1019 (N_1019,In_878,In_474);
and U1020 (N_1020,In_578,In_384);
nand U1021 (N_1021,In_749,In_209);
xor U1022 (N_1022,In_70,In_188);
and U1023 (N_1023,In_660,In_497);
nand U1024 (N_1024,In_939,In_217);
or U1025 (N_1025,In_409,In_668);
nand U1026 (N_1026,In_555,In_376);
nand U1027 (N_1027,In_177,In_739);
and U1028 (N_1028,In_164,In_690);
xnor U1029 (N_1029,In_528,In_35);
nand U1030 (N_1030,In_424,In_510);
nor U1031 (N_1031,In_283,In_931);
nand U1032 (N_1032,In_502,In_402);
and U1033 (N_1033,In_594,In_954);
and U1034 (N_1034,In_574,In_576);
or U1035 (N_1035,In_268,In_214);
nand U1036 (N_1036,In_189,In_819);
nor U1037 (N_1037,In_618,In_304);
nor U1038 (N_1038,In_504,In_656);
nand U1039 (N_1039,In_878,In_876);
and U1040 (N_1040,In_203,In_897);
nor U1041 (N_1041,In_427,In_489);
and U1042 (N_1042,In_505,In_34);
or U1043 (N_1043,In_855,In_148);
or U1044 (N_1044,In_495,In_372);
nand U1045 (N_1045,In_955,In_697);
and U1046 (N_1046,In_237,In_926);
nor U1047 (N_1047,In_478,In_232);
or U1048 (N_1048,In_814,In_433);
nand U1049 (N_1049,In_900,In_990);
and U1050 (N_1050,In_840,In_455);
or U1051 (N_1051,In_1,In_427);
nand U1052 (N_1052,In_917,In_866);
nor U1053 (N_1053,In_997,In_678);
and U1054 (N_1054,In_98,In_676);
and U1055 (N_1055,In_215,In_419);
and U1056 (N_1056,In_940,In_194);
xor U1057 (N_1057,In_445,In_946);
or U1058 (N_1058,In_70,In_123);
nor U1059 (N_1059,In_786,In_941);
or U1060 (N_1060,In_403,In_89);
nand U1061 (N_1061,In_646,In_653);
or U1062 (N_1062,In_758,In_811);
and U1063 (N_1063,In_579,In_267);
and U1064 (N_1064,In_933,In_69);
or U1065 (N_1065,In_497,In_945);
and U1066 (N_1066,In_165,In_906);
and U1067 (N_1067,In_760,In_751);
nor U1068 (N_1068,In_901,In_103);
nor U1069 (N_1069,In_299,In_758);
and U1070 (N_1070,In_553,In_957);
nor U1071 (N_1071,In_407,In_505);
or U1072 (N_1072,In_20,In_378);
nand U1073 (N_1073,In_278,In_551);
or U1074 (N_1074,In_384,In_454);
nor U1075 (N_1075,In_999,In_729);
and U1076 (N_1076,In_421,In_634);
and U1077 (N_1077,In_426,In_826);
or U1078 (N_1078,In_856,In_982);
and U1079 (N_1079,In_852,In_570);
xnor U1080 (N_1080,In_960,In_931);
nand U1081 (N_1081,In_112,In_968);
nand U1082 (N_1082,In_731,In_644);
and U1083 (N_1083,In_601,In_605);
nor U1084 (N_1084,In_81,In_462);
nand U1085 (N_1085,In_584,In_326);
xnor U1086 (N_1086,In_326,In_177);
or U1087 (N_1087,In_791,In_548);
or U1088 (N_1088,In_39,In_782);
and U1089 (N_1089,In_56,In_272);
nand U1090 (N_1090,In_905,In_985);
nand U1091 (N_1091,In_940,In_367);
nand U1092 (N_1092,In_755,In_609);
xnor U1093 (N_1093,In_203,In_528);
or U1094 (N_1094,In_265,In_510);
nor U1095 (N_1095,In_748,In_605);
or U1096 (N_1096,In_829,In_971);
or U1097 (N_1097,In_959,In_885);
nor U1098 (N_1098,In_166,In_219);
or U1099 (N_1099,In_461,In_199);
nand U1100 (N_1100,In_880,In_125);
or U1101 (N_1101,In_966,In_576);
nor U1102 (N_1102,In_294,In_159);
nor U1103 (N_1103,In_542,In_443);
nand U1104 (N_1104,In_83,In_960);
nand U1105 (N_1105,In_376,In_867);
nor U1106 (N_1106,In_419,In_354);
or U1107 (N_1107,In_347,In_339);
and U1108 (N_1108,In_761,In_110);
and U1109 (N_1109,In_796,In_840);
nor U1110 (N_1110,In_844,In_411);
nand U1111 (N_1111,In_389,In_703);
nor U1112 (N_1112,In_293,In_290);
nor U1113 (N_1113,In_320,In_222);
xor U1114 (N_1114,In_385,In_805);
nor U1115 (N_1115,In_145,In_494);
and U1116 (N_1116,In_962,In_994);
nand U1117 (N_1117,In_251,In_526);
or U1118 (N_1118,In_216,In_341);
nand U1119 (N_1119,In_474,In_312);
and U1120 (N_1120,In_2,In_395);
nor U1121 (N_1121,In_970,In_952);
nand U1122 (N_1122,In_204,In_704);
nor U1123 (N_1123,In_830,In_901);
and U1124 (N_1124,In_813,In_309);
and U1125 (N_1125,In_761,In_306);
or U1126 (N_1126,In_370,In_376);
nor U1127 (N_1127,In_772,In_717);
nor U1128 (N_1128,In_507,In_166);
nor U1129 (N_1129,In_720,In_112);
or U1130 (N_1130,In_335,In_78);
and U1131 (N_1131,In_198,In_457);
nor U1132 (N_1132,In_942,In_323);
nor U1133 (N_1133,In_979,In_962);
nor U1134 (N_1134,In_433,In_108);
and U1135 (N_1135,In_637,In_698);
and U1136 (N_1136,In_417,In_676);
and U1137 (N_1137,In_70,In_680);
nor U1138 (N_1138,In_53,In_616);
or U1139 (N_1139,In_693,In_80);
nor U1140 (N_1140,In_151,In_56);
or U1141 (N_1141,In_500,In_699);
or U1142 (N_1142,In_676,In_230);
or U1143 (N_1143,In_802,In_517);
and U1144 (N_1144,In_155,In_888);
or U1145 (N_1145,In_365,In_649);
or U1146 (N_1146,In_333,In_123);
xnor U1147 (N_1147,In_935,In_22);
nand U1148 (N_1148,In_553,In_789);
nor U1149 (N_1149,In_333,In_744);
or U1150 (N_1150,In_567,In_88);
or U1151 (N_1151,In_653,In_332);
and U1152 (N_1152,In_664,In_897);
and U1153 (N_1153,In_35,In_549);
and U1154 (N_1154,In_486,In_419);
and U1155 (N_1155,In_819,In_233);
nand U1156 (N_1156,In_653,In_399);
nor U1157 (N_1157,In_142,In_284);
nand U1158 (N_1158,In_729,In_91);
and U1159 (N_1159,In_782,In_689);
or U1160 (N_1160,In_85,In_859);
and U1161 (N_1161,In_553,In_400);
nor U1162 (N_1162,In_192,In_165);
nand U1163 (N_1163,In_164,In_727);
or U1164 (N_1164,In_598,In_730);
and U1165 (N_1165,In_481,In_482);
nor U1166 (N_1166,In_853,In_186);
nor U1167 (N_1167,In_998,In_674);
or U1168 (N_1168,In_296,In_319);
nand U1169 (N_1169,In_401,In_367);
nand U1170 (N_1170,In_274,In_941);
or U1171 (N_1171,In_535,In_240);
and U1172 (N_1172,In_693,In_42);
nor U1173 (N_1173,In_258,In_591);
nand U1174 (N_1174,In_344,In_488);
nor U1175 (N_1175,In_264,In_905);
nand U1176 (N_1176,In_736,In_382);
nor U1177 (N_1177,In_594,In_374);
or U1178 (N_1178,In_388,In_630);
nor U1179 (N_1179,In_3,In_840);
or U1180 (N_1180,In_574,In_429);
nand U1181 (N_1181,In_360,In_15);
and U1182 (N_1182,In_263,In_9);
or U1183 (N_1183,In_576,In_775);
nand U1184 (N_1184,In_579,In_182);
nand U1185 (N_1185,In_412,In_491);
and U1186 (N_1186,In_490,In_126);
nand U1187 (N_1187,In_294,In_962);
nor U1188 (N_1188,In_373,In_929);
xnor U1189 (N_1189,In_967,In_119);
or U1190 (N_1190,In_965,In_149);
nand U1191 (N_1191,In_112,In_141);
nor U1192 (N_1192,In_111,In_817);
or U1193 (N_1193,In_478,In_187);
or U1194 (N_1194,In_236,In_347);
xnor U1195 (N_1195,In_483,In_944);
nand U1196 (N_1196,In_985,In_125);
xor U1197 (N_1197,In_956,In_613);
nor U1198 (N_1198,In_435,In_529);
or U1199 (N_1199,In_198,In_810);
nand U1200 (N_1200,In_688,In_340);
or U1201 (N_1201,In_767,In_676);
nor U1202 (N_1202,In_741,In_349);
or U1203 (N_1203,In_779,In_115);
or U1204 (N_1204,In_487,In_457);
nor U1205 (N_1205,In_132,In_93);
and U1206 (N_1206,In_860,In_469);
and U1207 (N_1207,In_382,In_773);
nor U1208 (N_1208,In_388,In_789);
nand U1209 (N_1209,In_678,In_457);
nand U1210 (N_1210,In_85,In_305);
and U1211 (N_1211,In_211,In_334);
or U1212 (N_1212,In_139,In_590);
nor U1213 (N_1213,In_54,In_825);
and U1214 (N_1214,In_970,In_884);
or U1215 (N_1215,In_223,In_419);
and U1216 (N_1216,In_192,In_673);
nor U1217 (N_1217,In_836,In_668);
and U1218 (N_1218,In_106,In_570);
nor U1219 (N_1219,In_361,In_453);
and U1220 (N_1220,In_543,In_125);
xnor U1221 (N_1221,In_185,In_117);
and U1222 (N_1222,In_79,In_548);
nand U1223 (N_1223,In_199,In_130);
and U1224 (N_1224,In_192,In_122);
nand U1225 (N_1225,In_570,In_849);
nor U1226 (N_1226,In_588,In_383);
or U1227 (N_1227,In_823,In_921);
xnor U1228 (N_1228,In_410,In_948);
or U1229 (N_1229,In_741,In_573);
nand U1230 (N_1230,In_52,In_715);
and U1231 (N_1231,In_561,In_787);
or U1232 (N_1232,In_499,In_302);
and U1233 (N_1233,In_475,In_987);
or U1234 (N_1234,In_219,In_254);
xnor U1235 (N_1235,In_98,In_264);
xnor U1236 (N_1236,In_804,In_224);
nand U1237 (N_1237,In_602,In_293);
or U1238 (N_1238,In_197,In_736);
or U1239 (N_1239,In_181,In_617);
nor U1240 (N_1240,In_428,In_530);
nand U1241 (N_1241,In_956,In_885);
nand U1242 (N_1242,In_376,In_410);
nor U1243 (N_1243,In_586,In_465);
nand U1244 (N_1244,In_73,In_560);
nand U1245 (N_1245,In_752,In_596);
nand U1246 (N_1246,In_338,In_601);
or U1247 (N_1247,In_626,In_209);
xnor U1248 (N_1248,In_279,In_733);
and U1249 (N_1249,In_387,In_590);
nor U1250 (N_1250,In_4,In_94);
and U1251 (N_1251,In_446,In_140);
or U1252 (N_1252,In_146,In_901);
nor U1253 (N_1253,In_224,In_531);
or U1254 (N_1254,In_424,In_811);
or U1255 (N_1255,In_301,In_335);
and U1256 (N_1256,In_515,In_932);
or U1257 (N_1257,In_321,In_357);
nor U1258 (N_1258,In_85,In_475);
and U1259 (N_1259,In_75,In_998);
nand U1260 (N_1260,In_656,In_563);
nor U1261 (N_1261,In_477,In_668);
nand U1262 (N_1262,In_626,In_462);
or U1263 (N_1263,In_102,In_417);
or U1264 (N_1264,In_926,In_436);
and U1265 (N_1265,In_446,In_349);
nor U1266 (N_1266,In_484,In_781);
nand U1267 (N_1267,In_26,In_612);
or U1268 (N_1268,In_9,In_654);
nand U1269 (N_1269,In_987,In_724);
nand U1270 (N_1270,In_378,In_427);
nand U1271 (N_1271,In_76,In_21);
xnor U1272 (N_1272,In_272,In_168);
or U1273 (N_1273,In_955,In_522);
and U1274 (N_1274,In_405,In_743);
nand U1275 (N_1275,In_11,In_867);
and U1276 (N_1276,In_239,In_486);
and U1277 (N_1277,In_538,In_157);
nand U1278 (N_1278,In_121,In_475);
and U1279 (N_1279,In_487,In_573);
nor U1280 (N_1280,In_425,In_3);
and U1281 (N_1281,In_175,In_809);
nor U1282 (N_1282,In_423,In_608);
and U1283 (N_1283,In_719,In_170);
nor U1284 (N_1284,In_29,In_438);
nand U1285 (N_1285,In_879,In_813);
or U1286 (N_1286,In_353,In_328);
and U1287 (N_1287,In_396,In_794);
and U1288 (N_1288,In_906,In_507);
xnor U1289 (N_1289,In_770,In_119);
nor U1290 (N_1290,In_897,In_654);
and U1291 (N_1291,In_443,In_52);
or U1292 (N_1292,In_727,In_318);
nand U1293 (N_1293,In_273,In_487);
or U1294 (N_1294,In_366,In_100);
and U1295 (N_1295,In_419,In_450);
and U1296 (N_1296,In_687,In_224);
or U1297 (N_1297,In_935,In_883);
nand U1298 (N_1298,In_525,In_172);
nand U1299 (N_1299,In_362,In_176);
nor U1300 (N_1300,In_13,In_870);
nand U1301 (N_1301,In_627,In_100);
and U1302 (N_1302,In_299,In_934);
nand U1303 (N_1303,In_533,In_247);
or U1304 (N_1304,In_212,In_549);
or U1305 (N_1305,In_743,In_107);
nor U1306 (N_1306,In_463,In_266);
and U1307 (N_1307,In_478,In_359);
nand U1308 (N_1308,In_798,In_38);
nand U1309 (N_1309,In_20,In_589);
or U1310 (N_1310,In_201,In_1);
or U1311 (N_1311,In_902,In_310);
and U1312 (N_1312,In_830,In_305);
and U1313 (N_1313,In_843,In_336);
nor U1314 (N_1314,In_748,In_848);
nor U1315 (N_1315,In_925,In_518);
and U1316 (N_1316,In_147,In_949);
nand U1317 (N_1317,In_261,In_806);
or U1318 (N_1318,In_404,In_715);
nor U1319 (N_1319,In_296,In_736);
and U1320 (N_1320,In_303,In_441);
or U1321 (N_1321,In_468,In_678);
nor U1322 (N_1322,In_65,In_582);
nand U1323 (N_1323,In_809,In_484);
nor U1324 (N_1324,In_733,In_574);
nand U1325 (N_1325,In_226,In_559);
nor U1326 (N_1326,In_592,In_570);
nand U1327 (N_1327,In_313,In_738);
or U1328 (N_1328,In_609,In_451);
or U1329 (N_1329,In_814,In_693);
and U1330 (N_1330,In_795,In_818);
nor U1331 (N_1331,In_650,In_547);
nand U1332 (N_1332,In_487,In_14);
nand U1333 (N_1333,In_826,In_450);
nand U1334 (N_1334,In_905,In_956);
or U1335 (N_1335,In_757,In_542);
nand U1336 (N_1336,In_610,In_294);
xor U1337 (N_1337,In_130,In_81);
nor U1338 (N_1338,In_349,In_196);
nand U1339 (N_1339,In_900,In_889);
and U1340 (N_1340,In_450,In_882);
nand U1341 (N_1341,In_41,In_758);
and U1342 (N_1342,In_320,In_939);
nand U1343 (N_1343,In_981,In_302);
and U1344 (N_1344,In_186,In_802);
and U1345 (N_1345,In_66,In_152);
nand U1346 (N_1346,In_425,In_173);
or U1347 (N_1347,In_338,In_913);
or U1348 (N_1348,In_822,In_957);
and U1349 (N_1349,In_316,In_415);
or U1350 (N_1350,In_61,In_913);
nand U1351 (N_1351,In_157,In_84);
nor U1352 (N_1352,In_601,In_720);
and U1353 (N_1353,In_887,In_186);
or U1354 (N_1354,In_773,In_628);
or U1355 (N_1355,In_904,In_239);
nand U1356 (N_1356,In_861,In_329);
nor U1357 (N_1357,In_715,In_539);
and U1358 (N_1358,In_322,In_362);
nand U1359 (N_1359,In_514,In_717);
nor U1360 (N_1360,In_226,In_305);
and U1361 (N_1361,In_68,In_133);
or U1362 (N_1362,In_453,In_863);
nand U1363 (N_1363,In_375,In_10);
or U1364 (N_1364,In_470,In_404);
nand U1365 (N_1365,In_765,In_333);
nor U1366 (N_1366,In_644,In_234);
and U1367 (N_1367,In_274,In_297);
nand U1368 (N_1368,In_35,In_442);
nand U1369 (N_1369,In_134,In_390);
nor U1370 (N_1370,In_176,In_19);
nor U1371 (N_1371,In_791,In_683);
nor U1372 (N_1372,In_707,In_69);
or U1373 (N_1373,In_335,In_255);
nand U1374 (N_1374,In_633,In_283);
or U1375 (N_1375,In_412,In_106);
or U1376 (N_1376,In_266,In_664);
and U1377 (N_1377,In_768,In_741);
and U1378 (N_1378,In_68,In_930);
nor U1379 (N_1379,In_530,In_84);
nor U1380 (N_1380,In_797,In_175);
nand U1381 (N_1381,In_638,In_393);
or U1382 (N_1382,In_950,In_544);
and U1383 (N_1383,In_584,In_424);
or U1384 (N_1384,In_159,In_201);
nand U1385 (N_1385,In_593,In_266);
nor U1386 (N_1386,In_972,In_707);
nor U1387 (N_1387,In_101,In_172);
nand U1388 (N_1388,In_599,In_686);
and U1389 (N_1389,In_947,In_102);
and U1390 (N_1390,In_533,In_727);
nor U1391 (N_1391,In_364,In_998);
nand U1392 (N_1392,In_310,In_37);
xor U1393 (N_1393,In_441,In_268);
nor U1394 (N_1394,In_130,In_6);
nor U1395 (N_1395,In_184,In_213);
nor U1396 (N_1396,In_377,In_415);
or U1397 (N_1397,In_222,In_812);
nand U1398 (N_1398,In_456,In_529);
and U1399 (N_1399,In_746,In_17);
and U1400 (N_1400,In_706,In_967);
nand U1401 (N_1401,In_42,In_674);
nor U1402 (N_1402,In_420,In_111);
and U1403 (N_1403,In_456,In_290);
xor U1404 (N_1404,In_840,In_564);
or U1405 (N_1405,In_144,In_407);
or U1406 (N_1406,In_530,In_215);
and U1407 (N_1407,In_963,In_76);
or U1408 (N_1408,In_128,In_663);
xnor U1409 (N_1409,In_94,In_585);
nand U1410 (N_1410,In_345,In_489);
or U1411 (N_1411,In_610,In_50);
nor U1412 (N_1412,In_113,In_808);
nand U1413 (N_1413,In_721,In_402);
or U1414 (N_1414,In_325,In_88);
nand U1415 (N_1415,In_88,In_857);
and U1416 (N_1416,In_147,In_211);
nand U1417 (N_1417,In_875,In_891);
nand U1418 (N_1418,In_929,In_453);
nand U1419 (N_1419,In_500,In_364);
and U1420 (N_1420,In_140,In_812);
nand U1421 (N_1421,In_654,In_431);
or U1422 (N_1422,In_758,In_858);
nor U1423 (N_1423,In_379,In_765);
nor U1424 (N_1424,In_229,In_94);
nand U1425 (N_1425,In_758,In_820);
nand U1426 (N_1426,In_154,In_337);
and U1427 (N_1427,In_416,In_977);
or U1428 (N_1428,In_925,In_900);
and U1429 (N_1429,In_312,In_519);
nor U1430 (N_1430,In_575,In_554);
nor U1431 (N_1431,In_448,In_717);
nor U1432 (N_1432,In_192,In_820);
and U1433 (N_1433,In_820,In_694);
nand U1434 (N_1434,In_625,In_629);
and U1435 (N_1435,In_62,In_844);
and U1436 (N_1436,In_852,In_779);
or U1437 (N_1437,In_83,In_603);
nand U1438 (N_1438,In_178,In_634);
nand U1439 (N_1439,In_117,In_519);
or U1440 (N_1440,In_957,In_992);
nand U1441 (N_1441,In_721,In_220);
nand U1442 (N_1442,In_907,In_352);
nor U1443 (N_1443,In_960,In_811);
and U1444 (N_1444,In_2,In_765);
nand U1445 (N_1445,In_943,In_4);
xor U1446 (N_1446,In_459,In_210);
or U1447 (N_1447,In_106,In_28);
and U1448 (N_1448,In_818,In_513);
and U1449 (N_1449,In_231,In_964);
nor U1450 (N_1450,In_806,In_680);
nor U1451 (N_1451,In_996,In_620);
and U1452 (N_1452,In_315,In_843);
and U1453 (N_1453,In_971,In_330);
nand U1454 (N_1454,In_646,In_232);
nor U1455 (N_1455,In_852,In_666);
or U1456 (N_1456,In_484,In_568);
nand U1457 (N_1457,In_160,In_718);
nand U1458 (N_1458,In_480,In_451);
nor U1459 (N_1459,In_572,In_233);
nand U1460 (N_1460,In_486,In_785);
nand U1461 (N_1461,In_665,In_442);
nor U1462 (N_1462,In_626,In_84);
nand U1463 (N_1463,In_76,In_58);
nor U1464 (N_1464,In_599,In_718);
and U1465 (N_1465,In_695,In_879);
nor U1466 (N_1466,In_252,In_257);
nor U1467 (N_1467,In_375,In_285);
and U1468 (N_1468,In_513,In_424);
or U1469 (N_1469,In_482,In_507);
nor U1470 (N_1470,In_351,In_414);
or U1471 (N_1471,In_205,In_4);
nand U1472 (N_1472,In_862,In_101);
nor U1473 (N_1473,In_837,In_479);
and U1474 (N_1474,In_375,In_538);
nor U1475 (N_1475,In_549,In_727);
or U1476 (N_1476,In_117,In_104);
xnor U1477 (N_1477,In_823,In_561);
and U1478 (N_1478,In_830,In_135);
or U1479 (N_1479,In_831,In_345);
nor U1480 (N_1480,In_316,In_723);
and U1481 (N_1481,In_720,In_848);
and U1482 (N_1482,In_595,In_246);
nand U1483 (N_1483,In_491,In_456);
or U1484 (N_1484,In_451,In_370);
or U1485 (N_1485,In_496,In_728);
and U1486 (N_1486,In_933,In_975);
and U1487 (N_1487,In_271,In_422);
and U1488 (N_1488,In_932,In_912);
nor U1489 (N_1489,In_494,In_759);
and U1490 (N_1490,In_225,In_708);
or U1491 (N_1491,In_19,In_322);
nor U1492 (N_1492,In_433,In_279);
and U1493 (N_1493,In_413,In_193);
xor U1494 (N_1494,In_858,In_452);
nand U1495 (N_1495,In_955,In_407);
and U1496 (N_1496,In_994,In_194);
and U1497 (N_1497,In_522,In_831);
and U1498 (N_1498,In_841,In_619);
nand U1499 (N_1499,In_636,In_813);
nor U1500 (N_1500,In_681,In_589);
nor U1501 (N_1501,In_328,In_37);
nand U1502 (N_1502,In_230,In_423);
and U1503 (N_1503,In_456,In_682);
or U1504 (N_1504,In_716,In_393);
and U1505 (N_1505,In_465,In_601);
or U1506 (N_1506,In_837,In_817);
nand U1507 (N_1507,In_714,In_899);
or U1508 (N_1508,In_571,In_890);
and U1509 (N_1509,In_790,In_20);
nor U1510 (N_1510,In_513,In_872);
and U1511 (N_1511,In_810,In_11);
and U1512 (N_1512,In_305,In_516);
nor U1513 (N_1513,In_936,In_979);
or U1514 (N_1514,In_895,In_818);
and U1515 (N_1515,In_20,In_920);
and U1516 (N_1516,In_271,In_369);
and U1517 (N_1517,In_214,In_553);
nor U1518 (N_1518,In_529,In_520);
nand U1519 (N_1519,In_544,In_73);
and U1520 (N_1520,In_511,In_521);
nor U1521 (N_1521,In_964,In_76);
and U1522 (N_1522,In_508,In_63);
or U1523 (N_1523,In_74,In_572);
nand U1524 (N_1524,In_909,In_21);
nand U1525 (N_1525,In_883,In_107);
nor U1526 (N_1526,In_295,In_896);
or U1527 (N_1527,In_110,In_724);
or U1528 (N_1528,In_291,In_442);
nand U1529 (N_1529,In_995,In_727);
nand U1530 (N_1530,In_841,In_629);
nor U1531 (N_1531,In_608,In_614);
or U1532 (N_1532,In_875,In_772);
and U1533 (N_1533,In_481,In_290);
nand U1534 (N_1534,In_1,In_591);
or U1535 (N_1535,In_91,In_887);
nor U1536 (N_1536,In_35,In_582);
or U1537 (N_1537,In_759,In_595);
and U1538 (N_1538,In_928,In_654);
or U1539 (N_1539,In_241,In_138);
nand U1540 (N_1540,In_13,In_347);
nand U1541 (N_1541,In_360,In_687);
and U1542 (N_1542,In_509,In_230);
and U1543 (N_1543,In_540,In_898);
nand U1544 (N_1544,In_744,In_541);
nand U1545 (N_1545,In_378,In_341);
nor U1546 (N_1546,In_453,In_849);
or U1547 (N_1547,In_880,In_579);
xor U1548 (N_1548,In_995,In_268);
nand U1549 (N_1549,In_424,In_772);
or U1550 (N_1550,In_740,In_768);
and U1551 (N_1551,In_347,In_393);
nor U1552 (N_1552,In_163,In_461);
nor U1553 (N_1553,In_488,In_480);
and U1554 (N_1554,In_52,In_356);
or U1555 (N_1555,In_241,In_616);
nor U1556 (N_1556,In_830,In_872);
nand U1557 (N_1557,In_113,In_199);
nor U1558 (N_1558,In_205,In_98);
and U1559 (N_1559,In_557,In_488);
or U1560 (N_1560,In_893,In_784);
nand U1561 (N_1561,In_883,In_172);
nand U1562 (N_1562,In_453,In_772);
and U1563 (N_1563,In_188,In_25);
or U1564 (N_1564,In_549,In_717);
nand U1565 (N_1565,In_895,In_769);
nor U1566 (N_1566,In_7,In_154);
nand U1567 (N_1567,In_459,In_176);
nand U1568 (N_1568,In_946,In_238);
nand U1569 (N_1569,In_537,In_393);
or U1570 (N_1570,In_755,In_401);
and U1571 (N_1571,In_159,In_760);
nand U1572 (N_1572,In_835,In_672);
nor U1573 (N_1573,In_438,In_881);
or U1574 (N_1574,In_813,In_371);
xnor U1575 (N_1575,In_291,In_492);
or U1576 (N_1576,In_416,In_928);
nand U1577 (N_1577,In_77,In_830);
and U1578 (N_1578,In_582,In_609);
or U1579 (N_1579,In_665,In_632);
nand U1580 (N_1580,In_997,In_497);
xnor U1581 (N_1581,In_613,In_949);
nor U1582 (N_1582,In_301,In_707);
nor U1583 (N_1583,In_59,In_159);
nand U1584 (N_1584,In_85,In_409);
or U1585 (N_1585,In_177,In_646);
or U1586 (N_1586,In_203,In_933);
or U1587 (N_1587,In_908,In_554);
nand U1588 (N_1588,In_746,In_218);
nand U1589 (N_1589,In_857,In_668);
nor U1590 (N_1590,In_841,In_193);
nand U1591 (N_1591,In_42,In_321);
nor U1592 (N_1592,In_476,In_287);
nand U1593 (N_1593,In_481,In_690);
nor U1594 (N_1594,In_229,In_221);
nor U1595 (N_1595,In_196,In_742);
nor U1596 (N_1596,In_929,In_491);
or U1597 (N_1597,In_252,In_108);
nor U1598 (N_1598,In_581,In_508);
or U1599 (N_1599,In_11,In_632);
xnor U1600 (N_1600,In_360,In_785);
and U1601 (N_1601,In_730,In_716);
nor U1602 (N_1602,In_878,In_987);
and U1603 (N_1603,In_223,In_726);
or U1604 (N_1604,In_266,In_951);
nand U1605 (N_1605,In_824,In_935);
or U1606 (N_1606,In_838,In_22);
or U1607 (N_1607,In_621,In_801);
or U1608 (N_1608,In_328,In_754);
nand U1609 (N_1609,In_461,In_861);
nand U1610 (N_1610,In_4,In_911);
nand U1611 (N_1611,In_274,In_11);
or U1612 (N_1612,In_374,In_350);
nand U1613 (N_1613,In_324,In_354);
and U1614 (N_1614,In_480,In_269);
nand U1615 (N_1615,In_477,In_568);
nor U1616 (N_1616,In_345,In_247);
or U1617 (N_1617,In_438,In_162);
xnor U1618 (N_1618,In_534,In_826);
nand U1619 (N_1619,In_99,In_68);
nand U1620 (N_1620,In_373,In_564);
nor U1621 (N_1621,In_452,In_948);
or U1622 (N_1622,In_793,In_877);
nor U1623 (N_1623,In_725,In_844);
or U1624 (N_1624,In_303,In_68);
nor U1625 (N_1625,In_911,In_416);
and U1626 (N_1626,In_303,In_536);
or U1627 (N_1627,In_101,In_134);
nor U1628 (N_1628,In_75,In_651);
and U1629 (N_1629,In_755,In_866);
nor U1630 (N_1630,In_596,In_890);
or U1631 (N_1631,In_588,In_195);
or U1632 (N_1632,In_482,In_307);
and U1633 (N_1633,In_941,In_568);
nand U1634 (N_1634,In_373,In_279);
and U1635 (N_1635,In_54,In_736);
and U1636 (N_1636,In_900,In_863);
or U1637 (N_1637,In_72,In_943);
nor U1638 (N_1638,In_545,In_797);
nor U1639 (N_1639,In_515,In_626);
or U1640 (N_1640,In_64,In_329);
nand U1641 (N_1641,In_328,In_272);
nand U1642 (N_1642,In_888,In_80);
or U1643 (N_1643,In_505,In_462);
or U1644 (N_1644,In_464,In_444);
nor U1645 (N_1645,In_286,In_197);
or U1646 (N_1646,In_757,In_95);
or U1647 (N_1647,In_49,In_827);
and U1648 (N_1648,In_81,In_471);
or U1649 (N_1649,In_995,In_871);
and U1650 (N_1650,In_944,In_465);
and U1651 (N_1651,In_250,In_602);
or U1652 (N_1652,In_919,In_620);
and U1653 (N_1653,In_665,In_637);
nand U1654 (N_1654,In_373,In_800);
and U1655 (N_1655,In_820,In_560);
or U1656 (N_1656,In_70,In_65);
nand U1657 (N_1657,In_276,In_355);
nand U1658 (N_1658,In_943,In_467);
or U1659 (N_1659,In_821,In_563);
or U1660 (N_1660,In_579,In_655);
nor U1661 (N_1661,In_435,In_488);
and U1662 (N_1662,In_109,In_926);
nand U1663 (N_1663,In_356,In_998);
nor U1664 (N_1664,In_700,In_602);
nand U1665 (N_1665,In_199,In_983);
and U1666 (N_1666,In_529,In_467);
and U1667 (N_1667,In_319,In_267);
nand U1668 (N_1668,In_420,In_513);
or U1669 (N_1669,In_739,In_238);
and U1670 (N_1670,In_790,In_311);
or U1671 (N_1671,In_169,In_397);
and U1672 (N_1672,In_613,In_934);
nor U1673 (N_1673,In_931,In_620);
and U1674 (N_1674,In_423,In_139);
nor U1675 (N_1675,In_147,In_383);
nand U1676 (N_1676,In_955,In_894);
or U1677 (N_1677,In_50,In_574);
nand U1678 (N_1678,In_164,In_596);
and U1679 (N_1679,In_931,In_16);
nand U1680 (N_1680,In_870,In_921);
nand U1681 (N_1681,In_621,In_580);
and U1682 (N_1682,In_567,In_592);
nor U1683 (N_1683,In_716,In_949);
nand U1684 (N_1684,In_627,In_752);
nor U1685 (N_1685,In_20,In_435);
nand U1686 (N_1686,In_844,In_923);
or U1687 (N_1687,In_577,In_162);
or U1688 (N_1688,In_69,In_943);
nand U1689 (N_1689,In_462,In_688);
or U1690 (N_1690,In_223,In_347);
nand U1691 (N_1691,In_695,In_201);
nand U1692 (N_1692,In_89,In_619);
and U1693 (N_1693,In_185,In_875);
nand U1694 (N_1694,In_605,In_50);
nor U1695 (N_1695,In_198,In_473);
or U1696 (N_1696,In_109,In_860);
xor U1697 (N_1697,In_279,In_923);
or U1698 (N_1698,In_432,In_847);
and U1699 (N_1699,In_863,In_484);
and U1700 (N_1700,In_100,In_575);
nand U1701 (N_1701,In_446,In_289);
or U1702 (N_1702,In_192,In_732);
or U1703 (N_1703,In_473,In_706);
nand U1704 (N_1704,In_580,In_612);
nand U1705 (N_1705,In_959,In_874);
nand U1706 (N_1706,In_943,In_657);
or U1707 (N_1707,In_671,In_606);
or U1708 (N_1708,In_260,In_498);
and U1709 (N_1709,In_818,In_754);
and U1710 (N_1710,In_608,In_890);
and U1711 (N_1711,In_792,In_604);
nand U1712 (N_1712,In_934,In_562);
nand U1713 (N_1713,In_245,In_343);
or U1714 (N_1714,In_187,In_775);
nor U1715 (N_1715,In_862,In_688);
nand U1716 (N_1716,In_761,In_218);
nor U1717 (N_1717,In_967,In_770);
or U1718 (N_1718,In_812,In_300);
nor U1719 (N_1719,In_159,In_728);
or U1720 (N_1720,In_601,In_182);
and U1721 (N_1721,In_510,In_750);
and U1722 (N_1722,In_619,In_36);
and U1723 (N_1723,In_840,In_746);
and U1724 (N_1724,In_23,In_595);
and U1725 (N_1725,In_857,In_884);
and U1726 (N_1726,In_998,In_549);
and U1727 (N_1727,In_856,In_917);
nand U1728 (N_1728,In_324,In_518);
and U1729 (N_1729,In_268,In_607);
nor U1730 (N_1730,In_543,In_81);
and U1731 (N_1731,In_382,In_984);
nor U1732 (N_1732,In_336,In_400);
and U1733 (N_1733,In_795,In_74);
or U1734 (N_1734,In_84,In_615);
and U1735 (N_1735,In_951,In_622);
or U1736 (N_1736,In_259,In_675);
xnor U1737 (N_1737,In_321,In_7);
nand U1738 (N_1738,In_93,In_527);
and U1739 (N_1739,In_636,In_313);
nand U1740 (N_1740,In_874,In_616);
nor U1741 (N_1741,In_629,In_592);
nor U1742 (N_1742,In_962,In_511);
nor U1743 (N_1743,In_163,In_113);
or U1744 (N_1744,In_887,In_936);
nor U1745 (N_1745,In_74,In_622);
nor U1746 (N_1746,In_561,In_641);
nor U1747 (N_1747,In_308,In_783);
nor U1748 (N_1748,In_438,In_621);
and U1749 (N_1749,In_258,In_111);
and U1750 (N_1750,In_472,In_673);
nor U1751 (N_1751,In_966,In_391);
or U1752 (N_1752,In_12,In_854);
nand U1753 (N_1753,In_846,In_982);
and U1754 (N_1754,In_254,In_138);
nand U1755 (N_1755,In_698,In_691);
and U1756 (N_1756,In_38,In_259);
or U1757 (N_1757,In_136,In_401);
and U1758 (N_1758,In_440,In_932);
nand U1759 (N_1759,In_213,In_754);
nand U1760 (N_1760,In_243,In_373);
nand U1761 (N_1761,In_735,In_470);
or U1762 (N_1762,In_627,In_554);
nor U1763 (N_1763,In_130,In_783);
and U1764 (N_1764,In_205,In_39);
nand U1765 (N_1765,In_970,In_42);
and U1766 (N_1766,In_519,In_642);
nor U1767 (N_1767,In_71,In_438);
or U1768 (N_1768,In_164,In_756);
or U1769 (N_1769,In_809,In_102);
or U1770 (N_1770,In_20,In_80);
nand U1771 (N_1771,In_675,In_253);
and U1772 (N_1772,In_821,In_732);
nor U1773 (N_1773,In_953,In_628);
nor U1774 (N_1774,In_78,In_30);
or U1775 (N_1775,In_908,In_191);
and U1776 (N_1776,In_981,In_781);
or U1777 (N_1777,In_127,In_222);
or U1778 (N_1778,In_198,In_254);
xor U1779 (N_1779,In_689,In_30);
nor U1780 (N_1780,In_901,In_928);
nor U1781 (N_1781,In_262,In_876);
nand U1782 (N_1782,In_764,In_994);
or U1783 (N_1783,In_42,In_505);
nor U1784 (N_1784,In_142,In_968);
nor U1785 (N_1785,In_908,In_575);
xor U1786 (N_1786,In_294,In_842);
and U1787 (N_1787,In_552,In_470);
nand U1788 (N_1788,In_322,In_677);
or U1789 (N_1789,In_677,In_5);
nand U1790 (N_1790,In_680,In_848);
and U1791 (N_1791,In_904,In_928);
nand U1792 (N_1792,In_373,In_699);
and U1793 (N_1793,In_533,In_504);
or U1794 (N_1794,In_576,In_569);
or U1795 (N_1795,In_142,In_122);
nand U1796 (N_1796,In_136,In_363);
and U1797 (N_1797,In_904,In_486);
or U1798 (N_1798,In_106,In_887);
or U1799 (N_1799,In_862,In_349);
nor U1800 (N_1800,In_774,In_896);
nor U1801 (N_1801,In_965,In_126);
and U1802 (N_1802,In_503,In_185);
and U1803 (N_1803,In_676,In_602);
nor U1804 (N_1804,In_43,In_543);
xor U1805 (N_1805,In_28,In_249);
nor U1806 (N_1806,In_409,In_178);
and U1807 (N_1807,In_905,In_446);
and U1808 (N_1808,In_113,In_242);
and U1809 (N_1809,In_788,In_172);
and U1810 (N_1810,In_687,In_344);
nor U1811 (N_1811,In_127,In_95);
or U1812 (N_1812,In_943,In_412);
and U1813 (N_1813,In_871,In_796);
or U1814 (N_1814,In_327,In_220);
nor U1815 (N_1815,In_940,In_915);
nor U1816 (N_1816,In_977,In_7);
or U1817 (N_1817,In_463,In_959);
nand U1818 (N_1818,In_651,In_316);
nand U1819 (N_1819,In_885,In_483);
nor U1820 (N_1820,In_610,In_654);
and U1821 (N_1821,In_968,In_306);
or U1822 (N_1822,In_751,In_842);
and U1823 (N_1823,In_492,In_642);
and U1824 (N_1824,In_669,In_400);
and U1825 (N_1825,In_340,In_986);
and U1826 (N_1826,In_514,In_122);
nand U1827 (N_1827,In_950,In_204);
nand U1828 (N_1828,In_495,In_240);
nand U1829 (N_1829,In_731,In_335);
nand U1830 (N_1830,In_495,In_351);
nor U1831 (N_1831,In_615,In_917);
and U1832 (N_1832,In_897,In_171);
and U1833 (N_1833,In_274,In_216);
nand U1834 (N_1834,In_45,In_386);
or U1835 (N_1835,In_565,In_356);
or U1836 (N_1836,In_33,In_948);
or U1837 (N_1837,In_518,In_198);
xnor U1838 (N_1838,In_10,In_876);
xor U1839 (N_1839,In_759,In_744);
or U1840 (N_1840,In_115,In_890);
or U1841 (N_1841,In_341,In_961);
xor U1842 (N_1842,In_509,In_896);
or U1843 (N_1843,In_836,In_924);
nor U1844 (N_1844,In_694,In_399);
nor U1845 (N_1845,In_908,In_864);
nor U1846 (N_1846,In_463,In_361);
and U1847 (N_1847,In_816,In_626);
nand U1848 (N_1848,In_621,In_728);
and U1849 (N_1849,In_887,In_17);
nand U1850 (N_1850,In_665,In_656);
and U1851 (N_1851,In_279,In_267);
or U1852 (N_1852,In_865,In_501);
nand U1853 (N_1853,In_725,In_202);
nor U1854 (N_1854,In_845,In_226);
nand U1855 (N_1855,In_506,In_99);
and U1856 (N_1856,In_504,In_350);
and U1857 (N_1857,In_982,In_285);
or U1858 (N_1858,In_896,In_434);
nor U1859 (N_1859,In_436,In_226);
or U1860 (N_1860,In_425,In_30);
or U1861 (N_1861,In_943,In_658);
nand U1862 (N_1862,In_996,In_125);
nor U1863 (N_1863,In_743,In_944);
nand U1864 (N_1864,In_729,In_969);
or U1865 (N_1865,In_809,In_523);
and U1866 (N_1866,In_537,In_536);
and U1867 (N_1867,In_859,In_392);
nor U1868 (N_1868,In_73,In_787);
or U1869 (N_1869,In_785,In_126);
nand U1870 (N_1870,In_346,In_331);
xor U1871 (N_1871,In_769,In_739);
and U1872 (N_1872,In_309,In_257);
nor U1873 (N_1873,In_630,In_280);
nor U1874 (N_1874,In_203,In_29);
and U1875 (N_1875,In_887,In_532);
nor U1876 (N_1876,In_566,In_933);
nand U1877 (N_1877,In_191,In_723);
nand U1878 (N_1878,In_754,In_604);
nand U1879 (N_1879,In_421,In_303);
and U1880 (N_1880,In_385,In_451);
nor U1881 (N_1881,In_84,In_298);
and U1882 (N_1882,In_997,In_952);
nor U1883 (N_1883,In_851,In_907);
and U1884 (N_1884,In_667,In_346);
or U1885 (N_1885,In_244,In_328);
nand U1886 (N_1886,In_145,In_902);
nand U1887 (N_1887,In_376,In_726);
nand U1888 (N_1888,In_671,In_306);
nor U1889 (N_1889,In_746,In_300);
or U1890 (N_1890,In_245,In_568);
and U1891 (N_1891,In_50,In_793);
and U1892 (N_1892,In_529,In_547);
nor U1893 (N_1893,In_808,In_682);
nor U1894 (N_1894,In_812,In_117);
nor U1895 (N_1895,In_457,In_226);
and U1896 (N_1896,In_121,In_739);
nor U1897 (N_1897,In_226,In_920);
and U1898 (N_1898,In_747,In_404);
nand U1899 (N_1899,In_913,In_640);
and U1900 (N_1900,In_320,In_675);
nor U1901 (N_1901,In_944,In_858);
xor U1902 (N_1902,In_368,In_884);
nand U1903 (N_1903,In_935,In_762);
nand U1904 (N_1904,In_917,In_41);
nand U1905 (N_1905,In_350,In_395);
or U1906 (N_1906,In_26,In_225);
and U1907 (N_1907,In_209,In_775);
and U1908 (N_1908,In_758,In_190);
nor U1909 (N_1909,In_197,In_467);
and U1910 (N_1910,In_101,In_582);
and U1911 (N_1911,In_990,In_126);
nand U1912 (N_1912,In_579,In_726);
and U1913 (N_1913,In_8,In_985);
nor U1914 (N_1914,In_769,In_80);
nor U1915 (N_1915,In_842,In_306);
nand U1916 (N_1916,In_210,In_71);
nor U1917 (N_1917,In_292,In_971);
and U1918 (N_1918,In_722,In_669);
and U1919 (N_1919,In_661,In_316);
nand U1920 (N_1920,In_114,In_417);
and U1921 (N_1921,In_447,In_190);
or U1922 (N_1922,In_535,In_963);
nor U1923 (N_1923,In_821,In_152);
nor U1924 (N_1924,In_307,In_635);
nor U1925 (N_1925,In_994,In_487);
nor U1926 (N_1926,In_230,In_188);
or U1927 (N_1927,In_681,In_743);
and U1928 (N_1928,In_18,In_679);
and U1929 (N_1929,In_987,In_249);
or U1930 (N_1930,In_161,In_366);
nor U1931 (N_1931,In_459,In_146);
nand U1932 (N_1932,In_999,In_908);
nor U1933 (N_1933,In_764,In_630);
xnor U1934 (N_1934,In_40,In_450);
nand U1935 (N_1935,In_302,In_433);
and U1936 (N_1936,In_637,In_661);
nand U1937 (N_1937,In_807,In_698);
nor U1938 (N_1938,In_94,In_455);
or U1939 (N_1939,In_268,In_165);
or U1940 (N_1940,In_845,In_193);
nand U1941 (N_1941,In_657,In_519);
xnor U1942 (N_1942,In_126,In_120);
and U1943 (N_1943,In_40,In_837);
nand U1944 (N_1944,In_641,In_629);
nand U1945 (N_1945,In_132,In_355);
nor U1946 (N_1946,In_981,In_42);
or U1947 (N_1947,In_301,In_897);
nand U1948 (N_1948,In_703,In_575);
and U1949 (N_1949,In_55,In_462);
or U1950 (N_1950,In_718,In_197);
and U1951 (N_1951,In_0,In_243);
and U1952 (N_1952,In_887,In_401);
or U1953 (N_1953,In_43,In_7);
or U1954 (N_1954,In_194,In_204);
nor U1955 (N_1955,In_758,In_100);
nor U1956 (N_1956,In_376,In_646);
nor U1957 (N_1957,In_811,In_249);
xnor U1958 (N_1958,In_140,In_280);
and U1959 (N_1959,In_490,In_825);
or U1960 (N_1960,In_575,In_482);
nand U1961 (N_1961,In_724,In_382);
nand U1962 (N_1962,In_293,In_752);
nor U1963 (N_1963,In_752,In_898);
nor U1964 (N_1964,In_873,In_577);
nand U1965 (N_1965,In_478,In_925);
nand U1966 (N_1966,In_542,In_354);
or U1967 (N_1967,In_200,In_446);
or U1968 (N_1968,In_580,In_238);
or U1969 (N_1969,In_369,In_629);
and U1970 (N_1970,In_567,In_299);
and U1971 (N_1971,In_889,In_420);
nand U1972 (N_1972,In_227,In_827);
or U1973 (N_1973,In_569,In_941);
and U1974 (N_1974,In_415,In_357);
nand U1975 (N_1975,In_948,In_479);
and U1976 (N_1976,In_600,In_33);
and U1977 (N_1977,In_60,In_325);
and U1978 (N_1978,In_63,In_104);
nand U1979 (N_1979,In_173,In_548);
nand U1980 (N_1980,In_965,In_940);
nor U1981 (N_1981,In_259,In_627);
nor U1982 (N_1982,In_286,In_748);
or U1983 (N_1983,In_713,In_883);
or U1984 (N_1984,In_287,In_432);
or U1985 (N_1985,In_206,In_473);
xor U1986 (N_1986,In_692,In_72);
and U1987 (N_1987,In_842,In_668);
nand U1988 (N_1988,In_459,In_392);
nand U1989 (N_1989,In_540,In_138);
and U1990 (N_1990,In_332,In_216);
or U1991 (N_1991,In_807,In_715);
nor U1992 (N_1992,In_702,In_364);
nand U1993 (N_1993,In_441,In_715);
and U1994 (N_1994,In_793,In_895);
xnor U1995 (N_1995,In_478,In_990);
and U1996 (N_1996,In_692,In_17);
and U1997 (N_1997,In_71,In_932);
nand U1998 (N_1998,In_276,In_745);
nor U1999 (N_1999,In_996,In_508);
nand U2000 (N_2000,In_691,In_894);
nor U2001 (N_2001,In_187,In_872);
nand U2002 (N_2002,In_601,In_246);
nand U2003 (N_2003,In_433,In_315);
or U2004 (N_2004,In_21,In_691);
or U2005 (N_2005,In_518,In_266);
nand U2006 (N_2006,In_446,In_252);
or U2007 (N_2007,In_209,In_902);
nor U2008 (N_2008,In_72,In_353);
and U2009 (N_2009,In_954,In_889);
or U2010 (N_2010,In_405,In_359);
nor U2011 (N_2011,In_726,In_829);
nand U2012 (N_2012,In_845,In_584);
xor U2013 (N_2013,In_566,In_173);
or U2014 (N_2014,In_977,In_423);
and U2015 (N_2015,In_375,In_7);
and U2016 (N_2016,In_319,In_192);
and U2017 (N_2017,In_179,In_670);
nor U2018 (N_2018,In_580,In_190);
and U2019 (N_2019,In_279,In_200);
and U2020 (N_2020,In_411,In_651);
or U2021 (N_2021,In_160,In_61);
nand U2022 (N_2022,In_503,In_991);
nand U2023 (N_2023,In_45,In_211);
or U2024 (N_2024,In_438,In_994);
nand U2025 (N_2025,In_819,In_960);
or U2026 (N_2026,In_81,In_464);
and U2027 (N_2027,In_281,In_957);
or U2028 (N_2028,In_85,In_582);
nand U2029 (N_2029,In_949,In_963);
xor U2030 (N_2030,In_451,In_811);
or U2031 (N_2031,In_853,In_2);
or U2032 (N_2032,In_955,In_976);
and U2033 (N_2033,In_130,In_931);
and U2034 (N_2034,In_636,In_625);
and U2035 (N_2035,In_836,In_297);
nand U2036 (N_2036,In_71,In_709);
nor U2037 (N_2037,In_895,In_374);
or U2038 (N_2038,In_821,In_537);
or U2039 (N_2039,In_907,In_35);
or U2040 (N_2040,In_961,In_446);
nor U2041 (N_2041,In_24,In_903);
and U2042 (N_2042,In_695,In_916);
and U2043 (N_2043,In_953,In_434);
and U2044 (N_2044,In_730,In_57);
and U2045 (N_2045,In_395,In_110);
and U2046 (N_2046,In_13,In_828);
xor U2047 (N_2047,In_264,In_134);
or U2048 (N_2048,In_934,In_458);
and U2049 (N_2049,In_490,In_212);
nand U2050 (N_2050,In_370,In_296);
nand U2051 (N_2051,In_836,In_894);
nor U2052 (N_2052,In_733,In_580);
and U2053 (N_2053,In_812,In_800);
and U2054 (N_2054,In_185,In_161);
or U2055 (N_2055,In_784,In_460);
nor U2056 (N_2056,In_552,In_646);
or U2057 (N_2057,In_296,In_56);
nand U2058 (N_2058,In_590,In_979);
or U2059 (N_2059,In_8,In_909);
nor U2060 (N_2060,In_149,In_308);
and U2061 (N_2061,In_936,In_562);
or U2062 (N_2062,In_80,In_741);
and U2063 (N_2063,In_649,In_315);
nor U2064 (N_2064,In_701,In_885);
and U2065 (N_2065,In_838,In_30);
and U2066 (N_2066,In_889,In_998);
or U2067 (N_2067,In_605,In_76);
and U2068 (N_2068,In_163,In_390);
or U2069 (N_2069,In_84,In_104);
or U2070 (N_2070,In_874,In_288);
or U2071 (N_2071,In_504,In_810);
nand U2072 (N_2072,In_563,In_267);
nor U2073 (N_2073,In_618,In_116);
nor U2074 (N_2074,In_982,In_27);
nor U2075 (N_2075,In_420,In_587);
nor U2076 (N_2076,In_566,In_78);
nand U2077 (N_2077,In_430,In_667);
nor U2078 (N_2078,In_669,In_705);
or U2079 (N_2079,In_974,In_615);
or U2080 (N_2080,In_791,In_555);
nor U2081 (N_2081,In_236,In_711);
or U2082 (N_2082,In_490,In_921);
xnor U2083 (N_2083,In_300,In_903);
nand U2084 (N_2084,In_244,In_482);
nand U2085 (N_2085,In_514,In_982);
and U2086 (N_2086,In_341,In_912);
nand U2087 (N_2087,In_666,In_494);
or U2088 (N_2088,In_993,In_410);
or U2089 (N_2089,In_796,In_48);
nor U2090 (N_2090,In_594,In_534);
nor U2091 (N_2091,In_300,In_550);
and U2092 (N_2092,In_660,In_347);
nand U2093 (N_2093,In_718,In_985);
or U2094 (N_2094,In_690,In_692);
and U2095 (N_2095,In_847,In_770);
nor U2096 (N_2096,In_574,In_578);
nor U2097 (N_2097,In_256,In_550);
nor U2098 (N_2098,In_617,In_131);
nand U2099 (N_2099,In_787,In_197);
and U2100 (N_2100,In_559,In_449);
nand U2101 (N_2101,In_143,In_70);
and U2102 (N_2102,In_213,In_640);
nand U2103 (N_2103,In_210,In_328);
nand U2104 (N_2104,In_827,In_634);
xnor U2105 (N_2105,In_310,In_931);
or U2106 (N_2106,In_678,In_987);
nor U2107 (N_2107,In_249,In_370);
and U2108 (N_2108,In_320,In_466);
nand U2109 (N_2109,In_296,In_861);
or U2110 (N_2110,In_231,In_616);
nand U2111 (N_2111,In_327,In_899);
nor U2112 (N_2112,In_898,In_274);
nand U2113 (N_2113,In_342,In_451);
nor U2114 (N_2114,In_328,In_501);
and U2115 (N_2115,In_252,In_186);
or U2116 (N_2116,In_272,In_277);
or U2117 (N_2117,In_161,In_108);
and U2118 (N_2118,In_685,In_800);
and U2119 (N_2119,In_94,In_173);
nand U2120 (N_2120,In_731,In_346);
and U2121 (N_2121,In_627,In_885);
or U2122 (N_2122,In_306,In_461);
and U2123 (N_2123,In_138,In_72);
nor U2124 (N_2124,In_594,In_963);
nor U2125 (N_2125,In_684,In_790);
nand U2126 (N_2126,In_513,In_158);
nor U2127 (N_2127,In_721,In_363);
nor U2128 (N_2128,In_335,In_120);
xnor U2129 (N_2129,In_432,In_241);
nor U2130 (N_2130,In_917,In_225);
nand U2131 (N_2131,In_183,In_190);
or U2132 (N_2132,In_478,In_840);
and U2133 (N_2133,In_12,In_153);
and U2134 (N_2134,In_211,In_609);
nor U2135 (N_2135,In_859,In_319);
nor U2136 (N_2136,In_505,In_516);
or U2137 (N_2137,In_612,In_502);
nand U2138 (N_2138,In_370,In_552);
or U2139 (N_2139,In_560,In_334);
or U2140 (N_2140,In_852,In_438);
and U2141 (N_2141,In_223,In_768);
nor U2142 (N_2142,In_780,In_920);
and U2143 (N_2143,In_362,In_903);
or U2144 (N_2144,In_680,In_152);
and U2145 (N_2145,In_995,In_428);
nor U2146 (N_2146,In_988,In_549);
nand U2147 (N_2147,In_694,In_830);
or U2148 (N_2148,In_252,In_47);
nor U2149 (N_2149,In_110,In_831);
and U2150 (N_2150,In_559,In_937);
or U2151 (N_2151,In_603,In_509);
xor U2152 (N_2152,In_633,In_508);
nand U2153 (N_2153,In_932,In_655);
nor U2154 (N_2154,In_929,In_20);
nand U2155 (N_2155,In_967,In_870);
and U2156 (N_2156,In_894,In_155);
and U2157 (N_2157,In_326,In_577);
nand U2158 (N_2158,In_527,In_256);
and U2159 (N_2159,In_126,In_616);
nand U2160 (N_2160,In_832,In_915);
nor U2161 (N_2161,In_233,In_647);
nor U2162 (N_2162,In_350,In_855);
or U2163 (N_2163,In_333,In_352);
or U2164 (N_2164,In_192,In_10);
and U2165 (N_2165,In_734,In_111);
nor U2166 (N_2166,In_674,In_27);
or U2167 (N_2167,In_215,In_131);
nor U2168 (N_2168,In_760,In_2);
or U2169 (N_2169,In_465,In_573);
or U2170 (N_2170,In_686,In_512);
or U2171 (N_2171,In_195,In_642);
xor U2172 (N_2172,In_712,In_953);
and U2173 (N_2173,In_408,In_507);
and U2174 (N_2174,In_33,In_464);
or U2175 (N_2175,In_18,In_743);
xnor U2176 (N_2176,In_902,In_771);
and U2177 (N_2177,In_602,In_824);
xor U2178 (N_2178,In_12,In_860);
nand U2179 (N_2179,In_736,In_577);
nand U2180 (N_2180,In_364,In_752);
and U2181 (N_2181,In_227,In_26);
nand U2182 (N_2182,In_366,In_4);
nand U2183 (N_2183,In_850,In_448);
xor U2184 (N_2184,In_933,In_190);
nand U2185 (N_2185,In_597,In_236);
nand U2186 (N_2186,In_382,In_657);
nor U2187 (N_2187,In_429,In_79);
nand U2188 (N_2188,In_967,In_652);
nor U2189 (N_2189,In_578,In_416);
xor U2190 (N_2190,In_46,In_31);
nand U2191 (N_2191,In_694,In_174);
nand U2192 (N_2192,In_932,In_83);
and U2193 (N_2193,In_570,In_680);
and U2194 (N_2194,In_243,In_515);
or U2195 (N_2195,In_669,In_534);
nor U2196 (N_2196,In_630,In_501);
or U2197 (N_2197,In_173,In_769);
nand U2198 (N_2198,In_224,In_952);
xnor U2199 (N_2199,In_323,In_38);
and U2200 (N_2200,In_330,In_761);
nand U2201 (N_2201,In_964,In_73);
or U2202 (N_2202,In_573,In_777);
nor U2203 (N_2203,In_321,In_128);
and U2204 (N_2204,In_761,In_279);
and U2205 (N_2205,In_194,In_553);
and U2206 (N_2206,In_249,In_192);
nor U2207 (N_2207,In_38,In_575);
nand U2208 (N_2208,In_389,In_686);
nor U2209 (N_2209,In_361,In_973);
or U2210 (N_2210,In_106,In_323);
nand U2211 (N_2211,In_613,In_775);
nor U2212 (N_2212,In_558,In_441);
nor U2213 (N_2213,In_295,In_415);
or U2214 (N_2214,In_887,In_390);
nor U2215 (N_2215,In_945,In_704);
or U2216 (N_2216,In_322,In_732);
nand U2217 (N_2217,In_623,In_916);
and U2218 (N_2218,In_883,In_720);
or U2219 (N_2219,In_744,In_747);
nand U2220 (N_2220,In_756,In_162);
or U2221 (N_2221,In_234,In_777);
xor U2222 (N_2222,In_319,In_521);
and U2223 (N_2223,In_90,In_794);
nand U2224 (N_2224,In_921,In_872);
nand U2225 (N_2225,In_375,In_699);
and U2226 (N_2226,In_613,In_997);
nand U2227 (N_2227,In_439,In_999);
nand U2228 (N_2228,In_387,In_396);
and U2229 (N_2229,In_903,In_43);
nand U2230 (N_2230,In_596,In_677);
or U2231 (N_2231,In_286,In_352);
nor U2232 (N_2232,In_205,In_327);
nand U2233 (N_2233,In_220,In_243);
nand U2234 (N_2234,In_985,In_338);
xor U2235 (N_2235,In_127,In_172);
nand U2236 (N_2236,In_324,In_782);
nor U2237 (N_2237,In_526,In_260);
xnor U2238 (N_2238,In_686,In_290);
nor U2239 (N_2239,In_348,In_579);
or U2240 (N_2240,In_509,In_487);
and U2241 (N_2241,In_505,In_555);
or U2242 (N_2242,In_750,In_743);
nor U2243 (N_2243,In_79,In_33);
and U2244 (N_2244,In_244,In_442);
nand U2245 (N_2245,In_725,In_278);
xnor U2246 (N_2246,In_316,In_578);
and U2247 (N_2247,In_849,In_748);
and U2248 (N_2248,In_934,In_628);
or U2249 (N_2249,In_984,In_399);
or U2250 (N_2250,In_798,In_690);
or U2251 (N_2251,In_779,In_496);
nand U2252 (N_2252,In_962,In_748);
nor U2253 (N_2253,In_396,In_972);
or U2254 (N_2254,In_279,In_768);
or U2255 (N_2255,In_527,In_239);
and U2256 (N_2256,In_178,In_568);
and U2257 (N_2257,In_47,In_268);
nand U2258 (N_2258,In_150,In_808);
or U2259 (N_2259,In_809,In_697);
nor U2260 (N_2260,In_927,In_412);
nand U2261 (N_2261,In_978,In_945);
nand U2262 (N_2262,In_351,In_224);
nor U2263 (N_2263,In_247,In_529);
and U2264 (N_2264,In_175,In_867);
nor U2265 (N_2265,In_865,In_490);
nand U2266 (N_2266,In_991,In_70);
or U2267 (N_2267,In_456,In_371);
nand U2268 (N_2268,In_632,In_925);
or U2269 (N_2269,In_9,In_487);
nor U2270 (N_2270,In_872,In_772);
or U2271 (N_2271,In_76,In_229);
and U2272 (N_2272,In_565,In_382);
or U2273 (N_2273,In_797,In_361);
or U2274 (N_2274,In_173,In_516);
xnor U2275 (N_2275,In_632,In_442);
and U2276 (N_2276,In_148,In_932);
nand U2277 (N_2277,In_945,In_474);
nand U2278 (N_2278,In_696,In_612);
nor U2279 (N_2279,In_533,In_5);
and U2280 (N_2280,In_830,In_798);
or U2281 (N_2281,In_854,In_883);
nor U2282 (N_2282,In_122,In_360);
and U2283 (N_2283,In_746,In_322);
and U2284 (N_2284,In_259,In_492);
nor U2285 (N_2285,In_923,In_137);
or U2286 (N_2286,In_951,In_950);
nand U2287 (N_2287,In_407,In_796);
nand U2288 (N_2288,In_587,In_978);
and U2289 (N_2289,In_421,In_879);
nor U2290 (N_2290,In_582,In_996);
and U2291 (N_2291,In_796,In_867);
and U2292 (N_2292,In_496,In_294);
nor U2293 (N_2293,In_31,In_700);
nor U2294 (N_2294,In_25,In_550);
nand U2295 (N_2295,In_824,In_229);
nand U2296 (N_2296,In_974,In_296);
nor U2297 (N_2297,In_302,In_942);
nand U2298 (N_2298,In_172,In_800);
xnor U2299 (N_2299,In_10,In_50);
and U2300 (N_2300,In_171,In_62);
nand U2301 (N_2301,In_185,In_944);
nand U2302 (N_2302,In_857,In_531);
and U2303 (N_2303,In_120,In_437);
nor U2304 (N_2304,In_265,In_160);
nor U2305 (N_2305,In_634,In_966);
or U2306 (N_2306,In_815,In_899);
or U2307 (N_2307,In_937,In_307);
nand U2308 (N_2308,In_564,In_917);
or U2309 (N_2309,In_788,In_258);
nand U2310 (N_2310,In_557,In_185);
and U2311 (N_2311,In_759,In_463);
nand U2312 (N_2312,In_917,In_717);
and U2313 (N_2313,In_26,In_810);
nor U2314 (N_2314,In_980,In_217);
nor U2315 (N_2315,In_631,In_522);
nor U2316 (N_2316,In_102,In_90);
or U2317 (N_2317,In_38,In_369);
or U2318 (N_2318,In_976,In_722);
and U2319 (N_2319,In_666,In_324);
or U2320 (N_2320,In_577,In_420);
xnor U2321 (N_2321,In_896,In_321);
and U2322 (N_2322,In_489,In_774);
nand U2323 (N_2323,In_320,In_311);
nand U2324 (N_2324,In_255,In_585);
and U2325 (N_2325,In_742,In_374);
nand U2326 (N_2326,In_500,In_217);
nand U2327 (N_2327,In_937,In_570);
or U2328 (N_2328,In_546,In_659);
or U2329 (N_2329,In_384,In_606);
or U2330 (N_2330,In_606,In_320);
nor U2331 (N_2331,In_723,In_504);
and U2332 (N_2332,In_337,In_344);
and U2333 (N_2333,In_821,In_108);
or U2334 (N_2334,In_896,In_537);
nand U2335 (N_2335,In_133,In_356);
nor U2336 (N_2336,In_181,In_465);
nand U2337 (N_2337,In_293,In_367);
nand U2338 (N_2338,In_577,In_68);
nand U2339 (N_2339,In_80,In_465);
and U2340 (N_2340,In_268,In_275);
xnor U2341 (N_2341,In_174,In_539);
and U2342 (N_2342,In_676,In_178);
and U2343 (N_2343,In_428,In_495);
nand U2344 (N_2344,In_41,In_61);
and U2345 (N_2345,In_84,In_956);
nor U2346 (N_2346,In_206,In_657);
nor U2347 (N_2347,In_34,In_252);
nor U2348 (N_2348,In_989,In_339);
nor U2349 (N_2349,In_16,In_210);
and U2350 (N_2350,In_817,In_728);
or U2351 (N_2351,In_564,In_593);
and U2352 (N_2352,In_830,In_301);
and U2353 (N_2353,In_482,In_533);
or U2354 (N_2354,In_205,In_78);
nand U2355 (N_2355,In_109,In_147);
nand U2356 (N_2356,In_676,In_584);
nor U2357 (N_2357,In_871,In_110);
nor U2358 (N_2358,In_941,In_73);
or U2359 (N_2359,In_183,In_650);
or U2360 (N_2360,In_695,In_514);
and U2361 (N_2361,In_218,In_971);
xnor U2362 (N_2362,In_156,In_546);
nand U2363 (N_2363,In_172,In_730);
nand U2364 (N_2364,In_627,In_767);
nand U2365 (N_2365,In_978,In_146);
nor U2366 (N_2366,In_811,In_906);
nand U2367 (N_2367,In_466,In_362);
and U2368 (N_2368,In_652,In_692);
and U2369 (N_2369,In_49,In_115);
and U2370 (N_2370,In_752,In_747);
or U2371 (N_2371,In_121,In_403);
xor U2372 (N_2372,In_489,In_330);
and U2373 (N_2373,In_248,In_771);
nand U2374 (N_2374,In_627,In_864);
nand U2375 (N_2375,In_453,In_188);
nand U2376 (N_2376,In_706,In_257);
or U2377 (N_2377,In_507,In_324);
and U2378 (N_2378,In_729,In_301);
nor U2379 (N_2379,In_856,In_841);
and U2380 (N_2380,In_734,In_549);
nand U2381 (N_2381,In_286,In_755);
or U2382 (N_2382,In_616,In_560);
nor U2383 (N_2383,In_899,In_217);
or U2384 (N_2384,In_554,In_518);
nor U2385 (N_2385,In_551,In_256);
nor U2386 (N_2386,In_390,In_667);
and U2387 (N_2387,In_775,In_58);
or U2388 (N_2388,In_486,In_5);
or U2389 (N_2389,In_938,In_715);
nand U2390 (N_2390,In_354,In_207);
and U2391 (N_2391,In_166,In_692);
nand U2392 (N_2392,In_976,In_678);
nand U2393 (N_2393,In_860,In_810);
and U2394 (N_2394,In_844,In_791);
and U2395 (N_2395,In_620,In_348);
and U2396 (N_2396,In_481,In_23);
nand U2397 (N_2397,In_974,In_212);
nand U2398 (N_2398,In_758,In_294);
and U2399 (N_2399,In_883,In_633);
nand U2400 (N_2400,In_314,In_77);
or U2401 (N_2401,In_632,In_602);
or U2402 (N_2402,In_71,In_844);
and U2403 (N_2403,In_828,In_519);
nand U2404 (N_2404,In_9,In_997);
nor U2405 (N_2405,In_78,In_462);
and U2406 (N_2406,In_15,In_206);
or U2407 (N_2407,In_823,In_926);
and U2408 (N_2408,In_348,In_153);
nor U2409 (N_2409,In_881,In_706);
nor U2410 (N_2410,In_333,In_232);
nor U2411 (N_2411,In_239,In_75);
and U2412 (N_2412,In_882,In_243);
or U2413 (N_2413,In_975,In_728);
or U2414 (N_2414,In_547,In_612);
nand U2415 (N_2415,In_346,In_173);
nand U2416 (N_2416,In_911,In_136);
nor U2417 (N_2417,In_19,In_904);
nor U2418 (N_2418,In_455,In_576);
and U2419 (N_2419,In_153,In_479);
and U2420 (N_2420,In_137,In_293);
nand U2421 (N_2421,In_916,In_128);
nor U2422 (N_2422,In_296,In_729);
nand U2423 (N_2423,In_785,In_503);
nor U2424 (N_2424,In_62,In_142);
or U2425 (N_2425,In_434,In_279);
and U2426 (N_2426,In_136,In_819);
nand U2427 (N_2427,In_771,In_107);
nor U2428 (N_2428,In_778,In_563);
and U2429 (N_2429,In_650,In_9);
or U2430 (N_2430,In_30,In_114);
or U2431 (N_2431,In_57,In_668);
nand U2432 (N_2432,In_412,In_506);
nor U2433 (N_2433,In_186,In_116);
nand U2434 (N_2434,In_126,In_499);
or U2435 (N_2435,In_373,In_551);
and U2436 (N_2436,In_965,In_471);
or U2437 (N_2437,In_570,In_279);
nor U2438 (N_2438,In_407,In_167);
or U2439 (N_2439,In_61,In_142);
nor U2440 (N_2440,In_718,In_690);
and U2441 (N_2441,In_499,In_369);
nor U2442 (N_2442,In_849,In_388);
nand U2443 (N_2443,In_958,In_997);
nor U2444 (N_2444,In_879,In_338);
and U2445 (N_2445,In_275,In_793);
and U2446 (N_2446,In_914,In_701);
xnor U2447 (N_2447,In_448,In_316);
and U2448 (N_2448,In_963,In_798);
and U2449 (N_2449,In_560,In_153);
or U2450 (N_2450,In_71,In_901);
or U2451 (N_2451,In_857,In_373);
or U2452 (N_2452,In_157,In_970);
nor U2453 (N_2453,In_937,In_687);
or U2454 (N_2454,In_619,In_156);
and U2455 (N_2455,In_863,In_938);
or U2456 (N_2456,In_979,In_905);
or U2457 (N_2457,In_607,In_658);
and U2458 (N_2458,In_779,In_568);
and U2459 (N_2459,In_995,In_225);
nand U2460 (N_2460,In_505,In_224);
and U2461 (N_2461,In_122,In_427);
xor U2462 (N_2462,In_572,In_487);
nor U2463 (N_2463,In_57,In_760);
or U2464 (N_2464,In_945,In_800);
nor U2465 (N_2465,In_820,In_123);
nand U2466 (N_2466,In_890,In_690);
nand U2467 (N_2467,In_184,In_714);
or U2468 (N_2468,In_518,In_456);
and U2469 (N_2469,In_274,In_446);
nand U2470 (N_2470,In_722,In_908);
and U2471 (N_2471,In_141,In_994);
nor U2472 (N_2472,In_742,In_76);
and U2473 (N_2473,In_484,In_894);
nor U2474 (N_2474,In_138,In_921);
or U2475 (N_2475,In_103,In_805);
or U2476 (N_2476,In_352,In_155);
and U2477 (N_2477,In_62,In_972);
and U2478 (N_2478,In_253,In_530);
and U2479 (N_2479,In_768,In_38);
or U2480 (N_2480,In_601,In_813);
and U2481 (N_2481,In_972,In_880);
nor U2482 (N_2482,In_373,In_534);
nor U2483 (N_2483,In_975,In_209);
or U2484 (N_2484,In_727,In_238);
nor U2485 (N_2485,In_832,In_610);
and U2486 (N_2486,In_211,In_548);
nor U2487 (N_2487,In_684,In_30);
or U2488 (N_2488,In_101,In_213);
or U2489 (N_2489,In_867,In_617);
nor U2490 (N_2490,In_814,In_939);
xnor U2491 (N_2491,In_288,In_278);
nor U2492 (N_2492,In_972,In_481);
nand U2493 (N_2493,In_95,In_922);
nor U2494 (N_2494,In_62,In_499);
and U2495 (N_2495,In_697,In_398);
or U2496 (N_2496,In_56,In_329);
and U2497 (N_2497,In_921,In_311);
and U2498 (N_2498,In_461,In_74);
nor U2499 (N_2499,In_114,In_12);
nor U2500 (N_2500,In_190,In_916);
nor U2501 (N_2501,In_412,In_520);
and U2502 (N_2502,In_285,In_261);
or U2503 (N_2503,In_188,In_401);
nor U2504 (N_2504,In_457,In_907);
nand U2505 (N_2505,In_582,In_347);
nand U2506 (N_2506,In_417,In_736);
nand U2507 (N_2507,In_887,In_706);
and U2508 (N_2508,In_65,In_542);
nand U2509 (N_2509,In_905,In_241);
nor U2510 (N_2510,In_726,In_154);
nand U2511 (N_2511,In_244,In_983);
and U2512 (N_2512,In_260,In_557);
xnor U2513 (N_2513,In_885,In_643);
and U2514 (N_2514,In_903,In_238);
nor U2515 (N_2515,In_84,In_23);
nor U2516 (N_2516,In_627,In_212);
or U2517 (N_2517,In_943,In_868);
nor U2518 (N_2518,In_828,In_789);
nand U2519 (N_2519,In_153,In_816);
nor U2520 (N_2520,In_863,In_778);
and U2521 (N_2521,In_243,In_569);
nand U2522 (N_2522,In_186,In_174);
and U2523 (N_2523,In_147,In_881);
or U2524 (N_2524,In_423,In_543);
nor U2525 (N_2525,In_580,In_269);
and U2526 (N_2526,In_9,In_801);
nand U2527 (N_2527,In_282,In_498);
nor U2528 (N_2528,In_394,In_610);
nand U2529 (N_2529,In_909,In_173);
xor U2530 (N_2530,In_903,In_752);
or U2531 (N_2531,In_927,In_419);
or U2532 (N_2532,In_206,In_674);
nand U2533 (N_2533,In_222,In_736);
nor U2534 (N_2534,In_363,In_362);
and U2535 (N_2535,In_863,In_254);
and U2536 (N_2536,In_212,In_152);
nand U2537 (N_2537,In_799,In_242);
nand U2538 (N_2538,In_876,In_133);
or U2539 (N_2539,In_607,In_343);
nand U2540 (N_2540,In_353,In_991);
and U2541 (N_2541,In_253,In_564);
nor U2542 (N_2542,In_4,In_759);
nand U2543 (N_2543,In_650,In_999);
nand U2544 (N_2544,In_664,In_719);
xnor U2545 (N_2545,In_97,In_366);
nand U2546 (N_2546,In_300,In_578);
or U2547 (N_2547,In_704,In_480);
and U2548 (N_2548,In_172,In_293);
and U2549 (N_2549,In_540,In_844);
and U2550 (N_2550,In_390,In_337);
and U2551 (N_2551,In_982,In_611);
and U2552 (N_2552,In_957,In_302);
or U2553 (N_2553,In_375,In_257);
and U2554 (N_2554,In_417,In_960);
nor U2555 (N_2555,In_633,In_894);
or U2556 (N_2556,In_116,In_971);
and U2557 (N_2557,In_998,In_657);
nand U2558 (N_2558,In_188,In_837);
or U2559 (N_2559,In_981,In_289);
and U2560 (N_2560,In_826,In_504);
or U2561 (N_2561,In_999,In_119);
and U2562 (N_2562,In_855,In_857);
xnor U2563 (N_2563,In_500,In_941);
nand U2564 (N_2564,In_359,In_924);
nand U2565 (N_2565,In_456,In_125);
nor U2566 (N_2566,In_171,In_499);
or U2567 (N_2567,In_701,In_805);
or U2568 (N_2568,In_790,In_338);
or U2569 (N_2569,In_428,In_426);
nand U2570 (N_2570,In_828,In_958);
and U2571 (N_2571,In_171,In_714);
or U2572 (N_2572,In_354,In_370);
or U2573 (N_2573,In_462,In_669);
nand U2574 (N_2574,In_66,In_228);
and U2575 (N_2575,In_146,In_224);
nor U2576 (N_2576,In_35,In_695);
nor U2577 (N_2577,In_598,In_403);
xnor U2578 (N_2578,In_14,In_804);
and U2579 (N_2579,In_786,In_37);
and U2580 (N_2580,In_496,In_326);
and U2581 (N_2581,In_407,In_689);
nor U2582 (N_2582,In_444,In_174);
nor U2583 (N_2583,In_214,In_577);
and U2584 (N_2584,In_397,In_289);
nand U2585 (N_2585,In_380,In_220);
or U2586 (N_2586,In_534,In_194);
nand U2587 (N_2587,In_639,In_973);
nor U2588 (N_2588,In_768,In_104);
xor U2589 (N_2589,In_169,In_993);
or U2590 (N_2590,In_280,In_750);
or U2591 (N_2591,In_860,In_919);
nor U2592 (N_2592,In_559,In_125);
nand U2593 (N_2593,In_388,In_959);
and U2594 (N_2594,In_362,In_849);
and U2595 (N_2595,In_545,In_642);
or U2596 (N_2596,In_996,In_493);
xnor U2597 (N_2597,In_198,In_374);
nor U2598 (N_2598,In_641,In_396);
nor U2599 (N_2599,In_592,In_695);
or U2600 (N_2600,In_726,In_51);
or U2601 (N_2601,In_191,In_752);
and U2602 (N_2602,In_363,In_642);
nor U2603 (N_2603,In_398,In_556);
and U2604 (N_2604,In_178,In_223);
nor U2605 (N_2605,In_552,In_636);
nor U2606 (N_2606,In_898,In_325);
nor U2607 (N_2607,In_987,In_989);
nor U2608 (N_2608,In_741,In_388);
and U2609 (N_2609,In_456,In_525);
xor U2610 (N_2610,In_147,In_224);
nand U2611 (N_2611,In_543,In_446);
nand U2612 (N_2612,In_503,In_480);
nor U2613 (N_2613,In_771,In_633);
nor U2614 (N_2614,In_888,In_110);
or U2615 (N_2615,In_399,In_27);
xor U2616 (N_2616,In_633,In_189);
nor U2617 (N_2617,In_124,In_904);
and U2618 (N_2618,In_35,In_719);
nand U2619 (N_2619,In_962,In_573);
and U2620 (N_2620,In_424,In_667);
nor U2621 (N_2621,In_294,In_485);
and U2622 (N_2622,In_376,In_219);
or U2623 (N_2623,In_49,In_63);
or U2624 (N_2624,In_87,In_558);
nor U2625 (N_2625,In_462,In_602);
nand U2626 (N_2626,In_919,In_772);
xor U2627 (N_2627,In_675,In_662);
and U2628 (N_2628,In_543,In_776);
nor U2629 (N_2629,In_428,In_196);
nor U2630 (N_2630,In_552,In_136);
or U2631 (N_2631,In_651,In_322);
or U2632 (N_2632,In_935,In_455);
and U2633 (N_2633,In_12,In_327);
and U2634 (N_2634,In_93,In_922);
nor U2635 (N_2635,In_926,In_771);
nor U2636 (N_2636,In_692,In_150);
nand U2637 (N_2637,In_89,In_628);
nand U2638 (N_2638,In_14,In_277);
nand U2639 (N_2639,In_855,In_725);
and U2640 (N_2640,In_359,In_243);
or U2641 (N_2641,In_435,In_14);
or U2642 (N_2642,In_789,In_856);
nor U2643 (N_2643,In_150,In_504);
or U2644 (N_2644,In_236,In_408);
and U2645 (N_2645,In_782,In_832);
or U2646 (N_2646,In_252,In_143);
nand U2647 (N_2647,In_874,In_372);
or U2648 (N_2648,In_724,In_41);
or U2649 (N_2649,In_482,In_285);
and U2650 (N_2650,In_465,In_504);
nor U2651 (N_2651,In_456,In_482);
nand U2652 (N_2652,In_139,In_12);
or U2653 (N_2653,In_449,In_906);
or U2654 (N_2654,In_707,In_300);
nand U2655 (N_2655,In_639,In_697);
or U2656 (N_2656,In_921,In_376);
nor U2657 (N_2657,In_301,In_90);
nor U2658 (N_2658,In_191,In_76);
or U2659 (N_2659,In_180,In_375);
nor U2660 (N_2660,In_249,In_157);
nor U2661 (N_2661,In_219,In_10);
nor U2662 (N_2662,In_137,In_756);
nor U2663 (N_2663,In_796,In_945);
nand U2664 (N_2664,In_253,In_885);
and U2665 (N_2665,In_984,In_165);
nor U2666 (N_2666,In_157,In_282);
and U2667 (N_2667,In_727,In_45);
and U2668 (N_2668,In_391,In_954);
or U2669 (N_2669,In_626,In_799);
and U2670 (N_2670,In_890,In_673);
or U2671 (N_2671,In_769,In_206);
nand U2672 (N_2672,In_435,In_567);
or U2673 (N_2673,In_731,In_497);
nor U2674 (N_2674,In_686,In_308);
xnor U2675 (N_2675,In_675,In_126);
and U2676 (N_2676,In_854,In_591);
nor U2677 (N_2677,In_372,In_585);
nor U2678 (N_2678,In_652,In_636);
or U2679 (N_2679,In_753,In_915);
nand U2680 (N_2680,In_358,In_799);
nor U2681 (N_2681,In_793,In_392);
and U2682 (N_2682,In_109,In_909);
nor U2683 (N_2683,In_578,In_363);
nand U2684 (N_2684,In_17,In_510);
nor U2685 (N_2685,In_485,In_133);
nor U2686 (N_2686,In_104,In_815);
nand U2687 (N_2687,In_868,In_32);
or U2688 (N_2688,In_476,In_957);
and U2689 (N_2689,In_473,In_122);
nand U2690 (N_2690,In_921,In_682);
nor U2691 (N_2691,In_238,In_145);
nand U2692 (N_2692,In_358,In_280);
and U2693 (N_2693,In_385,In_242);
and U2694 (N_2694,In_800,In_264);
and U2695 (N_2695,In_593,In_26);
nand U2696 (N_2696,In_636,In_591);
nand U2697 (N_2697,In_949,In_843);
or U2698 (N_2698,In_569,In_220);
nor U2699 (N_2699,In_715,In_612);
nor U2700 (N_2700,In_136,In_536);
nand U2701 (N_2701,In_573,In_567);
and U2702 (N_2702,In_9,In_267);
and U2703 (N_2703,In_871,In_395);
nand U2704 (N_2704,In_397,In_90);
or U2705 (N_2705,In_326,In_304);
and U2706 (N_2706,In_475,In_692);
xnor U2707 (N_2707,In_807,In_468);
or U2708 (N_2708,In_742,In_566);
and U2709 (N_2709,In_443,In_287);
and U2710 (N_2710,In_712,In_683);
nor U2711 (N_2711,In_237,In_480);
nor U2712 (N_2712,In_640,In_869);
and U2713 (N_2713,In_403,In_239);
and U2714 (N_2714,In_611,In_231);
nor U2715 (N_2715,In_439,In_770);
or U2716 (N_2716,In_590,In_662);
and U2717 (N_2717,In_898,In_921);
nor U2718 (N_2718,In_225,In_67);
and U2719 (N_2719,In_477,In_806);
or U2720 (N_2720,In_624,In_412);
and U2721 (N_2721,In_979,In_430);
and U2722 (N_2722,In_430,In_784);
or U2723 (N_2723,In_282,In_663);
or U2724 (N_2724,In_182,In_875);
nor U2725 (N_2725,In_83,In_730);
nand U2726 (N_2726,In_576,In_876);
or U2727 (N_2727,In_542,In_746);
or U2728 (N_2728,In_80,In_841);
xor U2729 (N_2729,In_971,In_91);
and U2730 (N_2730,In_708,In_10);
nor U2731 (N_2731,In_5,In_420);
nand U2732 (N_2732,In_336,In_602);
nand U2733 (N_2733,In_314,In_323);
or U2734 (N_2734,In_55,In_69);
nand U2735 (N_2735,In_996,In_737);
nand U2736 (N_2736,In_992,In_328);
or U2737 (N_2737,In_22,In_168);
or U2738 (N_2738,In_483,In_472);
nand U2739 (N_2739,In_513,In_426);
nor U2740 (N_2740,In_935,In_207);
nor U2741 (N_2741,In_403,In_606);
or U2742 (N_2742,In_252,In_152);
nand U2743 (N_2743,In_170,In_580);
or U2744 (N_2744,In_248,In_50);
or U2745 (N_2745,In_200,In_963);
or U2746 (N_2746,In_575,In_644);
nand U2747 (N_2747,In_364,In_773);
or U2748 (N_2748,In_348,In_686);
nor U2749 (N_2749,In_928,In_762);
or U2750 (N_2750,In_974,In_926);
or U2751 (N_2751,In_933,In_458);
nand U2752 (N_2752,In_443,In_742);
nand U2753 (N_2753,In_145,In_821);
nand U2754 (N_2754,In_155,In_811);
or U2755 (N_2755,In_497,In_925);
nor U2756 (N_2756,In_655,In_385);
nor U2757 (N_2757,In_97,In_421);
nand U2758 (N_2758,In_409,In_998);
nor U2759 (N_2759,In_594,In_691);
or U2760 (N_2760,In_832,In_126);
nor U2761 (N_2761,In_861,In_654);
or U2762 (N_2762,In_499,In_149);
xor U2763 (N_2763,In_702,In_906);
or U2764 (N_2764,In_178,In_88);
xnor U2765 (N_2765,In_599,In_224);
or U2766 (N_2766,In_69,In_421);
nand U2767 (N_2767,In_360,In_42);
or U2768 (N_2768,In_154,In_888);
and U2769 (N_2769,In_87,In_242);
nor U2770 (N_2770,In_656,In_926);
or U2771 (N_2771,In_127,In_735);
and U2772 (N_2772,In_883,In_80);
and U2773 (N_2773,In_254,In_845);
or U2774 (N_2774,In_111,In_861);
or U2775 (N_2775,In_717,In_143);
and U2776 (N_2776,In_864,In_143);
nand U2777 (N_2777,In_622,In_511);
nand U2778 (N_2778,In_501,In_599);
nand U2779 (N_2779,In_890,In_851);
nand U2780 (N_2780,In_979,In_780);
and U2781 (N_2781,In_429,In_450);
nand U2782 (N_2782,In_937,In_638);
nor U2783 (N_2783,In_732,In_599);
nand U2784 (N_2784,In_554,In_250);
and U2785 (N_2785,In_538,In_507);
nand U2786 (N_2786,In_260,In_535);
and U2787 (N_2787,In_588,In_686);
xor U2788 (N_2788,In_421,In_795);
nor U2789 (N_2789,In_910,In_646);
nand U2790 (N_2790,In_318,In_648);
or U2791 (N_2791,In_549,In_859);
nand U2792 (N_2792,In_110,In_751);
nor U2793 (N_2793,In_279,In_249);
or U2794 (N_2794,In_836,In_39);
and U2795 (N_2795,In_233,In_628);
and U2796 (N_2796,In_179,In_475);
or U2797 (N_2797,In_256,In_824);
nor U2798 (N_2798,In_11,In_268);
xor U2799 (N_2799,In_496,In_283);
and U2800 (N_2800,In_733,In_806);
or U2801 (N_2801,In_149,In_915);
nor U2802 (N_2802,In_693,In_401);
nor U2803 (N_2803,In_154,In_664);
or U2804 (N_2804,In_961,In_651);
or U2805 (N_2805,In_637,In_340);
or U2806 (N_2806,In_976,In_843);
nand U2807 (N_2807,In_928,In_622);
nand U2808 (N_2808,In_175,In_929);
or U2809 (N_2809,In_545,In_115);
or U2810 (N_2810,In_978,In_18);
or U2811 (N_2811,In_336,In_242);
nand U2812 (N_2812,In_58,In_231);
and U2813 (N_2813,In_415,In_329);
nor U2814 (N_2814,In_129,In_237);
nand U2815 (N_2815,In_663,In_806);
or U2816 (N_2816,In_160,In_975);
and U2817 (N_2817,In_886,In_917);
nand U2818 (N_2818,In_378,In_303);
nor U2819 (N_2819,In_35,In_576);
and U2820 (N_2820,In_492,In_365);
xor U2821 (N_2821,In_818,In_380);
or U2822 (N_2822,In_972,In_42);
nand U2823 (N_2823,In_548,In_831);
nand U2824 (N_2824,In_622,In_177);
and U2825 (N_2825,In_152,In_682);
nand U2826 (N_2826,In_319,In_456);
nand U2827 (N_2827,In_809,In_534);
nand U2828 (N_2828,In_763,In_97);
or U2829 (N_2829,In_376,In_944);
or U2830 (N_2830,In_326,In_663);
or U2831 (N_2831,In_256,In_732);
nand U2832 (N_2832,In_597,In_502);
or U2833 (N_2833,In_443,In_478);
nand U2834 (N_2834,In_605,In_73);
nand U2835 (N_2835,In_73,In_535);
and U2836 (N_2836,In_943,In_74);
and U2837 (N_2837,In_625,In_688);
or U2838 (N_2838,In_464,In_579);
or U2839 (N_2839,In_240,In_304);
nand U2840 (N_2840,In_722,In_107);
nor U2841 (N_2841,In_778,In_432);
nor U2842 (N_2842,In_622,In_836);
nand U2843 (N_2843,In_512,In_681);
nor U2844 (N_2844,In_414,In_186);
nor U2845 (N_2845,In_664,In_486);
or U2846 (N_2846,In_122,In_590);
nor U2847 (N_2847,In_839,In_580);
nand U2848 (N_2848,In_200,In_448);
nor U2849 (N_2849,In_779,In_581);
and U2850 (N_2850,In_350,In_379);
and U2851 (N_2851,In_593,In_210);
nor U2852 (N_2852,In_510,In_944);
nand U2853 (N_2853,In_341,In_255);
nor U2854 (N_2854,In_544,In_5);
xor U2855 (N_2855,In_454,In_658);
or U2856 (N_2856,In_575,In_720);
nor U2857 (N_2857,In_695,In_525);
nand U2858 (N_2858,In_759,In_31);
and U2859 (N_2859,In_580,In_571);
nand U2860 (N_2860,In_407,In_323);
nor U2861 (N_2861,In_818,In_590);
and U2862 (N_2862,In_230,In_565);
and U2863 (N_2863,In_287,In_54);
and U2864 (N_2864,In_820,In_299);
and U2865 (N_2865,In_949,In_100);
nor U2866 (N_2866,In_882,In_733);
xor U2867 (N_2867,In_258,In_931);
or U2868 (N_2868,In_274,In_654);
or U2869 (N_2869,In_520,In_468);
nor U2870 (N_2870,In_540,In_320);
nand U2871 (N_2871,In_77,In_80);
and U2872 (N_2872,In_62,In_620);
nor U2873 (N_2873,In_254,In_758);
and U2874 (N_2874,In_985,In_385);
nor U2875 (N_2875,In_947,In_756);
or U2876 (N_2876,In_803,In_836);
nor U2877 (N_2877,In_160,In_450);
or U2878 (N_2878,In_791,In_685);
nand U2879 (N_2879,In_270,In_570);
nand U2880 (N_2880,In_18,In_941);
and U2881 (N_2881,In_851,In_866);
nand U2882 (N_2882,In_304,In_285);
nor U2883 (N_2883,In_23,In_982);
or U2884 (N_2884,In_129,In_397);
nor U2885 (N_2885,In_633,In_830);
or U2886 (N_2886,In_272,In_163);
nand U2887 (N_2887,In_620,In_339);
nor U2888 (N_2888,In_165,In_778);
and U2889 (N_2889,In_308,In_324);
nor U2890 (N_2890,In_458,In_588);
nand U2891 (N_2891,In_182,In_14);
xnor U2892 (N_2892,In_799,In_320);
and U2893 (N_2893,In_127,In_399);
and U2894 (N_2894,In_764,In_246);
and U2895 (N_2895,In_705,In_655);
or U2896 (N_2896,In_874,In_215);
nor U2897 (N_2897,In_953,In_200);
or U2898 (N_2898,In_228,In_912);
nor U2899 (N_2899,In_521,In_461);
nor U2900 (N_2900,In_558,In_317);
nand U2901 (N_2901,In_1,In_778);
nor U2902 (N_2902,In_3,In_185);
xor U2903 (N_2903,In_95,In_686);
or U2904 (N_2904,In_501,In_378);
and U2905 (N_2905,In_345,In_903);
and U2906 (N_2906,In_517,In_361);
and U2907 (N_2907,In_583,In_644);
or U2908 (N_2908,In_466,In_802);
nor U2909 (N_2909,In_493,In_85);
nand U2910 (N_2910,In_403,In_173);
nand U2911 (N_2911,In_27,In_569);
and U2912 (N_2912,In_8,In_924);
or U2913 (N_2913,In_891,In_403);
nor U2914 (N_2914,In_500,In_170);
nand U2915 (N_2915,In_215,In_996);
and U2916 (N_2916,In_618,In_203);
nor U2917 (N_2917,In_334,In_255);
nand U2918 (N_2918,In_152,In_692);
nor U2919 (N_2919,In_247,In_978);
nor U2920 (N_2920,In_674,In_745);
nor U2921 (N_2921,In_676,In_607);
xnor U2922 (N_2922,In_690,In_169);
nand U2923 (N_2923,In_6,In_311);
nand U2924 (N_2924,In_252,In_691);
nand U2925 (N_2925,In_965,In_556);
nor U2926 (N_2926,In_513,In_601);
xnor U2927 (N_2927,In_651,In_664);
or U2928 (N_2928,In_848,In_115);
or U2929 (N_2929,In_520,In_669);
nor U2930 (N_2930,In_903,In_687);
nand U2931 (N_2931,In_411,In_822);
and U2932 (N_2932,In_342,In_489);
nor U2933 (N_2933,In_779,In_654);
nand U2934 (N_2934,In_145,In_822);
or U2935 (N_2935,In_114,In_830);
nand U2936 (N_2936,In_215,In_545);
and U2937 (N_2937,In_564,In_227);
and U2938 (N_2938,In_782,In_346);
and U2939 (N_2939,In_772,In_681);
and U2940 (N_2940,In_486,In_772);
nand U2941 (N_2941,In_414,In_667);
and U2942 (N_2942,In_602,In_650);
or U2943 (N_2943,In_535,In_729);
or U2944 (N_2944,In_207,In_735);
or U2945 (N_2945,In_677,In_615);
nor U2946 (N_2946,In_831,In_942);
nor U2947 (N_2947,In_18,In_847);
or U2948 (N_2948,In_423,In_14);
or U2949 (N_2949,In_696,In_480);
or U2950 (N_2950,In_111,In_950);
nand U2951 (N_2951,In_504,In_313);
or U2952 (N_2952,In_503,In_745);
or U2953 (N_2953,In_687,In_78);
nand U2954 (N_2954,In_612,In_971);
nor U2955 (N_2955,In_356,In_759);
and U2956 (N_2956,In_92,In_533);
nor U2957 (N_2957,In_181,In_136);
xor U2958 (N_2958,In_826,In_528);
nand U2959 (N_2959,In_403,In_136);
nand U2960 (N_2960,In_43,In_990);
xor U2961 (N_2961,In_71,In_900);
nand U2962 (N_2962,In_17,In_965);
nand U2963 (N_2963,In_295,In_486);
nor U2964 (N_2964,In_424,In_209);
nand U2965 (N_2965,In_653,In_335);
nand U2966 (N_2966,In_4,In_511);
or U2967 (N_2967,In_238,In_196);
xor U2968 (N_2968,In_800,In_173);
or U2969 (N_2969,In_560,In_463);
and U2970 (N_2970,In_347,In_416);
and U2971 (N_2971,In_898,In_392);
or U2972 (N_2972,In_285,In_974);
nor U2973 (N_2973,In_604,In_433);
xnor U2974 (N_2974,In_956,In_276);
xnor U2975 (N_2975,In_940,In_715);
nor U2976 (N_2976,In_914,In_954);
nand U2977 (N_2977,In_425,In_854);
nand U2978 (N_2978,In_335,In_243);
nor U2979 (N_2979,In_812,In_910);
nor U2980 (N_2980,In_71,In_515);
or U2981 (N_2981,In_881,In_165);
and U2982 (N_2982,In_464,In_165);
or U2983 (N_2983,In_416,In_921);
or U2984 (N_2984,In_299,In_216);
or U2985 (N_2985,In_548,In_850);
and U2986 (N_2986,In_974,In_756);
xor U2987 (N_2987,In_244,In_727);
nor U2988 (N_2988,In_702,In_969);
nand U2989 (N_2989,In_552,In_296);
and U2990 (N_2990,In_386,In_404);
nor U2991 (N_2991,In_830,In_674);
or U2992 (N_2992,In_827,In_740);
or U2993 (N_2993,In_594,In_391);
or U2994 (N_2994,In_876,In_290);
or U2995 (N_2995,In_867,In_578);
nor U2996 (N_2996,In_400,In_716);
nand U2997 (N_2997,In_527,In_255);
nand U2998 (N_2998,In_554,In_547);
or U2999 (N_2999,In_13,In_358);
nor U3000 (N_3000,In_566,In_445);
xor U3001 (N_3001,In_456,In_743);
or U3002 (N_3002,In_446,In_192);
and U3003 (N_3003,In_859,In_411);
or U3004 (N_3004,In_944,In_832);
nand U3005 (N_3005,In_234,In_73);
or U3006 (N_3006,In_594,In_302);
or U3007 (N_3007,In_320,In_590);
nand U3008 (N_3008,In_131,In_15);
and U3009 (N_3009,In_504,In_729);
or U3010 (N_3010,In_785,In_211);
nand U3011 (N_3011,In_499,In_851);
or U3012 (N_3012,In_375,In_703);
nand U3013 (N_3013,In_428,In_966);
and U3014 (N_3014,In_954,In_744);
nor U3015 (N_3015,In_377,In_303);
nand U3016 (N_3016,In_2,In_461);
and U3017 (N_3017,In_863,In_366);
nor U3018 (N_3018,In_115,In_647);
xor U3019 (N_3019,In_266,In_154);
and U3020 (N_3020,In_256,In_360);
or U3021 (N_3021,In_620,In_694);
nor U3022 (N_3022,In_583,In_840);
and U3023 (N_3023,In_25,In_594);
or U3024 (N_3024,In_561,In_732);
and U3025 (N_3025,In_518,In_160);
xor U3026 (N_3026,In_803,In_565);
nand U3027 (N_3027,In_878,In_504);
or U3028 (N_3028,In_66,In_499);
nor U3029 (N_3029,In_811,In_99);
and U3030 (N_3030,In_551,In_17);
nand U3031 (N_3031,In_775,In_991);
nand U3032 (N_3032,In_319,In_310);
nand U3033 (N_3033,In_987,In_641);
nand U3034 (N_3034,In_361,In_997);
or U3035 (N_3035,In_418,In_927);
and U3036 (N_3036,In_354,In_165);
nor U3037 (N_3037,In_475,In_472);
xnor U3038 (N_3038,In_468,In_60);
nor U3039 (N_3039,In_911,In_640);
nand U3040 (N_3040,In_333,In_627);
nand U3041 (N_3041,In_31,In_971);
xor U3042 (N_3042,In_101,In_174);
nor U3043 (N_3043,In_320,In_583);
or U3044 (N_3044,In_962,In_922);
nor U3045 (N_3045,In_771,In_241);
nand U3046 (N_3046,In_419,In_994);
nor U3047 (N_3047,In_663,In_384);
nand U3048 (N_3048,In_688,In_490);
nand U3049 (N_3049,In_815,In_987);
nor U3050 (N_3050,In_25,In_873);
and U3051 (N_3051,In_69,In_987);
nor U3052 (N_3052,In_264,In_315);
or U3053 (N_3053,In_839,In_342);
nand U3054 (N_3054,In_586,In_864);
and U3055 (N_3055,In_826,In_515);
nor U3056 (N_3056,In_298,In_987);
nand U3057 (N_3057,In_589,In_274);
nand U3058 (N_3058,In_802,In_14);
and U3059 (N_3059,In_746,In_119);
and U3060 (N_3060,In_955,In_293);
and U3061 (N_3061,In_76,In_749);
nand U3062 (N_3062,In_958,In_848);
and U3063 (N_3063,In_28,In_547);
nand U3064 (N_3064,In_908,In_924);
or U3065 (N_3065,In_497,In_687);
nand U3066 (N_3066,In_408,In_109);
or U3067 (N_3067,In_323,In_864);
nand U3068 (N_3068,In_561,In_865);
and U3069 (N_3069,In_199,In_695);
or U3070 (N_3070,In_242,In_700);
and U3071 (N_3071,In_140,In_947);
nand U3072 (N_3072,In_980,In_598);
or U3073 (N_3073,In_263,In_412);
and U3074 (N_3074,In_684,In_948);
nand U3075 (N_3075,In_94,In_979);
or U3076 (N_3076,In_604,In_472);
nor U3077 (N_3077,In_751,In_457);
nor U3078 (N_3078,In_387,In_984);
xnor U3079 (N_3079,In_915,In_328);
nor U3080 (N_3080,In_53,In_673);
and U3081 (N_3081,In_564,In_631);
nand U3082 (N_3082,In_16,In_863);
or U3083 (N_3083,In_64,In_988);
or U3084 (N_3084,In_692,In_511);
nor U3085 (N_3085,In_1,In_680);
xnor U3086 (N_3086,In_954,In_766);
nor U3087 (N_3087,In_684,In_290);
and U3088 (N_3088,In_259,In_170);
and U3089 (N_3089,In_963,In_240);
and U3090 (N_3090,In_964,In_797);
xor U3091 (N_3091,In_190,In_458);
and U3092 (N_3092,In_954,In_4);
and U3093 (N_3093,In_450,In_144);
xnor U3094 (N_3094,In_241,In_86);
and U3095 (N_3095,In_605,In_757);
and U3096 (N_3096,In_295,In_461);
or U3097 (N_3097,In_345,In_536);
xor U3098 (N_3098,In_986,In_668);
nand U3099 (N_3099,In_645,In_519);
and U3100 (N_3100,In_518,In_32);
nor U3101 (N_3101,In_632,In_887);
nor U3102 (N_3102,In_415,In_512);
nor U3103 (N_3103,In_439,In_197);
or U3104 (N_3104,In_545,In_993);
nor U3105 (N_3105,In_846,In_831);
and U3106 (N_3106,In_446,In_904);
or U3107 (N_3107,In_49,In_299);
nor U3108 (N_3108,In_573,In_9);
nor U3109 (N_3109,In_654,In_833);
nor U3110 (N_3110,In_254,In_4);
and U3111 (N_3111,In_43,In_118);
or U3112 (N_3112,In_271,In_505);
nor U3113 (N_3113,In_311,In_658);
or U3114 (N_3114,In_278,In_259);
nor U3115 (N_3115,In_511,In_135);
nand U3116 (N_3116,In_809,In_406);
or U3117 (N_3117,In_735,In_427);
nor U3118 (N_3118,In_942,In_955);
or U3119 (N_3119,In_467,In_457);
and U3120 (N_3120,In_126,In_29);
nor U3121 (N_3121,In_553,In_924);
and U3122 (N_3122,In_310,In_674);
nor U3123 (N_3123,In_29,In_633);
and U3124 (N_3124,In_294,In_29);
and U3125 (N_3125,In_674,In_963);
nor U3126 (N_3126,In_597,In_228);
nor U3127 (N_3127,In_138,In_543);
nor U3128 (N_3128,In_764,In_650);
nand U3129 (N_3129,In_483,In_121);
or U3130 (N_3130,In_435,In_494);
or U3131 (N_3131,In_926,In_721);
or U3132 (N_3132,In_657,In_780);
and U3133 (N_3133,In_365,In_119);
and U3134 (N_3134,In_375,In_834);
and U3135 (N_3135,In_119,In_944);
nor U3136 (N_3136,In_557,In_499);
or U3137 (N_3137,In_368,In_92);
and U3138 (N_3138,In_291,In_66);
nand U3139 (N_3139,In_252,In_92);
nor U3140 (N_3140,In_844,In_114);
nor U3141 (N_3141,In_597,In_554);
or U3142 (N_3142,In_896,In_708);
xor U3143 (N_3143,In_592,In_982);
nand U3144 (N_3144,In_404,In_797);
xnor U3145 (N_3145,In_136,In_474);
nand U3146 (N_3146,In_914,In_465);
nor U3147 (N_3147,In_311,In_711);
nor U3148 (N_3148,In_55,In_142);
or U3149 (N_3149,In_876,In_790);
nor U3150 (N_3150,In_20,In_873);
and U3151 (N_3151,In_23,In_956);
nand U3152 (N_3152,In_685,In_519);
nor U3153 (N_3153,In_125,In_58);
xor U3154 (N_3154,In_378,In_875);
nand U3155 (N_3155,In_770,In_250);
and U3156 (N_3156,In_670,In_559);
nand U3157 (N_3157,In_565,In_685);
nand U3158 (N_3158,In_555,In_280);
or U3159 (N_3159,In_903,In_934);
nor U3160 (N_3160,In_972,In_574);
nand U3161 (N_3161,In_45,In_707);
or U3162 (N_3162,In_476,In_379);
or U3163 (N_3163,In_785,In_507);
and U3164 (N_3164,In_458,In_943);
nand U3165 (N_3165,In_691,In_218);
nand U3166 (N_3166,In_23,In_919);
and U3167 (N_3167,In_173,In_236);
nor U3168 (N_3168,In_210,In_939);
and U3169 (N_3169,In_498,In_878);
or U3170 (N_3170,In_686,In_227);
and U3171 (N_3171,In_911,In_942);
nor U3172 (N_3172,In_71,In_530);
nand U3173 (N_3173,In_868,In_138);
or U3174 (N_3174,In_43,In_264);
nor U3175 (N_3175,In_149,In_632);
or U3176 (N_3176,In_741,In_16);
nor U3177 (N_3177,In_746,In_511);
and U3178 (N_3178,In_501,In_969);
nor U3179 (N_3179,In_712,In_414);
nand U3180 (N_3180,In_926,In_63);
nor U3181 (N_3181,In_524,In_538);
and U3182 (N_3182,In_588,In_809);
and U3183 (N_3183,In_287,In_663);
and U3184 (N_3184,In_691,In_450);
nand U3185 (N_3185,In_656,In_529);
nand U3186 (N_3186,In_376,In_584);
xnor U3187 (N_3187,In_34,In_291);
nand U3188 (N_3188,In_924,In_802);
nand U3189 (N_3189,In_23,In_150);
nand U3190 (N_3190,In_570,In_899);
nor U3191 (N_3191,In_680,In_610);
or U3192 (N_3192,In_347,In_917);
and U3193 (N_3193,In_59,In_175);
and U3194 (N_3194,In_503,In_847);
nor U3195 (N_3195,In_129,In_7);
nand U3196 (N_3196,In_809,In_933);
and U3197 (N_3197,In_205,In_202);
and U3198 (N_3198,In_871,In_850);
nor U3199 (N_3199,In_335,In_849);
or U3200 (N_3200,In_118,In_851);
and U3201 (N_3201,In_801,In_579);
or U3202 (N_3202,In_778,In_23);
nand U3203 (N_3203,In_74,In_618);
and U3204 (N_3204,In_132,In_683);
nor U3205 (N_3205,In_756,In_246);
nand U3206 (N_3206,In_813,In_336);
or U3207 (N_3207,In_566,In_456);
nand U3208 (N_3208,In_74,In_85);
nor U3209 (N_3209,In_908,In_156);
nand U3210 (N_3210,In_321,In_440);
nand U3211 (N_3211,In_55,In_195);
nor U3212 (N_3212,In_814,In_564);
nand U3213 (N_3213,In_483,In_704);
nand U3214 (N_3214,In_456,In_304);
nand U3215 (N_3215,In_39,In_608);
or U3216 (N_3216,In_139,In_779);
or U3217 (N_3217,In_624,In_171);
nand U3218 (N_3218,In_614,In_907);
or U3219 (N_3219,In_722,In_561);
or U3220 (N_3220,In_560,In_321);
nor U3221 (N_3221,In_566,In_291);
nor U3222 (N_3222,In_987,In_905);
nand U3223 (N_3223,In_315,In_776);
nand U3224 (N_3224,In_973,In_655);
nor U3225 (N_3225,In_681,In_462);
or U3226 (N_3226,In_419,In_817);
xor U3227 (N_3227,In_339,In_955);
and U3228 (N_3228,In_63,In_444);
nand U3229 (N_3229,In_366,In_362);
xnor U3230 (N_3230,In_186,In_292);
and U3231 (N_3231,In_308,In_639);
xor U3232 (N_3232,In_619,In_216);
nor U3233 (N_3233,In_748,In_8);
nand U3234 (N_3234,In_392,In_469);
nand U3235 (N_3235,In_217,In_342);
and U3236 (N_3236,In_703,In_614);
or U3237 (N_3237,In_425,In_121);
nor U3238 (N_3238,In_837,In_810);
nand U3239 (N_3239,In_718,In_582);
nand U3240 (N_3240,In_725,In_835);
xnor U3241 (N_3241,In_914,In_198);
nand U3242 (N_3242,In_559,In_456);
and U3243 (N_3243,In_10,In_318);
nand U3244 (N_3244,In_211,In_379);
and U3245 (N_3245,In_665,In_24);
and U3246 (N_3246,In_763,In_38);
nor U3247 (N_3247,In_294,In_183);
and U3248 (N_3248,In_655,In_158);
nor U3249 (N_3249,In_268,In_699);
nor U3250 (N_3250,In_238,In_23);
nand U3251 (N_3251,In_55,In_43);
nand U3252 (N_3252,In_839,In_126);
and U3253 (N_3253,In_644,In_655);
nand U3254 (N_3254,In_992,In_751);
xor U3255 (N_3255,In_62,In_604);
nand U3256 (N_3256,In_403,In_753);
or U3257 (N_3257,In_499,In_43);
and U3258 (N_3258,In_928,In_40);
or U3259 (N_3259,In_309,In_802);
or U3260 (N_3260,In_360,In_985);
nand U3261 (N_3261,In_886,In_107);
or U3262 (N_3262,In_624,In_549);
and U3263 (N_3263,In_447,In_65);
or U3264 (N_3264,In_295,In_851);
and U3265 (N_3265,In_25,In_772);
nand U3266 (N_3266,In_349,In_601);
nor U3267 (N_3267,In_849,In_119);
or U3268 (N_3268,In_10,In_116);
or U3269 (N_3269,In_628,In_136);
nor U3270 (N_3270,In_170,In_290);
and U3271 (N_3271,In_797,In_180);
or U3272 (N_3272,In_892,In_275);
or U3273 (N_3273,In_280,In_375);
or U3274 (N_3274,In_162,In_625);
or U3275 (N_3275,In_393,In_660);
nor U3276 (N_3276,In_209,In_985);
and U3277 (N_3277,In_113,In_403);
nand U3278 (N_3278,In_781,In_486);
and U3279 (N_3279,In_543,In_544);
nor U3280 (N_3280,In_933,In_484);
and U3281 (N_3281,In_829,In_667);
nand U3282 (N_3282,In_164,In_361);
nand U3283 (N_3283,In_542,In_462);
and U3284 (N_3284,In_776,In_306);
nand U3285 (N_3285,In_130,In_502);
or U3286 (N_3286,In_870,In_159);
nor U3287 (N_3287,In_123,In_782);
nand U3288 (N_3288,In_119,In_874);
nand U3289 (N_3289,In_320,In_272);
or U3290 (N_3290,In_333,In_472);
and U3291 (N_3291,In_726,In_346);
or U3292 (N_3292,In_839,In_125);
nor U3293 (N_3293,In_531,In_505);
and U3294 (N_3294,In_178,In_670);
and U3295 (N_3295,In_953,In_554);
and U3296 (N_3296,In_342,In_632);
nor U3297 (N_3297,In_193,In_446);
nand U3298 (N_3298,In_941,In_132);
nand U3299 (N_3299,In_67,In_419);
nor U3300 (N_3300,In_549,In_690);
nor U3301 (N_3301,In_353,In_526);
or U3302 (N_3302,In_555,In_735);
nand U3303 (N_3303,In_934,In_423);
or U3304 (N_3304,In_203,In_444);
nor U3305 (N_3305,In_415,In_227);
and U3306 (N_3306,In_815,In_583);
nand U3307 (N_3307,In_745,In_918);
or U3308 (N_3308,In_431,In_728);
nand U3309 (N_3309,In_470,In_523);
nand U3310 (N_3310,In_979,In_999);
and U3311 (N_3311,In_995,In_143);
nand U3312 (N_3312,In_558,In_689);
nor U3313 (N_3313,In_248,In_330);
and U3314 (N_3314,In_762,In_567);
nand U3315 (N_3315,In_915,In_91);
nor U3316 (N_3316,In_315,In_163);
nand U3317 (N_3317,In_897,In_440);
nand U3318 (N_3318,In_81,In_553);
nor U3319 (N_3319,In_222,In_441);
or U3320 (N_3320,In_206,In_112);
and U3321 (N_3321,In_22,In_38);
and U3322 (N_3322,In_827,In_849);
or U3323 (N_3323,In_100,In_886);
nor U3324 (N_3324,In_517,In_459);
and U3325 (N_3325,In_472,In_949);
nand U3326 (N_3326,In_371,In_73);
and U3327 (N_3327,In_780,In_684);
or U3328 (N_3328,In_123,In_50);
or U3329 (N_3329,In_294,In_456);
or U3330 (N_3330,In_943,In_852);
xnor U3331 (N_3331,In_470,In_225);
and U3332 (N_3332,In_256,In_745);
or U3333 (N_3333,In_613,In_554);
nand U3334 (N_3334,In_857,In_107);
or U3335 (N_3335,In_46,In_641);
and U3336 (N_3336,In_970,In_587);
nor U3337 (N_3337,In_598,In_624);
nor U3338 (N_3338,In_879,In_719);
nand U3339 (N_3339,In_956,In_80);
nor U3340 (N_3340,In_141,In_772);
nor U3341 (N_3341,In_364,In_858);
and U3342 (N_3342,In_47,In_862);
nor U3343 (N_3343,In_89,In_279);
and U3344 (N_3344,In_414,In_945);
and U3345 (N_3345,In_426,In_836);
nand U3346 (N_3346,In_687,In_736);
or U3347 (N_3347,In_579,In_396);
nand U3348 (N_3348,In_213,In_994);
xor U3349 (N_3349,In_79,In_946);
nand U3350 (N_3350,In_932,In_314);
xor U3351 (N_3351,In_176,In_430);
nand U3352 (N_3352,In_898,In_890);
or U3353 (N_3353,In_986,In_756);
nand U3354 (N_3354,In_818,In_127);
or U3355 (N_3355,In_7,In_783);
nand U3356 (N_3356,In_647,In_738);
nor U3357 (N_3357,In_299,In_787);
or U3358 (N_3358,In_817,In_813);
and U3359 (N_3359,In_758,In_698);
or U3360 (N_3360,In_13,In_459);
and U3361 (N_3361,In_427,In_776);
nor U3362 (N_3362,In_271,In_872);
or U3363 (N_3363,In_675,In_26);
or U3364 (N_3364,In_802,In_456);
or U3365 (N_3365,In_146,In_421);
nand U3366 (N_3366,In_482,In_834);
nor U3367 (N_3367,In_400,In_602);
or U3368 (N_3368,In_834,In_690);
and U3369 (N_3369,In_185,In_647);
or U3370 (N_3370,In_924,In_642);
or U3371 (N_3371,In_388,In_68);
or U3372 (N_3372,In_943,In_665);
nor U3373 (N_3373,In_917,In_380);
nor U3374 (N_3374,In_322,In_972);
or U3375 (N_3375,In_439,In_435);
or U3376 (N_3376,In_49,In_393);
nand U3377 (N_3377,In_371,In_807);
nor U3378 (N_3378,In_382,In_808);
nand U3379 (N_3379,In_134,In_671);
nor U3380 (N_3380,In_747,In_867);
nand U3381 (N_3381,In_925,In_584);
and U3382 (N_3382,In_676,In_148);
nor U3383 (N_3383,In_747,In_956);
or U3384 (N_3384,In_618,In_751);
and U3385 (N_3385,In_716,In_27);
or U3386 (N_3386,In_449,In_345);
nor U3387 (N_3387,In_952,In_573);
nand U3388 (N_3388,In_56,In_701);
nor U3389 (N_3389,In_165,In_206);
nand U3390 (N_3390,In_114,In_348);
nand U3391 (N_3391,In_473,In_221);
or U3392 (N_3392,In_515,In_59);
or U3393 (N_3393,In_284,In_728);
nor U3394 (N_3394,In_381,In_50);
and U3395 (N_3395,In_408,In_349);
or U3396 (N_3396,In_994,In_70);
nor U3397 (N_3397,In_827,In_150);
or U3398 (N_3398,In_91,In_47);
and U3399 (N_3399,In_978,In_76);
nand U3400 (N_3400,In_314,In_190);
nor U3401 (N_3401,In_392,In_430);
or U3402 (N_3402,In_347,In_967);
or U3403 (N_3403,In_75,In_585);
and U3404 (N_3404,In_196,In_214);
nand U3405 (N_3405,In_158,In_339);
or U3406 (N_3406,In_243,In_771);
nor U3407 (N_3407,In_902,In_433);
nor U3408 (N_3408,In_10,In_359);
nand U3409 (N_3409,In_60,In_948);
nand U3410 (N_3410,In_421,In_42);
or U3411 (N_3411,In_972,In_684);
nor U3412 (N_3412,In_168,In_39);
or U3413 (N_3413,In_383,In_534);
nand U3414 (N_3414,In_505,In_139);
nor U3415 (N_3415,In_695,In_595);
and U3416 (N_3416,In_424,In_262);
or U3417 (N_3417,In_251,In_393);
nand U3418 (N_3418,In_801,In_901);
and U3419 (N_3419,In_486,In_532);
nor U3420 (N_3420,In_650,In_514);
or U3421 (N_3421,In_332,In_869);
and U3422 (N_3422,In_918,In_282);
or U3423 (N_3423,In_844,In_324);
nand U3424 (N_3424,In_788,In_227);
and U3425 (N_3425,In_170,In_343);
or U3426 (N_3426,In_311,In_293);
or U3427 (N_3427,In_916,In_512);
nor U3428 (N_3428,In_785,In_612);
nor U3429 (N_3429,In_244,In_105);
and U3430 (N_3430,In_407,In_890);
nand U3431 (N_3431,In_719,In_951);
or U3432 (N_3432,In_761,In_900);
and U3433 (N_3433,In_593,In_209);
nor U3434 (N_3434,In_961,In_870);
or U3435 (N_3435,In_750,In_225);
xnor U3436 (N_3436,In_436,In_201);
xnor U3437 (N_3437,In_205,In_195);
nand U3438 (N_3438,In_4,In_317);
or U3439 (N_3439,In_951,In_914);
and U3440 (N_3440,In_91,In_399);
nor U3441 (N_3441,In_290,In_401);
or U3442 (N_3442,In_957,In_723);
or U3443 (N_3443,In_465,In_333);
and U3444 (N_3444,In_123,In_262);
and U3445 (N_3445,In_386,In_896);
nand U3446 (N_3446,In_265,In_180);
nor U3447 (N_3447,In_931,In_372);
nand U3448 (N_3448,In_605,In_844);
nand U3449 (N_3449,In_69,In_132);
and U3450 (N_3450,In_257,In_203);
nor U3451 (N_3451,In_384,In_207);
nand U3452 (N_3452,In_451,In_266);
and U3453 (N_3453,In_682,In_669);
and U3454 (N_3454,In_405,In_749);
nand U3455 (N_3455,In_437,In_278);
and U3456 (N_3456,In_594,In_474);
nor U3457 (N_3457,In_267,In_796);
nor U3458 (N_3458,In_441,In_61);
or U3459 (N_3459,In_952,In_185);
and U3460 (N_3460,In_374,In_940);
nand U3461 (N_3461,In_870,In_992);
nand U3462 (N_3462,In_787,In_325);
nand U3463 (N_3463,In_999,In_706);
or U3464 (N_3464,In_630,In_668);
nor U3465 (N_3465,In_516,In_781);
nand U3466 (N_3466,In_341,In_307);
nor U3467 (N_3467,In_658,In_118);
and U3468 (N_3468,In_281,In_716);
or U3469 (N_3469,In_793,In_874);
and U3470 (N_3470,In_201,In_829);
nand U3471 (N_3471,In_179,In_2);
or U3472 (N_3472,In_873,In_961);
nand U3473 (N_3473,In_855,In_87);
and U3474 (N_3474,In_988,In_440);
nor U3475 (N_3475,In_398,In_348);
or U3476 (N_3476,In_691,In_795);
xnor U3477 (N_3477,In_573,In_988);
nand U3478 (N_3478,In_919,In_329);
nand U3479 (N_3479,In_791,In_335);
nor U3480 (N_3480,In_730,In_668);
or U3481 (N_3481,In_86,In_531);
xnor U3482 (N_3482,In_590,In_131);
nor U3483 (N_3483,In_72,In_380);
and U3484 (N_3484,In_110,In_387);
nor U3485 (N_3485,In_527,In_537);
nor U3486 (N_3486,In_617,In_440);
nor U3487 (N_3487,In_109,In_621);
and U3488 (N_3488,In_699,In_886);
nor U3489 (N_3489,In_21,In_728);
nor U3490 (N_3490,In_439,In_480);
nor U3491 (N_3491,In_263,In_538);
or U3492 (N_3492,In_365,In_183);
or U3493 (N_3493,In_405,In_446);
nand U3494 (N_3494,In_287,In_199);
nor U3495 (N_3495,In_906,In_8);
or U3496 (N_3496,In_64,In_248);
or U3497 (N_3497,In_355,In_271);
or U3498 (N_3498,In_998,In_860);
nand U3499 (N_3499,In_343,In_945);
and U3500 (N_3500,In_210,In_308);
nor U3501 (N_3501,In_320,In_862);
or U3502 (N_3502,In_552,In_671);
nand U3503 (N_3503,In_211,In_346);
nand U3504 (N_3504,In_311,In_368);
and U3505 (N_3505,In_371,In_297);
nor U3506 (N_3506,In_863,In_443);
or U3507 (N_3507,In_1,In_294);
and U3508 (N_3508,In_81,In_474);
nor U3509 (N_3509,In_461,In_850);
and U3510 (N_3510,In_552,In_430);
or U3511 (N_3511,In_705,In_993);
nor U3512 (N_3512,In_536,In_850);
nor U3513 (N_3513,In_958,In_932);
and U3514 (N_3514,In_728,In_94);
or U3515 (N_3515,In_760,In_673);
nand U3516 (N_3516,In_740,In_251);
and U3517 (N_3517,In_774,In_967);
or U3518 (N_3518,In_655,In_82);
and U3519 (N_3519,In_891,In_408);
nor U3520 (N_3520,In_396,In_994);
and U3521 (N_3521,In_452,In_450);
or U3522 (N_3522,In_23,In_724);
or U3523 (N_3523,In_669,In_212);
and U3524 (N_3524,In_391,In_604);
or U3525 (N_3525,In_304,In_319);
and U3526 (N_3526,In_893,In_864);
nand U3527 (N_3527,In_749,In_598);
nor U3528 (N_3528,In_293,In_802);
xor U3529 (N_3529,In_241,In_627);
or U3530 (N_3530,In_833,In_538);
nor U3531 (N_3531,In_755,In_575);
and U3532 (N_3532,In_931,In_446);
and U3533 (N_3533,In_204,In_293);
xnor U3534 (N_3534,In_205,In_937);
nand U3535 (N_3535,In_97,In_247);
nand U3536 (N_3536,In_237,In_764);
nand U3537 (N_3537,In_173,In_10);
nand U3538 (N_3538,In_562,In_134);
nor U3539 (N_3539,In_700,In_461);
nor U3540 (N_3540,In_662,In_416);
nor U3541 (N_3541,In_118,In_222);
nor U3542 (N_3542,In_280,In_632);
nor U3543 (N_3543,In_628,In_202);
and U3544 (N_3544,In_207,In_939);
and U3545 (N_3545,In_713,In_441);
and U3546 (N_3546,In_842,In_789);
nor U3547 (N_3547,In_985,In_40);
nand U3548 (N_3548,In_226,In_530);
xnor U3549 (N_3549,In_606,In_610);
and U3550 (N_3550,In_607,In_495);
or U3551 (N_3551,In_274,In_389);
nor U3552 (N_3552,In_477,In_911);
nand U3553 (N_3553,In_47,In_628);
or U3554 (N_3554,In_375,In_709);
or U3555 (N_3555,In_727,In_445);
nor U3556 (N_3556,In_292,In_236);
and U3557 (N_3557,In_54,In_503);
and U3558 (N_3558,In_10,In_376);
nor U3559 (N_3559,In_683,In_191);
or U3560 (N_3560,In_579,In_357);
or U3561 (N_3561,In_263,In_647);
and U3562 (N_3562,In_625,In_620);
nor U3563 (N_3563,In_925,In_574);
or U3564 (N_3564,In_147,In_452);
nand U3565 (N_3565,In_359,In_578);
nor U3566 (N_3566,In_977,In_690);
nand U3567 (N_3567,In_150,In_669);
or U3568 (N_3568,In_918,In_311);
nand U3569 (N_3569,In_515,In_835);
and U3570 (N_3570,In_764,In_57);
and U3571 (N_3571,In_505,In_709);
or U3572 (N_3572,In_442,In_292);
and U3573 (N_3573,In_716,In_551);
nor U3574 (N_3574,In_427,In_255);
nor U3575 (N_3575,In_608,In_261);
nand U3576 (N_3576,In_944,In_982);
or U3577 (N_3577,In_623,In_4);
nand U3578 (N_3578,In_642,In_204);
nor U3579 (N_3579,In_338,In_470);
or U3580 (N_3580,In_423,In_195);
and U3581 (N_3581,In_26,In_620);
and U3582 (N_3582,In_907,In_898);
or U3583 (N_3583,In_956,In_13);
or U3584 (N_3584,In_95,In_70);
or U3585 (N_3585,In_862,In_821);
nand U3586 (N_3586,In_646,In_362);
nand U3587 (N_3587,In_688,In_75);
nor U3588 (N_3588,In_431,In_142);
and U3589 (N_3589,In_363,In_517);
nand U3590 (N_3590,In_597,In_941);
nor U3591 (N_3591,In_478,In_179);
and U3592 (N_3592,In_477,In_986);
or U3593 (N_3593,In_113,In_500);
or U3594 (N_3594,In_79,In_793);
nor U3595 (N_3595,In_216,In_212);
xor U3596 (N_3596,In_108,In_586);
nor U3597 (N_3597,In_875,In_474);
xor U3598 (N_3598,In_319,In_678);
and U3599 (N_3599,In_969,In_543);
nand U3600 (N_3600,In_222,In_376);
nand U3601 (N_3601,In_868,In_618);
and U3602 (N_3602,In_791,In_737);
and U3603 (N_3603,In_489,In_25);
and U3604 (N_3604,In_67,In_763);
and U3605 (N_3605,In_22,In_506);
nand U3606 (N_3606,In_749,In_977);
nand U3607 (N_3607,In_792,In_945);
nand U3608 (N_3608,In_618,In_175);
and U3609 (N_3609,In_136,In_821);
or U3610 (N_3610,In_52,In_104);
or U3611 (N_3611,In_779,In_939);
or U3612 (N_3612,In_89,In_8);
xnor U3613 (N_3613,In_188,In_894);
nand U3614 (N_3614,In_988,In_995);
and U3615 (N_3615,In_884,In_716);
and U3616 (N_3616,In_858,In_328);
nor U3617 (N_3617,In_563,In_189);
nand U3618 (N_3618,In_945,In_651);
nand U3619 (N_3619,In_909,In_970);
nor U3620 (N_3620,In_181,In_542);
or U3621 (N_3621,In_657,In_821);
nand U3622 (N_3622,In_966,In_187);
nor U3623 (N_3623,In_847,In_425);
nand U3624 (N_3624,In_689,In_302);
nor U3625 (N_3625,In_928,In_461);
and U3626 (N_3626,In_580,In_537);
nor U3627 (N_3627,In_971,In_748);
nor U3628 (N_3628,In_433,In_99);
or U3629 (N_3629,In_97,In_936);
nor U3630 (N_3630,In_352,In_866);
nor U3631 (N_3631,In_376,In_939);
nor U3632 (N_3632,In_954,In_596);
nand U3633 (N_3633,In_556,In_505);
nand U3634 (N_3634,In_179,In_922);
and U3635 (N_3635,In_965,In_55);
nand U3636 (N_3636,In_785,In_445);
and U3637 (N_3637,In_772,In_928);
or U3638 (N_3638,In_132,In_514);
or U3639 (N_3639,In_313,In_493);
nand U3640 (N_3640,In_861,In_200);
and U3641 (N_3641,In_617,In_140);
and U3642 (N_3642,In_250,In_965);
nand U3643 (N_3643,In_179,In_403);
nand U3644 (N_3644,In_990,In_610);
nor U3645 (N_3645,In_839,In_232);
and U3646 (N_3646,In_585,In_531);
nand U3647 (N_3647,In_414,In_709);
and U3648 (N_3648,In_172,In_567);
nand U3649 (N_3649,In_975,In_363);
nand U3650 (N_3650,In_83,In_657);
xor U3651 (N_3651,In_203,In_786);
and U3652 (N_3652,In_962,In_371);
nand U3653 (N_3653,In_843,In_766);
nor U3654 (N_3654,In_800,In_129);
or U3655 (N_3655,In_968,In_691);
nand U3656 (N_3656,In_977,In_464);
nor U3657 (N_3657,In_897,In_352);
nand U3658 (N_3658,In_776,In_945);
nand U3659 (N_3659,In_972,In_854);
nor U3660 (N_3660,In_693,In_833);
and U3661 (N_3661,In_656,In_444);
nor U3662 (N_3662,In_311,In_401);
nand U3663 (N_3663,In_732,In_772);
and U3664 (N_3664,In_49,In_757);
and U3665 (N_3665,In_835,In_529);
nor U3666 (N_3666,In_588,In_204);
or U3667 (N_3667,In_599,In_774);
and U3668 (N_3668,In_519,In_885);
nand U3669 (N_3669,In_803,In_346);
or U3670 (N_3670,In_200,In_77);
or U3671 (N_3671,In_896,In_489);
and U3672 (N_3672,In_840,In_830);
nor U3673 (N_3673,In_459,In_804);
or U3674 (N_3674,In_849,In_316);
and U3675 (N_3675,In_608,In_231);
and U3676 (N_3676,In_42,In_373);
and U3677 (N_3677,In_774,In_597);
nor U3678 (N_3678,In_704,In_211);
nor U3679 (N_3679,In_430,In_740);
nor U3680 (N_3680,In_269,In_73);
nor U3681 (N_3681,In_351,In_959);
or U3682 (N_3682,In_809,In_220);
and U3683 (N_3683,In_684,In_83);
nor U3684 (N_3684,In_998,In_943);
or U3685 (N_3685,In_542,In_879);
or U3686 (N_3686,In_635,In_290);
xor U3687 (N_3687,In_65,In_803);
nor U3688 (N_3688,In_445,In_32);
and U3689 (N_3689,In_261,In_644);
nor U3690 (N_3690,In_930,In_571);
or U3691 (N_3691,In_298,In_172);
or U3692 (N_3692,In_767,In_594);
or U3693 (N_3693,In_607,In_781);
or U3694 (N_3694,In_58,In_462);
or U3695 (N_3695,In_309,In_648);
nand U3696 (N_3696,In_900,In_106);
or U3697 (N_3697,In_589,In_198);
nand U3698 (N_3698,In_908,In_295);
nand U3699 (N_3699,In_436,In_335);
or U3700 (N_3700,In_33,In_970);
and U3701 (N_3701,In_523,In_995);
nand U3702 (N_3702,In_638,In_769);
nand U3703 (N_3703,In_549,In_960);
nand U3704 (N_3704,In_732,In_157);
and U3705 (N_3705,In_538,In_726);
and U3706 (N_3706,In_285,In_369);
and U3707 (N_3707,In_583,In_91);
or U3708 (N_3708,In_840,In_586);
nor U3709 (N_3709,In_83,In_84);
nand U3710 (N_3710,In_312,In_791);
nor U3711 (N_3711,In_253,In_882);
nor U3712 (N_3712,In_970,In_695);
nand U3713 (N_3713,In_783,In_133);
nor U3714 (N_3714,In_405,In_360);
nand U3715 (N_3715,In_662,In_120);
nand U3716 (N_3716,In_385,In_857);
and U3717 (N_3717,In_916,In_47);
nand U3718 (N_3718,In_949,In_797);
nor U3719 (N_3719,In_789,In_427);
nand U3720 (N_3720,In_107,In_368);
and U3721 (N_3721,In_286,In_410);
nor U3722 (N_3722,In_366,In_508);
and U3723 (N_3723,In_500,In_362);
or U3724 (N_3724,In_192,In_188);
and U3725 (N_3725,In_71,In_672);
and U3726 (N_3726,In_30,In_49);
nor U3727 (N_3727,In_315,In_904);
or U3728 (N_3728,In_77,In_482);
nor U3729 (N_3729,In_636,In_555);
and U3730 (N_3730,In_622,In_181);
nor U3731 (N_3731,In_877,In_558);
nor U3732 (N_3732,In_399,In_974);
nor U3733 (N_3733,In_353,In_619);
or U3734 (N_3734,In_824,In_996);
or U3735 (N_3735,In_669,In_553);
nand U3736 (N_3736,In_814,In_33);
and U3737 (N_3737,In_968,In_494);
nor U3738 (N_3738,In_368,In_843);
nor U3739 (N_3739,In_484,In_952);
and U3740 (N_3740,In_744,In_466);
and U3741 (N_3741,In_862,In_698);
or U3742 (N_3742,In_451,In_150);
nor U3743 (N_3743,In_420,In_116);
nor U3744 (N_3744,In_392,In_526);
or U3745 (N_3745,In_545,In_427);
and U3746 (N_3746,In_590,In_866);
or U3747 (N_3747,In_19,In_885);
nor U3748 (N_3748,In_713,In_14);
and U3749 (N_3749,In_871,In_106);
nor U3750 (N_3750,In_236,In_504);
and U3751 (N_3751,In_394,In_61);
and U3752 (N_3752,In_116,In_868);
or U3753 (N_3753,In_336,In_339);
nand U3754 (N_3754,In_378,In_539);
nor U3755 (N_3755,In_710,In_800);
or U3756 (N_3756,In_929,In_706);
and U3757 (N_3757,In_246,In_57);
nor U3758 (N_3758,In_868,In_662);
and U3759 (N_3759,In_53,In_781);
nor U3760 (N_3760,In_672,In_271);
nand U3761 (N_3761,In_716,In_0);
nand U3762 (N_3762,In_375,In_785);
or U3763 (N_3763,In_700,In_638);
nor U3764 (N_3764,In_872,In_730);
and U3765 (N_3765,In_423,In_756);
and U3766 (N_3766,In_678,In_776);
nand U3767 (N_3767,In_226,In_690);
nor U3768 (N_3768,In_934,In_763);
or U3769 (N_3769,In_397,In_179);
or U3770 (N_3770,In_784,In_595);
or U3771 (N_3771,In_130,In_960);
nand U3772 (N_3772,In_51,In_388);
nand U3773 (N_3773,In_415,In_626);
nand U3774 (N_3774,In_597,In_863);
and U3775 (N_3775,In_504,In_912);
nor U3776 (N_3776,In_167,In_97);
nor U3777 (N_3777,In_357,In_476);
nand U3778 (N_3778,In_463,In_244);
or U3779 (N_3779,In_565,In_615);
nand U3780 (N_3780,In_843,In_184);
nand U3781 (N_3781,In_585,In_778);
and U3782 (N_3782,In_6,In_707);
nand U3783 (N_3783,In_431,In_959);
or U3784 (N_3784,In_913,In_931);
nand U3785 (N_3785,In_393,In_128);
and U3786 (N_3786,In_120,In_714);
nor U3787 (N_3787,In_482,In_746);
and U3788 (N_3788,In_48,In_391);
nand U3789 (N_3789,In_459,In_395);
nand U3790 (N_3790,In_686,In_900);
nand U3791 (N_3791,In_390,In_307);
or U3792 (N_3792,In_789,In_164);
or U3793 (N_3793,In_396,In_801);
and U3794 (N_3794,In_225,In_520);
or U3795 (N_3795,In_808,In_658);
and U3796 (N_3796,In_484,In_349);
or U3797 (N_3797,In_443,In_906);
or U3798 (N_3798,In_867,In_574);
xnor U3799 (N_3799,In_753,In_806);
nor U3800 (N_3800,In_934,In_384);
nor U3801 (N_3801,In_252,In_550);
nand U3802 (N_3802,In_83,In_592);
nor U3803 (N_3803,In_307,In_768);
and U3804 (N_3804,In_11,In_101);
or U3805 (N_3805,In_102,In_720);
nor U3806 (N_3806,In_260,In_52);
or U3807 (N_3807,In_519,In_810);
or U3808 (N_3808,In_163,In_800);
nor U3809 (N_3809,In_102,In_850);
nor U3810 (N_3810,In_954,In_143);
nand U3811 (N_3811,In_857,In_279);
and U3812 (N_3812,In_497,In_617);
or U3813 (N_3813,In_651,In_146);
nand U3814 (N_3814,In_840,In_735);
or U3815 (N_3815,In_456,In_549);
and U3816 (N_3816,In_22,In_64);
nand U3817 (N_3817,In_771,In_636);
and U3818 (N_3818,In_668,In_553);
or U3819 (N_3819,In_909,In_485);
or U3820 (N_3820,In_602,In_898);
and U3821 (N_3821,In_206,In_874);
nand U3822 (N_3822,In_192,In_534);
nand U3823 (N_3823,In_106,In_426);
or U3824 (N_3824,In_629,In_351);
and U3825 (N_3825,In_902,In_889);
nor U3826 (N_3826,In_16,In_385);
and U3827 (N_3827,In_825,In_983);
nor U3828 (N_3828,In_660,In_147);
nand U3829 (N_3829,In_618,In_160);
or U3830 (N_3830,In_730,In_679);
nor U3831 (N_3831,In_575,In_159);
or U3832 (N_3832,In_503,In_386);
or U3833 (N_3833,In_61,In_926);
or U3834 (N_3834,In_361,In_263);
nor U3835 (N_3835,In_20,In_12);
and U3836 (N_3836,In_56,In_820);
nor U3837 (N_3837,In_55,In_22);
nand U3838 (N_3838,In_760,In_657);
or U3839 (N_3839,In_838,In_890);
or U3840 (N_3840,In_255,In_64);
nor U3841 (N_3841,In_740,In_709);
or U3842 (N_3842,In_921,In_410);
and U3843 (N_3843,In_484,In_328);
nand U3844 (N_3844,In_151,In_809);
nor U3845 (N_3845,In_259,In_584);
nor U3846 (N_3846,In_679,In_503);
or U3847 (N_3847,In_583,In_930);
nand U3848 (N_3848,In_124,In_533);
nand U3849 (N_3849,In_478,In_594);
or U3850 (N_3850,In_131,In_192);
nor U3851 (N_3851,In_639,In_83);
nor U3852 (N_3852,In_247,In_671);
xor U3853 (N_3853,In_863,In_445);
nand U3854 (N_3854,In_725,In_135);
and U3855 (N_3855,In_735,In_63);
nor U3856 (N_3856,In_669,In_548);
or U3857 (N_3857,In_156,In_153);
nand U3858 (N_3858,In_972,In_325);
and U3859 (N_3859,In_68,In_188);
nand U3860 (N_3860,In_892,In_276);
or U3861 (N_3861,In_358,In_823);
nor U3862 (N_3862,In_350,In_301);
nor U3863 (N_3863,In_658,In_711);
nor U3864 (N_3864,In_536,In_199);
nand U3865 (N_3865,In_848,In_924);
nand U3866 (N_3866,In_722,In_718);
or U3867 (N_3867,In_507,In_646);
nand U3868 (N_3868,In_129,In_794);
or U3869 (N_3869,In_30,In_565);
and U3870 (N_3870,In_801,In_872);
or U3871 (N_3871,In_725,In_986);
or U3872 (N_3872,In_464,In_818);
nor U3873 (N_3873,In_898,In_875);
or U3874 (N_3874,In_408,In_338);
nor U3875 (N_3875,In_608,In_241);
nor U3876 (N_3876,In_148,In_252);
nor U3877 (N_3877,In_809,In_365);
nand U3878 (N_3878,In_774,In_173);
nand U3879 (N_3879,In_326,In_364);
and U3880 (N_3880,In_764,In_934);
and U3881 (N_3881,In_253,In_558);
nor U3882 (N_3882,In_759,In_258);
nor U3883 (N_3883,In_998,In_445);
nand U3884 (N_3884,In_760,In_757);
nand U3885 (N_3885,In_5,In_775);
nor U3886 (N_3886,In_121,In_971);
nor U3887 (N_3887,In_657,In_634);
nand U3888 (N_3888,In_750,In_648);
nor U3889 (N_3889,In_158,In_860);
or U3890 (N_3890,In_20,In_33);
nor U3891 (N_3891,In_98,In_408);
nor U3892 (N_3892,In_507,In_960);
nor U3893 (N_3893,In_305,In_339);
nand U3894 (N_3894,In_897,In_87);
xnor U3895 (N_3895,In_253,In_691);
nor U3896 (N_3896,In_637,In_815);
nand U3897 (N_3897,In_366,In_713);
and U3898 (N_3898,In_473,In_676);
nor U3899 (N_3899,In_290,In_194);
nor U3900 (N_3900,In_650,In_595);
and U3901 (N_3901,In_104,In_267);
or U3902 (N_3902,In_45,In_151);
nand U3903 (N_3903,In_575,In_369);
nor U3904 (N_3904,In_897,In_503);
nor U3905 (N_3905,In_607,In_559);
nor U3906 (N_3906,In_936,In_390);
nand U3907 (N_3907,In_720,In_196);
and U3908 (N_3908,In_660,In_470);
nor U3909 (N_3909,In_629,In_614);
nand U3910 (N_3910,In_16,In_27);
and U3911 (N_3911,In_818,In_665);
nand U3912 (N_3912,In_662,In_760);
or U3913 (N_3913,In_326,In_880);
nand U3914 (N_3914,In_615,In_824);
or U3915 (N_3915,In_448,In_967);
or U3916 (N_3916,In_294,In_445);
nand U3917 (N_3917,In_128,In_817);
or U3918 (N_3918,In_522,In_717);
and U3919 (N_3919,In_361,In_186);
xor U3920 (N_3920,In_82,In_195);
or U3921 (N_3921,In_144,In_158);
nor U3922 (N_3922,In_111,In_323);
nor U3923 (N_3923,In_121,In_280);
nor U3924 (N_3924,In_365,In_924);
nand U3925 (N_3925,In_346,In_822);
and U3926 (N_3926,In_399,In_763);
nand U3927 (N_3927,In_989,In_940);
or U3928 (N_3928,In_546,In_69);
nand U3929 (N_3929,In_185,In_566);
xnor U3930 (N_3930,In_701,In_167);
xor U3931 (N_3931,In_56,In_99);
and U3932 (N_3932,In_453,In_831);
nand U3933 (N_3933,In_850,In_452);
nand U3934 (N_3934,In_468,In_907);
or U3935 (N_3935,In_970,In_447);
nor U3936 (N_3936,In_175,In_406);
nand U3937 (N_3937,In_47,In_299);
nor U3938 (N_3938,In_339,In_837);
nor U3939 (N_3939,In_331,In_178);
or U3940 (N_3940,In_234,In_223);
nor U3941 (N_3941,In_825,In_454);
or U3942 (N_3942,In_74,In_922);
xor U3943 (N_3943,In_265,In_289);
or U3944 (N_3944,In_749,In_992);
and U3945 (N_3945,In_695,In_296);
nand U3946 (N_3946,In_38,In_446);
and U3947 (N_3947,In_625,In_948);
nand U3948 (N_3948,In_902,In_918);
nor U3949 (N_3949,In_71,In_894);
nand U3950 (N_3950,In_406,In_706);
nand U3951 (N_3951,In_386,In_329);
and U3952 (N_3952,In_689,In_480);
nand U3953 (N_3953,In_397,In_463);
nand U3954 (N_3954,In_812,In_123);
or U3955 (N_3955,In_121,In_422);
or U3956 (N_3956,In_889,In_507);
nor U3957 (N_3957,In_47,In_961);
nor U3958 (N_3958,In_755,In_27);
and U3959 (N_3959,In_372,In_207);
nand U3960 (N_3960,In_294,In_471);
and U3961 (N_3961,In_538,In_290);
nor U3962 (N_3962,In_229,In_680);
nand U3963 (N_3963,In_583,In_131);
or U3964 (N_3964,In_111,In_470);
xor U3965 (N_3965,In_401,In_322);
nor U3966 (N_3966,In_223,In_870);
nor U3967 (N_3967,In_438,In_295);
and U3968 (N_3968,In_614,In_814);
or U3969 (N_3969,In_394,In_737);
or U3970 (N_3970,In_614,In_991);
and U3971 (N_3971,In_857,In_707);
or U3972 (N_3972,In_904,In_827);
nand U3973 (N_3973,In_634,In_872);
and U3974 (N_3974,In_607,In_969);
and U3975 (N_3975,In_137,In_457);
nor U3976 (N_3976,In_365,In_273);
nand U3977 (N_3977,In_853,In_962);
or U3978 (N_3978,In_16,In_759);
nor U3979 (N_3979,In_507,In_229);
or U3980 (N_3980,In_558,In_212);
nor U3981 (N_3981,In_886,In_570);
or U3982 (N_3982,In_479,In_512);
nor U3983 (N_3983,In_445,In_689);
or U3984 (N_3984,In_255,In_881);
nand U3985 (N_3985,In_143,In_435);
nor U3986 (N_3986,In_6,In_916);
nand U3987 (N_3987,In_338,In_788);
and U3988 (N_3988,In_817,In_968);
nand U3989 (N_3989,In_139,In_976);
or U3990 (N_3990,In_59,In_544);
or U3991 (N_3991,In_930,In_564);
and U3992 (N_3992,In_516,In_951);
nand U3993 (N_3993,In_259,In_241);
or U3994 (N_3994,In_13,In_626);
nand U3995 (N_3995,In_278,In_301);
or U3996 (N_3996,In_673,In_707);
and U3997 (N_3997,In_90,In_546);
nor U3998 (N_3998,In_906,In_114);
nand U3999 (N_3999,In_998,In_757);
and U4000 (N_4000,In_997,In_48);
or U4001 (N_4001,In_19,In_509);
and U4002 (N_4002,In_145,In_716);
and U4003 (N_4003,In_590,In_552);
or U4004 (N_4004,In_822,In_27);
xnor U4005 (N_4005,In_714,In_825);
nand U4006 (N_4006,In_918,In_989);
nand U4007 (N_4007,In_875,In_194);
nand U4008 (N_4008,In_693,In_745);
and U4009 (N_4009,In_582,In_284);
nand U4010 (N_4010,In_19,In_83);
and U4011 (N_4011,In_860,In_31);
and U4012 (N_4012,In_980,In_604);
or U4013 (N_4013,In_737,In_172);
xnor U4014 (N_4014,In_769,In_372);
nor U4015 (N_4015,In_663,In_658);
nand U4016 (N_4016,In_290,In_58);
nor U4017 (N_4017,In_18,In_210);
and U4018 (N_4018,In_946,In_714);
nor U4019 (N_4019,In_453,In_809);
and U4020 (N_4020,In_197,In_772);
or U4021 (N_4021,In_876,In_390);
or U4022 (N_4022,In_79,In_698);
nand U4023 (N_4023,In_619,In_178);
and U4024 (N_4024,In_763,In_430);
nand U4025 (N_4025,In_884,In_999);
or U4026 (N_4026,In_922,In_177);
nor U4027 (N_4027,In_103,In_691);
nand U4028 (N_4028,In_595,In_103);
xnor U4029 (N_4029,In_852,In_426);
nand U4030 (N_4030,In_633,In_492);
or U4031 (N_4031,In_279,In_402);
or U4032 (N_4032,In_334,In_869);
nor U4033 (N_4033,In_391,In_526);
nand U4034 (N_4034,In_872,In_705);
nand U4035 (N_4035,In_937,In_281);
nor U4036 (N_4036,In_969,In_445);
and U4037 (N_4037,In_871,In_345);
or U4038 (N_4038,In_638,In_231);
nor U4039 (N_4039,In_994,In_931);
or U4040 (N_4040,In_793,In_112);
or U4041 (N_4041,In_505,In_828);
nand U4042 (N_4042,In_67,In_182);
nor U4043 (N_4043,In_65,In_272);
and U4044 (N_4044,In_242,In_536);
or U4045 (N_4045,In_964,In_662);
or U4046 (N_4046,In_590,In_423);
and U4047 (N_4047,In_394,In_467);
nor U4048 (N_4048,In_464,In_847);
and U4049 (N_4049,In_612,In_483);
and U4050 (N_4050,In_242,In_786);
or U4051 (N_4051,In_195,In_660);
and U4052 (N_4052,In_29,In_796);
or U4053 (N_4053,In_357,In_589);
nand U4054 (N_4054,In_808,In_325);
or U4055 (N_4055,In_873,In_40);
and U4056 (N_4056,In_266,In_532);
nand U4057 (N_4057,In_545,In_920);
and U4058 (N_4058,In_995,In_800);
nor U4059 (N_4059,In_518,In_206);
or U4060 (N_4060,In_805,In_152);
or U4061 (N_4061,In_980,In_434);
nand U4062 (N_4062,In_301,In_66);
nor U4063 (N_4063,In_417,In_84);
and U4064 (N_4064,In_951,In_146);
or U4065 (N_4065,In_437,In_603);
nand U4066 (N_4066,In_229,In_811);
and U4067 (N_4067,In_121,In_345);
or U4068 (N_4068,In_617,In_940);
or U4069 (N_4069,In_422,In_615);
nor U4070 (N_4070,In_519,In_898);
nor U4071 (N_4071,In_981,In_261);
nor U4072 (N_4072,In_577,In_509);
and U4073 (N_4073,In_591,In_665);
nand U4074 (N_4074,In_962,In_39);
nor U4075 (N_4075,In_223,In_664);
or U4076 (N_4076,In_384,In_395);
xnor U4077 (N_4077,In_376,In_581);
and U4078 (N_4078,In_979,In_440);
or U4079 (N_4079,In_802,In_850);
and U4080 (N_4080,In_620,In_316);
or U4081 (N_4081,In_593,In_863);
nand U4082 (N_4082,In_722,In_245);
and U4083 (N_4083,In_749,In_602);
or U4084 (N_4084,In_624,In_572);
and U4085 (N_4085,In_525,In_987);
xor U4086 (N_4086,In_987,In_870);
or U4087 (N_4087,In_159,In_715);
or U4088 (N_4088,In_607,In_81);
nand U4089 (N_4089,In_91,In_68);
nand U4090 (N_4090,In_286,In_440);
xnor U4091 (N_4091,In_575,In_999);
nand U4092 (N_4092,In_549,In_792);
or U4093 (N_4093,In_847,In_600);
nand U4094 (N_4094,In_752,In_591);
or U4095 (N_4095,In_34,In_681);
nor U4096 (N_4096,In_397,In_958);
nor U4097 (N_4097,In_769,In_760);
and U4098 (N_4098,In_993,In_187);
or U4099 (N_4099,In_21,In_969);
nor U4100 (N_4100,In_266,In_81);
nor U4101 (N_4101,In_842,In_787);
nor U4102 (N_4102,In_576,In_936);
or U4103 (N_4103,In_714,In_281);
nor U4104 (N_4104,In_495,In_621);
nand U4105 (N_4105,In_891,In_336);
and U4106 (N_4106,In_261,In_554);
or U4107 (N_4107,In_12,In_197);
nor U4108 (N_4108,In_161,In_421);
and U4109 (N_4109,In_130,In_195);
nand U4110 (N_4110,In_955,In_325);
xor U4111 (N_4111,In_455,In_820);
nand U4112 (N_4112,In_928,In_591);
xor U4113 (N_4113,In_945,In_817);
or U4114 (N_4114,In_687,In_942);
or U4115 (N_4115,In_341,In_123);
or U4116 (N_4116,In_736,In_801);
nor U4117 (N_4117,In_278,In_920);
or U4118 (N_4118,In_893,In_30);
and U4119 (N_4119,In_346,In_541);
nor U4120 (N_4120,In_754,In_557);
nand U4121 (N_4121,In_22,In_493);
nand U4122 (N_4122,In_385,In_401);
nor U4123 (N_4123,In_94,In_602);
nor U4124 (N_4124,In_341,In_209);
or U4125 (N_4125,In_88,In_243);
or U4126 (N_4126,In_410,In_148);
nand U4127 (N_4127,In_873,In_915);
nand U4128 (N_4128,In_549,In_529);
or U4129 (N_4129,In_171,In_957);
or U4130 (N_4130,In_670,In_455);
nand U4131 (N_4131,In_751,In_940);
or U4132 (N_4132,In_877,In_860);
or U4133 (N_4133,In_7,In_41);
or U4134 (N_4134,In_691,In_949);
or U4135 (N_4135,In_919,In_197);
or U4136 (N_4136,In_750,In_837);
or U4137 (N_4137,In_725,In_225);
and U4138 (N_4138,In_585,In_103);
nor U4139 (N_4139,In_192,In_785);
nor U4140 (N_4140,In_840,In_684);
and U4141 (N_4141,In_202,In_939);
or U4142 (N_4142,In_219,In_701);
nor U4143 (N_4143,In_774,In_749);
nor U4144 (N_4144,In_353,In_688);
and U4145 (N_4145,In_62,In_272);
nand U4146 (N_4146,In_279,In_774);
nor U4147 (N_4147,In_480,In_178);
nor U4148 (N_4148,In_692,In_405);
nand U4149 (N_4149,In_926,In_189);
and U4150 (N_4150,In_147,In_154);
or U4151 (N_4151,In_249,In_890);
nor U4152 (N_4152,In_621,In_930);
nor U4153 (N_4153,In_566,In_892);
nor U4154 (N_4154,In_872,In_690);
nor U4155 (N_4155,In_799,In_874);
nand U4156 (N_4156,In_89,In_560);
or U4157 (N_4157,In_238,In_318);
nand U4158 (N_4158,In_408,In_445);
xor U4159 (N_4159,In_535,In_437);
nor U4160 (N_4160,In_676,In_28);
or U4161 (N_4161,In_5,In_481);
or U4162 (N_4162,In_266,In_69);
nor U4163 (N_4163,In_111,In_16);
or U4164 (N_4164,In_710,In_838);
nand U4165 (N_4165,In_258,In_605);
nor U4166 (N_4166,In_363,In_179);
nor U4167 (N_4167,In_322,In_556);
nand U4168 (N_4168,In_274,In_678);
and U4169 (N_4169,In_265,In_791);
nor U4170 (N_4170,In_265,In_716);
nor U4171 (N_4171,In_560,In_620);
or U4172 (N_4172,In_292,In_299);
nor U4173 (N_4173,In_815,In_407);
or U4174 (N_4174,In_659,In_523);
nor U4175 (N_4175,In_971,In_77);
or U4176 (N_4176,In_951,In_121);
nor U4177 (N_4177,In_305,In_707);
and U4178 (N_4178,In_319,In_685);
and U4179 (N_4179,In_764,In_29);
nor U4180 (N_4180,In_127,In_424);
nor U4181 (N_4181,In_808,In_352);
or U4182 (N_4182,In_389,In_901);
or U4183 (N_4183,In_671,In_246);
or U4184 (N_4184,In_100,In_349);
nand U4185 (N_4185,In_606,In_515);
or U4186 (N_4186,In_622,In_616);
or U4187 (N_4187,In_825,In_365);
nand U4188 (N_4188,In_788,In_364);
nor U4189 (N_4189,In_963,In_135);
nand U4190 (N_4190,In_412,In_750);
or U4191 (N_4191,In_374,In_558);
nand U4192 (N_4192,In_923,In_680);
or U4193 (N_4193,In_624,In_594);
and U4194 (N_4194,In_256,In_454);
nand U4195 (N_4195,In_252,In_904);
nand U4196 (N_4196,In_362,In_489);
nand U4197 (N_4197,In_185,In_129);
nor U4198 (N_4198,In_299,In_598);
or U4199 (N_4199,In_546,In_543);
or U4200 (N_4200,In_246,In_210);
nor U4201 (N_4201,In_55,In_958);
nand U4202 (N_4202,In_585,In_141);
and U4203 (N_4203,In_552,In_309);
and U4204 (N_4204,In_885,In_354);
xnor U4205 (N_4205,In_400,In_286);
or U4206 (N_4206,In_691,In_825);
or U4207 (N_4207,In_774,In_298);
nor U4208 (N_4208,In_980,In_279);
and U4209 (N_4209,In_772,In_351);
nand U4210 (N_4210,In_157,In_875);
or U4211 (N_4211,In_545,In_45);
or U4212 (N_4212,In_750,In_103);
nand U4213 (N_4213,In_985,In_265);
xnor U4214 (N_4214,In_95,In_976);
and U4215 (N_4215,In_363,In_596);
or U4216 (N_4216,In_90,In_966);
nand U4217 (N_4217,In_208,In_901);
nand U4218 (N_4218,In_96,In_763);
nor U4219 (N_4219,In_629,In_637);
nor U4220 (N_4220,In_640,In_915);
and U4221 (N_4221,In_228,In_699);
nor U4222 (N_4222,In_428,In_311);
or U4223 (N_4223,In_565,In_297);
nand U4224 (N_4224,In_631,In_925);
nand U4225 (N_4225,In_440,In_912);
nand U4226 (N_4226,In_832,In_333);
nor U4227 (N_4227,In_261,In_747);
and U4228 (N_4228,In_38,In_702);
nand U4229 (N_4229,In_215,In_123);
nor U4230 (N_4230,In_489,In_151);
nor U4231 (N_4231,In_290,In_42);
nand U4232 (N_4232,In_706,In_305);
and U4233 (N_4233,In_576,In_492);
nor U4234 (N_4234,In_749,In_933);
nor U4235 (N_4235,In_328,In_867);
nand U4236 (N_4236,In_19,In_698);
and U4237 (N_4237,In_338,In_674);
and U4238 (N_4238,In_62,In_170);
or U4239 (N_4239,In_745,In_608);
nand U4240 (N_4240,In_23,In_268);
and U4241 (N_4241,In_397,In_508);
xor U4242 (N_4242,In_89,In_539);
nand U4243 (N_4243,In_931,In_623);
nor U4244 (N_4244,In_98,In_258);
nand U4245 (N_4245,In_461,In_499);
nand U4246 (N_4246,In_332,In_171);
or U4247 (N_4247,In_16,In_319);
nor U4248 (N_4248,In_4,In_491);
or U4249 (N_4249,In_157,In_861);
and U4250 (N_4250,In_766,In_375);
nand U4251 (N_4251,In_435,In_984);
nor U4252 (N_4252,In_886,In_26);
nand U4253 (N_4253,In_4,In_275);
nand U4254 (N_4254,In_530,In_595);
nand U4255 (N_4255,In_605,In_307);
and U4256 (N_4256,In_57,In_742);
or U4257 (N_4257,In_740,In_775);
and U4258 (N_4258,In_888,In_339);
or U4259 (N_4259,In_679,In_787);
nand U4260 (N_4260,In_956,In_44);
and U4261 (N_4261,In_288,In_86);
nor U4262 (N_4262,In_467,In_53);
and U4263 (N_4263,In_576,In_109);
nor U4264 (N_4264,In_851,In_988);
or U4265 (N_4265,In_595,In_608);
nor U4266 (N_4266,In_53,In_127);
nor U4267 (N_4267,In_796,In_890);
nand U4268 (N_4268,In_422,In_158);
and U4269 (N_4269,In_275,In_662);
nor U4270 (N_4270,In_388,In_704);
nor U4271 (N_4271,In_465,In_98);
or U4272 (N_4272,In_204,In_146);
and U4273 (N_4273,In_192,In_533);
or U4274 (N_4274,In_5,In_54);
nor U4275 (N_4275,In_659,In_153);
or U4276 (N_4276,In_358,In_464);
nand U4277 (N_4277,In_197,In_880);
nor U4278 (N_4278,In_817,In_293);
or U4279 (N_4279,In_156,In_822);
and U4280 (N_4280,In_507,In_907);
nor U4281 (N_4281,In_355,In_591);
nand U4282 (N_4282,In_955,In_110);
nand U4283 (N_4283,In_687,In_317);
and U4284 (N_4284,In_556,In_969);
nor U4285 (N_4285,In_620,In_188);
nand U4286 (N_4286,In_196,In_20);
nor U4287 (N_4287,In_242,In_16);
nand U4288 (N_4288,In_752,In_379);
nor U4289 (N_4289,In_141,In_693);
nand U4290 (N_4290,In_767,In_43);
and U4291 (N_4291,In_277,In_695);
and U4292 (N_4292,In_758,In_411);
nor U4293 (N_4293,In_362,In_154);
nand U4294 (N_4294,In_889,In_33);
or U4295 (N_4295,In_720,In_311);
or U4296 (N_4296,In_86,In_78);
and U4297 (N_4297,In_671,In_17);
nand U4298 (N_4298,In_731,In_987);
or U4299 (N_4299,In_818,In_908);
and U4300 (N_4300,In_851,In_592);
and U4301 (N_4301,In_697,In_9);
nand U4302 (N_4302,In_638,In_509);
nand U4303 (N_4303,In_592,In_588);
nand U4304 (N_4304,In_526,In_55);
nor U4305 (N_4305,In_760,In_588);
nand U4306 (N_4306,In_990,In_959);
and U4307 (N_4307,In_591,In_193);
and U4308 (N_4308,In_725,In_373);
and U4309 (N_4309,In_700,In_728);
or U4310 (N_4310,In_536,In_995);
nor U4311 (N_4311,In_534,In_279);
nand U4312 (N_4312,In_543,In_73);
or U4313 (N_4313,In_372,In_375);
and U4314 (N_4314,In_718,In_881);
nand U4315 (N_4315,In_434,In_327);
nand U4316 (N_4316,In_909,In_793);
nand U4317 (N_4317,In_375,In_209);
nor U4318 (N_4318,In_155,In_841);
nand U4319 (N_4319,In_427,In_494);
nand U4320 (N_4320,In_485,In_321);
or U4321 (N_4321,In_861,In_137);
nor U4322 (N_4322,In_213,In_643);
or U4323 (N_4323,In_359,In_950);
nor U4324 (N_4324,In_723,In_379);
and U4325 (N_4325,In_825,In_175);
nand U4326 (N_4326,In_763,In_829);
and U4327 (N_4327,In_843,In_314);
and U4328 (N_4328,In_307,In_869);
nor U4329 (N_4329,In_100,In_177);
or U4330 (N_4330,In_684,In_220);
and U4331 (N_4331,In_354,In_645);
xnor U4332 (N_4332,In_935,In_618);
nand U4333 (N_4333,In_440,In_217);
nor U4334 (N_4334,In_988,In_232);
nor U4335 (N_4335,In_406,In_508);
nand U4336 (N_4336,In_119,In_372);
and U4337 (N_4337,In_947,In_399);
nand U4338 (N_4338,In_20,In_971);
or U4339 (N_4339,In_806,In_821);
nor U4340 (N_4340,In_567,In_466);
or U4341 (N_4341,In_112,In_13);
or U4342 (N_4342,In_386,In_355);
or U4343 (N_4343,In_843,In_282);
nand U4344 (N_4344,In_145,In_369);
and U4345 (N_4345,In_153,In_171);
nand U4346 (N_4346,In_303,In_851);
or U4347 (N_4347,In_226,In_648);
and U4348 (N_4348,In_31,In_712);
and U4349 (N_4349,In_72,In_543);
or U4350 (N_4350,In_42,In_567);
nor U4351 (N_4351,In_701,In_162);
or U4352 (N_4352,In_79,In_91);
nand U4353 (N_4353,In_574,In_314);
or U4354 (N_4354,In_983,In_210);
and U4355 (N_4355,In_436,In_787);
or U4356 (N_4356,In_405,In_555);
and U4357 (N_4357,In_856,In_250);
nor U4358 (N_4358,In_261,In_351);
nand U4359 (N_4359,In_215,In_714);
and U4360 (N_4360,In_767,In_174);
and U4361 (N_4361,In_413,In_334);
and U4362 (N_4362,In_61,In_180);
nor U4363 (N_4363,In_391,In_98);
nor U4364 (N_4364,In_928,In_806);
and U4365 (N_4365,In_695,In_476);
nor U4366 (N_4366,In_20,In_464);
nand U4367 (N_4367,In_975,In_285);
nor U4368 (N_4368,In_384,In_726);
nor U4369 (N_4369,In_644,In_786);
nand U4370 (N_4370,In_622,In_583);
or U4371 (N_4371,In_834,In_930);
and U4372 (N_4372,In_0,In_398);
nor U4373 (N_4373,In_485,In_884);
nor U4374 (N_4374,In_913,In_382);
nor U4375 (N_4375,In_122,In_399);
xor U4376 (N_4376,In_483,In_274);
nand U4377 (N_4377,In_852,In_942);
nor U4378 (N_4378,In_701,In_468);
or U4379 (N_4379,In_123,In_933);
nand U4380 (N_4380,In_486,In_637);
and U4381 (N_4381,In_837,In_331);
nand U4382 (N_4382,In_602,In_850);
and U4383 (N_4383,In_262,In_367);
and U4384 (N_4384,In_110,In_352);
nor U4385 (N_4385,In_211,In_862);
nand U4386 (N_4386,In_468,In_240);
or U4387 (N_4387,In_18,In_260);
nor U4388 (N_4388,In_516,In_59);
and U4389 (N_4389,In_699,In_149);
or U4390 (N_4390,In_20,In_306);
nor U4391 (N_4391,In_289,In_262);
or U4392 (N_4392,In_158,In_608);
or U4393 (N_4393,In_308,In_693);
xnor U4394 (N_4394,In_12,In_719);
nand U4395 (N_4395,In_411,In_130);
and U4396 (N_4396,In_488,In_883);
nor U4397 (N_4397,In_228,In_636);
nor U4398 (N_4398,In_861,In_3);
nand U4399 (N_4399,In_564,In_200);
or U4400 (N_4400,In_614,In_47);
or U4401 (N_4401,In_758,In_285);
nand U4402 (N_4402,In_489,In_354);
nand U4403 (N_4403,In_609,In_525);
or U4404 (N_4404,In_634,In_692);
or U4405 (N_4405,In_369,In_25);
nand U4406 (N_4406,In_316,In_299);
or U4407 (N_4407,In_502,In_767);
nor U4408 (N_4408,In_89,In_714);
or U4409 (N_4409,In_589,In_74);
nand U4410 (N_4410,In_440,In_479);
nor U4411 (N_4411,In_660,In_380);
xor U4412 (N_4412,In_287,In_857);
or U4413 (N_4413,In_778,In_607);
and U4414 (N_4414,In_895,In_336);
nor U4415 (N_4415,In_718,In_312);
nor U4416 (N_4416,In_154,In_351);
and U4417 (N_4417,In_681,In_815);
or U4418 (N_4418,In_134,In_176);
or U4419 (N_4419,In_733,In_67);
nor U4420 (N_4420,In_982,In_887);
or U4421 (N_4421,In_476,In_186);
or U4422 (N_4422,In_813,In_434);
nor U4423 (N_4423,In_918,In_242);
nand U4424 (N_4424,In_230,In_267);
and U4425 (N_4425,In_180,In_99);
or U4426 (N_4426,In_965,In_165);
or U4427 (N_4427,In_328,In_839);
or U4428 (N_4428,In_903,In_174);
nor U4429 (N_4429,In_667,In_991);
nor U4430 (N_4430,In_939,In_878);
nor U4431 (N_4431,In_268,In_375);
nor U4432 (N_4432,In_170,In_739);
or U4433 (N_4433,In_234,In_473);
and U4434 (N_4434,In_8,In_912);
nor U4435 (N_4435,In_400,In_880);
and U4436 (N_4436,In_89,In_110);
nand U4437 (N_4437,In_807,In_664);
and U4438 (N_4438,In_320,In_919);
and U4439 (N_4439,In_71,In_446);
and U4440 (N_4440,In_125,In_132);
and U4441 (N_4441,In_196,In_900);
nand U4442 (N_4442,In_430,In_687);
nand U4443 (N_4443,In_713,In_648);
nor U4444 (N_4444,In_119,In_699);
nand U4445 (N_4445,In_154,In_466);
and U4446 (N_4446,In_209,In_140);
and U4447 (N_4447,In_645,In_315);
nor U4448 (N_4448,In_668,In_353);
nor U4449 (N_4449,In_533,In_79);
nand U4450 (N_4450,In_779,In_934);
nor U4451 (N_4451,In_652,In_277);
nor U4452 (N_4452,In_363,In_320);
nand U4453 (N_4453,In_353,In_672);
or U4454 (N_4454,In_914,In_329);
nor U4455 (N_4455,In_654,In_297);
nor U4456 (N_4456,In_746,In_332);
or U4457 (N_4457,In_892,In_932);
and U4458 (N_4458,In_455,In_457);
nor U4459 (N_4459,In_875,In_313);
nand U4460 (N_4460,In_647,In_236);
and U4461 (N_4461,In_272,In_696);
or U4462 (N_4462,In_666,In_654);
nand U4463 (N_4463,In_864,In_61);
nand U4464 (N_4464,In_902,In_718);
or U4465 (N_4465,In_214,In_928);
nand U4466 (N_4466,In_313,In_969);
or U4467 (N_4467,In_452,In_293);
nand U4468 (N_4468,In_279,In_436);
nand U4469 (N_4469,In_882,In_629);
nor U4470 (N_4470,In_563,In_839);
and U4471 (N_4471,In_268,In_201);
or U4472 (N_4472,In_642,In_468);
nand U4473 (N_4473,In_829,In_469);
or U4474 (N_4474,In_779,In_281);
and U4475 (N_4475,In_956,In_132);
or U4476 (N_4476,In_237,In_635);
nor U4477 (N_4477,In_40,In_370);
or U4478 (N_4478,In_620,In_943);
nor U4479 (N_4479,In_31,In_753);
and U4480 (N_4480,In_542,In_29);
nor U4481 (N_4481,In_104,In_8);
and U4482 (N_4482,In_317,In_616);
nand U4483 (N_4483,In_454,In_746);
nor U4484 (N_4484,In_181,In_990);
nand U4485 (N_4485,In_938,In_951);
nand U4486 (N_4486,In_742,In_117);
nor U4487 (N_4487,In_548,In_934);
xnor U4488 (N_4488,In_545,In_363);
xnor U4489 (N_4489,In_302,In_984);
nor U4490 (N_4490,In_729,In_566);
and U4491 (N_4491,In_438,In_148);
and U4492 (N_4492,In_920,In_75);
or U4493 (N_4493,In_92,In_847);
nor U4494 (N_4494,In_470,In_180);
nand U4495 (N_4495,In_704,In_553);
nor U4496 (N_4496,In_703,In_345);
or U4497 (N_4497,In_958,In_152);
and U4498 (N_4498,In_157,In_200);
nor U4499 (N_4499,In_173,In_473);
and U4500 (N_4500,In_213,In_938);
and U4501 (N_4501,In_229,In_492);
or U4502 (N_4502,In_68,In_348);
and U4503 (N_4503,In_558,In_605);
nor U4504 (N_4504,In_579,In_916);
and U4505 (N_4505,In_39,In_182);
and U4506 (N_4506,In_867,In_810);
xor U4507 (N_4507,In_326,In_530);
nand U4508 (N_4508,In_177,In_463);
xor U4509 (N_4509,In_819,In_18);
and U4510 (N_4510,In_259,In_779);
nor U4511 (N_4511,In_415,In_402);
nor U4512 (N_4512,In_968,In_587);
xnor U4513 (N_4513,In_225,In_220);
nor U4514 (N_4514,In_845,In_702);
nor U4515 (N_4515,In_388,In_577);
or U4516 (N_4516,In_566,In_400);
nor U4517 (N_4517,In_42,In_78);
nand U4518 (N_4518,In_486,In_102);
and U4519 (N_4519,In_200,In_810);
nand U4520 (N_4520,In_920,In_858);
and U4521 (N_4521,In_379,In_70);
nand U4522 (N_4522,In_470,In_779);
nor U4523 (N_4523,In_261,In_142);
nand U4524 (N_4524,In_942,In_873);
and U4525 (N_4525,In_501,In_890);
nor U4526 (N_4526,In_793,In_641);
nor U4527 (N_4527,In_134,In_44);
or U4528 (N_4528,In_220,In_972);
nand U4529 (N_4529,In_68,In_405);
nand U4530 (N_4530,In_431,In_473);
nand U4531 (N_4531,In_655,In_259);
nor U4532 (N_4532,In_274,In_335);
and U4533 (N_4533,In_253,In_656);
nor U4534 (N_4534,In_300,In_597);
nor U4535 (N_4535,In_18,In_21);
nand U4536 (N_4536,In_419,In_550);
xnor U4537 (N_4537,In_175,In_142);
nand U4538 (N_4538,In_449,In_910);
and U4539 (N_4539,In_126,In_995);
and U4540 (N_4540,In_558,In_223);
and U4541 (N_4541,In_805,In_515);
or U4542 (N_4542,In_63,In_423);
nor U4543 (N_4543,In_452,In_965);
or U4544 (N_4544,In_67,In_797);
nor U4545 (N_4545,In_550,In_510);
and U4546 (N_4546,In_336,In_38);
nor U4547 (N_4547,In_181,In_737);
or U4548 (N_4548,In_753,In_332);
nor U4549 (N_4549,In_318,In_606);
nor U4550 (N_4550,In_386,In_27);
and U4551 (N_4551,In_393,In_975);
nor U4552 (N_4552,In_518,In_233);
nand U4553 (N_4553,In_744,In_936);
or U4554 (N_4554,In_87,In_588);
or U4555 (N_4555,In_428,In_13);
or U4556 (N_4556,In_416,In_421);
and U4557 (N_4557,In_7,In_980);
or U4558 (N_4558,In_609,In_309);
nand U4559 (N_4559,In_827,In_759);
or U4560 (N_4560,In_881,In_926);
and U4561 (N_4561,In_85,In_624);
nor U4562 (N_4562,In_353,In_976);
nor U4563 (N_4563,In_693,In_344);
nor U4564 (N_4564,In_116,In_356);
nand U4565 (N_4565,In_1,In_231);
and U4566 (N_4566,In_99,In_363);
and U4567 (N_4567,In_56,In_937);
nand U4568 (N_4568,In_611,In_482);
and U4569 (N_4569,In_950,In_761);
or U4570 (N_4570,In_550,In_773);
nor U4571 (N_4571,In_986,In_847);
and U4572 (N_4572,In_647,In_21);
or U4573 (N_4573,In_880,In_376);
nand U4574 (N_4574,In_565,In_611);
nor U4575 (N_4575,In_59,In_165);
nor U4576 (N_4576,In_480,In_927);
or U4577 (N_4577,In_217,In_685);
nand U4578 (N_4578,In_279,In_586);
or U4579 (N_4579,In_572,In_640);
and U4580 (N_4580,In_521,In_70);
or U4581 (N_4581,In_149,In_844);
nor U4582 (N_4582,In_769,In_626);
nor U4583 (N_4583,In_839,In_273);
and U4584 (N_4584,In_500,In_457);
and U4585 (N_4585,In_551,In_637);
nor U4586 (N_4586,In_568,In_678);
or U4587 (N_4587,In_923,In_70);
or U4588 (N_4588,In_756,In_649);
nor U4589 (N_4589,In_589,In_756);
xor U4590 (N_4590,In_712,In_673);
nor U4591 (N_4591,In_503,In_250);
and U4592 (N_4592,In_553,In_391);
and U4593 (N_4593,In_560,In_472);
nand U4594 (N_4594,In_494,In_432);
xnor U4595 (N_4595,In_711,In_891);
nor U4596 (N_4596,In_8,In_244);
nor U4597 (N_4597,In_82,In_470);
xnor U4598 (N_4598,In_698,In_880);
nand U4599 (N_4599,In_754,In_469);
nor U4600 (N_4600,In_558,In_394);
or U4601 (N_4601,In_79,In_342);
nand U4602 (N_4602,In_590,In_447);
nor U4603 (N_4603,In_175,In_278);
nor U4604 (N_4604,In_592,In_385);
or U4605 (N_4605,In_760,In_386);
nor U4606 (N_4606,In_173,In_243);
and U4607 (N_4607,In_16,In_314);
and U4608 (N_4608,In_125,In_591);
nand U4609 (N_4609,In_193,In_813);
nand U4610 (N_4610,In_166,In_916);
nor U4611 (N_4611,In_580,In_937);
xnor U4612 (N_4612,In_59,In_566);
nor U4613 (N_4613,In_666,In_387);
or U4614 (N_4614,In_175,In_194);
xnor U4615 (N_4615,In_870,In_941);
nand U4616 (N_4616,In_733,In_883);
nand U4617 (N_4617,In_76,In_88);
nor U4618 (N_4618,In_540,In_874);
or U4619 (N_4619,In_830,In_571);
or U4620 (N_4620,In_846,In_808);
and U4621 (N_4621,In_146,In_604);
nor U4622 (N_4622,In_751,In_670);
nand U4623 (N_4623,In_848,In_493);
nor U4624 (N_4624,In_43,In_513);
nor U4625 (N_4625,In_690,In_228);
nand U4626 (N_4626,In_466,In_201);
nand U4627 (N_4627,In_893,In_9);
and U4628 (N_4628,In_391,In_81);
and U4629 (N_4629,In_836,In_808);
or U4630 (N_4630,In_832,In_429);
nand U4631 (N_4631,In_312,In_599);
or U4632 (N_4632,In_783,In_958);
or U4633 (N_4633,In_286,In_980);
and U4634 (N_4634,In_539,In_103);
nand U4635 (N_4635,In_741,In_310);
nand U4636 (N_4636,In_864,In_362);
or U4637 (N_4637,In_613,In_331);
nor U4638 (N_4638,In_160,In_582);
or U4639 (N_4639,In_913,In_621);
nor U4640 (N_4640,In_101,In_60);
nor U4641 (N_4641,In_841,In_97);
nor U4642 (N_4642,In_592,In_157);
and U4643 (N_4643,In_135,In_269);
or U4644 (N_4644,In_188,In_385);
nor U4645 (N_4645,In_134,In_237);
and U4646 (N_4646,In_731,In_864);
and U4647 (N_4647,In_799,In_752);
nand U4648 (N_4648,In_962,In_540);
nor U4649 (N_4649,In_91,In_457);
xor U4650 (N_4650,In_720,In_915);
nand U4651 (N_4651,In_922,In_791);
nor U4652 (N_4652,In_316,In_202);
or U4653 (N_4653,In_299,In_719);
nand U4654 (N_4654,In_622,In_880);
nor U4655 (N_4655,In_321,In_174);
or U4656 (N_4656,In_433,In_871);
and U4657 (N_4657,In_348,In_440);
and U4658 (N_4658,In_66,In_98);
nor U4659 (N_4659,In_276,In_875);
nor U4660 (N_4660,In_969,In_349);
or U4661 (N_4661,In_142,In_486);
nor U4662 (N_4662,In_939,In_122);
nand U4663 (N_4663,In_842,In_67);
and U4664 (N_4664,In_375,In_327);
or U4665 (N_4665,In_267,In_272);
nor U4666 (N_4666,In_625,In_159);
nor U4667 (N_4667,In_525,In_693);
nand U4668 (N_4668,In_766,In_963);
and U4669 (N_4669,In_992,In_958);
xnor U4670 (N_4670,In_850,In_155);
nand U4671 (N_4671,In_432,In_983);
nand U4672 (N_4672,In_35,In_357);
nor U4673 (N_4673,In_3,In_891);
and U4674 (N_4674,In_945,In_554);
or U4675 (N_4675,In_87,In_846);
or U4676 (N_4676,In_861,In_153);
nor U4677 (N_4677,In_340,In_442);
or U4678 (N_4678,In_258,In_561);
and U4679 (N_4679,In_556,In_114);
nand U4680 (N_4680,In_222,In_700);
and U4681 (N_4681,In_572,In_654);
and U4682 (N_4682,In_462,In_411);
and U4683 (N_4683,In_548,In_329);
or U4684 (N_4684,In_730,In_845);
or U4685 (N_4685,In_773,In_969);
nor U4686 (N_4686,In_373,In_424);
nor U4687 (N_4687,In_647,In_209);
nand U4688 (N_4688,In_697,In_222);
nand U4689 (N_4689,In_116,In_424);
or U4690 (N_4690,In_572,In_663);
nor U4691 (N_4691,In_7,In_999);
and U4692 (N_4692,In_386,In_209);
nand U4693 (N_4693,In_864,In_68);
or U4694 (N_4694,In_355,In_412);
nor U4695 (N_4695,In_368,In_252);
nor U4696 (N_4696,In_204,In_359);
or U4697 (N_4697,In_349,In_105);
or U4698 (N_4698,In_816,In_454);
and U4699 (N_4699,In_779,In_577);
and U4700 (N_4700,In_739,In_495);
nand U4701 (N_4701,In_381,In_8);
nor U4702 (N_4702,In_289,In_111);
or U4703 (N_4703,In_766,In_774);
and U4704 (N_4704,In_828,In_863);
or U4705 (N_4705,In_776,In_284);
xnor U4706 (N_4706,In_543,In_562);
nand U4707 (N_4707,In_333,In_772);
or U4708 (N_4708,In_70,In_172);
and U4709 (N_4709,In_880,In_564);
nand U4710 (N_4710,In_45,In_831);
and U4711 (N_4711,In_263,In_287);
nor U4712 (N_4712,In_12,In_950);
or U4713 (N_4713,In_198,In_32);
and U4714 (N_4714,In_91,In_604);
or U4715 (N_4715,In_895,In_442);
or U4716 (N_4716,In_30,In_675);
nand U4717 (N_4717,In_395,In_210);
or U4718 (N_4718,In_360,In_602);
nand U4719 (N_4719,In_548,In_208);
nand U4720 (N_4720,In_251,In_472);
nor U4721 (N_4721,In_357,In_145);
xor U4722 (N_4722,In_631,In_859);
nor U4723 (N_4723,In_304,In_90);
nor U4724 (N_4724,In_626,In_57);
or U4725 (N_4725,In_338,In_734);
nor U4726 (N_4726,In_850,In_927);
and U4727 (N_4727,In_597,In_855);
or U4728 (N_4728,In_487,In_520);
and U4729 (N_4729,In_149,In_178);
nand U4730 (N_4730,In_544,In_579);
and U4731 (N_4731,In_380,In_860);
or U4732 (N_4732,In_205,In_662);
and U4733 (N_4733,In_312,In_803);
and U4734 (N_4734,In_942,In_294);
nand U4735 (N_4735,In_939,In_463);
or U4736 (N_4736,In_172,In_478);
nor U4737 (N_4737,In_451,In_596);
nor U4738 (N_4738,In_777,In_771);
xor U4739 (N_4739,In_344,In_915);
and U4740 (N_4740,In_160,In_448);
nand U4741 (N_4741,In_109,In_178);
nand U4742 (N_4742,In_795,In_779);
nor U4743 (N_4743,In_707,In_271);
and U4744 (N_4744,In_683,In_430);
nor U4745 (N_4745,In_587,In_389);
nor U4746 (N_4746,In_56,In_476);
nand U4747 (N_4747,In_290,In_340);
or U4748 (N_4748,In_309,In_182);
nor U4749 (N_4749,In_676,In_770);
nor U4750 (N_4750,In_786,In_166);
nor U4751 (N_4751,In_870,In_653);
nand U4752 (N_4752,In_867,In_261);
nor U4753 (N_4753,In_943,In_927);
or U4754 (N_4754,In_765,In_33);
or U4755 (N_4755,In_308,In_446);
and U4756 (N_4756,In_568,In_160);
nand U4757 (N_4757,In_155,In_408);
and U4758 (N_4758,In_313,In_301);
xor U4759 (N_4759,In_42,In_342);
and U4760 (N_4760,In_471,In_121);
nand U4761 (N_4761,In_156,In_766);
or U4762 (N_4762,In_772,In_408);
nand U4763 (N_4763,In_603,In_727);
nor U4764 (N_4764,In_907,In_798);
nor U4765 (N_4765,In_741,In_45);
nand U4766 (N_4766,In_463,In_487);
or U4767 (N_4767,In_703,In_783);
or U4768 (N_4768,In_284,In_428);
nand U4769 (N_4769,In_318,In_194);
nand U4770 (N_4770,In_634,In_826);
nor U4771 (N_4771,In_881,In_755);
nand U4772 (N_4772,In_191,In_363);
and U4773 (N_4773,In_174,In_103);
xnor U4774 (N_4774,In_687,In_805);
nand U4775 (N_4775,In_4,In_66);
nand U4776 (N_4776,In_224,In_513);
nand U4777 (N_4777,In_551,In_579);
nor U4778 (N_4778,In_690,In_674);
or U4779 (N_4779,In_728,In_587);
nand U4780 (N_4780,In_304,In_101);
or U4781 (N_4781,In_506,In_748);
nand U4782 (N_4782,In_866,In_915);
or U4783 (N_4783,In_513,In_11);
nor U4784 (N_4784,In_5,In_220);
nor U4785 (N_4785,In_509,In_429);
nor U4786 (N_4786,In_370,In_95);
and U4787 (N_4787,In_290,In_887);
nand U4788 (N_4788,In_872,In_440);
nand U4789 (N_4789,In_810,In_855);
nor U4790 (N_4790,In_88,In_570);
nor U4791 (N_4791,In_651,In_428);
nor U4792 (N_4792,In_831,In_35);
and U4793 (N_4793,In_426,In_755);
or U4794 (N_4794,In_661,In_459);
or U4795 (N_4795,In_408,In_587);
nand U4796 (N_4796,In_256,In_252);
nor U4797 (N_4797,In_401,In_532);
nor U4798 (N_4798,In_963,In_67);
or U4799 (N_4799,In_209,In_880);
nand U4800 (N_4800,In_925,In_726);
or U4801 (N_4801,In_977,In_24);
nand U4802 (N_4802,In_4,In_76);
nor U4803 (N_4803,In_358,In_690);
and U4804 (N_4804,In_322,In_228);
nand U4805 (N_4805,In_858,In_691);
nor U4806 (N_4806,In_495,In_198);
nand U4807 (N_4807,In_709,In_759);
and U4808 (N_4808,In_325,In_215);
or U4809 (N_4809,In_880,In_385);
and U4810 (N_4810,In_879,In_884);
nor U4811 (N_4811,In_378,In_957);
nand U4812 (N_4812,In_375,In_654);
or U4813 (N_4813,In_421,In_792);
or U4814 (N_4814,In_765,In_116);
and U4815 (N_4815,In_342,In_502);
nand U4816 (N_4816,In_982,In_275);
and U4817 (N_4817,In_378,In_751);
nand U4818 (N_4818,In_478,In_100);
nor U4819 (N_4819,In_110,In_925);
and U4820 (N_4820,In_32,In_688);
or U4821 (N_4821,In_233,In_251);
or U4822 (N_4822,In_766,In_457);
or U4823 (N_4823,In_667,In_774);
nand U4824 (N_4824,In_478,In_866);
nor U4825 (N_4825,In_437,In_776);
nand U4826 (N_4826,In_303,In_810);
or U4827 (N_4827,In_922,In_229);
or U4828 (N_4828,In_534,In_79);
and U4829 (N_4829,In_692,In_462);
and U4830 (N_4830,In_140,In_196);
nor U4831 (N_4831,In_856,In_296);
and U4832 (N_4832,In_52,In_789);
or U4833 (N_4833,In_577,In_80);
and U4834 (N_4834,In_119,In_936);
nor U4835 (N_4835,In_139,In_384);
nand U4836 (N_4836,In_83,In_997);
or U4837 (N_4837,In_98,In_921);
nand U4838 (N_4838,In_670,In_404);
or U4839 (N_4839,In_208,In_789);
or U4840 (N_4840,In_100,In_194);
nor U4841 (N_4841,In_508,In_846);
nand U4842 (N_4842,In_65,In_967);
nand U4843 (N_4843,In_766,In_419);
nor U4844 (N_4844,In_797,In_11);
and U4845 (N_4845,In_846,In_531);
and U4846 (N_4846,In_643,In_122);
nand U4847 (N_4847,In_80,In_619);
or U4848 (N_4848,In_50,In_499);
nand U4849 (N_4849,In_390,In_836);
or U4850 (N_4850,In_667,In_613);
nor U4851 (N_4851,In_553,In_523);
and U4852 (N_4852,In_692,In_790);
nand U4853 (N_4853,In_316,In_105);
nor U4854 (N_4854,In_790,In_172);
or U4855 (N_4855,In_80,In_384);
nor U4856 (N_4856,In_359,In_535);
nor U4857 (N_4857,In_889,In_555);
or U4858 (N_4858,In_451,In_362);
nand U4859 (N_4859,In_980,In_350);
nor U4860 (N_4860,In_98,In_158);
and U4861 (N_4861,In_583,In_335);
nand U4862 (N_4862,In_929,In_646);
nor U4863 (N_4863,In_314,In_352);
xor U4864 (N_4864,In_610,In_518);
nor U4865 (N_4865,In_223,In_589);
nor U4866 (N_4866,In_700,In_612);
nand U4867 (N_4867,In_747,In_566);
and U4868 (N_4868,In_945,In_136);
nor U4869 (N_4869,In_477,In_817);
nand U4870 (N_4870,In_117,In_419);
nor U4871 (N_4871,In_9,In_751);
nand U4872 (N_4872,In_340,In_518);
and U4873 (N_4873,In_653,In_384);
nor U4874 (N_4874,In_85,In_250);
nor U4875 (N_4875,In_623,In_474);
nand U4876 (N_4876,In_148,In_691);
nor U4877 (N_4877,In_502,In_339);
or U4878 (N_4878,In_844,In_507);
nand U4879 (N_4879,In_731,In_718);
and U4880 (N_4880,In_166,In_50);
or U4881 (N_4881,In_303,In_23);
or U4882 (N_4882,In_854,In_20);
and U4883 (N_4883,In_474,In_289);
nand U4884 (N_4884,In_879,In_141);
or U4885 (N_4885,In_851,In_388);
nor U4886 (N_4886,In_545,In_724);
xnor U4887 (N_4887,In_464,In_454);
or U4888 (N_4888,In_149,In_476);
or U4889 (N_4889,In_847,In_649);
and U4890 (N_4890,In_751,In_631);
nor U4891 (N_4891,In_596,In_899);
nand U4892 (N_4892,In_137,In_349);
nand U4893 (N_4893,In_79,In_204);
nand U4894 (N_4894,In_144,In_495);
and U4895 (N_4895,In_709,In_779);
nor U4896 (N_4896,In_190,In_714);
and U4897 (N_4897,In_314,In_868);
or U4898 (N_4898,In_265,In_394);
and U4899 (N_4899,In_850,In_414);
and U4900 (N_4900,In_244,In_909);
nand U4901 (N_4901,In_598,In_648);
and U4902 (N_4902,In_992,In_890);
or U4903 (N_4903,In_8,In_327);
nand U4904 (N_4904,In_186,In_959);
nand U4905 (N_4905,In_4,In_417);
or U4906 (N_4906,In_933,In_505);
and U4907 (N_4907,In_568,In_935);
nand U4908 (N_4908,In_570,In_892);
nand U4909 (N_4909,In_197,In_97);
and U4910 (N_4910,In_161,In_477);
nor U4911 (N_4911,In_794,In_506);
and U4912 (N_4912,In_242,In_430);
nand U4913 (N_4913,In_634,In_270);
or U4914 (N_4914,In_212,In_521);
and U4915 (N_4915,In_406,In_916);
nor U4916 (N_4916,In_905,In_161);
and U4917 (N_4917,In_949,In_134);
and U4918 (N_4918,In_855,In_718);
nand U4919 (N_4919,In_891,In_124);
or U4920 (N_4920,In_286,In_763);
and U4921 (N_4921,In_974,In_689);
nor U4922 (N_4922,In_896,In_920);
xnor U4923 (N_4923,In_930,In_810);
and U4924 (N_4924,In_586,In_636);
or U4925 (N_4925,In_612,In_556);
or U4926 (N_4926,In_587,In_116);
or U4927 (N_4927,In_183,In_139);
or U4928 (N_4928,In_219,In_477);
nor U4929 (N_4929,In_876,In_739);
nand U4930 (N_4930,In_759,In_34);
nor U4931 (N_4931,In_184,In_995);
and U4932 (N_4932,In_639,In_243);
or U4933 (N_4933,In_546,In_874);
and U4934 (N_4934,In_149,In_545);
nand U4935 (N_4935,In_622,In_232);
nand U4936 (N_4936,In_134,In_768);
or U4937 (N_4937,In_216,In_237);
nand U4938 (N_4938,In_218,In_532);
or U4939 (N_4939,In_862,In_978);
or U4940 (N_4940,In_449,In_107);
and U4941 (N_4941,In_438,In_24);
nor U4942 (N_4942,In_747,In_354);
nand U4943 (N_4943,In_571,In_613);
nand U4944 (N_4944,In_792,In_851);
nor U4945 (N_4945,In_286,In_997);
nor U4946 (N_4946,In_111,In_696);
xnor U4947 (N_4947,In_166,In_566);
nand U4948 (N_4948,In_950,In_589);
or U4949 (N_4949,In_702,In_344);
nor U4950 (N_4950,In_898,In_983);
xnor U4951 (N_4951,In_924,In_93);
nand U4952 (N_4952,In_366,In_531);
nor U4953 (N_4953,In_648,In_909);
nor U4954 (N_4954,In_695,In_136);
or U4955 (N_4955,In_298,In_685);
nor U4956 (N_4956,In_189,In_861);
nor U4957 (N_4957,In_880,In_17);
and U4958 (N_4958,In_380,In_102);
or U4959 (N_4959,In_222,In_799);
nand U4960 (N_4960,In_354,In_549);
nor U4961 (N_4961,In_619,In_422);
or U4962 (N_4962,In_884,In_323);
and U4963 (N_4963,In_676,In_637);
or U4964 (N_4964,In_392,In_658);
and U4965 (N_4965,In_10,In_997);
nor U4966 (N_4966,In_508,In_15);
or U4967 (N_4967,In_311,In_556);
nand U4968 (N_4968,In_189,In_682);
nand U4969 (N_4969,In_891,In_938);
nor U4970 (N_4970,In_600,In_104);
nand U4971 (N_4971,In_647,In_548);
nor U4972 (N_4972,In_261,In_926);
or U4973 (N_4973,In_590,In_48);
nand U4974 (N_4974,In_834,In_593);
xnor U4975 (N_4975,In_792,In_351);
or U4976 (N_4976,In_901,In_47);
and U4977 (N_4977,In_731,In_836);
and U4978 (N_4978,In_389,In_84);
nand U4979 (N_4979,In_837,In_778);
xor U4980 (N_4980,In_49,In_654);
nor U4981 (N_4981,In_346,In_638);
nor U4982 (N_4982,In_918,In_497);
or U4983 (N_4983,In_222,In_678);
or U4984 (N_4984,In_908,In_571);
or U4985 (N_4985,In_143,In_431);
nor U4986 (N_4986,In_773,In_653);
and U4987 (N_4987,In_364,In_828);
or U4988 (N_4988,In_865,In_598);
and U4989 (N_4989,In_118,In_413);
nand U4990 (N_4990,In_654,In_469);
nand U4991 (N_4991,In_495,In_394);
or U4992 (N_4992,In_478,In_439);
nand U4993 (N_4993,In_917,In_605);
nand U4994 (N_4994,In_866,In_540);
nor U4995 (N_4995,In_37,In_319);
xor U4996 (N_4996,In_156,In_640);
and U4997 (N_4997,In_430,In_358);
nand U4998 (N_4998,In_781,In_514);
and U4999 (N_4999,In_874,In_325);
or U5000 (N_5000,N_323,N_4533);
nand U5001 (N_5001,N_2223,N_3971);
and U5002 (N_5002,N_1851,N_4395);
and U5003 (N_5003,N_4570,N_286);
nand U5004 (N_5004,N_3771,N_4610);
or U5005 (N_5005,N_1435,N_1193);
and U5006 (N_5006,N_3639,N_2291);
and U5007 (N_5007,N_766,N_4902);
and U5008 (N_5008,N_4816,N_538);
xor U5009 (N_5009,N_3592,N_4225);
and U5010 (N_5010,N_2415,N_652);
or U5011 (N_5011,N_2327,N_2626);
nor U5012 (N_5012,N_4964,N_3661);
nand U5013 (N_5013,N_3527,N_3922);
or U5014 (N_5014,N_2780,N_2219);
and U5015 (N_5015,N_759,N_680);
nand U5016 (N_5016,N_1198,N_2154);
nor U5017 (N_5017,N_172,N_3052);
nand U5018 (N_5018,N_3786,N_3295);
nand U5019 (N_5019,N_1544,N_1499);
nor U5020 (N_5020,N_902,N_712);
and U5021 (N_5021,N_3127,N_2323);
or U5022 (N_5022,N_3243,N_1052);
nor U5023 (N_5023,N_3921,N_825);
nor U5024 (N_5024,N_103,N_3703);
nand U5025 (N_5025,N_1809,N_4996);
nand U5026 (N_5026,N_4532,N_4763);
nor U5027 (N_5027,N_3718,N_986);
or U5028 (N_5028,N_1322,N_3851);
or U5029 (N_5029,N_3335,N_3100);
or U5030 (N_5030,N_4809,N_3827);
nand U5031 (N_5031,N_1192,N_1055);
and U5032 (N_5032,N_198,N_4681);
and U5033 (N_5033,N_581,N_2893);
nor U5034 (N_5034,N_4264,N_2143);
or U5035 (N_5035,N_2700,N_1961);
nor U5036 (N_5036,N_4486,N_2258);
nor U5037 (N_5037,N_266,N_3445);
nor U5038 (N_5038,N_2837,N_608);
nand U5039 (N_5039,N_3858,N_4590);
and U5040 (N_5040,N_4620,N_1229);
nand U5041 (N_5041,N_3466,N_2277);
nor U5042 (N_5042,N_350,N_1995);
nor U5043 (N_5043,N_301,N_456);
and U5044 (N_5044,N_1692,N_4981);
and U5045 (N_5045,N_3524,N_1076);
and U5046 (N_5046,N_2884,N_1420);
nor U5047 (N_5047,N_2553,N_2040);
nand U5048 (N_5048,N_10,N_3753);
nor U5049 (N_5049,N_522,N_158);
or U5050 (N_5050,N_4668,N_3382);
nor U5051 (N_5051,N_4934,N_4725);
or U5052 (N_5052,N_2688,N_3724);
nor U5053 (N_5053,N_3435,N_566);
nand U5054 (N_5054,N_838,N_3679);
nand U5055 (N_5055,N_104,N_1265);
and U5056 (N_5056,N_4276,N_3772);
and U5057 (N_5057,N_2345,N_1459);
or U5058 (N_5058,N_474,N_4596);
and U5059 (N_5059,N_720,N_46);
nor U5060 (N_5060,N_796,N_713);
and U5061 (N_5061,N_4552,N_3650);
or U5062 (N_5062,N_1138,N_4207);
nor U5063 (N_5063,N_130,N_2580);
or U5064 (N_5064,N_683,N_2081);
nor U5065 (N_5065,N_11,N_2481);
and U5066 (N_5066,N_1820,N_3239);
and U5067 (N_5067,N_917,N_2319);
or U5068 (N_5068,N_2589,N_2850);
nand U5069 (N_5069,N_4961,N_4321);
nor U5070 (N_5070,N_3627,N_2233);
or U5071 (N_5071,N_1136,N_2075);
and U5072 (N_5072,N_879,N_1253);
or U5073 (N_5073,N_3265,N_2925);
and U5074 (N_5074,N_1795,N_3492);
nor U5075 (N_5075,N_2887,N_2587);
or U5076 (N_5076,N_4257,N_3051);
and U5077 (N_5077,N_3220,N_189);
nand U5078 (N_5078,N_1838,N_3958);
or U5079 (N_5079,N_4699,N_4953);
nor U5080 (N_5080,N_1894,N_1911);
nor U5081 (N_5081,N_1555,N_4930);
nor U5082 (N_5082,N_2696,N_924);
and U5083 (N_5083,N_2875,N_1454);
nand U5084 (N_5084,N_3904,N_4513);
nor U5085 (N_5085,N_767,N_654);
or U5086 (N_5086,N_1977,N_963);
or U5087 (N_5087,N_3881,N_3934);
nand U5088 (N_5088,N_3636,N_386);
or U5089 (N_5089,N_578,N_2509);
nand U5090 (N_5090,N_4737,N_2866);
nand U5091 (N_5091,N_513,N_1205);
nand U5092 (N_5092,N_2654,N_3195);
and U5093 (N_5093,N_4982,N_1842);
and U5094 (N_5094,N_3874,N_2176);
and U5095 (N_5095,N_4866,N_3551);
nor U5096 (N_5096,N_75,N_3966);
and U5097 (N_5097,N_2982,N_2877);
or U5098 (N_5098,N_4020,N_131);
or U5099 (N_5099,N_3537,N_2769);
nor U5100 (N_5100,N_3652,N_2969);
and U5101 (N_5101,N_4447,N_1788);
nand U5102 (N_5102,N_2214,N_4634);
or U5103 (N_5103,N_1216,N_4550);
and U5104 (N_5104,N_1955,N_1509);
nand U5105 (N_5105,N_4506,N_2241);
and U5106 (N_5106,N_1108,N_157);
or U5107 (N_5107,N_4661,N_1690);
xor U5108 (N_5108,N_1916,N_4966);
nand U5109 (N_5109,N_1935,N_1092);
and U5110 (N_5110,N_4178,N_2380);
nor U5111 (N_5111,N_3436,N_2301);
or U5112 (N_5112,N_4925,N_3569);
and U5113 (N_5113,N_4921,N_912);
nor U5114 (N_5114,N_4038,N_1744);
and U5115 (N_5115,N_316,N_3873);
nor U5116 (N_5116,N_3259,N_4793);
and U5117 (N_5117,N_1739,N_4988);
nor U5118 (N_5118,N_1208,N_1080);
and U5119 (N_5119,N_1440,N_3326);
or U5120 (N_5120,N_3473,N_3043);
nand U5121 (N_5121,N_987,N_2104);
and U5122 (N_5122,N_3015,N_2604);
or U5123 (N_5123,N_641,N_1834);
or U5124 (N_5124,N_2201,N_251);
or U5125 (N_5125,N_2285,N_2934);
nand U5126 (N_5126,N_4086,N_2399);
nor U5127 (N_5127,N_1402,N_3993);
and U5128 (N_5128,N_2191,N_111);
nand U5129 (N_5129,N_4489,N_2713);
and U5130 (N_5130,N_1112,N_2039);
nand U5131 (N_5131,N_508,N_4161);
nor U5132 (N_5132,N_4419,N_1036);
nand U5133 (N_5133,N_3625,N_4567);
or U5134 (N_5134,N_4312,N_2076);
or U5135 (N_5135,N_1389,N_4108);
nor U5136 (N_5136,N_2365,N_592);
and U5137 (N_5137,N_3893,N_3228);
nor U5138 (N_5138,N_4865,N_109);
or U5139 (N_5139,N_660,N_4530);
nor U5140 (N_5140,N_1237,N_2245);
nor U5141 (N_5141,N_3684,N_2375);
or U5142 (N_5142,N_4787,N_3790);
or U5143 (N_5143,N_6,N_1829);
and U5144 (N_5144,N_1832,N_1156);
nand U5145 (N_5145,N_2976,N_3188);
nor U5146 (N_5146,N_4650,N_2111);
nand U5147 (N_5147,N_4526,N_2356);
nand U5148 (N_5148,N_4559,N_3321);
and U5149 (N_5149,N_3540,N_2647);
nand U5150 (N_5150,N_4114,N_1965);
or U5151 (N_5151,N_3235,N_848);
nor U5152 (N_5152,N_476,N_2282);
and U5153 (N_5153,N_2494,N_4511);
or U5154 (N_5154,N_1494,N_2648);
and U5155 (N_5155,N_3489,N_3419);
and U5156 (N_5156,N_4329,N_2435);
and U5157 (N_5157,N_2198,N_1094);
and U5158 (N_5158,N_2612,N_840);
nand U5159 (N_5159,N_2489,N_139);
nor U5160 (N_5160,N_1053,N_1316);
or U5161 (N_5161,N_1849,N_528);
and U5162 (N_5162,N_2359,N_2185);
and U5163 (N_5163,N_2159,N_1321);
xor U5164 (N_5164,N_971,N_145);
or U5165 (N_5165,N_2086,N_1817);
or U5166 (N_5166,N_404,N_588);
or U5167 (N_5167,N_2928,N_2473);
nor U5168 (N_5168,N_1147,N_1014);
and U5169 (N_5169,N_1644,N_2789);
nand U5170 (N_5170,N_3481,N_3504);
and U5171 (N_5171,N_2472,N_3111);
and U5172 (N_5172,N_3856,N_3078);
and U5173 (N_5173,N_1331,N_3596);
and U5174 (N_5174,N_4367,N_2361);
nor U5175 (N_5175,N_1275,N_2052);
and U5176 (N_5176,N_4818,N_2657);
or U5177 (N_5177,N_2635,N_4980);
nand U5178 (N_5178,N_1283,N_2243);
or U5179 (N_5179,N_471,N_579);
nand U5180 (N_5180,N_589,N_3460);
nand U5181 (N_5181,N_2994,N_3886);
nand U5182 (N_5182,N_4261,N_877);
and U5183 (N_5183,N_4602,N_320);
and U5184 (N_5184,N_4971,N_2582);
or U5185 (N_5185,N_1641,N_2265);
or U5186 (N_5186,N_1693,N_2448);
nand U5187 (N_5187,N_1179,N_2645);
and U5188 (N_5188,N_2715,N_485);
nand U5189 (N_5189,N_1380,N_3072);
nor U5190 (N_5190,N_1632,N_2339);
nor U5191 (N_5191,N_321,N_2248);
and U5192 (N_5192,N_4735,N_105);
nor U5193 (N_5193,N_1287,N_3119);
nor U5194 (N_5194,N_1490,N_3941);
nor U5195 (N_5195,N_3680,N_1844);
and U5196 (N_5196,N_2605,N_2961);
and U5197 (N_5197,N_858,N_1352);
or U5198 (N_5198,N_3096,N_3741);
nor U5199 (N_5199,N_752,N_3699);
and U5200 (N_5200,N_3142,N_4722);
or U5201 (N_5201,N_4515,N_3270);
or U5202 (N_5202,N_2337,N_4473);
nand U5203 (N_5203,N_1850,N_1363);
nand U5204 (N_5204,N_607,N_1586);
and U5205 (N_5205,N_4888,N_1706);
nand U5206 (N_5206,N_2406,N_3732);
nand U5207 (N_5207,N_1631,N_4327);
and U5208 (N_5208,N_1681,N_3638);
or U5209 (N_5209,N_2574,N_1127);
nor U5210 (N_5210,N_356,N_1449);
nor U5211 (N_5211,N_110,N_3773);
nand U5212 (N_5212,N_2662,N_3211);
or U5213 (N_5213,N_4783,N_1302);
nand U5214 (N_5214,N_2876,N_2712);
and U5215 (N_5215,N_951,N_4917);
nand U5216 (N_5216,N_1636,N_4767);
nor U5217 (N_5217,N_4652,N_3484);
or U5218 (N_5218,N_751,N_1379);
nor U5219 (N_5219,N_3510,N_4043);
and U5220 (N_5220,N_1304,N_1679);
nor U5221 (N_5221,N_3494,N_373);
nand U5222 (N_5222,N_2687,N_4179);
nor U5223 (N_5223,N_302,N_353);
and U5224 (N_5224,N_954,N_3044);
or U5225 (N_5225,N_4688,N_2240);
xor U5226 (N_5226,N_2911,N_3809);
and U5227 (N_5227,N_364,N_4854);
xor U5228 (N_5228,N_1333,N_4837);
nor U5229 (N_5229,N_1819,N_31);
or U5230 (N_5230,N_1174,N_1335);
nand U5231 (N_5231,N_1723,N_4910);
nor U5232 (N_5232,N_583,N_2121);
or U5233 (N_5233,N_4153,N_2409);
and U5234 (N_5234,N_996,N_3173);
nor U5235 (N_5235,N_4280,N_4840);
nor U5236 (N_5236,N_1295,N_2077);
or U5237 (N_5237,N_814,N_299);
and U5238 (N_5238,N_2331,N_3683);
nand U5239 (N_5239,N_3148,N_361);
xnor U5240 (N_5240,N_3869,N_453);
and U5241 (N_5241,N_257,N_775);
xnor U5242 (N_5242,N_3159,N_1922);
nand U5243 (N_5243,N_574,N_953);
nand U5244 (N_5244,N_4100,N_4899);
nand U5245 (N_5245,N_669,N_4549);
nor U5246 (N_5246,N_4831,N_1667);
and U5247 (N_5247,N_239,N_650);
nor U5248 (N_5248,N_362,N_4968);
nand U5249 (N_5249,N_406,N_154);
or U5250 (N_5250,N_290,N_2346);
nand U5251 (N_5251,N_3553,N_4868);
nand U5252 (N_5252,N_2905,N_3859);
or U5253 (N_5253,N_4090,N_4588);
and U5254 (N_5254,N_483,N_2002);
nor U5255 (N_5255,N_4702,N_212);
and U5256 (N_5256,N_2368,N_2396);
or U5257 (N_5257,N_1538,N_283);
nor U5258 (N_5258,N_1478,N_901);
and U5259 (N_5259,N_1529,N_494);
and U5260 (N_5260,N_423,N_211);
or U5261 (N_5261,N_4838,N_3758);
xor U5262 (N_5262,N_1060,N_1884);
or U5263 (N_5263,N_4449,N_2095);
or U5264 (N_5264,N_4617,N_4580);
nand U5265 (N_5265,N_2413,N_2089);
and U5266 (N_5266,N_2996,N_2990);
nand U5267 (N_5267,N_837,N_1178);
nor U5268 (N_5268,N_908,N_4605);
nand U5269 (N_5269,N_609,N_2617);
nor U5270 (N_5270,N_1516,N_4244);
and U5271 (N_5271,N_2385,N_3590);
and U5272 (N_5272,N_465,N_4524);
and U5273 (N_5273,N_2782,N_4529);
nor U5274 (N_5274,N_950,N_3544);
nor U5275 (N_5275,N_4879,N_4216);
nand U5276 (N_5276,N_1983,N_2513);
and U5277 (N_5277,N_401,N_4538);
and U5278 (N_5278,N_2535,N_2309);
nand U5279 (N_5279,N_761,N_533);
or U5280 (N_5280,N_2493,N_3244);
nor U5281 (N_5281,N_129,N_325);
nor U5282 (N_5282,N_3141,N_4135);
and U5283 (N_5283,N_454,N_3047);
nand U5284 (N_5284,N_3055,N_3765);
nand U5285 (N_5285,N_1040,N_3721);
and U5286 (N_5286,N_3775,N_4162);
and U5287 (N_5287,N_624,N_287);
and U5288 (N_5288,N_1135,N_3417);
nor U5289 (N_5289,N_1467,N_1642);
or U5290 (N_5290,N_2232,N_4006);
or U5291 (N_5291,N_1630,N_976);
nor U5292 (N_5292,N_3712,N_183);
or U5293 (N_5293,N_2844,N_4046);
nand U5294 (N_5294,N_155,N_3645);
and U5295 (N_5295,N_4491,N_4633);
nor U5296 (N_5296,N_584,N_2292);
or U5297 (N_5297,N_3898,N_3156);
or U5298 (N_5298,N_2998,N_3343);
or U5299 (N_5299,N_2175,N_1255);
nor U5300 (N_5300,N_4231,N_351);
and U5301 (N_5301,N_726,N_645);
and U5302 (N_5302,N_106,N_1541);
or U5303 (N_5303,N_3564,N_330);
and U5304 (N_5304,N_4670,N_1430);
nor U5305 (N_5305,N_206,N_2886);
or U5306 (N_5306,N_4527,N_1107);
nor U5307 (N_5307,N_4240,N_4846);
nand U5308 (N_5308,N_3969,N_3375);
or U5309 (N_5309,N_1896,N_4909);
nand U5310 (N_5310,N_101,N_696);
and U5311 (N_5311,N_2507,N_3810);
nand U5312 (N_5312,N_3012,N_2357);
nor U5313 (N_5313,N_3928,N_3023);
and U5314 (N_5314,N_4640,N_2296);
nor U5315 (N_5315,N_1220,N_3536);
nor U5316 (N_5316,N_4753,N_2078);
and U5317 (N_5317,N_572,N_787);
nand U5318 (N_5318,N_815,N_2314);
and U5319 (N_5319,N_506,N_2421);
or U5320 (N_5320,N_570,N_3013);
nand U5321 (N_5321,N_3065,N_4628);
nand U5322 (N_5322,N_3199,N_1370);
or U5323 (N_5323,N_4371,N_4101);
nand U5324 (N_5324,N_745,N_1292);
nor U5325 (N_5325,N_295,N_1562);
nand U5326 (N_5326,N_2907,N_3622);
nor U5327 (N_5327,N_1276,N_3629);
or U5328 (N_5328,N_3046,N_2006);
nand U5329 (N_5329,N_4305,N_399);
nand U5330 (N_5330,N_3264,N_2831);
nand U5331 (N_5331,N_4345,N_1900);
nor U5332 (N_5332,N_2788,N_1123);
xnor U5333 (N_5333,N_1593,N_2458);
and U5334 (N_5334,N_4998,N_4461);
nor U5335 (N_5335,N_276,N_1452);
and U5336 (N_5336,N_345,N_2622);
nor U5337 (N_5337,N_4779,N_582);
nand U5338 (N_5338,N_4476,N_892);
or U5339 (N_5339,N_4756,N_2817);
xor U5340 (N_5340,N_4875,N_4484);
nand U5341 (N_5341,N_419,N_2059);
xor U5342 (N_5342,N_2600,N_4587);
nand U5343 (N_5343,N_4102,N_383);
and U5344 (N_5344,N_4156,N_1155);
nand U5345 (N_5345,N_4245,N_4845);
xnor U5346 (N_5346,N_1421,N_1305);
or U5347 (N_5347,N_484,N_4521);
nor U5348 (N_5348,N_3694,N_4896);
nand U5349 (N_5349,N_4978,N_4157);
nor U5350 (N_5350,N_1576,N_1139);
nor U5351 (N_5351,N_1588,N_2678);
or U5352 (N_5352,N_2860,N_2354);
nand U5353 (N_5353,N_1129,N_3509);
and U5354 (N_5354,N_4855,N_1062);
or U5355 (N_5355,N_3177,N_4770);
nand U5356 (N_5356,N_3578,N_3942);
and U5357 (N_5357,N_2592,N_244);
and U5358 (N_5358,N_442,N_1406);
and U5359 (N_5359,N_2401,N_3533);
or U5360 (N_5360,N_121,N_1724);
or U5361 (N_5361,N_605,N_2461);
or U5362 (N_5362,N_3946,N_4184);
and U5363 (N_5363,N_2505,N_1584);
nor U5364 (N_5364,N_2315,N_2169);
nor U5365 (N_5365,N_1793,N_4174);
nor U5366 (N_5366,N_1514,N_190);
or U5367 (N_5367,N_3022,N_2366);
and U5368 (N_5368,N_236,N_2583);
and U5369 (N_5369,N_3085,N_2064);
nand U5370 (N_5370,N_4922,N_2390);
nand U5371 (N_5371,N_729,N_4457);
or U5372 (N_5372,N_870,N_4915);
or U5373 (N_5373,N_3833,N_4121);
nor U5374 (N_5374,N_2351,N_2548);
nor U5375 (N_5375,N_4347,N_2667);
nor U5376 (N_5376,N_4332,N_1273);
or U5377 (N_5377,N_2441,N_1749);
nand U5378 (N_5378,N_2872,N_3174);
nand U5379 (N_5379,N_2668,N_667);
and U5380 (N_5380,N_3550,N_2275);
nor U5381 (N_5381,N_4171,N_770);
or U5382 (N_5382,N_391,N_3296);
nor U5383 (N_5383,N_1117,N_4819);
and U5384 (N_5384,N_365,N_2839);
nor U5385 (N_5385,N_2773,N_1391);
or U5386 (N_5386,N_1807,N_4657);
or U5387 (N_5387,N_2761,N_2230);
nor U5388 (N_5388,N_2063,N_4301);
or U5389 (N_5389,N_3194,N_3572);
nor U5390 (N_5390,N_916,N_1968);
or U5391 (N_5391,N_4230,N_1225);
or U5392 (N_5392,N_1511,N_2312);
or U5393 (N_5393,N_3291,N_4897);
or U5394 (N_5394,N_3463,N_2332);
nor U5395 (N_5395,N_1912,N_396);
nand U5396 (N_5396,N_1470,N_4589);
nand U5397 (N_5397,N_3866,N_2974);
nor U5398 (N_5398,N_2829,N_740);
and U5399 (N_5399,N_4708,N_4166);
nand U5400 (N_5400,N_3108,N_3995);
nand U5401 (N_5401,N_4864,N_1007);
and U5402 (N_5402,N_4984,N_3181);
nor U5403 (N_5403,N_220,N_4732);
or U5404 (N_5404,N_615,N_4357);
nand U5405 (N_5405,N_1560,N_1134);
nor U5406 (N_5406,N_926,N_4124);
and U5407 (N_5407,N_2041,N_1589);
nor U5408 (N_5408,N_1564,N_4268);
nand U5409 (N_5409,N_3426,N_3031);
and U5410 (N_5410,N_899,N_1426);
and U5411 (N_5411,N_2335,N_1003);
nor U5412 (N_5412,N_4213,N_191);
nor U5413 (N_5413,N_4493,N_3021);
or U5414 (N_5414,N_1171,N_3113);
or U5415 (N_5415,N_644,N_448);
nor U5416 (N_5416,N_4409,N_990);
and U5417 (N_5417,N_1034,N_4727);
or U5418 (N_5418,N_4531,N_3899);
nand U5419 (N_5419,N_946,N_2074);
or U5420 (N_5420,N_4675,N_1557);
and U5421 (N_5421,N_1823,N_1072);
nand U5422 (N_5422,N_4678,N_1378);
nand U5423 (N_5423,N_4349,N_473);
nor U5424 (N_5424,N_4941,N_1468);
or U5425 (N_5425,N_3016,N_2062);
or U5426 (N_5426,N_468,N_784);
and U5427 (N_5427,N_4009,N_1340);
and U5428 (N_5428,N_2393,N_1689);
or U5429 (N_5429,N_1095,N_2695);
or U5430 (N_5430,N_59,N_4389);
and U5431 (N_5431,N_2950,N_2656);
nor U5432 (N_5432,N_2272,N_3954);
and U5433 (N_5433,N_4949,N_3777);
or U5434 (N_5434,N_2068,N_1732);
nand U5435 (N_5435,N_1387,N_3372);
or U5436 (N_5436,N_1802,N_2577);
and U5437 (N_5437,N_1424,N_2171);
and U5438 (N_5438,N_2707,N_2324);
nor U5439 (N_5439,N_3400,N_3011);
or U5440 (N_5440,N_3176,N_4458);
and U5441 (N_5441,N_2405,N_822);
or U5442 (N_5442,N_4674,N_3430);
or U5443 (N_5443,N_2593,N_2889);
and U5444 (N_5444,N_807,N_2871);
nor U5445 (N_5445,N_359,N_1567);
or U5446 (N_5446,N_50,N_1423);
nand U5447 (N_5447,N_3682,N_865);
nor U5448 (N_5448,N_972,N_467);
nor U5449 (N_5449,N_3449,N_4800);
nand U5450 (N_5450,N_2985,N_1745);
nand U5451 (N_5451,N_2578,N_2892);
and U5452 (N_5452,N_3088,N_1175);
nand U5453 (N_5453,N_1601,N_1290);
and U5454 (N_5454,N_1960,N_213);
nand U5455 (N_5455,N_4606,N_2417);
or U5456 (N_5456,N_2027,N_1608);
nor U5457 (N_5457,N_4739,N_492);
and U5458 (N_5458,N_3948,N_2910);
nand U5459 (N_5459,N_335,N_1358);
or U5460 (N_5460,N_3431,N_1778);
or U5461 (N_5461,N_1988,N_1569);
and U5462 (N_5462,N_1212,N_61);
nor U5463 (N_5463,N_2420,N_4133);
or U5464 (N_5464,N_1133,N_262);
nor U5465 (N_5465,N_3480,N_2038);
and U5466 (N_5466,N_4362,N_2188);
nor U5467 (N_5467,N_1224,N_1393);
nor U5468 (N_5468,N_2763,N_3709);
xnor U5469 (N_5469,N_2070,N_1978);
and U5470 (N_5470,N_3989,N_2200);
and U5471 (N_5471,N_3464,N_4907);
and U5472 (N_5472,N_2946,N_2597);
and U5473 (N_5473,N_4760,N_2128);
nand U5474 (N_5474,N_3266,N_4631);
and U5475 (N_5475,N_3618,N_2726);
and U5476 (N_5476,N_3428,N_1365);
and U5477 (N_5477,N_3249,N_161);
and U5478 (N_5478,N_2785,N_4612);
or U5479 (N_5479,N_510,N_3322);
and U5480 (N_5480,N_137,N_2845);
nor U5481 (N_5481,N_2491,N_4297);
or U5482 (N_5482,N_2503,N_2674);
and U5483 (N_5483,N_2757,N_2533);
or U5484 (N_5484,N_1130,N_3965);
or U5485 (N_5485,N_888,N_306);
nor U5486 (N_5486,N_3861,N_1185);
xnor U5487 (N_5487,N_2919,N_1312);
nor U5488 (N_5488,N_1323,N_3017);
or U5489 (N_5489,N_4940,N_4972);
or U5490 (N_5490,N_3956,N_2187);
nand U5491 (N_5491,N_3662,N_3062);
xnor U5492 (N_5492,N_1017,N_3277);
or U5493 (N_5493,N_4554,N_2897);
nand U5494 (N_5494,N_2774,N_3057);
nand U5495 (N_5495,N_4698,N_4481);
nor U5496 (N_5496,N_1417,N_1361);
or U5497 (N_5497,N_4499,N_3961);
nor U5498 (N_5498,N_1833,N_4169);
nand U5499 (N_5499,N_2289,N_670);
or U5500 (N_5500,N_202,N_2403);
nor U5501 (N_5501,N_3700,N_3045);
and U5502 (N_5502,N_4067,N_4561);
or U5503 (N_5503,N_2935,N_2815);
nand U5504 (N_5504,N_1513,N_1846);
nand U5505 (N_5505,N_4298,N_4711);
and U5506 (N_5506,N_4873,N_1585);
or U5507 (N_5507,N_3754,N_743);
nor U5508 (N_5508,N_3900,N_1750);
and U5509 (N_5509,N_1571,N_34);
and U5510 (N_5510,N_2975,N_417);
and U5511 (N_5511,N_2849,N_3325);
and U5512 (N_5512,N_1686,N_4065);
nand U5513 (N_5513,N_3929,N_4308);
or U5514 (N_5514,N_1448,N_478);
or U5515 (N_5515,N_1238,N_433);
and U5516 (N_5516,N_3496,N_547);
nor U5517 (N_5517,N_3102,N_3654);
or U5518 (N_5518,N_411,N_4403);
nand U5519 (N_5519,N_4189,N_974);
or U5520 (N_5520,N_343,N_3497);
or U5521 (N_5521,N_3482,N_117);
nor U5522 (N_5522,N_2960,N_1498);
nor U5523 (N_5523,N_3870,N_371);
nand U5524 (N_5524,N_4718,N_4959);
or U5525 (N_5525,N_2212,N_119);
nor U5526 (N_5526,N_1720,N_1103);
nand U5527 (N_5527,N_1675,N_1455);
nand U5528 (N_5528,N_2167,N_2449);
or U5529 (N_5529,N_4017,N_830);
and U5530 (N_5530,N_1969,N_4255);
nand U5531 (N_5531,N_2926,N_2521);
xor U5532 (N_5532,N_1051,N_4045);
nand U5533 (N_5533,N_3631,N_3548);
or U5534 (N_5534,N_918,N_2098);
nand U5535 (N_5535,N_1970,N_4049);
nor U5536 (N_5536,N_2488,N_760);
nor U5537 (N_5537,N_3788,N_4714);
nand U5538 (N_5538,N_3147,N_517);
or U5539 (N_5539,N_3744,N_1240);
nand U5540 (N_5540,N_2462,N_4285);
nand U5541 (N_5541,N_208,N_2463);
and U5542 (N_5542,N_2318,N_2023);
or U5543 (N_5543,N_4195,N_2701);
and U5544 (N_5544,N_764,N_2271);
or U5545 (N_5545,N_133,N_628);
nor U5546 (N_5546,N_2444,N_1396);
or U5547 (N_5547,N_836,N_2666);
nor U5548 (N_5548,N_721,N_3469);
nand U5549 (N_5549,N_3979,N_998);
nand U5550 (N_5550,N_2947,N_616);
or U5551 (N_5551,N_1432,N_2353);
xor U5552 (N_5552,N_832,N_2863);
and U5553 (N_5553,N_4600,N_1474);
or U5554 (N_5554,N_1554,N_2246);
or U5555 (N_5555,N_3443,N_461);
or U5556 (N_5556,N_493,N_1303);
or U5557 (N_5557,N_757,N_735);
nor U5558 (N_5558,N_4918,N_1187);
or U5559 (N_5559,N_540,N_1572);
and U5560 (N_5560,N_2754,N_4262);
and U5561 (N_5561,N_731,N_1518);
or U5562 (N_5562,N_4740,N_173);
and U5563 (N_5563,N_1372,N_1484);
nor U5564 (N_5564,N_868,N_671);
and U5565 (N_5565,N_1173,N_2534);
or U5566 (N_5566,N_587,N_748);
nand U5567 (N_5567,N_95,N_3158);
nor U5568 (N_5568,N_252,N_3232);
nor U5569 (N_5569,N_415,N_1451);
and U5570 (N_5570,N_4089,N_52);
nor U5571 (N_5571,N_1409,N_2793);
nor U5572 (N_5572,N_4762,N_30);
or U5573 (N_5573,N_3038,N_2014);
nand U5574 (N_5574,N_3319,N_4843);
nand U5575 (N_5575,N_613,N_68);
nand U5576 (N_5576,N_2652,N_1169);
nor U5577 (N_5577,N_2007,N_2705);
nand U5578 (N_5578,N_3075,N_3442);
nand U5579 (N_5579,N_3723,N_1716);
nor U5580 (N_5580,N_3283,N_1441);
and U5581 (N_5581,N_4785,N_2655);
nand U5582 (N_5582,N_4278,N_3454);
nor U5583 (N_5583,N_4097,N_529);
nand U5584 (N_5584,N_4051,N_834);
or U5585 (N_5585,N_962,N_2730);
and U5586 (N_5586,N_4,N_4111);
nand U5587 (N_5587,N_4397,N_4094);
and U5588 (N_5588,N_3799,N_3560);
nor U5589 (N_5589,N_1116,N_2954);
or U5590 (N_5590,N_717,N_3121);
xor U5591 (N_5591,N_3635,N_3475);
or U5592 (N_5592,N_1599,N_1839);
and U5593 (N_5593,N_1010,N_2195);
and U5594 (N_5594,N_440,N_1756);
or U5595 (N_5595,N_3289,N_618);
nor U5596 (N_5596,N_518,N_3425);
nor U5597 (N_5597,N_1531,N_369);
or U5598 (N_5598,N_1915,N_3290);
or U5599 (N_5599,N_4326,N_773);
nor U5600 (N_5600,N_1154,N_32);
nor U5601 (N_5601,N_867,N_2085);
nand U5602 (N_5602,N_754,N_1677);
or U5603 (N_5603,N_1759,N_3707);
nor U5604 (N_5604,N_3479,N_4754);
nand U5605 (N_5605,N_4542,N_1354);
nor U5606 (N_5606,N_1221,N_2790);
and U5607 (N_5607,N_758,N_2523);
nand U5608 (N_5608,N_1609,N_1157);
nor U5609 (N_5609,N_1835,N_324);
nor U5610 (N_5610,N_2407,N_1067);
or U5611 (N_5611,N_966,N_4242);
nor U5612 (N_5612,N_4342,N_4296);
nor U5613 (N_5613,N_4556,N_4713);
or U5614 (N_5614,N_563,N_4586);
nor U5615 (N_5615,N_2942,N_3915);
or U5616 (N_5616,N_4019,N_1923);
and U5617 (N_5617,N_2722,N_1122);
nand U5618 (N_5618,N_3233,N_3160);
and U5619 (N_5619,N_3186,N_3365);
nand U5620 (N_5620,N_4050,N_4435);
and U5621 (N_5621,N_2364,N_4175);
nand U5622 (N_5622,N_4647,N_2288);
nand U5623 (N_5623,N_1289,N_3151);
and U5624 (N_5624,N_2336,N_968);
nor U5625 (N_5625,N_2854,N_604);
or U5626 (N_5626,N_4537,N_1056);
nor U5627 (N_5627,N_1326,N_2226);
and U5628 (N_5628,N_3913,N_835);
or U5629 (N_5629,N_3844,N_496);
and U5630 (N_5630,N_4394,N_2970);
nand U5631 (N_5631,N_3378,N_1465);
nand U5632 (N_5632,N_2870,N_3923);
nor U5633 (N_5633,N_1114,N_3747);
xnor U5634 (N_5634,N_3669,N_1903);
nor U5635 (N_5635,N_4126,N_2962);
or U5636 (N_5636,N_3397,N_3513);
nor U5637 (N_5637,N_4286,N_3814);
nand U5638 (N_5638,N_408,N_3672);
nand U5639 (N_5639,N_2846,N_4503);
and U5640 (N_5640,N_4813,N_2644);
nor U5641 (N_5641,N_3191,N_3685);
or U5642 (N_5642,N_3376,N_26);
nand U5643 (N_5643,N_4683,N_2181);
nand U5644 (N_5644,N_3617,N_1942);
and U5645 (N_5645,N_446,N_4113);
and U5646 (N_5646,N_2832,N_3568);
nand U5647 (N_5647,N_363,N_519);
or U5648 (N_5648,N_1574,N_1497);
and U5649 (N_5649,N_2620,N_2218);
or U5650 (N_5650,N_1073,N_1867);
nand U5651 (N_5651,N_4035,N_4096);
nand U5652 (N_5652,N_4354,N_2123);
nand U5653 (N_5653,N_3600,N_2260);
and U5654 (N_5654,N_4891,N_3920);
and U5655 (N_5655,N_4939,N_3697);
or U5656 (N_5656,N_3642,N_2504);
and U5657 (N_5657,N_4350,N_39);
nand U5658 (N_5658,N_2333,N_3668);
nor U5659 (N_5659,N_2018,N_1740);
nor U5660 (N_5660,N_2882,N_1652);
or U5661 (N_5661,N_2009,N_4877);
nand U5662 (N_5662,N_1899,N_682);
nor U5663 (N_5663,N_3304,N_424);
or U5664 (N_5664,N_4393,N_3751);
or U5665 (N_5665,N_2692,N_1628);
or U5666 (N_5666,N_3458,N_1770);
nand U5667 (N_5667,N_1729,N_3838);
and U5668 (N_5668,N_2908,N_3812);
nor U5669 (N_5669,N_1493,N_1500);
or U5670 (N_5670,N_3344,N_1929);
and U5671 (N_5671,N_1747,N_486);
and U5672 (N_5672,N_3865,N_4624);
or U5673 (N_5673,N_4103,N_542);
nor U5674 (N_5674,N_4534,N_2071);
nor U5675 (N_5675,N_4584,N_384);
nor U5676 (N_5676,N_1011,N_2968);
or U5677 (N_5677,N_4212,N_2640);
and U5678 (N_5678,N_3502,N_3105);
nor U5679 (N_5679,N_1926,N_25);
or U5680 (N_5680,N_4830,N_4116);
or U5681 (N_5681,N_2771,N_2160);
or U5682 (N_5682,N_4468,N_4220);
nand U5683 (N_5683,N_4098,N_4523);
or U5684 (N_5684,N_2728,N_3752);
and U5685 (N_5685,N_594,N_2115);
and U5686 (N_5686,N_3099,N_4892);
nand U5687 (N_5687,N_2270,N_2084);
nor U5688 (N_5688,N_3756,N_1704);
nand U5689 (N_5689,N_3150,N_1620);
and U5690 (N_5690,N_1429,N_3357);
nor U5691 (N_5691,N_4052,N_4565);
nand U5692 (N_5692,N_2178,N_3577);
or U5693 (N_5693,N_2302,N_1043);
nand U5694 (N_5694,N_3840,N_3717);
nand U5695 (N_5695,N_631,N_2221);
nand U5696 (N_5696,N_813,N_2727);
nor U5697 (N_5697,N_4238,N_434);
nand U5698 (N_5698,N_1443,N_952);
and U5699 (N_5699,N_4127,N_268);
nand U5700 (N_5700,N_3381,N_395);
nor U5701 (N_5701,N_995,N_1075);
and U5702 (N_5702,N_4168,N_1368);
or U5703 (N_5703,N_3888,N_4236);
nor U5704 (N_5704,N_3586,N_438);
or U5705 (N_5705,N_790,N_4495);
or U5706 (N_5706,N_2146,N_4270);
and U5707 (N_5707,N_802,N_3408);
nor U5708 (N_5708,N_1951,N_246);
or U5709 (N_5709,N_2051,N_3395);
nand U5710 (N_5710,N_3125,N_3988);
and U5711 (N_5711,N_1748,N_2290);
nor U5712 (N_5712,N_2102,N_3835);
nand U5713 (N_5713,N_4851,N_4558);
xor U5714 (N_5714,N_2234,N_2940);
nor U5715 (N_5715,N_1825,N_2239);
and U5716 (N_5716,N_2569,N_1830);
or U5717 (N_5717,N_4248,N_3010);
nand U5718 (N_5718,N_4804,N_4356);
nor U5719 (N_5719,N_354,N_3602);
or U5720 (N_5720,N_2980,N_2561);
and U5721 (N_5721,N_1543,N_3260);
xor U5722 (N_5722,N_2841,N_327);
xor U5723 (N_5723,N_3839,N_3167);
and U5724 (N_5724,N_2279,N_1733);
nor U5725 (N_5725,N_3559,N_4139);
nor U5726 (N_5726,N_1217,N_171);
and U5727 (N_5727,N_3770,N_2474);
nand U5728 (N_5728,N_308,N_303);
nor U5729 (N_5729,N_4333,N_3049);
nand U5730 (N_5730,N_1113,N_2294);
nand U5731 (N_5731,N_2865,N_4071);
and U5732 (N_5732,N_4316,N_2414);
and U5733 (N_5733,N_2216,N_4376);
and U5734 (N_5734,N_1731,N_3185);
nor U5735 (N_5735,N_2161,N_4512);
nor U5736 (N_5736,N_114,N_1891);
or U5737 (N_5737,N_270,N_3109);
and U5738 (N_5738,N_1551,N_4834);
and U5739 (N_5739,N_2297,N_2634);
and U5740 (N_5740,N_2723,N_4932);
or U5741 (N_5741,N_4562,N_1808);
nor U5742 (N_5742,N_2710,N_4200);
or U5743 (N_5743,N_2711,N_4627);
and U5744 (N_5744,N_2512,N_3581);
and U5745 (N_5745,N_1311,N_3077);
or U5746 (N_5746,N_1547,N_282);
nor U5747 (N_5747,N_3446,N_564);
and U5748 (N_5748,N_44,N_3330);
nor U5749 (N_5749,N_585,N_338);
nand U5750 (N_5750,N_937,N_3002);
nor U5751 (N_5751,N_936,N_4583);
nor U5752 (N_5752,N_2196,N_3006);
nand U5753 (N_5753,N_2963,N_907);
nor U5754 (N_5754,N_3128,N_2519);
or U5755 (N_5755,N_1013,N_2464);
nor U5756 (N_5756,N_1994,N_1317);
xor U5757 (N_5757,N_1866,N_3252);
or U5758 (N_5758,N_2029,N_1438);
and U5759 (N_5759,N_1142,N_1299);
and U5760 (N_5760,N_1125,N_1327);
or U5761 (N_5761,N_147,N_3517);
nand U5762 (N_5762,N_1919,N_265);
and U5763 (N_5763,N_1115,N_4811);
or U5764 (N_5764,N_3665,N_4223);
or U5765 (N_5765,N_1374,N_4411);
and U5766 (N_5766,N_2979,N_2552);
nand U5767 (N_5767,N_74,N_2642);
nor U5768 (N_5768,N_100,N_2244);
or U5769 (N_5769,N_3124,N_2651);
nand U5770 (N_5770,N_2186,N_3867);
nor U5771 (N_5771,N_1872,N_1460);
and U5772 (N_5772,N_1712,N_2693);
and U5773 (N_5773,N_3501,N_3019);
and U5774 (N_5774,N_2680,N_4025);
nand U5775 (N_5775,N_422,N_2807);
nand U5776 (N_5776,N_2856,N_3864);
or U5777 (N_5777,N_2308,N_2608);
and U5778 (N_5778,N_2042,N_1700);
nor U5779 (N_5779,N_1860,N_4319);
nand U5780 (N_5780,N_2932,N_710);
or U5781 (N_5781,N_1206,N_750);
nor U5782 (N_5782,N_808,N_151);
nor U5783 (N_5783,N_1902,N_2611);
or U5784 (N_5784,N_4547,N_4933);
nand U5785 (N_5785,N_1313,N_4744);
nor U5786 (N_5786,N_33,N_2781);
nor U5787 (N_5787,N_4081,N_248);
or U5788 (N_5788,N_4814,N_3183);
or U5789 (N_5789,N_4869,N_2902);
or U5790 (N_5790,N_4410,N_2510);
nor U5791 (N_5791,N_4796,N_909);
nand U5792 (N_5792,N_3599,N_2322);
nor U5793 (N_5793,N_931,N_2697);
nor U5794 (N_5794,N_3209,N_3286);
or U5795 (N_5795,N_2400,N_3912);
nand U5796 (N_5796,N_3757,N_4082);
nor U5797 (N_5797,N_1124,N_2391);
or U5798 (N_5798,N_3349,N_3452);
xnor U5799 (N_5799,N_4894,N_614);
and U5800 (N_5800,N_168,N_4163);
and U5801 (N_5801,N_3691,N_3164);
and U5802 (N_5802,N_3522,N_3710);
or U5803 (N_5803,N_1162,N_4390);
nand U5804 (N_5804,N_3053,N_3523);
or U5805 (N_5805,N_2885,N_2686);
nor U5806 (N_5806,N_3285,N_242);
nor U5807 (N_5807,N_3530,N_2055);
nor U5808 (N_5808,N_3354,N_3896);
or U5809 (N_5809,N_1779,N_2514);
and U5810 (N_5810,N_1385,N_3837);
nor U5811 (N_5811,N_3616,N_3555);
or U5812 (N_5812,N_944,N_1697);
and U5813 (N_5813,N_2412,N_2779);
nand U5814 (N_5814,N_4073,N_96);
or U5815 (N_5815,N_3033,N_795);
or U5816 (N_5816,N_1843,N_4222);
nand U5817 (N_5817,N_933,N_4791);
and U5818 (N_5818,N_1102,N_1996);
or U5819 (N_5819,N_1024,N_4365);
or U5820 (N_5820,N_4505,N_855);
or U5821 (N_5821,N_3307,N_69);
nor U5822 (N_5822,N_3807,N_1375);
nand U5823 (N_5823,N_1765,N_357);
nand U5824 (N_5824,N_2304,N_2207);
nand U5825 (N_5825,N_2768,N_3585);
or U5826 (N_5826,N_1286,N_4622);
nor U5827 (N_5827,N_1875,N_4719);
nand U5828 (N_5828,N_3410,N_2929);
nand U5829 (N_5829,N_1647,N_956);
and U5830 (N_5830,N_3977,N_2613);
xor U5831 (N_5831,N_298,N_3029);
xnor U5832 (N_5832,N_4204,N_2813);
and U5833 (N_5833,N_2659,N_499);
nand U5834 (N_5834,N_842,N_4720);
or U5835 (N_5835,N_3632,N_1726);
and U5836 (N_5836,N_1863,N_4428);
nand U5837 (N_5837,N_112,N_1106);
nand U5838 (N_5838,N_2061,N_73);
or U5839 (N_5839,N_4798,N_4769);
xnor U5840 (N_5840,N_3145,N_1751);
nand U5841 (N_5841,N_1132,N_2136);
nand U5842 (N_5842,N_2134,N_4249);
and U5843 (N_5843,N_4192,N_2810);
xnor U5844 (N_5844,N_3042,N_1758);
nor U5845 (N_5845,N_4801,N_1254);
xnor U5846 (N_5846,N_4022,N_1083);
nor U5847 (N_5847,N_175,N_736);
and U5848 (N_5848,N_4619,N_3880);
and U5849 (N_5849,N_4825,N_502);
nor U5850 (N_5850,N_1044,N_2470);
and U5851 (N_5851,N_1079,N_2895);
nor U5852 (N_5852,N_1635,N_1654);
or U5853 (N_5853,N_1434,N_2132);
or U5854 (N_5854,N_1066,N_771);
and U5855 (N_5855,N_4271,N_1359);
nand U5856 (N_5856,N_1721,N_3139);
nand U5857 (N_5857,N_4734,N_3110);
nor U5858 (N_5858,N_375,N_4149);
and U5859 (N_5859,N_1214,N_475);
or U5860 (N_5860,N_4581,N_3216);
or U5861 (N_5861,N_3413,N_1722);
or U5862 (N_5862,N_2579,N_3800);
xor U5863 (N_5863,N_4508,N_1319);
nand U5864 (N_5864,N_2820,N_2822);
nand U5865 (N_5865,N_1403,N_3279);
nand U5866 (N_5866,N_2430,N_3926);
nand U5867 (N_5867,N_1618,N_4485);
xor U5868 (N_5868,N_4856,N_1624);
nor U5869 (N_5869,N_1592,N_4076);
nand U5870 (N_5870,N_3447,N_1371);
or U5871 (N_5871,N_3388,N_2222);
nor U5872 (N_5872,N_1264,N_3626);
nor U5873 (N_5873,N_3238,N_3315);
nand U5874 (N_5874,N_132,N_4504);
or U5875 (N_5875,N_3508,N_226);
nand U5876 (N_5876,N_3890,N_58);
xnor U5877 (N_5877,N_4666,N_3037);
nand U5878 (N_5878,N_1845,N_2453);
and U5879 (N_5879,N_3634,N_1471);
nand U5880 (N_5880,N_629,N_2958);
nand U5881 (N_5881,N_2545,N_3313);
or U5882 (N_5882,N_272,N_3841);
and U5883 (N_5883,N_4044,N_4836);
nor U5884 (N_5884,N_48,N_3182);
nor U5885 (N_5885,N_2484,N_991);
and U5886 (N_5886,N_3336,N_2165);
nand U5887 (N_5887,N_4545,N_1263);
or U5888 (N_5888,N_3287,N_4187);
nand U5889 (N_5889,N_3056,N_2032);
nand U5890 (N_5890,N_149,N_3486);
nand U5891 (N_5891,N_51,N_1710);
and U5892 (N_5892,N_2468,N_4252);
nand U5893 (N_5893,N_2426,N_3556);
or U5894 (N_5894,N_3653,N_1109);
or U5895 (N_5895,N_3308,N_2487);
xor U5896 (N_5896,N_3660,N_4426);
nor U5897 (N_5897,N_1246,N_4284);
and U5898 (N_5898,N_1627,N_4574);
nor U5899 (N_5899,N_2251,N_3892);
or U5900 (N_5900,N_700,N_3906);
or U5901 (N_5901,N_1218,N_692);
nor U5902 (N_5902,N_2284,N_863);
and U5903 (N_5903,N_3580,N_2193);
or U5904 (N_5904,N_3387,N_3562);
and U5905 (N_5905,N_4364,N_4160);
and U5906 (N_5906,N_2100,N_2972);
nor U5907 (N_5907,N_76,N_4654);
and U5908 (N_5908,N_4137,N_4214);
nor U5909 (N_5909,N_1614,N_4794);
nand U5910 (N_5910,N_215,N_2162);
nand U5911 (N_5911,N_1797,N_3225);
and U5912 (N_5912,N_3152,N_4423);
xnor U5913 (N_5913,N_900,N_1949);
nand U5914 (N_5914,N_3597,N_469);
or U5915 (N_5915,N_636,N_1840);
nand U5916 (N_5916,N_2675,N_1172);
nor U5917 (N_5917,N_13,N_3755);
nor U5918 (N_5918,N_1230,N_4446);
nand U5919 (N_5919,N_4150,N_4012);
nand U5920 (N_5920,N_4924,N_3223);
nand U5921 (N_5921,N_2606,N_549);
and U5922 (N_5922,N_3104,N_3930);
nand U5923 (N_5923,N_521,N_2163);
nor U5924 (N_5924,N_394,N_455);
or U5925 (N_5925,N_3061,N_250);
nand U5926 (N_5926,N_1783,N_231);
nand U5927 (N_5927,N_3571,N_3933);
or U5928 (N_5928,N_1633,N_4406);
or U5929 (N_5929,N_4416,N_1999);
or U5930 (N_5930,N_4876,N_3352);
nand U5931 (N_5931,N_3229,N_2498);
nor U5932 (N_5932,N_859,N_843);
or U5933 (N_5933,N_3227,N_4817);
or U5934 (N_5934,N_4201,N_192);
or U5935 (N_5935,N_1655,N_4066);
nor U5936 (N_5936,N_3711,N_1388);
or U5937 (N_5937,N_544,N_558);
nor U5938 (N_5938,N_4679,N_1473);
nor U5939 (N_5939,N_1353,N_4243);
and U5940 (N_5940,N_3557,N_945);
and U5941 (N_5941,N_45,N_524);
and U5942 (N_5942,N_4808,N_3776);
nand U5943 (N_5943,N_2679,N_3212);
nand U5944 (N_5944,N_4464,N_3853);
nand U5945 (N_5945,N_797,N_2818);
or U5946 (N_5946,N_3695,N_187);
nand U5947 (N_5947,N_4075,N_4273);
nor U5948 (N_5948,N_3123,N_2433);
and U5949 (N_5949,N_4310,N_794);
and U5950 (N_5950,N_289,N_1776);
or U5951 (N_5951,N_718,N_1530);
or U5952 (N_5952,N_4293,N_1407);
or U5953 (N_5953,N_445,N_630);
and U5954 (N_5954,N_2362,N_3323);
or U5955 (N_5955,N_3623,N_2802);
and U5956 (N_5956,N_2862,N_4265);
or U5957 (N_5957,N_4715,N_3520);
or U5958 (N_5958,N_2340,N_253);
or U5959 (N_5959,N_3761,N_3589);
nor U5960 (N_5960,N_2012,N_2522);
and U5961 (N_5961,N_4374,N_4898);
nand U5962 (N_5962,N_1963,N_319);
nand U5963 (N_5963,N_2527,N_3782);
nor U5964 (N_5964,N_4250,N_4842);
and U5965 (N_5965,N_3944,N_2546);
nand U5966 (N_5966,N_1284,N_2045);
or U5967 (N_5967,N_2883,N_179);
and U5968 (N_5968,N_3131,N_1041);
nor U5969 (N_5969,N_1794,N_1);
or U5970 (N_5970,N_1537,N_4259);
and U5971 (N_5971,N_3316,N_70);
and U5972 (N_5972,N_3297,N_307);
nand U5973 (N_5973,N_2868,N_1268);
nor U5974 (N_5974,N_397,N_4004);
nand U5975 (N_5975,N_238,N_205);
nand U5976 (N_5976,N_1989,N_4931);
xnor U5977 (N_5977,N_2217,N_1738);
nor U5978 (N_5978,N_1110,N_2283);
and U5979 (N_5979,N_3367,N_2765);
nand U5980 (N_5980,N_988,N_957);
nor U5981 (N_5981,N_4414,N_561);
nor U5982 (N_5982,N_3779,N_3878);
and U5983 (N_5983,N_3457,N_4314);
nand U5984 (N_5984,N_1757,N_4405);
and U5985 (N_5985,N_747,N_4330);
nor U5986 (N_5986,N_1251,N_753);
and U5987 (N_5987,N_3917,N_2048);
nor U5988 (N_5988,N_1243,N_4470);
or U5989 (N_5989,N_2274,N_1694);
nand U5990 (N_5990,N_4181,N_3162);
nor U5991 (N_5991,N_803,N_2452);
nor U5992 (N_5992,N_853,N_1369);
nand U5993 (N_5993,N_1262,N_378);
nand U5994 (N_5994,N_3483,N_4690);
nand U5995 (N_5995,N_2973,N_1821);
nor U5996 (N_5996,N_1660,N_3692);
and U5997 (N_5997,N_398,N_393);
nor U5998 (N_5998,N_977,N_331);
and U5999 (N_5999,N_1065,N_2673);
nor U6000 (N_6000,N_1597,N_2037);
nor U6001 (N_6001,N_3498,N_124);
xor U6002 (N_6002,N_1550,N_3648);
or U6003 (N_6003,N_329,N_188);
xor U6004 (N_6004,N_3927,N_4145);
or U6005 (N_6005,N_3702,N_2511);
nand U6006 (N_6006,N_2777,N_4673);
and U6007 (N_6007,N_4987,N_4692);
and U6008 (N_6008,N_2157,N_1086);
and U6009 (N_6009,N_648,N_1933);
and U6010 (N_6010,N_2914,N_418);
nor U6011 (N_6011,N_821,N_214);
and U6012 (N_6012,N_1657,N_2716);
nor U6013 (N_6013,N_4300,N_1713);
or U6014 (N_6014,N_4593,N_1018);
and U6015 (N_6015,N_4383,N_2704);
or U6016 (N_6016,N_3024,N_1167);
or U6017 (N_6017,N_3385,N_1741);
and U6018 (N_6018,N_204,N_4867);
nand U6019 (N_6019,N_1878,N_360);
nor U6020 (N_6020,N_2355,N_1545);
and U6021 (N_6021,N_281,N_2901);
nor U6022 (N_6022,N_3664,N_3180);
and U6023 (N_6023,N_913,N_887);
and U6024 (N_6024,N_4709,N_4950);
nor U6025 (N_6025,N_3728,N_3163);
and U6026 (N_6026,N_99,N_4522);
or U6027 (N_6027,N_2804,N_4595);
and U6028 (N_6028,N_1855,N_2563);
or U6029 (N_6029,N_3819,N_2010);
and U6030 (N_6030,N_2900,N_4141);
nand U6031 (N_6031,N_716,N_1806);
or U6032 (N_6032,N_4553,N_783);
and U6033 (N_6033,N_2502,N_254);
and U6034 (N_6034,N_2717,N_1170);
nand U6035 (N_6035,N_1105,N_2653);
and U6036 (N_6036,N_799,N_2694);
nand U6037 (N_6037,N_3936,N_4448);
nor U6038 (N_6038,N_4663,N_3619);
nand U6039 (N_6039,N_3738,N_2567);
or U6040 (N_6040,N_3939,N_1924);
nor U6041 (N_6041,N_2859,N_1501);
or U6042 (N_6042,N_3461,N_184);
and U6043 (N_6043,N_134,N_340);
and U6044 (N_6044,N_3998,N_4014);
nand U6045 (N_6045,N_2938,N_2457);
nor U6046 (N_6046,N_1649,N_449);
nor U6047 (N_6047,N_3644,N_1145);
or U6048 (N_6048,N_1097,N_1427);
nand U6049 (N_6049,N_1785,N_516);
and U6050 (N_6050,N_2508,N_4920);
nand U6051 (N_6051,N_3666,N_3902);
nor U6052 (N_6052,N_4781,N_4764);
nand U6053 (N_6053,N_2602,N_2341);
or U6054 (N_6054,N_3842,N_511);
nand U6055 (N_6055,N_1824,N_3472);
nand U6056 (N_6056,N_3453,N_2650);
nand U6057 (N_6057,N_4823,N_727);
nand U6058 (N_6058,N_2377,N_146);
nand U6059 (N_6059,N_1573,N_1242);
nor U6060 (N_6060,N_38,N_3916);
and U6061 (N_6061,N_4062,N_3549);
nor U6062 (N_6062,N_277,N_3237);
and U6063 (N_6063,N_777,N_1796);
nand U6064 (N_6064,N_3610,N_2661);
nor U6065 (N_6065,N_626,N_4277);
nor U6066 (N_6066,N_545,N_1021);
nor U6067 (N_6067,N_2764,N_3637);
nand U6068 (N_6068,N_1482,N_334);
and U6069 (N_6069,N_1071,N_2261);
or U6070 (N_6070,N_3379,N_4696);
and U6071 (N_6071,N_4462,N_1288);
nand U6072 (N_6072,N_2603,N_3907);
nor U6073 (N_6073,N_2703,N_80);
and U6074 (N_6074,N_3720,N_4916);
or U6075 (N_6075,N_4281,N_140);
or U6076 (N_6076,N_4118,N_1665);
or U6077 (N_6077,N_3135,N_4000);
and U6078 (N_6078,N_4418,N_2460);
nor U6079 (N_6079,N_3346,N_3005);
or U6080 (N_6080,N_2130,N_3877);
or U6081 (N_6081,N_939,N_3201);
nor U6082 (N_6082,N_3369,N_4790);
xnor U6083 (N_6083,N_2177,N_4662);
nand U6084 (N_6084,N_4986,N_1377);
or U6085 (N_6085,N_3911,N_4889);
or U6086 (N_6086,N_1874,N_4377);
or U6087 (N_6087,N_4289,N_1639);
or U6088 (N_6088,N_4563,N_4079);
or U6089 (N_6089,N_691,N_1025);
nor U6090 (N_6090,N_1826,N_4438);
and U6091 (N_6091,N_885,N_2011);
or U6092 (N_6092,N_457,N_4085);
nand U6093 (N_6093,N_3444,N_2066);
nand U6094 (N_6094,N_1841,N_4741);
nand U6095 (N_6095,N_4324,N_1160);
or U6096 (N_6096,N_4215,N_1278);
or U6097 (N_6097,N_1643,N_4440);
or U6098 (N_6098,N_1350,N_1280);
nor U6099 (N_6099,N_4355,N_3529);
and U6100 (N_6100,N_2702,N_3871);
and U6101 (N_6101,N_4591,N_3515);
or U6102 (N_6102,N_2987,N_2445);
and U6103 (N_6103,N_55,N_706);
xor U6104 (N_6104,N_2370,N_778);
or U6105 (N_6105,N_3331,N_505);
nand U6106 (N_6106,N_3137,N_405);
or U6107 (N_6107,N_3740,N_4784);
nand U6108 (N_6108,N_2117,N_3894);
nand U6109 (N_6109,N_3884,N_2276);
or U6110 (N_6110,N_601,N_3716);
or U6111 (N_6111,N_210,N_2383);
or U6112 (N_6112,N_1945,N_4193);
nand U6113 (N_6113,N_413,N_2455);
and U6114 (N_6114,N_2685,N_2751);
nand U6115 (N_6115,N_4454,N_235);
nand U6116 (N_6116,N_3284,N_317);
and U6117 (N_6117,N_3975,N_3924);
or U6118 (N_6118,N_2663,N_1616);
nand U6119 (N_6119,N_4490,N_2016);
xnor U6120 (N_6120,N_5,N_3465);
and U6121 (N_6121,N_1883,N_1486);
and U6122 (N_6122,N_3166,N_2965);
nand U6123 (N_6123,N_2480,N_4860);
and U6124 (N_6124,N_1329,N_3804);
or U6125 (N_6125,N_1517,N_4246);
or U6126 (N_6126,N_997,N_543);
nand U6127 (N_6127,N_3745,N_3604);
nor U6128 (N_6128,N_1857,N_2964);
nor U6129 (N_6129,N_994,N_590);
or U6130 (N_6130,N_2286,N_1004);
or U6131 (N_6131,N_2293,N_1301);
xnor U6132 (N_6132,N_2747,N_2906);
or U6133 (N_6133,N_2515,N_3491);
nand U6134 (N_6134,N_4235,N_4313);
nand U6135 (N_6135,N_4693,N_2909);
and U6136 (N_6136,N_1266,N_4442);
nor U6137 (N_6137,N_1542,N_3686);
nor U6138 (N_6138,N_3149,N_2824);
and U6139 (N_6139,N_2273,N_2550);
nor U6140 (N_6140,N_1985,N_3434);
and U6141 (N_6141,N_17,N_961);
nand U6142 (N_6142,N_2255,N_649);
nand U6143 (N_6143,N_1799,N_1966);
nor U6144 (N_6144,N_2395,N_4519);
or U6145 (N_6145,N_1247,N_1400);
and U6146 (N_6146,N_1762,N_999);
and U6147 (N_6147,N_1528,N_1773);
nand U6148 (N_6148,N_3143,N_3130);
or U6149 (N_6149,N_4477,N_54);
nor U6150 (N_6150,N_1445,N_1921);
nor U6151 (N_6151,N_450,N_3688);
nand U6152 (N_6152,N_1549,N_4061);
nand U6153 (N_6153,N_1099,N_2803);
or U6154 (N_6154,N_1858,N_94);
nor U6155 (N_6155,N_1957,N_4198);
nor U6156 (N_6156,N_1153,N_2772);
and U6157 (N_6157,N_256,N_3000);
and U6158 (N_6158,N_2110,N_3704);
or U6159 (N_6159,N_4748,N_4516);
nor U6160 (N_6160,N_4901,N_3620);
nor U6161 (N_6161,N_1746,N_3887);
nand U6162 (N_6162,N_1296,N_3516);
nand U6163 (N_6163,N_269,N_2287);
and U6164 (N_6164,N_4288,N_2796);
nor U6165 (N_6165,N_1207,N_2639);
or U6166 (N_6166,N_1462,N_347);
nor U6167 (N_6167,N_707,N_1737);
and U6168 (N_6168,N_818,N_3311);
nand U6169 (N_6169,N_3314,N_431);
nor U6170 (N_6170,N_2172,N_4645);
nor U6171 (N_6171,N_3791,N_3997);
and U6172 (N_6172,N_97,N_4517);
nand U6173 (N_6173,N_3854,N_1906);
nor U6174 (N_6174,N_4155,N_1771);
nor U6175 (N_6175,N_2748,N_1002);
and U6176 (N_6176,N_1792,N_3247);
or U6177 (N_6177,N_91,N_1672);
nand U6178 (N_6178,N_2000,N_678);
nand U6179 (N_6179,N_935,N_2630);
nand U6180 (N_6180,N_2898,N_1717);
nand U6181 (N_6181,N_4055,N_1381);
and U6182 (N_6182,N_3353,N_1104);
and U6183 (N_6183,N_223,N_2404);
or U6184 (N_6184,N_426,N_3671);
xor U6185 (N_6185,N_4942,N_3696);
nand U6186 (N_6186,N_2734,N_4611);
nand U6187 (N_6187,N_3324,N_1087);
or U6188 (N_6188,N_1611,N_2328);
nor U6189 (N_6189,N_1563,N_2209);
and U6190 (N_6190,N_1774,N_3221);
nor U6191 (N_6191,N_2798,N_1815);
nor U6192 (N_6192,N_1991,N_3068);
and U6193 (N_6193,N_4381,N_765);
nor U6194 (N_6194,N_4958,N_3767);
nand U6195 (N_6195,N_2190,N_344);
nor U6196 (N_6196,N_4033,N_1580);
nor U6197 (N_6197,N_4576,N_3905);
and U6198 (N_6198,N_3360,N_4541);
nor U6199 (N_6199,N_3302,N_1535);
or U6200 (N_6200,N_400,N_4269);
and U6201 (N_6201,N_3432,N_3106);
and U6202 (N_6202,N_3918,N_2033);
nand U6203 (N_6203,N_4027,N_1324);
nor U6204 (N_6204,N_1476,N_1950);
nand U6205 (N_6205,N_3748,N_3563);
and U6206 (N_6206,N_3439,N_2933);
xnor U6207 (N_6207,N_1553,N_1507);
and U6208 (N_6208,N_1488,N_4578);
nor U6209 (N_6209,N_4757,N_622);
nand U6210 (N_6210,N_732,N_4815);
and U6211 (N_6211,N_3984,N_358);
xnor U6212 (N_6212,N_4256,N_3785);
nor U6213 (N_6213,N_294,N_2381);
and U6214 (N_6214,N_1461,N_4375);
or U6215 (N_6215,N_463,N_4358);
nor U6216 (N_6216,N_1143,N_2913);
nor U6217 (N_6217,N_2495,N_296);
and U6218 (N_6218,N_4407,N_597);
nor U6219 (N_6219,N_3850,N_2506);
nand U6220 (N_6220,N_1615,N_3415);
nor U6221 (N_6221,N_903,N_1715);
nor U6222 (N_6222,N_2194,N_2069);
nand U6223 (N_6223,N_4147,N_3575);
and U6224 (N_6224,N_2402,N_3834);
nor U6225 (N_6225,N_625,N_3674);
and U6226 (N_6226,N_4159,N_2378);
or U6227 (N_6227,N_4036,N_1920);
nand U6228 (N_6228,N_19,N_4074);
nor U6229 (N_6229,N_60,N_1761);
nor U6230 (N_6230,N_2855,N_278);
nand U6231 (N_6231,N_1568,N_4164);
nand U6232 (N_6232,N_3054,N_593);
nor U6233 (N_6233,N_1787,N_1905);
nor U6234 (N_6234,N_1118,N_4536);
or U6235 (N_6235,N_240,N_705);
nand U6236 (N_6236,N_655,N_576);
nor U6237 (N_6237,N_1742,N_4728);
nand U6238 (N_6238,N_1766,N_4638);
and U6239 (N_6239,N_4859,N_1121);
and U6240 (N_6240,N_3749,N_2745);
nor U6241 (N_6241,N_2416,N_376);
and U6242 (N_6242,N_3254,N_2348);
nor U6243 (N_6243,N_3621,N_4960);
and U6244 (N_6244,N_195,N_4820);
nand U6245 (N_6245,N_2382,N_1646);
and U6246 (N_6246,N_4776,N_403);
or U6247 (N_6247,N_274,N_3412);
nor U6248 (N_6248,N_1784,N_3950);
nor U6249 (N_6249,N_3086,N_1199);
or U6250 (N_6250,N_3404,N_915);
and U6251 (N_6251,N_2158,N_2912);
nand U6252 (N_6252,N_4717,N_3427);
nand U6253 (N_6253,N_894,N_2590);
nor U6254 (N_6254,N_2739,N_1189);
xnor U6255 (N_6255,N_4177,N_1604);
xnor U6256 (N_6256,N_3624,N_1077);
or U6257 (N_6257,N_1578,N_3609);
or U6258 (N_6258,N_1603,N_2709);
and U6259 (N_6259,N_2689,N_4107);
or U6260 (N_6260,N_1688,N_1049);
and U6261 (N_6261,N_4822,N_4976);
or U6262 (N_6262,N_2821,N_2795);
nand U6263 (N_6263,N_314,N_4385);
nor U6264 (N_6264,N_981,N_4459);
nor U6265 (N_6265,N_4003,N_4777);
nor U6266 (N_6266,N_4771,N_435);
nor U6267 (N_6267,N_3421,N_3215);
and U6268 (N_6268,N_2801,N_2767);
nor U6269 (N_6269,N_3872,N_428);
nand U6270 (N_6270,N_2632,N_1028);
nor U6271 (N_6271,N_828,N_4040);
nand U6272 (N_6272,N_739,N_150);
nor U6273 (N_6273,N_1195,N_4015);
nand U6274 (N_6274,N_3860,N_2334);
and U6275 (N_6275,N_3089,N_3994);
or U6276 (N_6276,N_209,N_3192);
and U6277 (N_6277,N_2141,N_676);
or U6278 (N_6278,N_387,N_3558);
or U6279 (N_6279,N_4745,N_2492);
nor U6280 (N_6280,N_3050,N_1581);
nor U6281 (N_6281,N_2389,N_3170);
nand U6282 (N_6282,N_3968,N_1444);
nand U6283 (N_6283,N_4850,N_633);
or U6284 (N_6284,N_3972,N_4130);
nor U6285 (N_6285,N_617,N_1093);
nor U6286 (N_6286,N_1090,N_4539);
and U6287 (N_6287,N_850,N_1082);
nor U6288 (N_6288,N_1927,N_3281);
nor U6289 (N_6289,N_1910,N_4436);
nor U6290 (N_6290,N_1959,N_728);
xnor U6291 (N_6291,N_1781,N_2993);
nand U6292 (N_6292,N_2746,N_4707);
or U6293 (N_6293,N_3440,N_2316);
and U6294 (N_6294,N_2082,N_1625);
or U6295 (N_6295,N_1798,N_1469);
nand U6296 (N_6296,N_2373,N_2584);
nor U6297 (N_6297,N_4425,N_4543);
or U6298 (N_6298,N_1425,N_662);
xor U6299 (N_6299,N_2439,N_788);
and U6300 (N_6300,N_4343,N_288);
and U6301 (N_6301,N_904,N_143);
nand U6302 (N_6302,N_1366,N_925);
or U6303 (N_6303,N_3722,N_1800);
nand U6304 (N_6304,N_185,N_2953);
or U6305 (N_6305,N_816,N_4323);
or U6306 (N_6306,N_4500,N_113);
nand U6307 (N_6307,N_975,N_2714);
xnor U6308 (N_6308,N_3500,N_2073);
and U6309 (N_6309,N_4598,N_2637);
and U6310 (N_6310,N_491,N_1873);
and U6311 (N_6311,N_3026,N_3983);
nand U6312 (N_6312,N_218,N_714);
nor U6313 (N_6313,N_1408,N_4799);
and U6314 (N_6314,N_4597,N_3112);
nand U6315 (N_6315,N_2459,N_1962);
and U6316 (N_6316,N_3200,N_3826);
nor U6317 (N_6317,N_632,N_4194);
nand U6318 (N_6318,N_3750,N_3306);
nor U6319 (N_6319,N_4945,N_1297);
nand U6320 (N_6320,N_1394,N_3155);
nor U6321 (N_6321,N_3230,N_2440);
nor U6322 (N_6322,N_4059,N_4582);
and U6323 (N_6323,N_36,N_4482);
nand U6324 (N_6324,N_42,N_2482);
nor U6325 (N_6325,N_4750,N_3069);
nand U6326 (N_6326,N_72,N_3734);
nand U6327 (N_6327,N_1158,N_4412);
nand U6328 (N_6328,N_738,N_4032);
nor U6329 (N_6329,N_2020,N_4387);
nand U6330 (N_6330,N_643,N_3565);
nor U6331 (N_6331,N_459,N_4507);
and U6332 (N_6332,N_4603,N_619);
nor U6333 (N_6333,N_1939,N_1489);
and U6334 (N_6334,N_2148,N_410);
nand U6335 (N_6335,N_4721,N_2305);
or U6336 (N_6336,N_3815,N_2374);
nand U6337 (N_6337,N_460,N_580);
xor U6338 (N_6338,N_416,N_1376);
or U6339 (N_6339,N_4380,N_4363);
nand U6340 (N_6340,N_500,N_1450);
and U6341 (N_6341,N_4430,N_2537);
or U6342 (N_6342,N_1211,N_846);
nor U6343 (N_6343,N_3783,N_1577);
or U6344 (N_6344,N_3101,N_1479);
or U6345 (N_6345,N_2269,N_755);
xnor U6346 (N_6346,N_2496,N_4789);
and U6347 (N_6347,N_2899,N_3806);
nor U6348 (N_6348,N_3366,N_2528);
nor U6349 (N_6349,N_3122,N_4686);
or U6350 (N_6350,N_1334,N_1256);
nand U6351 (N_6351,N_1870,N_1257);
and U6352 (N_6352,N_1399,N_441);
or U6353 (N_6353,N_1001,N_3766);
nor U6354 (N_6354,N_1645,N_123);
nor U6355 (N_6355,N_1805,N_826);
and U6356 (N_6356,N_2105,N_772);
or U6357 (N_6357,N_4023,N_3503);
nand U6358 (N_6358,N_4417,N_573);
and U6359 (N_6359,N_2437,N_1786);
and U6360 (N_6360,N_844,N_224);
or U6361 (N_6361,N_4369,N_199);
and U6362 (N_6362,N_653,N_4979);
nand U6363 (N_6363,N_1974,N_860);
or U6364 (N_6364,N_1892,N_1204);
nand U6365 (N_6365,N_1267,N_4983);
nand U6366 (N_6366,N_2878,N_4434);
or U6367 (N_6367,N_1546,N_2551);
and U6368 (N_6368,N_2329,N_1565);
nand U6369 (N_6369,N_2150,N_1235);
and U6370 (N_6370,N_3960,N_1418);
nor U6371 (N_6371,N_144,N_2731);
nand U6372 (N_6372,N_1314,N_3855);
xnor U6373 (N_6373,N_3949,N_4893);
nand U6374 (N_6374,N_1341,N_1755);
xor U6375 (N_6375,N_4487,N_3584);
nor U6376 (N_6376,N_1209,N_1952);
or U6377 (N_6377,N_864,N_2683);
or U6378 (N_6378,N_525,N_697);
nand U6379 (N_6379,N_3066,N_3603);
nor U6380 (N_6380,N_4047,N_1678);
nand U6381 (N_6381,N_82,N_552);
or U6382 (N_6382,N_1405,N_2471);
nor U6383 (N_6383,N_1658,N_3193);
nand U6384 (N_6384,N_1854,N_2369);
nand U6385 (N_6385,N_4560,N_3393);
nand U6386 (N_6386,N_2360,N_108);
and U6387 (N_6387,N_3157,N_1670);
nor U6388 (N_6388,N_539,N_3593);
or U6389 (N_6389,N_3175,N_2257);
nor U6390 (N_6390,N_3126,N_81);
nand U6391 (N_6391,N_2392,N_2156);
xnor U6392 (N_6392,N_2093,N_4382);
nand U6393 (N_6393,N_4290,N_4119);
or U6394 (N_6394,N_3655,N_3242);
and U6395 (N_6395,N_4755,N_1801);
nor U6396 (N_6396,N_2152,N_3063);
or U6397 (N_6397,N_1691,N_4956);
nand U6398 (N_6398,N_3251,N_1727);
or U6399 (N_6399,N_2623,N_3802);
and U6400 (N_6400,N_2828,N_1383);
and U6401 (N_6401,N_973,N_2049);
nand U6402 (N_6402,N_2447,N_4947);
nor U6403 (N_6403,N_4217,N_4039);
xnor U6404 (N_6404,N_4465,N_4579);
or U6405 (N_6405,N_1666,N_3705);
nand U6406 (N_6406,N_4601,N_3409);
and U6407 (N_6407,N_4710,N_1520);
and U6408 (N_6408,N_3278,N_3093);
nand U6409 (N_6409,N_4807,N_1386);
and U6410 (N_6410,N_1472,N_4287);
nor U6411 (N_6411,N_64,N_1767);
nand U6412 (N_6412,N_782,N_4378);
and U6413 (N_6413,N_1126,N_180);
xnor U6414 (N_6414,N_4197,N_4660);
xor U6415 (N_6415,N_3274,N_4173);
nand U6416 (N_6416,N_3025,N_4026);
nand U6417 (N_6417,N_4165,N_526);
nor U6418 (N_6418,N_3630,N_194);
and U6419 (N_6419,N_4723,N_3094);
nor U6420 (N_6420,N_2670,N_4926);
or U6421 (N_6421,N_3852,N_4648);
and U6422 (N_6422,N_4546,N_421);
or U6423 (N_6423,N_4937,N_934);
or U6424 (N_6424,N_3895,N_1871);
nor U6425 (N_6425,N_65,N_1575);
or U6426 (N_6426,N_2740,N_2627);
nand U6427 (N_6427,N_4203,N_2140);
nor U6428 (N_6428,N_4653,N_2083);
nand U6429 (N_6429,N_1954,N_1483);
and U6430 (N_6430,N_4571,N_160);
and U6431 (N_6431,N_4540,N_3020);
and U6432 (N_6432,N_2281,N_4483);
or U6433 (N_6433,N_896,N_2857);
or U6434 (N_6434,N_122,N_3735);
xnor U6435 (N_6435,N_1027,N_1344);
or U6436 (N_6436,N_1098,N_4795);
nand U6437 (N_6437,N_4335,N_3541);
xnor U6438 (N_6438,N_4989,N_4928);
or U6439 (N_6439,N_989,N_1987);
or U6440 (N_6440,N_546,N_2560);
and U6441 (N_6441,N_4724,N_3312);
xnor U6442 (N_6442,N_3140,N_3073);
xor U6443 (N_6443,N_4990,N_309);
or U6444 (N_6444,N_1913,N_4402);
and U6445 (N_6445,N_2477,N_3240);
or U6446 (N_6446,N_3467,N_1610);
and U6447 (N_6447,N_2699,N_4691);
nor U6448 (N_6448,N_3305,N_4384);
nand U6449 (N_6449,N_3514,N_464);
nor U6450 (N_6450,N_2429,N_2805);
and U6451 (N_6451,N_2065,N_3437);
and U6452 (N_6452,N_3456,N_2682);
nand U6453 (N_6453,N_708,N_2690);
nor U6454 (N_6454,N_2619,N_292);
or U6455 (N_6455,N_857,N_1270);
nor U6456 (N_6456,N_2598,N_2915);
nor U6457 (N_6457,N_4731,N_4752);
nor U6458 (N_6458,N_4975,N_4758);
and U6459 (N_6459,N_569,N_1526);
and U6460 (N_6460,N_2138,N_1763);
or U6461 (N_6461,N_3407,N_551);
xor U6462 (N_6462,N_77,N_4253);
xor U6463 (N_6463,N_1022,N_3820);
and U6464 (N_6464,N_3245,N_4643);
and U6465 (N_6465,N_3208,N_4344);
nor U6466 (N_6466,N_228,N_2120);
or U6467 (N_6467,N_4954,N_1534);
and U6468 (N_6468,N_4460,N_1760);
and U6469 (N_6469,N_480,N_1422);
and U6470 (N_6470,N_2615,N_3999);
and U6471 (N_6471,N_313,N_4874);
or U6472 (N_6472,N_3293,N_1882);
or U6473 (N_6473,N_2997,N_437);
or U6474 (N_6474,N_2544,N_4366);
nor U6475 (N_6475,N_2501,N_695);
nor U6476 (N_6476,N_3760,N_4307);
and U6477 (N_6477,N_2681,N_1510);
or U6478 (N_6478,N_1128,N_4704);
xnor U6479 (N_6479,N_79,N_742);
nor U6480 (N_6480,N_87,N_532);
xnor U6481 (N_6481,N_4274,N_1780);
or U6482 (N_6482,N_2625,N_809);
or U6483 (N_6483,N_1525,N_4535);
nand U6484 (N_6484,N_3499,N_2096);
nor U6485 (N_6485,N_2880,N_1702);
nand U6486 (N_6486,N_4969,N_1590);
or U6487 (N_6487,N_2989,N_2008);
nor U6488 (N_6488,N_3014,N_2806);
or U6489 (N_6489,N_2784,N_3231);
nor U6490 (N_6490,N_895,N_3370);
and U6491 (N_6491,N_4616,N_4400);
nand U6492 (N_6492,N_623,N_479);
nor U6493 (N_6493,N_2153,N_2808);
nor U6494 (N_6494,N_3813,N_851);
nor U6495 (N_6495,N_664,N_2056);
and U6496 (N_6496,N_3996,N_1973);
or U6497 (N_6497,N_4420,N_3909);
nor U6498 (N_6498,N_4520,N_3340);
and U6499 (N_6499,N_4229,N_1046);
xnor U6500 (N_6500,N_2556,N_481);
nand U6501 (N_6501,N_3727,N_3687);
nand U6502 (N_6502,N_4115,N_135);
nand U6503 (N_6503,N_16,N_820);
nor U6504 (N_6504,N_2559,N_14);
nor U6505 (N_6505,N_2665,N_2432);
nand U6506 (N_6506,N_1023,N_984);
or U6507 (N_6507,N_4592,N_249);
nand U6508 (N_6508,N_4439,N_3236);
nor U6509 (N_6509,N_4453,N_3332);
and U6510 (N_6510,N_1600,N_839);
nand U6511 (N_6511,N_3601,N_4226);
and U6512 (N_6512,N_534,N_1260);
nand U6513 (N_6513,N_4013,N_88);
or U6514 (N_6514,N_845,N_4502);
or U6515 (N_6515,N_1149,N_3891);
nand U6516 (N_6516,N_3831,N_219);
nand U6517 (N_6517,N_4258,N_4694);
and U6518 (N_6518,N_2053,N_2313);
nand U6519 (N_6519,N_2762,N_1466);
and U6520 (N_6520,N_1241,N_1944);
or U6521 (N_6521,N_1310,N_2759);
nor U6522 (N_6522,N_4644,N_1932);
nor U6523 (N_6523,N_3333,N_3576);
nor U6524 (N_6524,N_849,N_1285);
or U6525 (N_6525,N_3811,N_2142);
and U6526 (N_6526,N_2220,N_4148);
nand U6527 (N_6527,N_2616,N_3830);
nor U6528 (N_6528,N_4544,N_1946);
nand U6529 (N_6529,N_1941,N_4341);
nand U6530 (N_6530,N_4852,N_1274);
or U6531 (N_6531,N_2646,N_377);
or U6532 (N_6532,N_2575,N_2684);
xor U6533 (N_6533,N_3418,N_221);
or U6534 (N_6534,N_1428,N_3943);
and U6535 (N_6535,N_2418,N_2454);
or U6536 (N_6536,N_2981,N_1699);
or U6537 (N_6537,N_562,N_4182);
or U6538 (N_6538,N_4944,N_2833);
nor U6539 (N_6539,N_793,N_4224);
nand U6540 (N_6540,N_4233,N_3261);
nor U6541 (N_6541,N_638,N_2999);
or U6542 (N_6542,N_3250,N_3080);
nand U6543 (N_6543,N_2259,N_992);
nand U6544 (N_6544,N_1522,N_1623);
nand U6545 (N_6545,N_666,N_4669);
nand U6546 (N_6546,N_1515,N_702);
nor U6547 (N_6547,N_746,N_4935);
or U6548 (N_6548,N_948,N_4824);
and U6549 (N_6549,N_3931,N_2267);
nor U6550 (N_6550,N_2300,N_148);
and U6551 (N_6551,N_3422,N_955);
or U6552 (N_6552,N_923,N_3725);
and U6553 (N_6553,N_2151,N_4849);
or U6554 (N_6554,N_1918,N_3083);
and U6555 (N_6555,N_3561,N_4862);
or U6556 (N_6556,N_332,N_4923);
nor U6557 (N_6557,N_2428,N_2830);
nor U6558 (N_6558,N_4572,N_4072);
nor U6559 (N_6559,N_4452,N_388);
nor U6560 (N_6560,N_4351,N_1355);
nand U6561 (N_6561,N_4396,N_2708);
xnor U6562 (N_6562,N_2298,N_4677);
or U6563 (N_6563,N_2572,N_889);
and U6564 (N_6564,N_2756,N_3248);
and U6565 (N_6565,N_2183,N_304);
nor U6566 (N_6566,N_3798,N_3470);
and U6567 (N_6567,N_4829,N_789);
nand U6568 (N_6568,N_3009,N_4005);
nand U6569 (N_6569,N_3546,N_1606);
or U6570 (N_6570,N_1909,N_3172);
and U6571 (N_6571,N_2278,N_3764);
nand U6572 (N_6572,N_2215,N_2479);
or U6573 (N_6573,N_554,N_164);
or U6574 (N_6574,N_2601,N_2864);
or U6575 (N_6575,N_3384,N_2423);
or U6576 (N_6576,N_3423,N_4379);
or U6577 (N_6577,N_4239,N_2568);
or U6578 (N_6578,N_3925,N_1888);
nand U6579 (N_6579,N_4883,N_1120);
or U6580 (N_6580,N_4404,N_1059);
or U6581 (N_6581,N_824,N_230);
or U6582 (N_6582,N_4398,N_1852);
or U6583 (N_6583,N_737,N_3628);
nand U6584 (N_6584,N_4123,N_3932);
nor U6585 (N_6585,N_779,N_2080);
and U6586 (N_6586,N_4788,N_2799);
or U6587 (N_6587,N_3914,N_3028);
nand U6588 (N_6588,N_4695,N_2778);
or U6589 (N_6589,N_3059,N_3060);
nor U6590 (N_6590,N_4303,N_3411);
nor U6591 (N_6591,N_3134,N_557);
nor U6592 (N_6592,N_3300,N_4881);
and U6593 (N_6593,N_3808,N_3876);
and U6594 (N_6594,N_3611,N_3386);
and U6595 (N_6595,N_297,N_965);
nand U6596 (N_6596,N_201,N_3448);
or U6597 (N_6597,N_4870,N_4712);
nand U6598 (N_6598,N_2483,N_2179);
and U6599 (N_6599,N_2536,N_1346);
nor U6600 (N_6600,N_4774,N_722);
nor U6601 (N_6601,N_2001,N_4701);
nand U6602 (N_6602,N_4206,N_3288);
nor U6603 (N_6603,N_3506,N_3903);
or U6604 (N_6604,N_498,N_4266);
nor U6605 (N_6605,N_2450,N_4315);
and U6606 (N_6606,N_3543,N_4080);
or U6607 (N_6607,N_4128,N_603);
and U6608 (N_6608,N_4370,N_2792);
nor U6609 (N_6609,N_4729,N_4970);
nor U6610 (N_6610,N_2797,N_263);
nand U6611 (N_6611,N_882,N_1990);
and U6612 (N_6612,N_2192,N_2811);
or U6613 (N_6613,N_967,N_2629);
nor U6614 (N_6614,N_4768,N_4144);
and U6615 (N_6615,N_611,N_4142);
nand U6616 (N_6616,N_4228,N_3762);
nand U6617 (N_6617,N_4455,N_685);
nand U6618 (N_6618,N_4241,N_3606);
or U6619 (N_6619,N_891,N_427);
nor U6620 (N_6620,N_1345,N_3823);
nand U6621 (N_6621,N_197,N_2848);
and U6622 (N_6622,N_4957,N_4615);
nand U6623 (N_6623,N_3737,N_2931);
or U6624 (N_6624,N_1045,N_2753);
nand U6625 (N_6625,N_3318,N_1146);
nand U6626 (N_6626,N_1447,N_4974);
and U6627 (N_6627,N_436,N_530);
nor U6628 (N_6628,N_4138,N_2549);
and U6629 (N_6629,N_3214,N_4625);
nor U6630 (N_6630,N_4093,N_1210);
and U6631 (N_6631,N_4642,N_1395);
nor U6632 (N_6632,N_3084,N_4388);
or U6633 (N_6633,N_3528,N_78);
nand U6634 (N_6634,N_2469,N_1879);
or U6635 (N_6635,N_3992,N_2943);
and U6636 (N_6636,N_3985,N_4525);
nand U6637 (N_6637,N_1433,N_4992);
nand U6638 (N_6638,N_4422,N_3246);
nand U6639 (N_6639,N_1728,N_1775);
and U6640 (N_6640,N_1881,N_634);
xnor U6641 (N_6641,N_1318,N_3778);
nand U6642 (N_6642,N_1019,N_2719);
nor U6643 (N_6643,N_4068,N_3945);
and U6644 (N_6644,N_1769,N_2526);
nor U6645 (N_6645,N_1349,N_339);
or U6646 (N_6646,N_812,N_4185);
and U6647 (N_6647,N_2497,N_447);
or U6648 (N_6648,N_4911,N_1475);
nand U6649 (N_6649,N_3739,N_1325);
nand U6650 (N_6650,N_1674,N_927);
nor U6651 (N_6651,N_827,N_3794);
nand U6652 (N_6652,N_2766,N_4858);
nand U6653 (N_6653,N_3526,N_681);
and U6654 (N_6654,N_1937,N_1698);
nor U6655 (N_6655,N_2921,N_2858);
nand U6656 (N_6656,N_3394,N_701);
or U6657 (N_6657,N_3328,N_768);
nor U6658 (N_6658,N_3351,N_2573);
nor U6659 (N_6659,N_2208,N_3701);
nand U6660 (N_6660,N_4621,N_2129);
nand U6661 (N_6661,N_310,N_2894);
and U6662 (N_6662,N_1272,N_8);
nand U6663 (N_6663,N_3262,N_2122);
and U6664 (N_6664,N_4180,N_661);
nand U6665 (N_6665,N_2419,N_4812);
or U6666 (N_6666,N_1150,N_2721);
nand U6667 (N_6667,N_1148,N_4821);
or U6668 (N_6668,N_3485,N_1818);
nor U6669 (N_6669,N_693,N_2164);
nor U6670 (N_6670,N_2320,N_2197);
or U6671 (N_6671,N_4999,N_4056);
and U6672 (N_6672,N_3420,N_4806);
nor U6673 (N_6673,N_315,N_138);
or U6674 (N_6674,N_640,N_3468);
nand U6675 (N_6675,N_1487,N_495);
and U6676 (N_6676,N_2524,N_3079);
nor U6677 (N_6677,N_4943,N_2738);
and U6678 (N_6678,N_4733,N_4810);
or U6679 (N_6679,N_4608,N_4995);
nor U6680 (N_6680,N_3957,N_537);
or U6681 (N_6681,N_4146,N_780);
nand U6682 (N_6682,N_2955,N_207);
nand U6683 (N_6683,N_1184,N_4948);
or U6684 (N_6684,N_2896,N_3862);
nor U6685 (N_6685,N_4929,N_1886);
and U6686 (N_6686,N_979,N_2621);
nor U6687 (N_6687,N_4176,N_1416);
and U6688 (N_6688,N_174,N_2936);
and U6689 (N_6689,N_2939,N_4131);
nor U6690 (N_6690,N_501,N_374);
or U6691 (N_6691,N_2306,N_3910);
or U6692 (N_6692,N_1640,N_4091);
nor U6693 (N_6693,N_1596,N_3818);
nand U6694 (N_6694,N_2342,N_769);
and U6695 (N_6695,N_4906,N_1348);
nand U6696 (N_6696,N_1908,N_2017);
and U6697 (N_6697,N_1790,N_2599);
nand U6698 (N_6698,N_3380,N_1404);
nor U6699 (N_6699,N_3845,N_2109);
or U6700 (N_6700,N_4963,N_928);
or U6701 (N_6701,N_2022,N_255);
and U6702 (N_6702,N_4993,N_2247);
xnor U6703 (N_6703,N_2531,N_1413);
nor U6704 (N_6704,N_791,N_3614);
and U6705 (N_6705,N_1822,N_3202);
nor U6706 (N_6706,N_3976,N_452);
and U6707 (N_6707,N_2967,N_800);
nor U6708 (N_6708,N_3595,N_763);
nor U6709 (N_6709,N_1812,N_3329);
and U6710 (N_6710,N_2791,N_4689);
or U6711 (N_6711,N_3795,N_2166);
or U6712 (N_6712,N_2959,N_2825);
or U6713 (N_6713,N_3294,N_1457);
nand U6714 (N_6714,N_1979,N_2638);
nor U6715 (N_6715,N_2917,N_2676);
and U6716 (N_6716,N_4041,N_2015);
or U6717 (N_6717,N_169,N_1188);
xnor U6718 (N_6718,N_1653,N_3074);
nand U6719 (N_6719,N_2317,N_4053);
or U6720 (N_6720,N_3301,N_1695);
nand U6721 (N_6721,N_4002,N_577);
nor U6722 (N_6722,N_2794,N_2103);
and U6723 (N_6723,N_4132,N_1012);
or U6724 (N_6724,N_2031,N_938);
or U6725 (N_6725,N_3863,N_1736);
or U6726 (N_6726,N_4635,N_831);
and U6727 (N_6727,N_3171,N_2490);
or U6728 (N_6728,N_982,N_4805);
and U6729 (N_6729,N_1570,N_57);
nor U6730 (N_6730,N_3708,N_3768);
or U6731 (N_6731,N_2724,N_4994);
nor U6732 (N_6732,N_1227,N_639);
or U6733 (N_6733,N_642,N_1789);
nor U6734 (N_6734,N_2114,N_2026);
and U6735 (N_6735,N_2596,N_3161);
xor U6736 (N_6736,N_2918,N_684);
nand U6737 (N_6737,N_1931,N_98);
nor U6738 (N_6738,N_3429,N_4302);
and U6739 (N_6739,N_273,N_3035);
and U6740 (N_6740,N_4437,N_128);
nor U6741 (N_6741,N_4247,N_541);
or U6742 (N_6742,N_20,N_162);
nand U6743 (N_6743,N_2087,N_2379);
nor U6744 (N_6744,N_724,N_2809);
and U6745 (N_6745,N_2922,N_4441);
nor U6746 (N_6746,N_1626,N_4386);
nand U6747 (N_6747,N_3759,N_3769);
nand U6748 (N_6748,N_4210,N_2252);
or U6749 (N_6749,N_4514,N_3184);
nand U6750 (N_6750,N_2202,N_258);
nand U6751 (N_6751,N_3197,N_3981);
and U6752 (N_6752,N_3937,N_3612);
nor U6753 (N_6753,N_3282,N_4991);
nor U6754 (N_6754,N_3276,N_719);
and U6755 (N_6755,N_2486,N_1308);
nor U6756 (N_6756,N_2236,N_2542);
and U6757 (N_6757,N_1998,N_4637);
or U6758 (N_6758,N_267,N_3070);
and U6759 (N_6759,N_4279,N_4847);
and U6760 (N_6760,N_3383,N_2013);
nor U6761 (N_6761,N_3226,N_2310);
nor U6762 (N_6762,N_1163,N_1351);
nand U6763 (N_6763,N_2387,N_3257);
or U6764 (N_6764,N_3218,N_1030);
nand U6765 (N_6765,N_1561,N_233);
nor U6766 (N_6766,N_3836,N_1164);
or U6767 (N_6767,N_3144,N_4967);
and U6768 (N_6768,N_4904,N_93);
nand U6769 (N_6769,N_1101,N_3849);
and U6770 (N_6770,N_4551,N_2749);
nor U6771 (N_6771,N_3505,N_2107);
and U6772 (N_6772,N_4659,N_2398);
and U6773 (N_6773,N_3146,N_3847);
nand U6774 (N_6774,N_1975,N_3901);
or U6775 (N_6775,N_4391,N_3405);
or U6776 (N_6776,N_1061,N_420);
or U6777 (N_6777,N_385,N_366);
nand U6778 (N_6778,N_571,N_341);
nand U6779 (N_6779,N_305,N_4368);
or U6780 (N_6780,N_1063,N_2628);
nand U6781 (N_6781,N_2924,N_3071);
nand U6782 (N_6782,N_2036,N_2564);
and U6783 (N_6783,N_876,N_621);
or U6784 (N_6784,N_2408,N_3477);
nor U6785 (N_6785,N_1183,N_3299);
nand U6786 (N_6786,N_1725,N_4890);
nand U6787 (N_6787,N_2610,N_2570);
and U6788 (N_6788,N_4154,N_949);
nor U6789 (N_6789,N_4282,N_620);
or U6790 (N_6790,N_3780,N_2624);
and U6791 (N_6791,N_4498,N_3309);
and U6792 (N_6792,N_4431,N_4835);
or U6793 (N_6793,N_1020,N_3271);
nand U6794 (N_6794,N_2633,N_3399);
nand U6795 (N_6795,N_1159,N_3817);
nor U6796 (N_6796,N_4751,N_3545);
nand U6797 (N_6797,N_4221,N_880);
nand U6798 (N_6798,N_4475,N_871);
nand U6799 (N_6799,N_390,N_2873);
nor U6800 (N_6800,N_3607,N_3962);
nand U6801 (N_6801,N_2732,N_811);
and U6802 (N_6802,N_1245,N_3255);
and U6803 (N_6803,N_1971,N_4078);
nor U6804 (N_6804,N_4317,N_3613);
nor U6805 (N_6805,N_1250,N_4331);
and U6806 (N_6806,N_3681,N_3987);
and U6807 (N_6807,N_1249,N_3120);
nand U6808 (N_6808,N_1373,N_3272);
or U6809 (N_6809,N_1876,N_1085);
nand U6810 (N_6810,N_817,N_3356);
and U6811 (N_6811,N_2204,N_4938);
or U6812 (N_6812,N_1269,N_3222);
nor U6813 (N_6813,N_2263,N_4191);
and U6814 (N_6814,N_379,N_4170);
and U6815 (N_6815,N_1186,N_4946);
and U6816 (N_6816,N_1607,N_4011);
nand U6817 (N_6817,N_2,N_2384);
xor U6818 (N_6818,N_1015,N_4749);
or U6819 (N_6819,N_3310,N_1558);
and U6820 (N_6820,N_852,N_1032);
nor U6821 (N_6821,N_1993,N_1481);
nor U6822 (N_6822,N_3263,N_1078);
and U6823 (N_6823,N_4687,N_1521);
or U6824 (N_6824,N_237,N_126);
nand U6825 (N_6825,N_3647,N_4095);
nor U6826 (N_6826,N_1202,N_1068);
nand U6827 (N_6827,N_1539,N_2742);
nand U6828 (N_6828,N_786,N_2170);
and U6829 (N_6829,N_3424,N_1992);
or U6830 (N_6830,N_3736,N_3774);
and U6831 (N_6831,N_3897,N_595);
xnor U6832 (N_6832,N_2852,N_4594);
xor U6833 (N_6833,N_2986,N_4433);
and U6834 (N_6834,N_1415,N_462);
or U6835 (N_6835,N_4833,N_1048);
or U6836 (N_6836,N_1356,N_1081);
and U6837 (N_6837,N_1598,N_4480);
nor U6838 (N_6838,N_1782,N_409);
nor U6839 (N_6839,N_2737,N_1981);
or U6840 (N_6840,N_3640,N_3743);
nand U6841 (N_6841,N_4919,N_2736);
nor U6842 (N_6842,N_3,N_3973);
or U6843 (N_6843,N_1339,N_2636);
nand U6844 (N_6844,N_4700,N_1527);
xnor U6845 (N_6845,N_3535,N_3570);
or U6846 (N_6846,N_675,N_3392);
nand U6847 (N_6847,N_565,N_43);
or U6848 (N_6848,N_1309,N_3107);
nor U6849 (N_6849,N_4451,N_3138);
nor U6850 (N_6850,N_2025,N_3115);
or U6851 (N_6851,N_2091,N_4880);
nand U6852 (N_6852,N_3403,N_4884);
nand U6853 (N_6853,N_711,N_1503);
and U6854 (N_6854,N_3511,N_4844);
nand U6855 (N_6855,N_1613,N_1244);
or U6856 (N_6856,N_3269,N_3179);
nand U6857 (N_6857,N_4092,N_3007);
nor U6858 (N_6858,N_2184,N_2213);
nor U6859 (N_6859,N_1685,N_4614);
nor U6860 (N_6860,N_9,N_3258);
and U6861 (N_6861,N_4566,N_4291);
nand U6862 (N_6862,N_4632,N_3646);
nor U6863 (N_6863,N_504,N_1074);
nand U6864 (N_6864,N_1621,N_2113);
nor U6865 (N_6865,N_1261,N_120);
and U6866 (N_6866,N_1764,N_3676);
nand U6867 (N_6867,N_2530,N_3347);
or U6868 (N_6868,N_1533,N_2787);
and U6869 (N_6869,N_40,N_4575);
or U6870 (N_6870,N_3462,N_2090);
and U6871 (N_6871,N_1836,N_2698);
nand U6872 (N_6872,N_2203,N_3731);
nand U6873 (N_6873,N_4802,N_1054);
nand U6874 (N_6874,N_4997,N_2847);
xor U6875 (N_6875,N_3154,N_1412);
nor U6876 (N_6876,N_1258,N_4120);
or U6877 (N_6877,N_4908,N_2614);
and U6878 (N_6878,N_600,N_4887);
nand U6879 (N_6879,N_4322,N_1827);
nor U6880 (N_6880,N_2475,N_1463);
nand U6881 (N_6881,N_1536,N_275);
nand U6882 (N_6882,N_4962,N_177);
or U6883 (N_6883,N_4773,N_1166);
or U6884 (N_6884,N_3970,N_1804);
nor U6885 (N_6885,N_3117,N_756);
and U6886 (N_6886,N_1984,N_430);
nand U6887 (N_6887,N_4129,N_3713);
nor U6888 (N_6888,N_959,N_1006);
and U6889 (N_6889,N_1248,N_1140);
and U6890 (N_6890,N_2525,N_1008);
nand U6891 (N_6891,N_4973,N_4427);
nor U6892 (N_6892,N_1458,N_3608);
nand U6893 (N_6893,N_311,N_2422);
or U6894 (N_6894,N_4528,N_1831);
nor U6895 (N_6895,N_3064,N_4682);
nand U6896 (N_6896,N_1191,N_1980);
xor U6897 (N_6897,N_4334,N_225);
and U6898 (N_6898,N_886,N_1219);
nand U6899 (N_6899,N_4604,N_4736);
and U6900 (N_6900,N_4501,N_4339);
and U6901 (N_6901,N_1131,N_41);
nor U6902 (N_6902,N_4492,N_15);
and U6903 (N_6903,N_1029,N_3103);
xor U6904 (N_6904,N_3253,N_3168);
xor U6905 (N_6905,N_166,N_4106);
and U6906 (N_6906,N_2199,N_285);
or U6907 (N_6907,N_781,N_1300);
or U6908 (N_6908,N_1231,N_3196);
or U6909 (N_6909,N_116,N_1893);
and U6910 (N_6910,N_2952,N_3534);
nor U6911 (N_6911,N_4034,N_1194);
or U6912 (N_6912,N_823,N_1602);
nand U6913 (N_6913,N_801,N_2227);
nor U6914 (N_6914,N_2984,N_1901);
nor U6915 (N_6915,N_715,N_4172);
nor U6916 (N_6916,N_1684,N_2729);
and U6917 (N_6917,N_4008,N_1837);
and U6918 (N_6918,N_3187,N_602);
nor U6919 (N_6919,N_2326,N_3118);
nor U6920 (N_6920,N_792,N_4054);
nor U6921 (N_6921,N_2760,N_1233);
and U6922 (N_6922,N_1050,N_2750);
or U6923 (N_6923,N_322,N_3338);
or U6924 (N_6924,N_3030,N_1651);
xor U6925 (N_6925,N_125,N_906);
or U6926 (N_6926,N_535,N_1161);
nand U6927 (N_6927,N_2585,N_657);
or U6928 (N_6928,N_3781,N_3241);
nand U6929 (N_6929,N_1320,N_3091);
or U6930 (N_6930,N_4716,N_200);
or U6931 (N_6931,N_4353,N_4895);
nand U6932 (N_6932,N_4496,N_3359);
nand U6933 (N_6933,N_2571,N_531);
nor U6934 (N_6934,N_3406,N_1176);
and U6935 (N_6935,N_3224,N_3507);
nor U6936 (N_6936,N_28,N_4283);
and U6937 (N_6937,N_2983,N_439);
and U6938 (N_6938,N_3451,N_247);
or U6939 (N_6939,N_3951,N_749);
or U6940 (N_6940,N_2770,N_854);
and U6941 (N_6941,N_4125,N_4569);
nand U6942 (N_6942,N_1437,N_1180);
and U6943 (N_6943,N_2516,N_2649);
or U6944 (N_6944,N_4218,N_2034);
or U6945 (N_6945,N_1343,N_3334);
and U6946 (N_6946,N_2853,N_4024);
or U6947 (N_6947,N_4706,N_4186);
and U6948 (N_6948,N_4730,N_1828);
xor U6949 (N_6949,N_4069,N_3803);
nor U6950 (N_6950,N_4030,N_2500);
and U6951 (N_6951,N_559,N_2812);
or U6952 (N_6952,N_942,N_241);
nor U6953 (N_6953,N_0,N_2058);
nor U6954 (N_6954,N_1671,N_1398);
or U6955 (N_6955,N_4705,N_2072);
and U6956 (N_6956,N_4913,N_1070);
or U6957 (N_6957,N_1986,N_785);
nor U6958 (N_6958,N_4413,N_1519);
and U6959 (N_6959,N_1856,N_1234);
and U6960 (N_6960,N_3641,N_1940);
or U6961 (N_6961,N_318,N_1031);
or U6962 (N_6962,N_312,N_1236);
or U6963 (N_6963,N_4853,N_4325);
or U6964 (N_6964,N_637,N_4058);
and U6965 (N_6965,N_85,N_489);
and U6966 (N_6966,N_3374,N_1401);
and U6967 (N_6967,N_960,N_1508);
nand U6968 (N_6968,N_1904,N_49);
and U6969 (N_6969,N_1917,N_1661);
or U6970 (N_6970,N_4188,N_1676);
nand U6971 (N_6971,N_4759,N_847);
or U6972 (N_6972,N_4636,N_3495);
or U6973 (N_6973,N_883,N_3317);
nor U6974 (N_6974,N_3210,N_2499);
or U6975 (N_6975,N_1436,N_2618);
or U6976 (N_6976,N_3234,N_861);
and U6977 (N_6977,N_2003,N_4117);
or U6978 (N_6978,N_4360,N_3488);
or U6979 (N_6979,N_874,N_3327);
or U6980 (N_6980,N_1064,N_490);
and U6981 (N_6981,N_1495,N_3114);
nor U6982 (N_6982,N_873,N_1887);
nand U6983 (N_6983,N_4294,N_1037);
and U6984 (N_6984,N_555,N_4912);
nor U6985 (N_6985,N_4031,N_4861);
or U6986 (N_6986,N_3698,N_1587);
nand U6987 (N_6987,N_2237,N_264);
and U6988 (N_6988,N_2949,N_3401);
and U6989 (N_6989,N_964,N_4738);
xor U6990 (N_6990,N_1754,N_2371);
nor U6991 (N_6991,N_1703,N_2144);
nand U6992 (N_6992,N_2869,N_3875);
nand U6993 (N_6993,N_3742,N_3039);
or U6994 (N_6994,N_2307,N_536);
nand U6995 (N_6995,N_352,N_3132);
nor U6996 (N_6996,N_443,N_3967);
nand U6997 (N_6997,N_690,N_734);
nor U6998 (N_6998,N_4479,N_1419);
or U6999 (N_6999,N_18,N_869);
xor U7000 (N_7000,N_3371,N_1556);
or U7001 (N_7001,N_1390,N_890);
or U7002 (N_7002,N_2566,N_2930);
or U7003 (N_7003,N_1439,N_62);
nor U7004 (N_7004,N_1637,N_3746);
and U7005 (N_7005,N_805,N_3377);
or U7006 (N_7006,N_1735,N_1026);
nand U7007 (N_7007,N_1814,N_2658);
nor U7008 (N_7008,N_3574,N_227);
nor U7009 (N_7009,N_4338,N_679);
and U7010 (N_7010,N_4914,N_4857);
or U7011 (N_7011,N_470,N_3368);
or U7012 (N_7012,N_810,N_930);
nand U7013 (N_7013,N_2643,N_3036);
and U7014 (N_7014,N_1595,N_3978);
nand U7015 (N_7015,N_3087,N_741);
and U7016 (N_7016,N_2891,N_3829);
nand U7017 (N_7017,N_1392,N_367);
xor U7018 (N_7018,N_1360,N_2108);
nand U7019 (N_7019,N_372,N_2718);
nand U7020 (N_7020,N_4703,N_723);
or U7021 (N_7021,N_1151,N_1259);
or U7022 (N_7022,N_2046,N_2101);
nor U7023 (N_7023,N_1914,N_3868);
or U7024 (N_7024,N_1165,N_3787);
nor U7025 (N_7025,N_3363,N_2147);
nor U7026 (N_7026,N_932,N_2543);
nand U7027 (N_7027,N_2540,N_929);
nand U7028 (N_7028,N_651,N_1650);
or U7029 (N_7029,N_3169,N_4007);
nor U7030 (N_7030,N_2838,N_1431);
and U7031 (N_7031,N_1005,N_429);
and U7032 (N_7032,N_2937,N_4306);
and U7033 (N_7033,N_2280,N_1743);
nand U7034 (N_7034,N_3116,N_3982);
or U7035 (N_7035,N_3587,N_4658);
nand U7036 (N_7036,N_3796,N_659);
and U7037 (N_7037,N_1294,N_2977);
nand U7038 (N_7038,N_3092,N_2956);
and U7039 (N_7039,N_163,N_1972);
nand U7040 (N_7040,N_686,N_2054);
nor U7041 (N_7041,N_730,N_3204);
or U7042 (N_7042,N_3715,N_1496);
and U7043 (N_7043,N_326,N_4432);
nor U7044 (N_7044,N_56,N_1622);
nor U7045 (N_7045,N_3615,N_1141);
nor U7046 (N_7046,N_776,N_4016);
and U7047 (N_7047,N_610,N_1446);
nor U7048 (N_7048,N_4775,N_1152);
or U7049 (N_7049,N_3633,N_2067);
and U7050 (N_7050,N_2920,N_560);
and U7051 (N_7051,N_920,N_2562);
nand U7052 (N_7052,N_2372,N_3554);
and U7053 (N_7053,N_3219,N_2456);
or U7054 (N_7054,N_4112,N_1281);
and U7055 (N_7055,N_1928,N_3656);
nand U7056 (N_7056,N_89,N_4209);
or U7057 (N_7057,N_978,N_3706);
nor U7058 (N_7058,N_4318,N_2660);
nor U7059 (N_7059,N_1315,N_3693);
nor U7060 (N_7060,N_1384,N_1228);
and U7061 (N_7061,N_4336,N_1411);
or U7062 (N_7062,N_4122,N_3008);
and U7063 (N_7063,N_4029,N_2607);
or U7064 (N_7064,N_1506,N_4985);
nand U7065 (N_7065,N_3689,N_548);
and U7066 (N_7066,N_389,N_4443);
and U7067 (N_7067,N_4272,N_3345);
nand U7068 (N_7068,N_2376,N_2311);
and U7069 (N_7069,N_47,N_3882);
and U7070 (N_7070,N_12,N_1347);
and U7071 (N_7071,N_3797,N_86);
nand U7072 (N_7072,N_2434,N_4509);
nor U7073 (N_7073,N_3081,N_1934);
nand U7074 (N_7074,N_466,N_4346);
nor U7075 (N_7075,N_2004,N_4028);
nand U7076 (N_7076,N_4680,N_804);
or U7077 (N_7077,N_3659,N_3189);
and U7078 (N_7078,N_4237,N_1663);
nand U7079 (N_7079,N_1033,N_21);
or U7080 (N_7080,N_3373,N_2595);
nand U7081 (N_7081,N_3566,N_1091);
or U7082 (N_7082,N_1505,N_2520);
nand U7083 (N_7083,N_4060,N_2137);
or U7084 (N_7084,N_3032,N_658);
xor U7085 (N_7085,N_4373,N_4190);
or U7086 (N_7086,N_3990,N_4445);
nor U7087 (N_7087,N_4196,N_2325);
nor U7088 (N_7088,N_152,N_4630);
nand U7089 (N_7089,N_3542,N_1088);
nand U7090 (N_7090,N_2888,N_646);
nand U7091 (N_7091,N_4456,N_4905);
nand U7092 (N_7092,N_167,N_229);
nand U7093 (N_7093,N_4564,N_293);
xnor U7094 (N_7094,N_1659,N_596);
nand U7095 (N_7095,N_2669,N_4656);
or U7096 (N_7096,N_196,N_4685);
nor U7097 (N_7097,N_1307,N_1512);
nor U7098 (N_7098,N_1552,N_243);
or U7099 (N_7099,N_392,N_3726);
nand U7100 (N_7100,N_4424,N_2944);
or U7101 (N_7101,N_2927,N_2581);
and U7102 (N_7102,N_333,N_37);
nor U7103 (N_7103,N_488,N_3889);
nand U7104 (N_7104,N_514,N_568);
nor U7105 (N_7105,N_4152,N_4555);
and U7106 (N_7106,N_216,N_1009);
nor U7107 (N_7107,N_2189,N_53);
nand U7108 (N_7108,N_280,N_1634);
or U7109 (N_7109,N_1683,N_346);
and U7110 (N_7110,N_2995,N_2478);
nor U7111 (N_7111,N_1540,N_3588);
nand U7112 (N_7112,N_1364,N_4109);
nand U7113 (N_7113,N_910,N_1203);
or U7114 (N_7114,N_3206,N_2397);
xnor U7115 (N_7115,N_3090,N_2097);
and U7116 (N_7116,N_515,N_3433);
or U7117 (N_7117,N_4087,N_3991);
and U7118 (N_7118,N_4471,N_2229);
nor U7119 (N_7119,N_2529,N_668);
nor U7120 (N_7120,N_4885,N_2127);
nand U7121 (N_7121,N_4839,N_2256);
nand U7122 (N_7122,N_4585,N_3095);
nor U7123 (N_7123,N_2836,N_4965);
or U7124 (N_7124,N_153,N_3583);
or U7125 (N_7125,N_2443,N_507);
nor U7126 (N_7126,N_4136,N_3519);
nor U7127 (N_7127,N_1201,N_3348);
or U7128 (N_7128,N_672,N_2205);
and U7129 (N_7129,N_1696,N_665);
or U7130 (N_7130,N_4639,N_2211);
and U7131 (N_7131,N_2867,N_2586);
nor U7132 (N_7132,N_1791,N_2126);
and U7133 (N_7133,N_4110,N_985);
nand U7134 (N_7134,N_3801,N_4219);
nand U7135 (N_7135,N_1485,N_1714);
nor U7136 (N_7136,N_2641,N_4372);
and U7137 (N_7137,N_3832,N_4474);
nand U7138 (N_7138,N_694,N_4747);
and U7139 (N_7139,N_4466,N_2238);
and U7140 (N_7140,N_2425,N_1656);
or U7141 (N_7141,N_2047,N_674);
and U7142 (N_7142,N_4878,N_3040);
and U7143 (N_7143,N_2438,N_4882);
or U7144 (N_7144,N_4337,N_4260);
nor U7145 (N_7145,N_2411,N_2733);
or U7146 (N_7146,N_349,N_3677);
or U7147 (N_7147,N_4429,N_3547);
nor U7148 (N_7148,N_1548,N_2118);
or U7149 (N_7149,N_3848,N_2044);
or U7150 (N_7150,N_414,N_947);
and U7151 (N_7151,N_3675,N_4408);
nor U7152 (N_7152,N_4001,N_232);
and U7153 (N_7153,N_3822,N_2268);
xnor U7154 (N_7154,N_4167,N_3667);
or U7155 (N_7155,N_1709,N_673);
and U7156 (N_7156,N_4697,N_7);
nor U7157 (N_7157,N_627,N_2424);
nor U7158 (N_7158,N_3450,N_1752);
nor U7159 (N_7159,N_1442,N_1362);
or U7160 (N_7160,N_2631,N_4792);
or U7161 (N_7161,N_4672,N_245);
or U7162 (N_7162,N_1777,N_84);
nor U7163 (N_7163,N_3538,N_2262);
and U7164 (N_7164,N_1492,N_4977);
nor U7165 (N_7165,N_3320,N_1936);
and U7166 (N_7166,N_2028,N_2367);
or U7167 (N_7167,N_3963,N_4450);
xor U7168 (N_7168,N_4063,N_3136);
nor U7169 (N_7169,N_3512,N_3658);
nor U7170 (N_7170,N_3730,N_1938);
nor U7171 (N_7171,N_1907,N_4444);
or U7172 (N_7172,N_1861,N_2363);
nor U7173 (N_7173,N_342,N_3441);
nand U7174 (N_7174,N_2436,N_4927);
and U7175 (N_7175,N_4251,N_2783);
nor U7176 (N_7176,N_3789,N_3531);
nor U7177 (N_7177,N_527,N_2266);
or U7178 (N_7178,N_3358,N_4607);
nor U7179 (N_7179,N_3879,N_3337);
or U7180 (N_7180,N_2842,N_4573);
and U7181 (N_7181,N_3004,N_878);
or U7182 (N_7182,N_2834,N_1084);
nor U7183 (N_7183,N_3203,N_1456);
or U7184 (N_7184,N_4421,N_4311);
nand U7185 (N_7185,N_2173,N_4018);
nor U7186 (N_7186,N_4211,N_2541);
nor U7187 (N_7187,N_3098,N_4472);
nor U7188 (N_7188,N_4048,N_2125);
and U7189 (N_7189,N_993,N_4295);
or U7190 (N_7190,N_2099,N_4952);
or U7191 (N_7191,N_1701,N_922);
nand U7192 (N_7192,N_762,N_3952);
or U7193 (N_7193,N_1591,N_4320);
nor U7194 (N_7194,N_300,N_2538);
and U7195 (N_7195,N_4401,N_3048);
nand U7196 (N_7196,N_1719,N_2035);
nand U7197 (N_7197,N_1853,N_4467);
nand U7198 (N_7198,N_3003,N_4641);
nand U7199 (N_7199,N_3908,N_1705);
nor U7200 (N_7200,N_4299,N_677);
nand U7201 (N_7201,N_1953,N_2338);
or U7202 (N_7202,N_893,N_1816);
and U7203 (N_7203,N_2992,N_2343);
nor U7204 (N_7204,N_1982,N_2344);
and U7205 (N_7205,N_2030,N_1502);
and U7206 (N_7206,N_2224,N_1813);
nand U7207 (N_7207,N_1708,N_2060);
nand U7208 (N_7208,N_688,N_1865);
nand U7209 (N_7209,N_2843,N_1898);
and U7210 (N_7210,N_2819,N_2916);
or U7211 (N_7211,N_1414,N_1480);
and U7212 (N_7212,N_1213,N_3129);
or U7213 (N_7213,N_1328,N_1196);
nor U7214 (N_7214,N_4803,N_2119);
and U7215 (N_7215,N_291,N_1997);
and U7216 (N_7216,N_2352,N_2948);
and U7217 (N_7217,N_2180,N_833);
and U7218 (N_7218,N_856,N_4208);
nand U7219 (N_7219,N_1504,N_1925);
nor U7220 (N_7220,N_970,N_261);
nor U7221 (N_7221,N_487,N_1730);
or U7222 (N_7222,N_1718,N_3178);
or U7223 (N_7223,N_1223,N_1648);
or U7224 (N_7224,N_234,N_4037);
nand U7225 (N_7225,N_1226,N_3598);
or U7226 (N_7226,N_911,N_612);
and U7227 (N_7227,N_1197,N_1000);
or U7228 (N_7228,N_1864,N_1222);
nand U7229 (N_7229,N_2210,N_2941);
nand U7230 (N_7230,N_4292,N_1711);
nor U7231 (N_7231,N_1895,N_2092);
nor U7232 (N_7232,N_3217,N_1337);
nor U7233 (N_7233,N_90,N_3001);
or U7234 (N_7234,N_699,N_27);
or U7235 (N_7235,N_4361,N_1869);
nand U7236 (N_7236,N_222,N_4655);
nor U7237 (N_7237,N_4105,N_3487);
and U7238 (N_7238,N_2131,N_337);
nor U7239 (N_7239,N_1669,N_4263);
nor U7240 (N_7240,N_914,N_2816);
nor U7241 (N_7241,N_382,N_4227);
nor U7242 (N_7242,N_4104,N_1976);
nor U7243 (N_7243,N_3573,N_2295);
nor U7244 (N_7244,N_2835,N_1803);
nand U7245 (N_7245,N_3292,N_4084);
and U7246 (N_7246,N_3058,N_2758);
nor U7247 (N_7247,N_3076,N_1847);
nor U7248 (N_7248,N_24,N_67);
or U7249 (N_7249,N_170,N_2951);
and U7250 (N_7250,N_4780,N_4826);
nor U7251 (N_7251,N_477,N_3198);
nor U7252 (N_7252,N_4646,N_1594);
or U7253 (N_7253,N_444,N_4463);
xor U7254 (N_7254,N_4951,N_29);
or U7255 (N_7255,N_1137,N_4328);
and U7256 (N_7256,N_841,N_368);
and U7257 (N_7257,N_2021,N_3298);
nor U7258 (N_7258,N_458,N_3389);
nand U7259 (N_7259,N_136,N_3273);
nor U7260 (N_7260,N_3784,N_3986);
and U7261 (N_7261,N_2823,N_2235);
and U7262 (N_7262,N_1239,N_2079);
or U7263 (N_7263,N_1047,N_4151);
nor U7264 (N_7264,N_3398,N_897);
nand U7265 (N_7265,N_3034,N_866);
or U7266 (N_7266,N_3525,N_1332);
and U7267 (N_7267,N_3493,N_1177);
nor U7268 (N_7268,N_941,N_3303);
nor U7269 (N_7269,N_4202,N_3396);
nand U7270 (N_7270,N_1397,N_2057);
or U7271 (N_7271,N_260,N_2431);
nand U7272 (N_7272,N_4140,N_2874);
or U7273 (N_7273,N_550,N_4021);
xnor U7274 (N_7274,N_3280,N_512);
nand U7275 (N_7275,N_4232,N_2024);
or U7276 (N_7276,N_141,N_3341);
and U7277 (N_7277,N_943,N_284);
and U7278 (N_7278,N_1707,N_3471);
and U7279 (N_7279,N_586,N_4766);
nor U7280 (N_7280,N_3663,N_2725);
or U7281 (N_7281,N_503,N_178);
nor U7282 (N_7282,N_1058,N_1958);
and U7283 (N_7283,N_2752,N_176);
or U7284 (N_7284,N_4626,N_2168);
nor U7285 (N_7285,N_1862,N_575);
xnor U7286 (N_7286,N_1144,N_4936);
nand U7287 (N_7287,N_4183,N_3821);
or U7288 (N_7288,N_875,N_4134);
nand U7289 (N_7289,N_3605,N_3955);
and U7290 (N_7290,N_4548,N_2881);
xnor U7291 (N_7291,N_4772,N_3959);
and U7292 (N_7292,N_3763,N_142);
nand U7293 (N_7293,N_472,N_983);
nand U7294 (N_7294,N_919,N_1848);
and U7295 (N_7295,N_1662,N_1890);
and U7296 (N_7296,N_2124,N_279);
and U7297 (N_7297,N_1168,N_4577);
nor U7298 (N_7298,N_3552,N_2476);
and U7299 (N_7299,N_567,N_217);
or U7300 (N_7300,N_3733,N_4903);
and U7301 (N_7301,N_1582,N_2465);
or U7302 (N_7302,N_2228,N_4651);
nor U7303 (N_7303,N_3857,N_2741);
nor U7304 (N_7304,N_4746,N_635);
and U7305 (N_7305,N_704,N_881);
or U7306 (N_7306,N_2112,N_1111);
nor U7307 (N_7307,N_862,N_3474);
or U7308 (N_7308,N_4828,N_3438);
and U7309 (N_7309,N_1682,N_2517);
nor U7310 (N_7310,N_4871,N_4199);
and U7311 (N_7311,N_3213,N_4765);
nand U7312 (N_7312,N_1532,N_1182);
nand U7313 (N_7313,N_3651,N_4676);
nor U7314 (N_7314,N_3883,N_1252);
nand U7315 (N_7315,N_66,N_2923);
nor U7316 (N_7316,N_2094,N_4629);
nand U7317 (N_7317,N_3190,N_3714);
and U7318 (N_7318,N_1298,N_4494);
xor U7319 (N_7319,N_1566,N_509);
nand U7320 (N_7320,N_4070,N_523);
nand U7321 (N_7321,N_3792,N_4392);
nand U7322 (N_7322,N_4088,N_4099);
nand U7323 (N_7323,N_698,N_2957);
and U7324 (N_7324,N_3567,N_3532);
or U7325 (N_7325,N_3805,N_3391);
nor U7326 (N_7326,N_3518,N_1096);
nand U7327 (N_7327,N_1523,N_2264);
and U7328 (N_7328,N_2050,N_2840);
nor U7329 (N_7329,N_598,N_3591);
or U7330 (N_7330,N_3673,N_4352);
or U7331 (N_7331,N_2249,N_1069);
and U7332 (N_7332,N_2386,N_2945);
nand U7333 (N_7333,N_2321,N_3919);
and U7334 (N_7334,N_4649,N_4205);
or U7335 (N_7335,N_2743,N_2451);
nor U7336 (N_7336,N_4497,N_2254);
nor U7337 (N_7337,N_3153,N_3018);
or U7338 (N_7338,N_2557,N_1524);
nand U7339 (N_7339,N_656,N_2349);
or U7340 (N_7340,N_4900,N_4399);
nand U7341 (N_7341,N_4518,N_4664);
nand U7342 (N_7342,N_1859,N_689);
and U7343 (N_7343,N_4510,N_1477);
nor U7344 (N_7344,N_3935,N_2861);
nor U7345 (N_7345,N_2576,N_2558);
nand U7346 (N_7346,N_4599,N_4010);
nand U7347 (N_7347,N_4064,N_2609);
xnor U7348 (N_7348,N_4671,N_3097);
nand U7349 (N_7349,N_4832,N_3355);
and U7350 (N_7350,N_2427,N_1877);
nand U7351 (N_7351,N_1664,N_2890);
xor U7352 (N_7352,N_1617,N_425);
nor U7353 (N_7353,N_4665,N_3207);
and U7354 (N_7354,N_355,N_3361);
nor U7355 (N_7355,N_3670,N_4309);
nand U7356 (N_7356,N_4955,N_2554);
and U7357 (N_7357,N_647,N_2145);
nor U7358 (N_7358,N_4761,N_4469);
nand U7359 (N_7359,N_2088,N_1200);
nor U7360 (N_7360,N_35,N_3974);
and U7361 (N_7361,N_4778,N_3953);
and U7362 (N_7362,N_2744,N_1619);
nor U7363 (N_7363,N_107,N_4254);
nor U7364 (N_7364,N_4234,N_2532);
nor U7365 (N_7365,N_4348,N_4359);
and U7366 (N_7366,N_905,N_1868);
nor U7367 (N_7367,N_3478,N_3825);
or U7368 (N_7368,N_1038,N_83);
nor U7369 (N_7369,N_412,N_2971);
xor U7370 (N_7370,N_3067,N_1016);
and U7371 (N_7371,N_4797,N_2358);
nor U7372 (N_7372,N_4267,N_2776);
and U7373 (N_7373,N_1410,N_2851);
nor U7374 (N_7374,N_1605,N_3690);
or U7375 (N_7375,N_1673,N_2786);
or U7376 (N_7376,N_606,N_663);
nor U7377 (N_7377,N_4143,N_2135);
nand U7378 (N_7378,N_4827,N_709);
or U7379 (N_7379,N_482,N_1734);
and U7380 (N_7380,N_3539,N_2394);
or U7381 (N_7381,N_1367,N_407);
and U7382 (N_7382,N_2671,N_2720);
and U7383 (N_7383,N_1680,N_2706);
nor U7384 (N_7384,N_2206,N_165);
and U7385 (N_7385,N_3719,N_3350);
or U7386 (N_7386,N_2691,N_4742);
or U7387 (N_7387,N_127,N_829);
or U7388 (N_7388,N_3455,N_1947);
nand U7389 (N_7389,N_2735,N_203);
and U7390 (N_7390,N_2299,N_2814);
nand U7391 (N_7391,N_2518,N_2149);
nand U7392 (N_7392,N_186,N_3657);
or U7393 (N_7393,N_599,N_3256);
and U7394 (N_7394,N_1768,N_4077);
nor U7395 (N_7395,N_2903,N_4726);
or U7396 (N_7396,N_380,N_1057);
and U7397 (N_7397,N_370,N_520);
nand U7398 (N_7398,N_4667,N_819);
or U7399 (N_7399,N_3643,N_1943);
nand U7400 (N_7400,N_4340,N_328);
nor U7401 (N_7401,N_3824,N_884);
or U7402 (N_7402,N_3267,N_4304);
or U7403 (N_7403,N_744,N_3268);
and U7404 (N_7404,N_2775,N_4618);
and U7405 (N_7405,N_4158,N_3579);
nor U7406 (N_7406,N_2182,N_3459);
nand U7407 (N_7407,N_159,N_3082);
and U7408 (N_7408,N_2139,N_1277);
nor U7409 (N_7409,N_1100,N_725);
xnor U7410 (N_7410,N_4886,N_969);
nor U7411 (N_7411,N_432,N_2133);
and U7412 (N_7412,N_2800,N_3521);
nand U7413 (N_7413,N_1382,N_2225);
nor U7414 (N_7414,N_2466,N_2966);
or U7415 (N_7415,N_4415,N_1271);
nor U7416 (N_7416,N_2594,N_193);
nor U7417 (N_7417,N_4848,N_2755);
xnor U7418 (N_7418,N_381,N_958);
and U7419 (N_7419,N_3885,N_774);
and U7420 (N_7420,N_1232,N_2991);
nor U7421 (N_7421,N_3402,N_2978);
and U7422 (N_7422,N_497,N_4782);
nor U7423 (N_7423,N_3793,N_3947);
nand U7424 (N_7424,N_1491,N_4743);
or U7425 (N_7425,N_1948,N_4623);
nand U7426 (N_7426,N_2826,N_556);
and U7427 (N_7427,N_1880,N_3342);
or U7428 (N_7428,N_2043,N_2155);
and U7429 (N_7429,N_2005,N_3027);
nor U7430 (N_7430,N_4872,N_156);
nor U7431 (N_7431,N_1338,N_1579);
or U7432 (N_7432,N_3414,N_2253);
nor U7433 (N_7433,N_3649,N_2588);
or U7434 (N_7434,N_2485,N_2677);
and U7435 (N_7435,N_1035,N_71);
nand U7436 (N_7436,N_687,N_2827);
or U7437 (N_7437,N_63,N_2250);
and U7438 (N_7438,N_1772,N_3416);
and U7439 (N_7439,N_1687,N_1810);
nand U7440 (N_7440,N_4557,N_1089);
nor U7441 (N_7441,N_259,N_2242);
and U7442 (N_7442,N_872,N_3594);
or U7443 (N_7443,N_4275,N_3339);
nor U7444 (N_7444,N_2879,N_4488);
or U7445 (N_7445,N_921,N_1583);
and U7446 (N_7446,N_1559,N_1930);
and U7447 (N_7447,N_2565,N_2174);
and U7448 (N_7448,N_1215,N_2303);
and U7449 (N_7449,N_4684,N_3938);
or U7450 (N_7450,N_1282,N_2442);
and U7451 (N_7451,N_3816,N_3364);
or U7452 (N_7452,N_1279,N_3843);
and U7453 (N_7453,N_2446,N_3846);
or U7454 (N_7454,N_1342,N_2547);
or U7455 (N_7455,N_980,N_2231);
nor U7456 (N_7456,N_1967,N_553);
nor U7457 (N_7457,N_1897,N_2988);
and U7458 (N_7458,N_1964,N_1811);
nor U7459 (N_7459,N_4786,N_4057);
nor U7460 (N_7460,N_1629,N_3165);
nor U7461 (N_7461,N_591,N_115);
and U7462 (N_7462,N_1330,N_1956);
and U7463 (N_7463,N_22,N_2388);
and U7464 (N_7464,N_2672,N_23);
nor U7465 (N_7465,N_118,N_1306);
nor U7466 (N_7466,N_3729,N_181);
and U7467 (N_7467,N_4083,N_3582);
nor U7468 (N_7468,N_1119,N_940);
nand U7469 (N_7469,N_3964,N_336);
nor U7470 (N_7470,N_1042,N_3940);
or U7471 (N_7471,N_1181,N_1885);
nor U7472 (N_7472,N_1889,N_4863);
nand U7473 (N_7473,N_2019,N_3490);
or U7474 (N_7474,N_703,N_1357);
nor U7475 (N_7475,N_4478,N_2664);
and U7476 (N_7476,N_3275,N_3390);
and U7477 (N_7477,N_451,N_2410);
and U7478 (N_7478,N_1753,N_2106);
and U7479 (N_7479,N_4613,N_3476);
or U7480 (N_7480,N_182,N_2591);
or U7481 (N_7481,N_2347,N_3828);
and U7482 (N_7482,N_271,N_2904);
or U7483 (N_7483,N_3980,N_3133);
nor U7484 (N_7484,N_1638,N_1039);
or U7485 (N_7485,N_3205,N_4042);
or U7486 (N_7486,N_4841,N_348);
or U7487 (N_7487,N_1612,N_3362);
and U7488 (N_7488,N_2350,N_2555);
nand U7489 (N_7489,N_1190,N_806);
or U7490 (N_7490,N_2467,N_4609);
and U7491 (N_7491,N_1293,N_1336);
or U7492 (N_7492,N_1668,N_798);
nand U7493 (N_7493,N_2116,N_1464);
nand U7494 (N_7494,N_102,N_402);
nand U7495 (N_7495,N_2330,N_733);
or U7496 (N_7496,N_1291,N_1453);
nor U7497 (N_7497,N_2539,N_92);
and U7498 (N_7498,N_4568,N_898);
nand U7499 (N_7499,N_3041,N_3678);
nor U7500 (N_7500,N_1100,N_4652);
or U7501 (N_7501,N_4008,N_2281);
or U7502 (N_7502,N_4905,N_2093);
and U7503 (N_7503,N_4477,N_4202);
nand U7504 (N_7504,N_962,N_2554);
and U7505 (N_7505,N_2373,N_133);
and U7506 (N_7506,N_271,N_2137);
or U7507 (N_7507,N_2148,N_88);
nand U7508 (N_7508,N_4755,N_1530);
or U7509 (N_7509,N_2110,N_1424);
or U7510 (N_7510,N_4177,N_2766);
and U7511 (N_7511,N_4773,N_2235);
nor U7512 (N_7512,N_663,N_1053);
nor U7513 (N_7513,N_3794,N_2311);
or U7514 (N_7514,N_2341,N_3540);
or U7515 (N_7515,N_77,N_2328);
nand U7516 (N_7516,N_3369,N_3855);
or U7517 (N_7517,N_2575,N_1570);
nor U7518 (N_7518,N_1527,N_1475);
or U7519 (N_7519,N_3896,N_251);
nand U7520 (N_7520,N_781,N_4606);
nand U7521 (N_7521,N_3810,N_3594);
or U7522 (N_7522,N_3296,N_1464);
and U7523 (N_7523,N_766,N_2993);
and U7524 (N_7524,N_1364,N_3688);
and U7525 (N_7525,N_2212,N_1589);
nand U7526 (N_7526,N_574,N_1041);
nand U7527 (N_7527,N_2136,N_305);
or U7528 (N_7528,N_3031,N_1173);
or U7529 (N_7529,N_512,N_4470);
nand U7530 (N_7530,N_2686,N_4375);
nor U7531 (N_7531,N_1433,N_659);
nand U7532 (N_7532,N_3475,N_3331);
or U7533 (N_7533,N_4617,N_4648);
nand U7534 (N_7534,N_393,N_2638);
or U7535 (N_7535,N_4068,N_3790);
or U7536 (N_7536,N_208,N_3052);
or U7537 (N_7537,N_3774,N_4927);
or U7538 (N_7538,N_153,N_2782);
nand U7539 (N_7539,N_1748,N_1011);
nor U7540 (N_7540,N_2323,N_1004);
and U7541 (N_7541,N_100,N_644);
nand U7542 (N_7542,N_1891,N_2720);
nor U7543 (N_7543,N_3158,N_609);
nor U7544 (N_7544,N_1394,N_2776);
and U7545 (N_7545,N_326,N_2904);
xnor U7546 (N_7546,N_1045,N_234);
and U7547 (N_7547,N_4653,N_2404);
nand U7548 (N_7548,N_599,N_3720);
or U7549 (N_7549,N_189,N_3463);
nand U7550 (N_7550,N_4096,N_110);
nand U7551 (N_7551,N_4227,N_12);
nand U7552 (N_7552,N_3374,N_577);
and U7553 (N_7553,N_3265,N_1698);
nor U7554 (N_7554,N_2676,N_589);
and U7555 (N_7555,N_513,N_1605);
and U7556 (N_7556,N_3409,N_1390);
nor U7557 (N_7557,N_2717,N_536);
nand U7558 (N_7558,N_243,N_2184);
or U7559 (N_7559,N_3271,N_3811);
and U7560 (N_7560,N_4117,N_2108);
and U7561 (N_7561,N_4597,N_127);
xnor U7562 (N_7562,N_877,N_4392);
nor U7563 (N_7563,N_745,N_3033);
nand U7564 (N_7564,N_2808,N_3428);
or U7565 (N_7565,N_1185,N_4840);
nor U7566 (N_7566,N_3886,N_1694);
and U7567 (N_7567,N_4234,N_3182);
xor U7568 (N_7568,N_128,N_2677);
and U7569 (N_7569,N_666,N_2366);
and U7570 (N_7570,N_2597,N_351);
and U7571 (N_7571,N_3448,N_2577);
nor U7572 (N_7572,N_486,N_2301);
or U7573 (N_7573,N_1211,N_3016);
nor U7574 (N_7574,N_4199,N_2878);
nor U7575 (N_7575,N_793,N_4454);
and U7576 (N_7576,N_2804,N_1712);
and U7577 (N_7577,N_4023,N_29);
nand U7578 (N_7578,N_4314,N_270);
nand U7579 (N_7579,N_2134,N_2510);
or U7580 (N_7580,N_2895,N_4799);
xnor U7581 (N_7581,N_3291,N_1582);
or U7582 (N_7582,N_267,N_3942);
nor U7583 (N_7583,N_2351,N_2831);
nand U7584 (N_7584,N_3664,N_1360);
nand U7585 (N_7585,N_1551,N_1445);
nor U7586 (N_7586,N_3383,N_1355);
nand U7587 (N_7587,N_2475,N_4734);
nand U7588 (N_7588,N_2565,N_451);
or U7589 (N_7589,N_2988,N_1298);
nand U7590 (N_7590,N_3850,N_1780);
or U7591 (N_7591,N_2705,N_121);
and U7592 (N_7592,N_1294,N_798);
nor U7593 (N_7593,N_4102,N_4403);
nand U7594 (N_7594,N_3625,N_489);
or U7595 (N_7595,N_2311,N_4644);
or U7596 (N_7596,N_2766,N_2439);
or U7597 (N_7597,N_1891,N_3330);
or U7598 (N_7598,N_3647,N_627);
and U7599 (N_7599,N_3255,N_3502);
or U7600 (N_7600,N_1708,N_1402);
or U7601 (N_7601,N_4289,N_3770);
xor U7602 (N_7602,N_2522,N_1742);
xnor U7603 (N_7603,N_4352,N_4697);
and U7604 (N_7604,N_2882,N_1800);
and U7605 (N_7605,N_4291,N_3016);
or U7606 (N_7606,N_775,N_2251);
nand U7607 (N_7607,N_4538,N_284);
or U7608 (N_7608,N_4274,N_1620);
nand U7609 (N_7609,N_828,N_1973);
and U7610 (N_7610,N_1207,N_2053);
and U7611 (N_7611,N_2657,N_3011);
and U7612 (N_7612,N_311,N_2156);
nand U7613 (N_7613,N_2444,N_2962);
nand U7614 (N_7614,N_1929,N_1144);
and U7615 (N_7615,N_4038,N_2661);
nor U7616 (N_7616,N_4846,N_3740);
and U7617 (N_7617,N_4734,N_4133);
nand U7618 (N_7618,N_2801,N_3293);
nand U7619 (N_7619,N_3363,N_520);
and U7620 (N_7620,N_260,N_3191);
or U7621 (N_7621,N_2493,N_2595);
nand U7622 (N_7622,N_2091,N_1403);
or U7623 (N_7623,N_4110,N_3107);
nand U7624 (N_7624,N_2390,N_355);
nand U7625 (N_7625,N_2894,N_3988);
nand U7626 (N_7626,N_95,N_189);
nor U7627 (N_7627,N_2788,N_4395);
nand U7628 (N_7628,N_42,N_455);
nor U7629 (N_7629,N_165,N_2191);
nor U7630 (N_7630,N_2329,N_761);
or U7631 (N_7631,N_2458,N_3328);
and U7632 (N_7632,N_4854,N_377);
nand U7633 (N_7633,N_2757,N_2497);
and U7634 (N_7634,N_3751,N_3797);
or U7635 (N_7635,N_3369,N_134);
and U7636 (N_7636,N_1120,N_3152);
nand U7637 (N_7637,N_865,N_4564);
xor U7638 (N_7638,N_2243,N_1012);
or U7639 (N_7639,N_4578,N_958);
or U7640 (N_7640,N_3397,N_2669);
nand U7641 (N_7641,N_3810,N_2891);
and U7642 (N_7642,N_1415,N_1998);
or U7643 (N_7643,N_4098,N_3396);
nor U7644 (N_7644,N_4106,N_2252);
nor U7645 (N_7645,N_718,N_4409);
and U7646 (N_7646,N_4949,N_329);
and U7647 (N_7647,N_2875,N_4551);
and U7648 (N_7648,N_4087,N_3841);
or U7649 (N_7649,N_1252,N_1570);
and U7650 (N_7650,N_528,N_4750);
nand U7651 (N_7651,N_1070,N_1746);
or U7652 (N_7652,N_1252,N_4084);
xnor U7653 (N_7653,N_1032,N_190);
or U7654 (N_7654,N_2905,N_4055);
or U7655 (N_7655,N_3796,N_1742);
nor U7656 (N_7656,N_2342,N_3973);
or U7657 (N_7657,N_1763,N_4744);
or U7658 (N_7658,N_3517,N_1352);
and U7659 (N_7659,N_2877,N_2964);
nor U7660 (N_7660,N_1955,N_2477);
and U7661 (N_7661,N_263,N_1997);
or U7662 (N_7662,N_725,N_2445);
and U7663 (N_7663,N_2184,N_1327);
nand U7664 (N_7664,N_2515,N_3322);
nor U7665 (N_7665,N_3616,N_1290);
and U7666 (N_7666,N_930,N_2447);
or U7667 (N_7667,N_4967,N_4518);
nor U7668 (N_7668,N_2893,N_1869);
nand U7669 (N_7669,N_3465,N_4448);
or U7670 (N_7670,N_1075,N_4782);
nand U7671 (N_7671,N_2751,N_2624);
or U7672 (N_7672,N_2668,N_1402);
and U7673 (N_7673,N_576,N_2496);
or U7674 (N_7674,N_2658,N_4187);
or U7675 (N_7675,N_4657,N_3825);
or U7676 (N_7676,N_1017,N_970);
and U7677 (N_7677,N_4697,N_3288);
nor U7678 (N_7678,N_1675,N_4483);
xor U7679 (N_7679,N_3684,N_1907);
xor U7680 (N_7680,N_1765,N_4983);
and U7681 (N_7681,N_488,N_4763);
or U7682 (N_7682,N_821,N_2915);
nand U7683 (N_7683,N_1776,N_4581);
nor U7684 (N_7684,N_3503,N_3476);
xor U7685 (N_7685,N_352,N_1896);
nor U7686 (N_7686,N_2356,N_1072);
nand U7687 (N_7687,N_1825,N_1201);
and U7688 (N_7688,N_2841,N_4527);
nand U7689 (N_7689,N_1262,N_1679);
or U7690 (N_7690,N_4799,N_4702);
or U7691 (N_7691,N_1404,N_1255);
nor U7692 (N_7692,N_4312,N_1220);
or U7693 (N_7693,N_1549,N_4961);
or U7694 (N_7694,N_135,N_1231);
nand U7695 (N_7695,N_2364,N_1003);
or U7696 (N_7696,N_4145,N_4783);
nand U7697 (N_7697,N_4987,N_3027);
nand U7698 (N_7698,N_2094,N_681);
nand U7699 (N_7699,N_3413,N_4661);
nand U7700 (N_7700,N_1822,N_1419);
or U7701 (N_7701,N_2508,N_4134);
or U7702 (N_7702,N_2500,N_2728);
nor U7703 (N_7703,N_2354,N_2668);
nor U7704 (N_7704,N_2753,N_3564);
and U7705 (N_7705,N_3522,N_4780);
nor U7706 (N_7706,N_439,N_1263);
nor U7707 (N_7707,N_1605,N_4223);
nor U7708 (N_7708,N_1931,N_1502);
and U7709 (N_7709,N_1001,N_2871);
nor U7710 (N_7710,N_4335,N_4994);
nor U7711 (N_7711,N_1195,N_3218);
or U7712 (N_7712,N_4285,N_2089);
xor U7713 (N_7713,N_4142,N_2442);
or U7714 (N_7714,N_866,N_4755);
or U7715 (N_7715,N_3209,N_3788);
nor U7716 (N_7716,N_2993,N_1741);
nor U7717 (N_7717,N_3715,N_3607);
or U7718 (N_7718,N_1833,N_4638);
and U7719 (N_7719,N_1148,N_1092);
nor U7720 (N_7720,N_4788,N_787);
nand U7721 (N_7721,N_4890,N_3034);
nand U7722 (N_7722,N_4066,N_4031);
nor U7723 (N_7723,N_3413,N_4410);
nor U7724 (N_7724,N_2591,N_2885);
or U7725 (N_7725,N_336,N_4308);
or U7726 (N_7726,N_2174,N_4238);
and U7727 (N_7727,N_190,N_1356);
xnor U7728 (N_7728,N_436,N_1033);
nand U7729 (N_7729,N_4532,N_2091);
nor U7730 (N_7730,N_4204,N_1560);
nand U7731 (N_7731,N_3289,N_4121);
or U7732 (N_7732,N_4277,N_2830);
and U7733 (N_7733,N_4251,N_4195);
nand U7734 (N_7734,N_107,N_2580);
nor U7735 (N_7735,N_1515,N_4783);
nand U7736 (N_7736,N_3197,N_3043);
nand U7737 (N_7737,N_3953,N_4785);
nor U7738 (N_7738,N_3170,N_649);
nand U7739 (N_7739,N_2608,N_4396);
and U7740 (N_7740,N_99,N_4316);
and U7741 (N_7741,N_3088,N_2747);
and U7742 (N_7742,N_2242,N_4011);
nand U7743 (N_7743,N_1077,N_4183);
and U7744 (N_7744,N_3153,N_2615);
nand U7745 (N_7745,N_1914,N_386);
and U7746 (N_7746,N_2587,N_1563);
nor U7747 (N_7747,N_4407,N_3614);
nand U7748 (N_7748,N_3822,N_2433);
nor U7749 (N_7749,N_4777,N_4321);
nand U7750 (N_7750,N_3585,N_1679);
or U7751 (N_7751,N_1478,N_3475);
and U7752 (N_7752,N_3680,N_3235);
or U7753 (N_7753,N_4057,N_4761);
and U7754 (N_7754,N_1460,N_4978);
nand U7755 (N_7755,N_436,N_4449);
nand U7756 (N_7756,N_2522,N_4615);
nor U7757 (N_7757,N_3700,N_1097);
and U7758 (N_7758,N_1282,N_2584);
nand U7759 (N_7759,N_1466,N_4625);
and U7760 (N_7760,N_2654,N_2012);
nand U7761 (N_7761,N_3895,N_3257);
and U7762 (N_7762,N_1533,N_3568);
xnor U7763 (N_7763,N_3434,N_1451);
nor U7764 (N_7764,N_2143,N_1374);
nor U7765 (N_7765,N_800,N_3441);
or U7766 (N_7766,N_862,N_4528);
xor U7767 (N_7767,N_2890,N_1971);
and U7768 (N_7768,N_300,N_2920);
nand U7769 (N_7769,N_4613,N_1356);
and U7770 (N_7770,N_739,N_3168);
or U7771 (N_7771,N_3102,N_4191);
xor U7772 (N_7772,N_985,N_805);
nor U7773 (N_7773,N_1010,N_4163);
and U7774 (N_7774,N_934,N_2538);
xnor U7775 (N_7775,N_1754,N_3137);
nor U7776 (N_7776,N_1922,N_4984);
nand U7777 (N_7777,N_1689,N_89);
nor U7778 (N_7778,N_4797,N_1270);
nand U7779 (N_7779,N_2241,N_3619);
or U7780 (N_7780,N_3753,N_417);
or U7781 (N_7781,N_2267,N_4088);
nor U7782 (N_7782,N_4335,N_3307);
nand U7783 (N_7783,N_607,N_3603);
nand U7784 (N_7784,N_3521,N_2620);
and U7785 (N_7785,N_1914,N_1787);
nand U7786 (N_7786,N_1445,N_1739);
nor U7787 (N_7787,N_2426,N_4507);
or U7788 (N_7788,N_2800,N_78);
and U7789 (N_7789,N_2263,N_2132);
nor U7790 (N_7790,N_552,N_3092);
nand U7791 (N_7791,N_4144,N_2816);
and U7792 (N_7792,N_3508,N_4305);
nand U7793 (N_7793,N_1349,N_2603);
and U7794 (N_7794,N_4022,N_397);
and U7795 (N_7795,N_3697,N_801);
nor U7796 (N_7796,N_4472,N_2826);
and U7797 (N_7797,N_44,N_3253);
nand U7798 (N_7798,N_280,N_2518);
and U7799 (N_7799,N_3847,N_1598);
and U7800 (N_7800,N_1727,N_4617);
nand U7801 (N_7801,N_155,N_161);
and U7802 (N_7802,N_1862,N_2956);
nand U7803 (N_7803,N_4088,N_1321);
and U7804 (N_7804,N_2389,N_1086);
and U7805 (N_7805,N_1078,N_2);
and U7806 (N_7806,N_3553,N_2108);
and U7807 (N_7807,N_4019,N_3741);
or U7808 (N_7808,N_3263,N_1628);
and U7809 (N_7809,N_3067,N_4435);
and U7810 (N_7810,N_4353,N_2025);
nand U7811 (N_7811,N_1882,N_2786);
and U7812 (N_7812,N_886,N_1303);
or U7813 (N_7813,N_3642,N_1878);
and U7814 (N_7814,N_4729,N_1220);
and U7815 (N_7815,N_563,N_1694);
nor U7816 (N_7816,N_4196,N_192);
or U7817 (N_7817,N_3547,N_1568);
or U7818 (N_7818,N_905,N_355);
nand U7819 (N_7819,N_863,N_4144);
or U7820 (N_7820,N_4523,N_4093);
nor U7821 (N_7821,N_4384,N_295);
and U7822 (N_7822,N_4019,N_1441);
nand U7823 (N_7823,N_3883,N_3349);
xor U7824 (N_7824,N_1860,N_921);
or U7825 (N_7825,N_666,N_1267);
and U7826 (N_7826,N_2887,N_523);
and U7827 (N_7827,N_266,N_2063);
nor U7828 (N_7828,N_1163,N_1868);
nand U7829 (N_7829,N_3655,N_2877);
and U7830 (N_7830,N_2191,N_3223);
nand U7831 (N_7831,N_4237,N_64);
nand U7832 (N_7832,N_865,N_2753);
or U7833 (N_7833,N_2602,N_1204);
and U7834 (N_7834,N_3886,N_819);
and U7835 (N_7835,N_3331,N_1223);
nor U7836 (N_7836,N_4618,N_3825);
nand U7837 (N_7837,N_2426,N_2261);
or U7838 (N_7838,N_4819,N_1621);
nand U7839 (N_7839,N_3225,N_989);
nor U7840 (N_7840,N_2996,N_651);
nor U7841 (N_7841,N_656,N_2240);
or U7842 (N_7842,N_4885,N_4446);
nor U7843 (N_7843,N_2698,N_693);
nor U7844 (N_7844,N_1040,N_3221);
nand U7845 (N_7845,N_1674,N_3702);
xnor U7846 (N_7846,N_3390,N_2414);
nor U7847 (N_7847,N_3611,N_4865);
nor U7848 (N_7848,N_2164,N_2188);
nor U7849 (N_7849,N_692,N_3745);
or U7850 (N_7850,N_3248,N_2827);
nor U7851 (N_7851,N_3611,N_878);
nand U7852 (N_7852,N_4074,N_4168);
and U7853 (N_7853,N_582,N_2098);
nor U7854 (N_7854,N_3775,N_3239);
nor U7855 (N_7855,N_2496,N_1404);
and U7856 (N_7856,N_3128,N_4812);
nand U7857 (N_7857,N_1726,N_3269);
nor U7858 (N_7858,N_2379,N_2483);
nor U7859 (N_7859,N_3168,N_1991);
nand U7860 (N_7860,N_4874,N_3090);
nor U7861 (N_7861,N_2230,N_1128);
or U7862 (N_7862,N_437,N_2136);
nand U7863 (N_7863,N_3511,N_4022);
nor U7864 (N_7864,N_808,N_4255);
and U7865 (N_7865,N_3037,N_2367);
or U7866 (N_7866,N_320,N_1934);
or U7867 (N_7867,N_229,N_2832);
or U7868 (N_7868,N_4666,N_153);
and U7869 (N_7869,N_3188,N_4693);
and U7870 (N_7870,N_1141,N_660);
xnor U7871 (N_7871,N_2004,N_1517);
or U7872 (N_7872,N_1280,N_820);
or U7873 (N_7873,N_4567,N_109);
and U7874 (N_7874,N_4350,N_104);
or U7875 (N_7875,N_914,N_2520);
nand U7876 (N_7876,N_4509,N_2230);
or U7877 (N_7877,N_4809,N_283);
nor U7878 (N_7878,N_4293,N_1055);
or U7879 (N_7879,N_1016,N_189);
nor U7880 (N_7880,N_648,N_4214);
and U7881 (N_7881,N_351,N_1354);
xnor U7882 (N_7882,N_3088,N_1206);
nand U7883 (N_7883,N_326,N_834);
nor U7884 (N_7884,N_491,N_2308);
nor U7885 (N_7885,N_963,N_2112);
or U7886 (N_7886,N_3729,N_839);
and U7887 (N_7887,N_2290,N_3028);
nand U7888 (N_7888,N_4229,N_2208);
nor U7889 (N_7889,N_3398,N_4436);
or U7890 (N_7890,N_4914,N_1642);
nand U7891 (N_7891,N_4082,N_4586);
or U7892 (N_7892,N_2206,N_4034);
nor U7893 (N_7893,N_3671,N_3543);
or U7894 (N_7894,N_2129,N_3000);
nand U7895 (N_7895,N_1068,N_4086);
or U7896 (N_7896,N_3022,N_1597);
or U7897 (N_7897,N_4047,N_53);
nor U7898 (N_7898,N_1270,N_775);
nand U7899 (N_7899,N_1188,N_142);
nand U7900 (N_7900,N_2558,N_2108);
and U7901 (N_7901,N_2920,N_1328);
and U7902 (N_7902,N_1864,N_1415);
and U7903 (N_7903,N_1278,N_1865);
and U7904 (N_7904,N_615,N_2358);
nand U7905 (N_7905,N_2179,N_1384);
and U7906 (N_7906,N_3787,N_787);
nor U7907 (N_7907,N_2860,N_1745);
or U7908 (N_7908,N_3940,N_4605);
and U7909 (N_7909,N_1885,N_1841);
nand U7910 (N_7910,N_3624,N_2936);
nor U7911 (N_7911,N_4539,N_747);
or U7912 (N_7912,N_3618,N_988);
and U7913 (N_7913,N_2816,N_1599);
nor U7914 (N_7914,N_947,N_4909);
nand U7915 (N_7915,N_4152,N_2125);
xnor U7916 (N_7916,N_2645,N_1846);
nand U7917 (N_7917,N_364,N_4058);
nand U7918 (N_7918,N_791,N_2699);
nand U7919 (N_7919,N_3853,N_735);
nor U7920 (N_7920,N_4522,N_1357);
or U7921 (N_7921,N_2450,N_893);
nor U7922 (N_7922,N_363,N_3420);
nor U7923 (N_7923,N_2877,N_16);
nor U7924 (N_7924,N_571,N_3085);
or U7925 (N_7925,N_4215,N_2672);
xnor U7926 (N_7926,N_2205,N_3462);
nand U7927 (N_7927,N_1545,N_853);
nand U7928 (N_7928,N_4793,N_2470);
nand U7929 (N_7929,N_4117,N_3867);
and U7930 (N_7930,N_4746,N_1062);
nor U7931 (N_7931,N_1089,N_3848);
or U7932 (N_7932,N_232,N_4282);
nor U7933 (N_7933,N_2724,N_4615);
or U7934 (N_7934,N_2853,N_118);
and U7935 (N_7935,N_2996,N_54);
and U7936 (N_7936,N_4135,N_3752);
nand U7937 (N_7937,N_903,N_4086);
or U7938 (N_7938,N_3498,N_860);
nand U7939 (N_7939,N_33,N_3344);
and U7940 (N_7940,N_4571,N_2616);
nor U7941 (N_7941,N_699,N_2542);
or U7942 (N_7942,N_2085,N_1466);
xnor U7943 (N_7943,N_4264,N_3058);
nor U7944 (N_7944,N_2832,N_2731);
and U7945 (N_7945,N_4174,N_4479);
nor U7946 (N_7946,N_3724,N_7);
or U7947 (N_7947,N_704,N_11);
and U7948 (N_7948,N_2971,N_4544);
nor U7949 (N_7949,N_954,N_1635);
nor U7950 (N_7950,N_763,N_1188);
xnor U7951 (N_7951,N_3401,N_2361);
or U7952 (N_7952,N_2617,N_1255);
nor U7953 (N_7953,N_291,N_4196);
and U7954 (N_7954,N_420,N_1619);
and U7955 (N_7955,N_3758,N_1069);
nor U7956 (N_7956,N_1969,N_41);
xor U7957 (N_7957,N_4537,N_1654);
and U7958 (N_7958,N_3271,N_798);
and U7959 (N_7959,N_174,N_3346);
nand U7960 (N_7960,N_3800,N_2306);
and U7961 (N_7961,N_553,N_3280);
nand U7962 (N_7962,N_3436,N_3841);
or U7963 (N_7963,N_3377,N_3613);
nand U7964 (N_7964,N_4797,N_2418);
nor U7965 (N_7965,N_3558,N_1669);
and U7966 (N_7966,N_701,N_2254);
nor U7967 (N_7967,N_10,N_1345);
or U7968 (N_7968,N_2623,N_354);
and U7969 (N_7969,N_3141,N_4900);
nand U7970 (N_7970,N_4974,N_1886);
nand U7971 (N_7971,N_61,N_4438);
nand U7972 (N_7972,N_4440,N_2376);
nor U7973 (N_7973,N_1292,N_3204);
nand U7974 (N_7974,N_4487,N_441);
nor U7975 (N_7975,N_259,N_3928);
nand U7976 (N_7976,N_693,N_894);
and U7977 (N_7977,N_954,N_2369);
nor U7978 (N_7978,N_1316,N_3752);
nor U7979 (N_7979,N_721,N_3351);
or U7980 (N_7980,N_4104,N_2693);
or U7981 (N_7981,N_2824,N_3125);
nor U7982 (N_7982,N_4829,N_4855);
xnor U7983 (N_7983,N_647,N_1087);
and U7984 (N_7984,N_4605,N_1185);
nor U7985 (N_7985,N_279,N_2770);
or U7986 (N_7986,N_3049,N_269);
nor U7987 (N_7987,N_4024,N_4403);
or U7988 (N_7988,N_2689,N_1366);
nand U7989 (N_7989,N_3977,N_3154);
nor U7990 (N_7990,N_127,N_145);
or U7991 (N_7991,N_3942,N_16);
or U7992 (N_7992,N_1669,N_1524);
or U7993 (N_7993,N_1700,N_1914);
nand U7994 (N_7994,N_1572,N_2546);
nand U7995 (N_7995,N_3429,N_780);
or U7996 (N_7996,N_3779,N_3077);
nor U7997 (N_7997,N_3360,N_4023);
and U7998 (N_7998,N_3317,N_4701);
nand U7999 (N_7999,N_235,N_1946);
nand U8000 (N_8000,N_4627,N_1077);
and U8001 (N_8001,N_679,N_2479);
nor U8002 (N_8002,N_4850,N_814);
nor U8003 (N_8003,N_167,N_4753);
or U8004 (N_8004,N_1471,N_3760);
nand U8005 (N_8005,N_1996,N_4903);
nor U8006 (N_8006,N_2124,N_3106);
or U8007 (N_8007,N_2211,N_2878);
xnor U8008 (N_8008,N_4762,N_4999);
and U8009 (N_8009,N_796,N_4644);
xnor U8010 (N_8010,N_3158,N_523);
xnor U8011 (N_8011,N_2812,N_1765);
nor U8012 (N_8012,N_2304,N_3166);
nor U8013 (N_8013,N_960,N_2239);
or U8014 (N_8014,N_4687,N_4801);
nor U8015 (N_8015,N_4778,N_2778);
or U8016 (N_8016,N_2616,N_231);
nand U8017 (N_8017,N_595,N_4923);
and U8018 (N_8018,N_4488,N_2667);
nand U8019 (N_8019,N_3955,N_2539);
or U8020 (N_8020,N_3799,N_4028);
and U8021 (N_8021,N_3266,N_1781);
or U8022 (N_8022,N_4764,N_4156);
and U8023 (N_8023,N_2630,N_3218);
or U8024 (N_8024,N_2179,N_277);
nor U8025 (N_8025,N_3641,N_878);
nand U8026 (N_8026,N_119,N_3702);
nand U8027 (N_8027,N_3046,N_2695);
and U8028 (N_8028,N_4287,N_4334);
or U8029 (N_8029,N_1667,N_1673);
and U8030 (N_8030,N_15,N_1059);
or U8031 (N_8031,N_2973,N_2992);
nand U8032 (N_8032,N_130,N_4408);
nor U8033 (N_8033,N_1350,N_885);
nor U8034 (N_8034,N_142,N_3526);
or U8035 (N_8035,N_1659,N_1760);
and U8036 (N_8036,N_309,N_2066);
nand U8037 (N_8037,N_711,N_974);
nand U8038 (N_8038,N_2444,N_4486);
and U8039 (N_8039,N_1604,N_3804);
nand U8040 (N_8040,N_4523,N_3081);
or U8041 (N_8041,N_1934,N_1456);
xor U8042 (N_8042,N_1145,N_4232);
nor U8043 (N_8043,N_1267,N_4069);
and U8044 (N_8044,N_1807,N_3626);
xor U8045 (N_8045,N_2270,N_3027);
nor U8046 (N_8046,N_787,N_2569);
and U8047 (N_8047,N_466,N_4104);
nor U8048 (N_8048,N_1386,N_2067);
or U8049 (N_8049,N_324,N_2842);
or U8050 (N_8050,N_1958,N_554);
and U8051 (N_8051,N_46,N_2810);
or U8052 (N_8052,N_1991,N_533);
and U8053 (N_8053,N_1957,N_4686);
nor U8054 (N_8054,N_2388,N_569);
nor U8055 (N_8055,N_3646,N_1515);
and U8056 (N_8056,N_2925,N_3725);
nand U8057 (N_8057,N_4492,N_3533);
or U8058 (N_8058,N_4392,N_4294);
and U8059 (N_8059,N_4148,N_2632);
and U8060 (N_8060,N_4077,N_204);
nand U8061 (N_8061,N_2535,N_4379);
nor U8062 (N_8062,N_4227,N_1881);
nor U8063 (N_8063,N_2273,N_1351);
nor U8064 (N_8064,N_1162,N_16);
nand U8065 (N_8065,N_4240,N_4957);
nand U8066 (N_8066,N_2191,N_2867);
nand U8067 (N_8067,N_4554,N_3511);
and U8068 (N_8068,N_2695,N_273);
and U8069 (N_8069,N_3520,N_1039);
or U8070 (N_8070,N_560,N_3193);
and U8071 (N_8071,N_2757,N_2054);
and U8072 (N_8072,N_2305,N_4630);
or U8073 (N_8073,N_6,N_2356);
xnor U8074 (N_8074,N_1597,N_593);
xor U8075 (N_8075,N_1646,N_1252);
nor U8076 (N_8076,N_4335,N_4468);
nor U8077 (N_8077,N_4105,N_163);
and U8078 (N_8078,N_4802,N_4606);
and U8079 (N_8079,N_447,N_2224);
or U8080 (N_8080,N_2431,N_2114);
or U8081 (N_8081,N_2124,N_4010);
nand U8082 (N_8082,N_4590,N_3670);
nor U8083 (N_8083,N_3769,N_91);
nor U8084 (N_8084,N_1865,N_3284);
or U8085 (N_8085,N_1128,N_2185);
nor U8086 (N_8086,N_4021,N_2842);
or U8087 (N_8087,N_2052,N_4992);
nand U8088 (N_8088,N_1219,N_2409);
and U8089 (N_8089,N_1607,N_4816);
and U8090 (N_8090,N_3364,N_2788);
nor U8091 (N_8091,N_3272,N_1454);
or U8092 (N_8092,N_4044,N_4034);
and U8093 (N_8093,N_4129,N_3572);
and U8094 (N_8094,N_2429,N_1678);
nand U8095 (N_8095,N_1507,N_2931);
nand U8096 (N_8096,N_3419,N_1145);
xor U8097 (N_8097,N_4323,N_688);
nor U8098 (N_8098,N_2610,N_4187);
and U8099 (N_8099,N_3657,N_3679);
or U8100 (N_8100,N_1236,N_2896);
nor U8101 (N_8101,N_1377,N_1785);
nand U8102 (N_8102,N_950,N_1344);
or U8103 (N_8103,N_533,N_2628);
nor U8104 (N_8104,N_669,N_2722);
nand U8105 (N_8105,N_4661,N_472);
and U8106 (N_8106,N_859,N_3052);
nand U8107 (N_8107,N_2349,N_3337);
nor U8108 (N_8108,N_4392,N_3370);
nand U8109 (N_8109,N_2404,N_2658);
nor U8110 (N_8110,N_1647,N_2);
or U8111 (N_8111,N_1438,N_2276);
nor U8112 (N_8112,N_317,N_1241);
and U8113 (N_8113,N_2303,N_4925);
or U8114 (N_8114,N_3762,N_4557);
nand U8115 (N_8115,N_3872,N_1381);
nor U8116 (N_8116,N_2449,N_3541);
and U8117 (N_8117,N_3626,N_4869);
or U8118 (N_8118,N_4747,N_3544);
and U8119 (N_8119,N_2082,N_1696);
or U8120 (N_8120,N_4212,N_3067);
nand U8121 (N_8121,N_13,N_1586);
and U8122 (N_8122,N_4252,N_251);
nor U8123 (N_8123,N_2793,N_1447);
or U8124 (N_8124,N_1289,N_1593);
xnor U8125 (N_8125,N_460,N_1270);
and U8126 (N_8126,N_133,N_1048);
and U8127 (N_8127,N_108,N_3327);
nand U8128 (N_8128,N_1403,N_1846);
or U8129 (N_8129,N_2692,N_1799);
nand U8130 (N_8130,N_3477,N_2801);
nor U8131 (N_8131,N_926,N_89);
and U8132 (N_8132,N_2017,N_1222);
or U8133 (N_8133,N_2210,N_4238);
nand U8134 (N_8134,N_197,N_3287);
xor U8135 (N_8135,N_1814,N_4104);
or U8136 (N_8136,N_1654,N_820);
nor U8137 (N_8137,N_4579,N_1887);
nor U8138 (N_8138,N_1280,N_3752);
or U8139 (N_8139,N_3040,N_1637);
or U8140 (N_8140,N_1575,N_4774);
xor U8141 (N_8141,N_1887,N_4530);
and U8142 (N_8142,N_2547,N_4348);
and U8143 (N_8143,N_699,N_643);
and U8144 (N_8144,N_3706,N_4790);
and U8145 (N_8145,N_2785,N_4018);
nor U8146 (N_8146,N_260,N_3611);
nor U8147 (N_8147,N_4426,N_60);
nor U8148 (N_8148,N_4806,N_2672);
and U8149 (N_8149,N_1430,N_918);
and U8150 (N_8150,N_4676,N_1740);
xor U8151 (N_8151,N_3120,N_1240);
nor U8152 (N_8152,N_2261,N_3296);
and U8153 (N_8153,N_959,N_4986);
nand U8154 (N_8154,N_4371,N_3847);
or U8155 (N_8155,N_1332,N_437);
or U8156 (N_8156,N_138,N_3843);
nand U8157 (N_8157,N_4615,N_1969);
nor U8158 (N_8158,N_78,N_1019);
or U8159 (N_8159,N_4308,N_357);
nand U8160 (N_8160,N_2826,N_3950);
and U8161 (N_8161,N_2965,N_624);
xor U8162 (N_8162,N_0,N_3884);
and U8163 (N_8163,N_106,N_691);
or U8164 (N_8164,N_2768,N_4655);
and U8165 (N_8165,N_3418,N_3493);
nand U8166 (N_8166,N_2736,N_315);
or U8167 (N_8167,N_4540,N_1066);
or U8168 (N_8168,N_1016,N_2642);
and U8169 (N_8169,N_1049,N_3357);
or U8170 (N_8170,N_3161,N_4980);
xor U8171 (N_8171,N_203,N_2328);
nand U8172 (N_8172,N_531,N_1443);
and U8173 (N_8173,N_196,N_1480);
and U8174 (N_8174,N_2655,N_767);
or U8175 (N_8175,N_4556,N_4073);
nand U8176 (N_8176,N_0,N_3400);
nor U8177 (N_8177,N_1376,N_3748);
nand U8178 (N_8178,N_2460,N_2559);
and U8179 (N_8179,N_1802,N_4326);
nand U8180 (N_8180,N_1272,N_2683);
nand U8181 (N_8181,N_3835,N_3739);
or U8182 (N_8182,N_1712,N_2839);
or U8183 (N_8183,N_3298,N_3460);
nor U8184 (N_8184,N_3989,N_2884);
and U8185 (N_8185,N_4572,N_3974);
nor U8186 (N_8186,N_342,N_415);
nor U8187 (N_8187,N_244,N_87);
and U8188 (N_8188,N_352,N_3031);
nand U8189 (N_8189,N_4129,N_3021);
and U8190 (N_8190,N_4651,N_844);
nand U8191 (N_8191,N_2114,N_64);
nand U8192 (N_8192,N_1144,N_3816);
and U8193 (N_8193,N_79,N_23);
and U8194 (N_8194,N_4157,N_2589);
or U8195 (N_8195,N_1379,N_1216);
or U8196 (N_8196,N_2243,N_2915);
or U8197 (N_8197,N_725,N_692);
or U8198 (N_8198,N_2362,N_793);
or U8199 (N_8199,N_3748,N_2082);
nand U8200 (N_8200,N_3566,N_498);
and U8201 (N_8201,N_2226,N_2316);
nor U8202 (N_8202,N_63,N_405);
nand U8203 (N_8203,N_2353,N_3523);
nand U8204 (N_8204,N_1329,N_2576);
nor U8205 (N_8205,N_4098,N_2640);
nor U8206 (N_8206,N_483,N_3158);
or U8207 (N_8207,N_2812,N_839);
and U8208 (N_8208,N_1583,N_2645);
and U8209 (N_8209,N_933,N_3908);
nor U8210 (N_8210,N_1515,N_3000);
nor U8211 (N_8211,N_1806,N_3902);
nor U8212 (N_8212,N_3745,N_3574);
nand U8213 (N_8213,N_4115,N_3849);
nor U8214 (N_8214,N_4766,N_952);
and U8215 (N_8215,N_4377,N_732);
and U8216 (N_8216,N_4931,N_3480);
nand U8217 (N_8217,N_4199,N_3744);
nand U8218 (N_8218,N_3921,N_2821);
and U8219 (N_8219,N_869,N_3936);
nand U8220 (N_8220,N_4087,N_2472);
nand U8221 (N_8221,N_1639,N_867);
and U8222 (N_8222,N_2345,N_1831);
and U8223 (N_8223,N_4701,N_4857);
nor U8224 (N_8224,N_309,N_4413);
nand U8225 (N_8225,N_3194,N_4951);
nor U8226 (N_8226,N_174,N_3629);
or U8227 (N_8227,N_858,N_142);
xor U8228 (N_8228,N_602,N_4024);
and U8229 (N_8229,N_3320,N_418);
nand U8230 (N_8230,N_775,N_1680);
or U8231 (N_8231,N_2639,N_948);
and U8232 (N_8232,N_3839,N_2252);
nor U8233 (N_8233,N_2810,N_3984);
or U8234 (N_8234,N_4003,N_4948);
nand U8235 (N_8235,N_94,N_4011);
nand U8236 (N_8236,N_1616,N_4895);
and U8237 (N_8237,N_147,N_1983);
nor U8238 (N_8238,N_4145,N_3836);
nor U8239 (N_8239,N_836,N_2342);
or U8240 (N_8240,N_4253,N_2464);
nor U8241 (N_8241,N_1407,N_2369);
nor U8242 (N_8242,N_705,N_4838);
or U8243 (N_8243,N_793,N_1985);
nor U8244 (N_8244,N_1098,N_4826);
and U8245 (N_8245,N_4802,N_1835);
and U8246 (N_8246,N_3276,N_1235);
or U8247 (N_8247,N_1207,N_1641);
or U8248 (N_8248,N_4652,N_371);
nor U8249 (N_8249,N_4918,N_1838);
nor U8250 (N_8250,N_173,N_231);
and U8251 (N_8251,N_3721,N_2535);
nand U8252 (N_8252,N_4983,N_135);
or U8253 (N_8253,N_290,N_3416);
and U8254 (N_8254,N_3738,N_3984);
and U8255 (N_8255,N_1427,N_2403);
and U8256 (N_8256,N_1621,N_2462);
or U8257 (N_8257,N_2571,N_4339);
nand U8258 (N_8258,N_1997,N_1565);
and U8259 (N_8259,N_4688,N_4739);
xnor U8260 (N_8260,N_1282,N_4527);
nand U8261 (N_8261,N_3451,N_1689);
nand U8262 (N_8262,N_2747,N_4781);
or U8263 (N_8263,N_4377,N_1681);
nand U8264 (N_8264,N_3913,N_3365);
nand U8265 (N_8265,N_2798,N_316);
and U8266 (N_8266,N_3221,N_3674);
nor U8267 (N_8267,N_4006,N_726);
nor U8268 (N_8268,N_4497,N_2990);
or U8269 (N_8269,N_472,N_3560);
and U8270 (N_8270,N_4014,N_637);
and U8271 (N_8271,N_3868,N_4391);
nor U8272 (N_8272,N_32,N_2499);
nand U8273 (N_8273,N_196,N_1275);
xnor U8274 (N_8274,N_1851,N_556);
and U8275 (N_8275,N_1986,N_4499);
nor U8276 (N_8276,N_4023,N_4813);
nor U8277 (N_8277,N_3511,N_2660);
nand U8278 (N_8278,N_2023,N_1078);
nand U8279 (N_8279,N_1733,N_3090);
nor U8280 (N_8280,N_3562,N_818);
or U8281 (N_8281,N_4997,N_3667);
nor U8282 (N_8282,N_3519,N_4822);
nand U8283 (N_8283,N_270,N_1731);
and U8284 (N_8284,N_265,N_1588);
and U8285 (N_8285,N_1149,N_2776);
nand U8286 (N_8286,N_3271,N_474);
or U8287 (N_8287,N_1648,N_1890);
nand U8288 (N_8288,N_2185,N_213);
nor U8289 (N_8289,N_3185,N_4250);
and U8290 (N_8290,N_2547,N_462);
or U8291 (N_8291,N_4952,N_4027);
nor U8292 (N_8292,N_4829,N_2389);
and U8293 (N_8293,N_2449,N_2228);
nor U8294 (N_8294,N_4153,N_192);
nor U8295 (N_8295,N_3977,N_190);
nor U8296 (N_8296,N_3196,N_3089);
or U8297 (N_8297,N_863,N_3375);
and U8298 (N_8298,N_2149,N_512);
or U8299 (N_8299,N_1613,N_2750);
nor U8300 (N_8300,N_2042,N_2511);
nand U8301 (N_8301,N_4872,N_4955);
or U8302 (N_8302,N_3073,N_4707);
and U8303 (N_8303,N_4392,N_4120);
and U8304 (N_8304,N_3036,N_4164);
nand U8305 (N_8305,N_2816,N_3240);
and U8306 (N_8306,N_312,N_2693);
nor U8307 (N_8307,N_4624,N_4722);
nor U8308 (N_8308,N_911,N_1284);
nand U8309 (N_8309,N_639,N_3482);
or U8310 (N_8310,N_3711,N_1920);
or U8311 (N_8311,N_1214,N_2464);
or U8312 (N_8312,N_439,N_2817);
and U8313 (N_8313,N_3063,N_1215);
or U8314 (N_8314,N_1151,N_155);
nor U8315 (N_8315,N_3438,N_3854);
nor U8316 (N_8316,N_4632,N_2686);
and U8317 (N_8317,N_4261,N_2733);
nand U8318 (N_8318,N_4357,N_2170);
or U8319 (N_8319,N_3150,N_255);
nor U8320 (N_8320,N_1023,N_1135);
nand U8321 (N_8321,N_2538,N_597);
and U8322 (N_8322,N_2638,N_4328);
nand U8323 (N_8323,N_4827,N_2132);
and U8324 (N_8324,N_1652,N_2817);
and U8325 (N_8325,N_879,N_3835);
nand U8326 (N_8326,N_1129,N_2155);
and U8327 (N_8327,N_956,N_2668);
or U8328 (N_8328,N_4727,N_3862);
nor U8329 (N_8329,N_2188,N_4661);
and U8330 (N_8330,N_4744,N_82);
and U8331 (N_8331,N_4591,N_48);
nor U8332 (N_8332,N_562,N_2891);
and U8333 (N_8333,N_3530,N_3657);
nor U8334 (N_8334,N_2233,N_256);
nor U8335 (N_8335,N_2777,N_3709);
and U8336 (N_8336,N_2558,N_3361);
or U8337 (N_8337,N_3532,N_1119);
or U8338 (N_8338,N_4620,N_4158);
nor U8339 (N_8339,N_3541,N_4565);
nand U8340 (N_8340,N_4300,N_3387);
and U8341 (N_8341,N_4461,N_97);
and U8342 (N_8342,N_889,N_3766);
and U8343 (N_8343,N_4247,N_3573);
or U8344 (N_8344,N_281,N_3501);
and U8345 (N_8345,N_4088,N_389);
or U8346 (N_8346,N_189,N_4060);
xnor U8347 (N_8347,N_4560,N_2428);
nor U8348 (N_8348,N_3217,N_2802);
or U8349 (N_8349,N_4209,N_992);
and U8350 (N_8350,N_1798,N_487);
nor U8351 (N_8351,N_2953,N_4461);
nand U8352 (N_8352,N_3330,N_4325);
or U8353 (N_8353,N_1055,N_1936);
nor U8354 (N_8354,N_1830,N_2723);
xnor U8355 (N_8355,N_3034,N_4593);
and U8356 (N_8356,N_1199,N_414);
or U8357 (N_8357,N_148,N_3228);
and U8358 (N_8358,N_1861,N_723);
and U8359 (N_8359,N_2200,N_1815);
nand U8360 (N_8360,N_2679,N_3610);
and U8361 (N_8361,N_4245,N_3394);
nor U8362 (N_8362,N_4135,N_1430);
nor U8363 (N_8363,N_2403,N_1305);
and U8364 (N_8364,N_1827,N_4621);
nand U8365 (N_8365,N_337,N_2569);
or U8366 (N_8366,N_4163,N_626);
nand U8367 (N_8367,N_84,N_1770);
nand U8368 (N_8368,N_1199,N_3151);
nand U8369 (N_8369,N_2865,N_1989);
nand U8370 (N_8370,N_2649,N_100);
nand U8371 (N_8371,N_2406,N_3085);
or U8372 (N_8372,N_2724,N_3813);
or U8373 (N_8373,N_1519,N_546);
nand U8374 (N_8374,N_448,N_604);
and U8375 (N_8375,N_464,N_4192);
and U8376 (N_8376,N_3952,N_910);
and U8377 (N_8377,N_887,N_2363);
nor U8378 (N_8378,N_488,N_2114);
and U8379 (N_8379,N_3192,N_562);
nor U8380 (N_8380,N_4120,N_3671);
and U8381 (N_8381,N_3157,N_3712);
nand U8382 (N_8382,N_300,N_2089);
or U8383 (N_8383,N_838,N_3417);
and U8384 (N_8384,N_3703,N_1219);
or U8385 (N_8385,N_752,N_2675);
nor U8386 (N_8386,N_1534,N_130);
nand U8387 (N_8387,N_2155,N_2306);
and U8388 (N_8388,N_4112,N_1935);
and U8389 (N_8389,N_2540,N_4240);
nand U8390 (N_8390,N_2165,N_802);
nor U8391 (N_8391,N_169,N_4211);
nand U8392 (N_8392,N_1452,N_3582);
nor U8393 (N_8393,N_4178,N_965);
and U8394 (N_8394,N_670,N_1504);
or U8395 (N_8395,N_2707,N_837);
and U8396 (N_8396,N_2871,N_3764);
nand U8397 (N_8397,N_124,N_1422);
or U8398 (N_8398,N_2464,N_3027);
or U8399 (N_8399,N_1755,N_860);
nand U8400 (N_8400,N_2367,N_3708);
nor U8401 (N_8401,N_1792,N_475);
or U8402 (N_8402,N_3532,N_2355);
nor U8403 (N_8403,N_2532,N_2649);
or U8404 (N_8404,N_4448,N_1927);
and U8405 (N_8405,N_2690,N_643);
and U8406 (N_8406,N_4460,N_1433);
nand U8407 (N_8407,N_3060,N_3507);
and U8408 (N_8408,N_2973,N_2226);
and U8409 (N_8409,N_526,N_145);
and U8410 (N_8410,N_3035,N_3327);
nor U8411 (N_8411,N_3990,N_3656);
and U8412 (N_8412,N_4433,N_458);
nand U8413 (N_8413,N_1759,N_1041);
or U8414 (N_8414,N_4685,N_3400);
nor U8415 (N_8415,N_4237,N_183);
and U8416 (N_8416,N_1097,N_4371);
or U8417 (N_8417,N_2845,N_4241);
nor U8418 (N_8418,N_2124,N_1321);
nor U8419 (N_8419,N_631,N_4304);
and U8420 (N_8420,N_1636,N_3592);
or U8421 (N_8421,N_3293,N_1158);
nor U8422 (N_8422,N_1820,N_3411);
nor U8423 (N_8423,N_940,N_3131);
and U8424 (N_8424,N_2976,N_533);
nor U8425 (N_8425,N_3806,N_1008);
and U8426 (N_8426,N_3820,N_2534);
or U8427 (N_8427,N_2923,N_1397);
and U8428 (N_8428,N_2026,N_4680);
nor U8429 (N_8429,N_3199,N_3685);
or U8430 (N_8430,N_3657,N_91);
nand U8431 (N_8431,N_2257,N_2704);
nand U8432 (N_8432,N_2263,N_1719);
or U8433 (N_8433,N_4171,N_1799);
nor U8434 (N_8434,N_1553,N_4122);
xnor U8435 (N_8435,N_408,N_4400);
nand U8436 (N_8436,N_4868,N_917);
or U8437 (N_8437,N_2960,N_977);
nand U8438 (N_8438,N_4482,N_4902);
nand U8439 (N_8439,N_4127,N_4620);
and U8440 (N_8440,N_3073,N_1546);
and U8441 (N_8441,N_1924,N_3780);
nand U8442 (N_8442,N_4296,N_2516);
or U8443 (N_8443,N_620,N_1358);
nand U8444 (N_8444,N_1299,N_2645);
or U8445 (N_8445,N_19,N_3774);
or U8446 (N_8446,N_1579,N_3102);
or U8447 (N_8447,N_4231,N_2792);
or U8448 (N_8448,N_3794,N_2301);
nand U8449 (N_8449,N_612,N_997);
and U8450 (N_8450,N_1464,N_2988);
nand U8451 (N_8451,N_4037,N_2714);
and U8452 (N_8452,N_2504,N_4355);
or U8453 (N_8453,N_3545,N_2832);
nand U8454 (N_8454,N_672,N_1275);
or U8455 (N_8455,N_3476,N_1857);
nand U8456 (N_8456,N_1762,N_2642);
and U8457 (N_8457,N_4767,N_4964);
nor U8458 (N_8458,N_975,N_4017);
and U8459 (N_8459,N_3387,N_4009);
or U8460 (N_8460,N_382,N_2218);
nor U8461 (N_8461,N_4846,N_1525);
or U8462 (N_8462,N_2554,N_4601);
nand U8463 (N_8463,N_3964,N_303);
nand U8464 (N_8464,N_2022,N_985);
nor U8465 (N_8465,N_3494,N_4275);
nand U8466 (N_8466,N_3897,N_4214);
nand U8467 (N_8467,N_3724,N_2813);
and U8468 (N_8468,N_2978,N_1305);
and U8469 (N_8469,N_4476,N_4480);
and U8470 (N_8470,N_1343,N_3135);
nand U8471 (N_8471,N_5,N_1231);
and U8472 (N_8472,N_2796,N_442);
and U8473 (N_8473,N_2482,N_995);
or U8474 (N_8474,N_4187,N_2229);
nand U8475 (N_8475,N_1633,N_1929);
nand U8476 (N_8476,N_3343,N_4426);
nor U8477 (N_8477,N_812,N_1331);
or U8478 (N_8478,N_4992,N_4443);
or U8479 (N_8479,N_2449,N_3406);
nand U8480 (N_8480,N_766,N_4394);
nand U8481 (N_8481,N_2072,N_1592);
and U8482 (N_8482,N_3159,N_2481);
and U8483 (N_8483,N_4990,N_1294);
or U8484 (N_8484,N_54,N_2951);
and U8485 (N_8485,N_531,N_4126);
or U8486 (N_8486,N_3107,N_1260);
xnor U8487 (N_8487,N_4192,N_3394);
nand U8488 (N_8488,N_1586,N_4024);
or U8489 (N_8489,N_3986,N_1631);
nand U8490 (N_8490,N_1572,N_2740);
nand U8491 (N_8491,N_399,N_515);
and U8492 (N_8492,N_1060,N_2741);
nor U8493 (N_8493,N_3607,N_55);
and U8494 (N_8494,N_632,N_3355);
or U8495 (N_8495,N_1313,N_658);
nor U8496 (N_8496,N_4333,N_1212);
nand U8497 (N_8497,N_681,N_460);
nor U8498 (N_8498,N_2160,N_394);
nand U8499 (N_8499,N_4807,N_3031);
or U8500 (N_8500,N_1198,N_4291);
or U8501 (N_8501,N_1930,N_839);
and U8502 (N_8502,N_752,N_3646);
and U8503 (N_8503,N_3900,N_3024);
or U8504 (N_8504,N_4970,N_2905);
nand U8505 (N_8505,N_3358,N_4178);
and U8506 (N_8506,N_1117,N_594);
and U8507 (N_8507,N_4611,N_2591);
and U8508 (N_8508,N_2082,N_1864);
and U8509 (N_8509,N_2992,N_911);
nor U8510 (N_8510,N_1967,N_1130);
nand U8511 (N_8511,N_773,N_4247);
and U8512 (N_8512,N_3695,N_941);
nor U8513 (N_8513,N_4430,N_4322);
nor U8514 (N_8514,N_175,N_2182);
nand U8515 (N_8515,N_1455,N_826);
or U8516 (N_8516,N_4177,N_3489);
nor U8517 (N_8517,N_1328,N_1857);
nor U8518 (N_8518,N_252,N_4698);
and U8519 (N_8519,N_4981,N_1919);
nand U8520 (N_8520,N_2751,N_1948);
nor U8521 (N_8521,N_594,N_1187);
nor U8522 (N_8522,N_1760,N_2549);
nand U8523 (N_8523,N_2472,N_1999);
or U8524 (N_8524,N_1149,N_3734);
nand U8525 (N_8525,N_1471,N_2176);
nor U8526 (N_8526,N_3722,N_603);
and U8527 (N_8527,N_3045,N_1267);
nand U8528 (N_8528,N_1,N_4882);
or U8529 (N_8529,N_275,N_3279);
nand U8530 (N_8530,N_474,N_4429);
or U8531 (N_8531,N_2282,N_4547);
nand U8532 (N_8532,N_1738,N_2097);
nor U8533 (N_8533,N_4858,N_4641);
nor U8534 (N_8534,N_3976,N_2093);
nand U8535 (N_8535,N_4921,N_2273);
nor U8536 (N_8536,N_3063,N_1208);
and U8537 (N_8537,N_2387,N_2016);
nand U8538 (N_8538,N_2527,N_2419);
nand U8539 (N_8539,N_2535,N_697);
nor U8540 (N_8540,N_2610,N_3222);
or U8541 (N_8541,N_1187,N_343);
and U8542 (N_8542,N_4949,N_1732);
and U8543 (N_8543,N_152,N_3438);
nand U8544 (N_8544,N_3620,N_1967);
or U8545 (N_8545,N_2842,N_3329);
nand U8546 (N_8546,N_2915,N_1373);
nand U8547 (N_8547,N_2389,N_2763);
and U8548 (N_8548,N_1643,N_1380);
nor U8549 (N_8549,N_400,N_2781);
or U8550 (N_8550,N_4382,N_1006);
nand U8551 (N_8551,N_1400,N_3879);
and U8552 (N_8552,N_2339,N_4673);
xnor U8553 (N_8553,N_135,N_3576);
nor U8554 (N_8554,N_1003,N_516);
or U8555 (N_8555,N_817,N_3832);
nand U8556 (N_8556,N_1215,N_1159);
and U8557 (N_8557,N_3744,N_1165);
nor U8558 (N_8558,N_1478,N_3523);
or U8559 (N_8559,N_2432,N_529);
and U8560 (N_8560,N_207,N_1420);
and U8561 (N_8561,N_3683,N_4352);
nand U8562 (N_8562,N_2457,N_1548);
nor U8563 (N_8563,N_3551,N_4745);
xor U8564 (N_8564,N_3995,N_2059);
nand U8565 (N_8565,N_3391,N_1749);
nand U8566 (N_8566,N_1267,N_843);
nand U8567 (N_8567,N_3960,N_3920);
or U8568 (N_8568,N_381,N_3796);
nand U8569 (N_8569,N_3317,N_2036);
nand U8570 (N_8570,N_3005,N_1217);
and U8571 (N_8571,N_866,N_3763);
nor U8572 (N_8572,N_4398,N_2699);
nor U8573 (N_8573,N_4274,N_2056);
or U8574 (N_8574,N_165,N_4265);
nor U8575 (N_8575,N_2893,N_3041);
and U8576 (N_8576,N_48,N_4913);
or U8577 (N_8577,N_4798,N_570);
nor U8578 (N_8578,N_92,N_1897);
or U8579 (N_8579,N_1697,N_683);
or U8580 (N_8580,N_1885,N_2137);
and U8581 (N_8581,N_3165,N_3715);
nor U8582 (N_8582,N_2200,N_3221);
and U8583 (N_8583,N_2415,N_361);
nor U8584 (N_8584,N_2688,N_1690);
nand U8585 (N_8585,N_2749,N_3614);
nand U8586 (N_8586,N_1793,N_1694);
nand U8587 (N_8587,N_895,N_2755);
nand U8588 (N_8588,N_4525,N_249);
xor U8589 (N_8589,N_4899,N_3894);
and U8590 (N_8590,N_3197,N_2172);
or U8591 (N_8591,N_1263,N_758);
nand U8592 (N_8592,N_1614,N_3329);
nor U8593 (N_8593,N_4274,N_2526);
or U8594 (N_8594,N_4106,N_4286);
and U8595 (N_8595,N_960,N_105);
xor U8596 (N_8596,N_4328,N_4590);
or U8597 (N_8597,N_1370,N_3134);
and U8598 (N_8598,N_1404,N_3917);
nor U8599 (N_8599,N_1568,N_4506);
or U8600 (N_8600,N_2802,N_2371);
nand U8601 (N_8601,N_275,N_4885);
and U8602 (N_8602,N_2726,N_3107);
and U8603 (N_8603,N_755,N_4365);
and U8604 (N_8604,N_4755,N_2563);
or U8605 (N_8605,N_4172,N_3276);
or U8606 (N_8606,N_2454,N_3476);
or U8607 (N_8607,N_3088,N_3370);
nand U8608 (N_8608,N_2969,N_2125);
nand U8609 (N_8609,N_3765,N_3468);
nand U8610 (N_8610,N_4454,N_4653);
or U8611 (N_8611,N_4183,N_2690);
nand U8612 (N_8612,N_950,N_2530);
or U8613 (N_8613,N_2831,N_3563);
and U8614 (N_8614,N_2838,N_4052);
or U8615 (N_8615,N_230,N_553);
or U8616 (N_8616,N_4293,N_1269);
nor U8617 (N_8617,N_1569,N_120);
or U8618 (N_8618,N_1086,N_3386);
nand U8619 (N_8619,N_4216,N_3997);
or U8620 (N_8620,N_2913,N_436);
and U8621 (N_8621,N_4605,N_4800);
and U8622 (N_8622,N_1891,N_4848);
or U8623 (N_8623,N_2546,N_743);
nor U8624 (N_8624,N_2390,N_3729);
nor U8625 (N_8625,N_3670,N_1304);
nand U8626 (N_8626,N_3551,N_3456);
nor U8627 (N_8627,N_1432,N_4656);
nand U8628 (N_8628,N_1569,N_769);
or U8629 (N_8629,N_3724,N_4799);
or U8630 (N_8630,N_4266,N_745);
nand U8631 (N_8631,N_3554,N_2975);
nor U8632 (N_8632,N_4782,N_4137);
or U8633 (N_8633,N_2537,N_1791);
and U8634 (N_8634,N_284,N_4398);
or U8635 (N_8635,N_3910,N_3510);
nor U8636 (N_8636,N_1855,N_2090);
or U8637 (N_8637,N_648,N_227);
or U8638 (N_8638,N_2991,N_2330);
xnor U8639 (N_8639,N_1948,N_4952);
nor U8640 (N_8640,N_2139,N_2138);
or U8641 (N_8641,N_686,N_3670);
or U8642 (N_8642,N_4222,N_4095);
nor U8643 (N_8643,N_625,N_1491);
or U8644 (N_8644,N_1813,N_686);
nor U8645 (N_8645,N_1273,N_2148);
and U8646 (N_8646,N_1200,N_47);
nand U8647 (N_8647,N_1052,N_4043);
or U8648 (N_8648,N_3568,N_446);
and U8649 (N_8649,N_2277,N_247);
or U8650 (N_8650,N_4839,N_3969);
nand U8651 (N_8651,N_1700,N_671);
nor U8652 (N_8652,N_3520,N_4647);
xor U8653 (N_8653,N_1414,N_2853);
xor U8654 (N_8654,N_2596,N_3588);
or U8655 (N_8655,N_4100,N_1903);
nor U8656 (N_8656,N_87,N_988);
nor U8657 (N_8657,N_4955,N_3716);
or U8658 (N_8658,N_3721,N_3873);
nand U8659 (N_8659,N_3740,N_3317);
and U8660 (N_8660,N_4746,N_371);
nand U8661 (N_8661,N_3447,N_3237);
and U8662 (N_8662,N_614,N_4101);
and U8663 (N_8663,N_1907,N_4834);
and U8664 (N_8664,N_4375,N_536);
nand U8665 (N_8665,N_2633,N_3345);
nor U8666 (N_8666,N_1062,N_4602);
or U8667 (N_8667,N_1312,N_3966);
or U8668 (N_8668,N_3161,N_2773);
nand U8669 (N_8669,N_2469,N_3919);
and U8670 (N_8670,N_372,N_4554);
nand U8671 (N_8671,N_1928,N_3503);
nor U8672 (N_8672,N_1578,N_4749);
and U8673 (N_8673,N_3309,N_394);
and U8674 (N_8674,N_1542,N_3647);
or U8675 (N_8675,N_4517,N_3875);
nor U8676 (N_8676,N_1620,N_3948);
nand U8677 (N_8677,N_106,N_1375);
or U8678 (N_8678,N_494,N_1945);
or U8679 (N_8679,N_2250,N_2127);
nand U8680 (N_8680,N_1858,N_371);
nor U8681 (N_8681,N_3463,N_3023);
and U8682 (N_8682,N_4040,N_3511);
and U8683 (N_8683,N_364,N_1420);
nand U8684 (N_8684,N_3638,N_2974);
or U8685 (N_8685,N_4003,N_4929);
nor U8686 (N_8686,N_463,N_1716);
and U8687 (N_8687,N_57,N_4215);
nand U8688 (N_8688,N_3359,N_1418);
nand U8689 (N_8689,N_4896,N_3235);
nand U8690 (N_8690,N_2414,N_6);
nand U8691 (N_8691,N_1241,N_4980);
and U8692 (N_8692,N_676,N_4519);
or U8693 (N_8693,N_537,N_2479);
and U8694 (N_8694,N_4833,N_1726);
nor U8695 (N_8695,N_3966,N_2337);
nor U8696 (N_8696,N_2214,N_830);
nor U8697 (N_8697,N_4746,N_3811);
nor U8698 (N_8698,N_4853,N_3744);
and U8699 (N_8699,N_2827,N_2094);
nor U8700 (N_8700,N_4653,N_2554);
nand U8701 (N_8701,N_1601,N_2717);
nor U8702 (N_8702,N_1828,N_1793);
or U8703 (N_8703,N_1158,N_3763);
nand U8704 (N_8704,N_868,N_230);
or U8705 (N_8705,N_2014,N_1665);
and U8706 (N_8706,N_107,N_222);
nand U8707 (N_8707,N_640,N_1384);
nand U8708 (N_8708,N_234,N_3838);
nor U8709 (N_8709,N_3800,N_3369);
or U8710 (N_8710,N_812,N_695);
nand U8711 (N_8711,N_3435,N_3647);
nor U8712 (N_8712,N_690,N_4486);
or U8713 (N_8713,N_4505,N_4513);
nor U8714 (N_8714,N_1986,N_685);
and U8715 (N_8715,N_4164,N_920);
and U8716 (N_8716,N_3414,N_1490);
nand U8717 (N_8717,N_4350,N_3690);
nor U8718 (N_8718,N_4367,N_2208);
or U8719 (N_8719,N_1473,N_3512);
nand U8720 (N_8720,N_542,N_4747);
nand U8721 (N_8721,N_3785,N_1341);
or U8722 (N_8722,N_917,N_4420);
nand U8723 (N_8723,N_2824,N_3284);
or U8724 (N_8724,N_2706,N_2393);
nand U8725 (N_8725,N_4209,N_864);
nand U8726 (N_8726,N_170,N_4252);
nor U8727 (N_8727,N_4325,N_2062);
and U8728 (N_8728,N_1958,N_3549);
or U8729 (N_8729,N_1712,N_3469);
or U8730 (N_8730,N_251,N_1916);
or U8731 (N_8731,N_4180,N_1430);
nand U8732 (N_8732,N_3041,N_900);
nand U8733 (N_8733,N_2045,N_1448);
and U8734 (N_8734,N_3909,N_3294);
or U8735 (N_8735,N_787,N_1124);
and U8736 (N_8736,N_566,N_1000);
nand U8737 (N_8737,N_1708,N_4691);
or U8738 (N_8738,N_186,N_1540);
or U8739 (N_8739,N_3721,N_4539);
or U8740 (N_8740,N_2222,N_986);
xor U8741 (N_8741,N_1286,N_757);
and U8742 (N_8742,N_3041,N_325);
and U8743 (N_8743,N_2412,N_1306);
nor U8744 (N_8744,N_3608,N_1806);
nor U8745 (N_8745,N_2084,N_3717);
or U8746 (N_8746,N_1857,N_3792);
nor U8747 (N_8747,N_1136,N_4891);
or U8748 (N_8748,N_306,N_2119);
nand U8749 (N_8749,N_765,N_772);
and U8750 (N_8750,N_3166,N_3311);
and U8751 (N_8751,N_3313,N_1786);
and U8752 (N_8752,N_1824,N_2369);
nand U8753 (N_8753,N_4742,N_4900);
or U8754 (N_8754,N_4350,N_1807);
nand U8755 (N_8755,N_622,N_4342);
or U8756 (N_8756,N_4882,N_4748);
nor U8757 (N_8757,N_3262,N_3591);
nor U8758 (N_8758,N_4289,N_2599);
and U8759 (N_8759,N_3383,N_4744);
nor U8760 (N_8760,N_2636,N_2815);
nor U8761 (N_8761,N_2659,N_1736);
and U8762 (N_8762,N_3217,N_4130);
or U8763 (N_8763,N_3585,N_3052);
or U8764 (N_8764,N_27,N_954);
nand U8765 (N_8765,N_2029,N_3354);
nor U8766 (N_8766,N_2488,N_2213);
nand U8767 (N_8767,N_2171,N_1421);
nand U8768 (N_8768,N_3643,N_4775);
nor U8769 (N_8769,N_1144,N_2805);
or U8770 (N_8770,N_4038,N_1628);
and U8771 (N_8771,N_3967,N_4769);
or U8772 (N_8772,N_3507,N_251);
nand U8773 (N_8773,N_4724,N_1053);
or U8774 (N_8774,N_2348,N_1128);
nand U8775 (N_8775,N_4944,N_783);
xnor U8776 (N_8776,N_4022,N_2138);
nand U8777 (N_8777,N_929,N_4676);
xor U8778 (N_8778,N_2418,N_4546);
xnor U8779 (N_8779,N_2354,N_3583);
nand U8780 (N_8780,N_3080,N_1076);
nor U8781 (N_8781,N_179,N_4448);
nand U8782 (N_8782,N_856,N_4314);
nor U8783 (N_8783,N_2919,N_967);
nor U8784 (N_8784,N_1051,N_2873);
nor U8785 (N_8785,N_2368,N_2778);
nand U8786 (N_8786,N_1496,N_3328);
nor U8787 (N_8787,N_3724,N_3308);
nor U8788 (N_8788,N_2725,N_2843);
nand U8789 (N_8789,N_745,N_580);
nor U8790 (N_8790,N_4157,N_1714);
nor U8791 (N_8791,N_4793,N_104);
nand U8792 (N_8792,N_712,N_3363);
or U8793 (N_8793,N_345,N_2685);
nor U8794 (N_8794,N_384,N_1959);
nor U8795 (N_8795,N_1772,N_4287);
nand U8796 (N_8796,N_4967,N_1168);
nand U8797 (N_8797,N_4050,N_1638);
nand U8798 (N_8798,N_4800,N_1329);
nand U8799 (N_8799,N_298,N_2316);
nand U8800 (N_8800,N_4397,N_2011);
nand U8801 (N_8801,N_2451,N_4590);
xnor U8802 (N_8802,N_4961,N_4763);
xnor U8803 (N_8803,N_2822,N_4668);
nand U8804 (N_8804,N_4329,N_3193);
nand U8805 (N_8805,N_762,N_4802);
nand U8806 (N_8806,N_56,N_210);
nor U8807 (N_8807,N_3879,N_597);
or U8808 (N_8808,N_3363,N_3236);
and U8809 (N_8809,N_1534,N_1077);
or U8810 (N_8810,N_2352,N_2240);
nor U8811 (N_8811,N_4035,N_4800);
and U8812 (N_8812,N_443,N_3500);
or U8813 (N_8813,N_329,N_868);
nand U8814 (N_8814,N_3680,N_1273);
and U8815 (N_8815,N_4296,N_729);
or U8816 (N_8816,N_1261,N_841);
and U8817 (N_8817,N_4264,N_2083);
nor U8818 (N_8818,N_1703,N_2196);
or U8819 (N_8819,N_895,N_3799);
and U8820 (N_8820,N_64,N_2439);
nand U8821 (N_8821,N_2279,N_102);
or U8822 (N_8822,N_1685,N_3242);
nand U8823 (N_8823,N_4818,N_2153);
or U8824 (N_8824,N_1367,N_2419);
nor U8825 (N_8825,N_2494,N_3995);
or U8826 (N_8826,N_505,N_2404);
xnor U8827 (N_8827,N_4614,N_3859);
nand U8828 (N_8828,N_2025,N_3591);
or U8829 (N_8829,N_3914,N_2656);
and U8830 (N_8830,N_3232,N_2280);
xnor U8831 (N_8831,N_3909,N_2015);
and U8832 (N_8832,N_3426,N_1150);
or U8833 (N_8833,N_3020,N_1963);
and U8834 (N_8834,N_841,N_4227);
nand U8835 (N_8835,N_3534,N_2477);
and U8836 (N_8836,N_785,N_4570);
and U8837 (N_8837,N_1684,N_3167);
nor U8838 (N_8838,N_333,N_2668);
or U8839 (N_8839,N_2406,N_4319);
and U8840 (N_8840,N_1564,N_1786);
nand U8841 (N_8841,N_1270,N_2659);
and U8842 (N_8842,N_80,N_3395);
nand U8843 (N_8843,N_4139,N_2941);
and U8844 (N_8844,N_1348,N_532);
nor U8845 (N_8845,N_2717,N_2018);
or U8846 (N_8846,N_3519,N_4836);
nor U8847 (N_8847,N_4072,N_4734);
or U8848 (N_8848,N_3434,N_566);
and U8849 (N_8849,N_4164,N_3210);
nor U8850 (N_8850,N_566,N_2640);
nand U8851 (N_8851,N_3542,N_627);
or U8852 (N_8852,N_4342,N_4640);
nand U8853 (N_8853,N_1800,N_3257);
or U8854 (N_8854,N_2186,N_4207);
nor U8855 (N_8855,N_3354,N_2229);
nor U8856 (N_8856,N_4704,N_2495);
and U8857 (N_8857,N_829,N_131);
or U8858 (N_8858,N_3078,N_4308);
or U8859 (N_8859,N_2811,N_3518);
and U8860 (N_8860,N_4145,N_3145);
nor U8861 (N_8861,N_2749,N_2089);
xnor U8862 (N_8862,N_2666,N_581);
or U8863 (N_8863,N_345,N_950);
and U8864 (N_8864,N_1975,N_914);
xnor U8865 (N_8865,N_4644,N_2494);
and U8866 (N_8866,N_3803,N_4820);
nand U8867 (N_8867,N_1570,N_3209);
nand U8868 (N_8868,N_4043,N_448);
nand U8869 (N_8869,N_2291,N_3230);
nand U8870 (N_8870,N_902,N_1739);
or U8871 (N_8871,N_3124,N_2109);
and U8872 (N_8872,N_1069,N_395);
nand U8873 (N_8873,N_3886,N_877);
and U8874 (N_8874,N_4589,N_4231);
or U8875 (N_8875,N_3152,N_1222);
and U8876 (N_8876,N_4968,N_2848);
and U8877 (N_8877,N_2055,N_2660);
and U8878 (N_8878,N_4324,N_2172);
or U8879 (N_8879,N_1535,N_284);
nor U8880 (N_8880,N_2500,N_1996);
nand U8881 (N_8881,N_2726,N_1456);
and U8882 (N_8882,N_1173,N_1480);
nand U8883 (N_8883,N_995,N_1053);
nor U8884 (N_8884,N_3507,N_949);
nand U8885 (N_8885,N_3137,N_1101);
nand U8886 (N_8886,N_4919,N_409);
nand U8887 (N_8887,N_1840,N_1364);
and U8888 (N_8888,N_4120,N_3056);
and U8889 (N_8889,N_3342,N_247);
nand U8890 (N_8890,N_3984,N_1620);
nand U8891 (N_8891,N_4436,N_3973);
and U8892 (N_8892,N_2900,N_437);
and U8893 (N_8893,N_2712,N_516);
or U8894 (N_8894,N_1613,N_4620);
or U8895 (N_8895,N_1547,N_4103);
nand U8896 (N_8896,N_2687,N_2344);
and U8897 (N_8897,N_2552,N_735);
nor U8898 (N_8898,N_3730,N_1470);
nand U8899 (N_8899,N_1347,N_417);
nand U8900 (N_8900,N_1085,N_458);
and U8901 (N_8901,N_509,N_4715);
nor U8902 (N_8902,N_1929,N_1670);
nand U8903 (N_8903,N_2297,N_1100);
and U8904 (N_8904,N_37,N_2208);
or U8905 (N_8905,N_3416,N_1493);
nand U8906 (N_8906,N_3080,N_4937);
nor U8907 (N_8907,N_2533,N_2996);
nor U8908 (N_8908,N_2900,N_4912);
nand U8909 (N_8909,N_3824,N_650);
and U8910 (N_8910,N_2483,N_2155);
nand U8911 (N_8911,N_2762,N_3043);
or U8912 (N_8912,N_584,N_3716);
nor U8913 (N_8913,N_3237,N_1886);
nand U8914 (N_8914,N_559,N_3762);
or U8915 (N_8915,N_3495,N_3406);
or U8916 (N_8916,N_2816,N_2383);
nand U8917 (N_8917,N_3378,N_2196);
or U8918 (N_8918,N_537,N_2775);
nand U8919 (N_8919,N_646,N_1928);
or U8920 (N_8920,N_3877,N_3775);
and U8921 (N_8921,N_1324,N_4186);
and U8922 (N_8922,N_3874,N_2659);
or U8923 (N_8923,N_82,N_2262);
nand U8924 (N_8924,N_2494,N_4438);
and U8925 (N_8925,N_920,N_879);
xnor U8926 (N_8926,N_2171,N_94);
nor U8927 (N_8927,N_2409,N_3019);
and U8928 (N_8928,N_3576,N_3261);
or U8929 (N_8929,N_248,N_310);
or U8930 (N_8930,N_132,N_1529);
nand U8931 (N_8931,N_1908,N_1422);
nor U8932 (N_8932,N_24,N_2182);
nor U8933 (N_8933,N_2481,N_2813);
nor U8934 (N_8934,N_1717,N_2966);
and U8935 (N_8935,N_4686,N_4363);
and U8936 (N_8936,N_1157,N_3004);
and U8937 (N_8937,N_1639,N_2029);
nand U8938 (N_8938,N_1057,N_2864);
or U8939 (N_8939,N_2707,N_1670);
or U8940 (N_8940,N_1942,N_3669);
nor U8941 (N_8941,N_2937,N_4816);
nor U8942 (N_8942,N_2135,N_1188);
nand U8943 (N_8943,N_4671,N_4424);
and U8944 (N_8944,N_1850,N_4592);
nand U8945 (N_8945,N_2754,N_2179);
and U8946 (N_8946,N_4153,N_3453);
or U8947 (N_8947,N_1241,N_3912);
and U8948 (N_8948,N_191,N_252);
xor U8949 (N_8949,N_2733,N_2507);
nand U8950 (N_8950,N_529,N_1815);
and U8951 (N_8951,N_826,N_2898);
or U8952 (N_8952,N_866,N_2333);
nor U8953 (N_8953,N_1040,N_2424);
nand U8954 (N_8954,N_3541,N_1463);
and U8955 (N_8955,N_3651,N_590);
or U8956 (N_8956,N_2090,N_4518);
nand U8957 (N_8957,N_3486,N_4155);
nor U8958 (N_8958,N_2566,N_3991);
and U8959 (N_8959,N_1548,N_110);
nand U8960 (N_8960,N_4150,N_2944);
nor U8961 (N_8961,N_4920,N_293);
or U8962 (N_8962,N_1797,N_232);
and U8963 (N_8963,N_1294,N_4314);
and U8964 (N_8964,N_959,N_3929);
nand U8965 (N_8965,N_4102,N_2485);
or U8966 (N_8966,N_4248,N_2922);
or U8967 (N_8967,N_557,N_1897);
xnor U8968 (N_8968,N_4127,N_3942);
nor U8969 (N_8969,N_663,N_192);
or U8970 (N_8970,N_2790,N_4895);
or U8971 (N_8971,N_1013,N_2948);
or U8972 (N_8972,N_4857,N_3190);
or U8973 (N_8973,N_2262,N_375);
nand U8974 (N_8974,N_1614,N_229);
nand U8975 (N_8975,N_4234,N_2877);
nand U8976 (N_8976,N_2938,N_1601);
or U8977 (N_8977,N_1460,N_4670);
nand U8978 (N_8978,N_1647,N_2266);
nor U8979 (N_8979,N_1704,N_95);
or U8980 (N_8980,N_2753,N_1945);
and U8981 (N_8981,N_4675,N_314);
and U8982 (N_8982,N_3050,N_854);
and U8983 (N_8983,N_264,N_2040);
and U8984 (N_8984,N_2727,N_486);
nand U8985 (N_8985,N_4248,N_3698);
nand U8986 (N_8986,N_290,N_3873);
or U8987 (N_8987,N_3122,N_4518);
or U8988 (N_8988,N_2034,N_4707);
or U8989 (N_8989,N_132,N_234);
nor U8990 (N_8990,N_3339,N_3675);
and U8991 (N_8991,N_1007,N_668);
nand U8992 (N_8992,N_3848,N_1754);
nand U8993 (N_8993,N_2770,N_2172);
nand U8994 (N_8994,N_3779,N_4334);
or U8995 (N_8995,N_4530,N_3144);
or U8996 (N_8996,N_4053,N_4744);
nor U8997 (N_8997,N_1720,N_1099);
and U8998 (N_8998,N_4867,N_1544);
nor U8999 (N_8999,N_1078,N_4867);
or U9000 (N_9000,N_4038,N_2465);
nand U9001 (N_9001,N_3109,N_4544);
nor U9002 (N_9002,N_1354,N_4821);
nor U9003 (N_9003,N_3432,N_3351);
nor U9004 (N_9004,N_2517,N_4177);
nor U9005 (N_9005,N_160,N_3187);
nor U9006 (N_9006,N_834,N_2692);
nor U9007 (N_9007,N_1523,N_577);
nor U9008 (N_9008,N_1374,N_3220);
and U9009 (N_9009,N_2634,N_1817);
xor U9010 (N_9010,N_304,N_1212);
nor U9011 (N_9011,N_1370,N_1341);
nor U9012 (N_9012,N_1892,N_820);
and U9013 (N_9013,N_698,N_593);
and U9014 (N_9014,N_4183,N_3265);
and U9015 (N_9015,N_4568,N_4046);
nand U9016 (N_9016,N_551,N_3307);
and U9017 (N_9017,N_2092,N_3511);
or U9018 (N_9018,N_136,N_2661);
or U9019 (N_9019,N_802,N_4889);
nor U9020 (N_9020,N_3770,N_972);
or U9021 (N_9021,N_4658,N_1816);
nand U9022 (N_9022,N_4540,N_1456);
nor U9023 (N_9023,N_751,N_4632);
and U9024 (N_9024,N_1581,N_2354);
or U9025 (N_9025,N_4251,N_1042);
and U9026 (N_9026,N_1823,N_1507);
nand U9027 (N_9027,N_4150,N_403);
nor U9028 (N_9028,N_15,N_4544);
nand U9029 (N_9029,N_1459,N_3187);
nor U9030 (N_9030,N_192,N_2234);
nor U9031 (N_9031,N_4422,N_1017);
nor U9032 (N_9032,N_133,N_1310);
nand U9033 (N_9033,N_4189,N_109);
nand U9034 (N_9034,N_106,N_1578);
nor U9035 (N_9035,N_3894,N_3454);
and U9036 (N_9036,N_4510,N_2112);
nor U9037 (N_9037,N_4899,N_4611);
and U9038 (N_9038,N_4908,N_3443);
and U9039 (N_9039,N_1936,N_3598);
nand U9040 (N_9040,N_449,N_3791);
or U9041 (N_9041,N_2518,N_606);
and U9042 (N_9042,N_4106,N_2869);
and U9043 (N_9043,N_654,N_3364);
and U9044 (N_9044,N_1458,N_4214);
nor U9045 (N_9045,N_1077,N_3724);
nor U9046 (N_9046,N_4119,N_2934);
nor U9047 (N_9047,N_4430,N_4494);
nor U9048 (N_9048,N_3767,N_3301);
or U9049 (N_9049,N_1232,N_2848);
or U9050 (N_9050,N_4293,N_959);
nor U9051 (N_9051,N_386,N_29);
or U9052 (N_9052,N_1061,N_3651);
nor U9053 (N_9053,N_4706,N_1189);
and U9054 (N_9054,N_4828,N_1012);
nor U9055 (N_9055,N_2203,N_220);
or U9056 (N_9056,N_4726,N_4860);
nand U9057 (N_9057,N_4553,N_1611);
nand U9058 (N_9058,N_1807,N_2334);
and U9059 (N_9059,N_1243,N_2581);
or U9060 (N_9060,N_4810,N_979);
or U9061 (N_9061,N_4758,N_3659);
nand U9062 (N_9062,N_2238,N_3823);
nor U9063 (N_9063,N_4749,N_2450);
and U9064 (N_9064,N_1005,N_3904);
nand U9065 (N_9065,N_2022,N_3663);
or U9066 (N_9066,N_3478,N_3254);
nor U9067 (N_9067,N_1862,N_3449);
nor U9068 (N_9068,N_3444,N_4089);
or U9069 (N_9069,N_4331,N_1909);
or U9070 (N_9070,N_623,N_845);
nor U9071 (N_9071,N_2716,N_4680);
xnor U9072 (N_9072,N_4756,N_99);
nor U9073 (N_9073,N_713,N_4981);
xnor U9074 (N_9074,N_2230,N_267);
nor U9075 (N_9075,N_1428,N_467);
nand U9076 (N_9076,N_2527,N_3736);
and U9077 (N_9077,N_388,N_2613);
nor U9078 (N_9078,N_3200,N_4333);
and U9079 (N_9079,N_4225,N_3429);
and U9080 (N_9080,N_4259,N_2959);
nor U9081 (N_9081,N_4439,N_2209);
nand U9082 (N_9082,N_3324,N_4440);
nor U9083 (N_9083,N_387,N_4197);
and U9084 (N_9084,N_493,N_4232);
nand U9085 (N_9085,N_2125,N_3985);
nor U9086 (N_9086,N_686,N_1871);
or U9087 (N_9087,N_3742,N_3765);
or U9088 (N_9088,N_2417,N_2187);
nand U9089 (N_9089,N_2550,N_2590);
nor U9090 (N_9090,N_972,N_495);
or U9091 (N_9091,N_4340,N_2041);
or U9092 (N_9092,N_1994,N_2723);
xnor U9093 (N_9093,N_4900,N_3713);
and U9094 (N_9094,N_2872,N_135);
nor U9095 (N_9095,N_2784,N_4140);
nand U9096 (N_9096,N_2934,N_4894);
nand U9097 (N_9097,N_771,N_3416);
or U9098 (N_9098,N_1474,N_229);
or U9099 (N_9099,N_1510,N_1811);
and U9100 (N_9100,N_3780,N_1140);
or U9101 (N_9101,N_2405,N_3207);
and U9102 (N_9102,N_1909,N_4297);
nand U9103 (N_9103,N_2851,N_1366);
nor U9104 (N_9104,N_2711,N_1359);
nand U9105 (N_9105,N_935,N_2430);
nand U9106 (N_9106,N_3841,N_1185);
nand U9107 (N_9107,N_1311,N_3614);
or U9108 (N_9108,N_1761,N_1425);
nand U9109 (N_9109,N_1851,N_4587);
nor U9110 (N_9110,N_4678,N_866);
nand U9111 (N_9111,N_4725,N_2166);
and U9112 (N_9112,N_3812,N_972);
nor U9113 (N_9113,N_612,N_671);
or U9114 (N_9114,N_1393,N_3267);
or U9115 (N_9115,N_1065,N_3032);
and U9116 (N_9116,N_693,N_1974);
nor U9117 (N_9117,N_4053,N_1232);
nor U9118 (N_9118,N_4156,N_3620);
and U9119 (N_9119,N_2422,N_217);
or U9120 (N_9120,N_4009,N_4584);
or U9121 (N_9121,N_1896,N_2061);
nor U9122 (N_9122,N_305,N_687);
and U9123 (N_9123,N_769,N_2499);
nand U9124 (N_9124,N_1834,N_1654);
nand U9125 (N_9125,N_4566,N_1475);
nand U9126 (N_9126,N_930,N_1820);
nor U9127 (N_9127,N_2024,N_2565);
nand U9128 (N_9128,N_1697,N_4415);
nor U9129 (N_9129,N_1683,N_4468);
or U9130 (N_9130,N_3399,N_2848);
and U9131 (N_9131,N_2980,N_4893);
or U9132 (N_9132,N_326,N_993);
nand U9133 (N_9133,N_4948,N_2254);
nor U9134 (N_9134,N_2851,N_356);
or U9135 (N_9135,N_4615,N_4761);
nand U9136 (N_9136,N_738,N_1442);
and U9137 (N_9137,N_25,N_1979);
nand U9138 (N_9138,N_4333,N_1092);
or U9139 (N_9139,N_2237,N_3281);
and U9140 (N_9140,N_2581,N_371);
or U9141 (N_9141,N_3204,N_4585);
and U9142 (N_9142,N_1732,N_3715);
and U9143 (N_9143,N_4480,N_3728);
or U9144 (N_9144,N_2688,N_4212);
nor U9145 (N_9145,N_1914,N_2753);
nor U9146 (N_9146,N_3950,N_149);
and U9147 (N_9147,N_3729,N_3721);
and U9148 (N_9148,N_1993,N_464);
or U9149 (N_9149,N_1511,N_175);
nor U9150 (N_9150,N_4996,N_3997);
nand U9151 (N_9151,N_1375,N_1508);
nand U9152 (N_9152,N_4359,N_492);
nand U9153 (N_9153,N_3402,N_1520);
nor U9154 (N_9154,N_1315,N_2838);
xor U9155 (N_9155,N_1642,N_4519);
nand U9156 (N_9156,N_2678,N_3854);
nand U9157 (N_9157,N_3439,N_2072);
nor U9158 (N_9158,N_3534,N_3732);
and U9159 (N_9159,N_1004,N_2114);
or U9160 (N_9160,N_1396,N_4272);
nor U9161 (N_9161,N_2134,N_3501);
or U9162 (N_9162,N_1804,N_1736);
nor U9163 (N_9163,N_356,N_3710);
or U9164 (N_9164,N_1351,N_4986);
and U9165 (N_9165,N_1559,N_777);
or U9166 (N_9166,N_4170,N_4931);
or U9167 (N_9167,N_4170,N_3455);
xnor U9168 (N_9168,N_4498,N_4620);
nand U9169 (N_9169,N_1053,N_4459);
or U9170 (N_9170,N_59,N_1202);
nor U9171 (N_9171,N_2204,N_3909);
or U9172 (N_9172,N_3829,N_2243);
and U9173 (N_9173,N_4632,N_3508);
nand U9174 (N_9174,N_1021,N_2158);
nor U9175 (N_9175,N_1925,N_2044);
and U9176 (N_9176,N_2064,N_2718);
or U9177 (N_9177,N_564,N_1433);
or U9178 (N_9178,N_404,N_1938);
nand U9179 (N_9179,N_4717,N_765);
xor U9180 (N_9180,N_3625,N_2465);
nor U9181 (N_9181,N_1205,N_1920);
nor U9182 (N_9182,N_4444,N_3674);
nand U9183 (N_9183,N_1880,N_4042);
nor U9184 (N_9184,N_1293,N_4643);
or U9185 (N_9185,N_193,N_2136);
and U9186 (N_9186,N_4189,N_4486);
nor U9187 (N_9187,N_744,N_597);
or U9188 (N_9188,N_4501,N_230);
nand U9189 (N_9189,N_3045,N_2784);
nand U9190 (N_9190,N_172,N_4959);
and U9191 (N_9191,N_1663,N_3352);
and U9192 (N_9192,N_3342,N_76);
nor U9193 (N_9193,N_3607,N_3472);
nor U9194 (N_9194,N_630,N_3110);
nor U9195 (N_9195,N_3126,N_584);
or U9196 (N_9196,N_686,N_1420);
or U9197 (N_9197,N_855,N_934);
nand U9198 (N_9198,N_4854,N_4882);
nor U9199 (N_9199,N_2199,N_3400);
nor U9200 (N_9200,N_1980,N_4607);
nor U9201 (N_9201,N_4122,N_4393);
nor U9202 (N_9202,N_295,N_4962);
and U9203 (N_9203,N_4468,N_4256);
or U9204 (N_9204,N_2188,N_1144);
or U9205 (N_9205,N_1170,N_2463);
nor U9206 (N_9206,N_4888,N_1608);
nor U9207 (N_9207,N_4488,N_2951);
nand U9208 (N_9208,N_4279,N_3918);
nor U9209 (N_9209,N_4261,N_3950);
or U9210 (N_9210,N_800,N_2510);
nand U9211 (N_9211,N_2238,N_4699);
and U9212 (N_9212,N_822,N_798);
or U9213 (N_9213,N_373,N_1387);
nor U9214 (N_9214,N_2254,N_3673);
nand U9215 (N_9215,N_3488,N_122);
or U9216 (N_9216,N_4601,N_2818);
and U9217 (N_9217,N_3703,N_4559);
and U9218 (N_9218,N_683,N_1563);
nand U9219 (N_9219,N_2527,N_322);
nor U9220 (N_9220,N_3505,N_3518);
nor U9221 (N_9221,N_2827,N_2942);
nand U9222 (N_9222,N_71,N_3006);
nand U9223 (N_9223,N_3002,N_648);
nand U9224 (N_9224,N_107,N_4052);
nor U9225 (N_9225,N_4138,N_4108);
and U9226 (N_9226,N_708,N_1790);
and U9227 (N_9227,N_477,N_124);
nor U9228 (N_9228,N_1092,N_2975);
and U9229 (N_9229,N_4489,N_4635);
nor U9230 (N_9230,N_267,N_2828);
and U9231 (N_9231,N_4351,N_306);
nand U9232 (N_9232,N_2243,N_2432);
nor U9233 (N_9233,N_1463,N_3878);
nand U9234 (N_9234,N_1870,N_3529);
xor U9235 (N_9235,N_2674,N_1887);
nor U9236 (N_9236,N_3231,N_1413);
or U9237 (N_9237,N_3493,N_462);
nand U9238 (N_9238,N_3254,N_2007);
nand U9239 (N_9239,N_1471,N_4647);
or U9240 (N_9240,N_305,N_2157);
and U9241 (N_9241,N_3590,N_2167);
nor U9242 (N_9242,N_227,N_4555);
or U9243 (N_9243,N_3739,N_4261);
and U9244 (N_9244,N_2062,N_3330);
and U9245 (N_9245,N_1688,N_2231);
nand U9246 (N_9246,N_2016,N_995);
or U9247 (N_9247,N_1732,N_1151);
or U9248 (N_9248,N_628,N_1195);
nand U9249 (N_9249,N_1824,N_4514);
and U9250 (N_9250,N_688,N_2131);
nand U9251 (N_9251,N_3845,N_193);
or U9252 (N_9252,N_1891,N_3528);
nor U9253 (N_9253,N_1413,N_515);
and U9254 (N_9254,N_3854,N_1723);
and U9255 (N_9255,N_1602,N_868);
nand U9256 (N_9256,N_2211,N_1179);
and U9257 (N_9257,N_3744,N_3774);
and U9258 (N_9258,N_1671,N_655);
and U9259 (N_9259,N_4111,N_4530);
nor U9260 (N_9260,N_3174,N_1217);
nor U9261 (N_9261,N_2137,N_4540);
or U9262 (N_9262,N_4063,N_2402);
nor U9263 (N_9263,N_2370,N_1680);
or U9264 (N_9264,N_3619,N_4258);
and U9265 (N_9265,N_1187,N_3817);
nor U9266 (N_9266,N_4085,N_1772);
nand U9267 (N_9267,N_2795,N_1678);
nor U9268 (N_9268,N_88,N_4037);
or U9269 (N_9269,N_320,N_3973);
nor U9270 (N_9270,N_4009,N_3716);
or U9271 (N_9271,N_2257,N_1104);
nand U9272 (N_9272,N_1424,N_637);
nor U9273 (N_9273,N_2633,N_4013);
xor U9274 (N_9274,N_2609,N_825);
nand U9275 (N_9275,N_2802,N_3255);
or U9276 (N_9276,N_4570,N_3324);
nand U9277 (N_9277,N_1908,N_2056);
nor U9278 (N_9278,N_453,N_2384);
nor U9279 (N_9279,N_3597,N_4675);
xor U9280 (N_9280,N_163,N_946);
and U9281 (N_9281,N_2032,N_3304);
and U9282 (N_9282,N_1323,N_1884);
and U9283 (N_9283,N_1786,N_3340);
and U9284 (N_9284,N_4547,N_58);
or U9285 (N_9285,N_3585,N_2633);
nand U9286 (N_9286,N_2921,N_3568);
or U9287 (N_9287,N_3540,N_1973);
or U9288 (N_9288,N_1402,N_4971);
nor U9289 (N_9289,N_4816,N_734);
or U9290 (N_9290,N_4521,N_4071);
or U9291 (N_9291,N_2614,N_1671);
or U9292 (N_9292,N_473,N_1642);
nor U9293 (N_9293,N_2563,N_577);
and U9294 (N_9294,N_3463,N_2079);
or U9295 (N_9295,N_4688,N_2064);
and U9296 (N_9296,N_225,N_2809);
and U9297 (N_9297,N_3623,N_4510);
nand U9298 (N_9298,N_2619,N_1433);
or U9299 (N_9299,N_362,N_400);
and U9300 (N_9300,N_4242,N_4310);
and U9301 (N_9301,N_1430,N_3678);
nand U9302 (N_9302,N_3192,N_3440);
nand U9303 (N_9303,N_2974,N_3644);
and U9304 (N_9304,N_2801,N_4583);
nand U9305 (N_9305,N_1958,N_4100);
nand U9306 (N_9306,N_1287,N_164);
nand U9307 (N_9307,N_3772,N_423);
nand U9308 (N_9308,N_1183,N_2769);
nand U9309 (N_9309,N_3422,N_281);
nand U9310 (N_9310,N_3567,N_4969);
nor U9311 (N_9311,N_273,N_4738);
or U9312 (N_9312,N_1440,N_4051);
nor U9313 (N_9313,N_21,N_1970);
or U9314 (N_9314,N_22,N_2006);
nor U9315 (N_9315,N_1408,N_3671);
and U9316 (N_9316,N_4399,N_4549);
nor U9317 (N_9317,N_4731,N_3868);
nand U9318 (N_9318,N_120,N_3231);
nand U9319 (N_9319,N_1307,N_2023);
and U9320 (N_9320,N_427,N_2365);
nor U9321 (N_9321,N_981,N_2714);
and U9322 (N_9322,N_1447,N_63);
or U9323 (N_9323,N_143,N_1076);
nor U9324 (N_9324,N_1671,N_4037);
nor U9325 (N_9325,N_2513,N_160);
xor U9326 (N_9326,N_1964,N_2824);
and U9327 (N_9327,N_4027,N_1851);
and U9328 (N_9328,N_3512,N_4285);
nor U9329 (N_9329,N_4560,N_2570);
or U9330 (N_9330,N_4077,N_4598);
nor U9331 (N_9331,N_2708,N_113);
or U9332 (N_9332,N_1757,N_4462);
nor U9333 (N_9333,N_3668,N_1707);
or U9334 (N_9334,N_2219,N_2408);
and U9335 (N_9335,N_3938,N_962);
or U9336 (N_9336,N_666,N_478);
or U9337 (N_9337,N_1154,N_4322);
nor U9338 (N_9338,N_3911,N_1963);
nand U9339 (N_9339,N_3719,N_754);
and U9340 (N_9340,N_4172,N_833);
nand U9341 (N_9341,N_1805,N_1581);
or U9342 (N_9342,N_3987,N_4110);
or U9343 (N_9343,N_1741,N_2085);
and U9344 (N_9344,N_4684,N_3086);
nand U9345 (N_9345,N_4535,N_2630);
nor U9346 (N_9346,N_1492,N_4808);
nand U9347 (N_9347,N_3589,N_1068);
nand U9348 (N_9348,N_635,N_2228);
nand U9349 (N_9349,N_4909,N_493);
or U9350 (N_9350,N_904,N_274);
and U9351 (N_9351,N_3187,N_1175);
nor U9352 (N_9352,N_212,N_2040);
nor U9353 (N_9353,N_728,N_2530);
and U9354 (N_9354,N_2443,N_335);
and U9355 (N_9355,N_1790,N_4516);
or U9356 (N_9356,N_1202,N_3299);
nand U9357 (N_9357,N_4259,N_713);
or U9358 (N_9358,N_768,N_2204);
or U9359 (N_9359,N_1490,N_658);
nand U9360 (N_9360,N_1037,N_94);
nand U9361 (N_9361,N_1443,N_4999);
nor U9362 (N_9362,N_2983,N_4864);
nor U9363 (N_9363,N_4699,N_2122);
nand U9364 (N_9364,N_2611,N_2721);
and U9365 (N_9365,N_204,N_919);
and U9366 (N_9366,N_857,N_2044);
nand U9367 (N_9367,N_186,N_3598);
or U9368 (N_9368,N_3565,N_3216);
or U9369 (N_9369,N_2247,N_2471);
or U9370 (N_9370,N_2705,N_4253);
and U9371 (N_9371,N_3318,N_4087);
and U9372 (N_9372,N_56,N_2011);
and U9373 (N_9373,N_3243,N_4408);
and U9374 (N_9374,N_1350,N_2607);
nor U9375 (N_9375,N_3783,N_2695);
nor U9376 (N_9376,N_232,N_121);
nor U9377 (N_9377,N_3028,N_4437);
xnor U9378 (N_9378,N_4006,N_811);
nand U9379 (N_9379,N_1225,N_2046);
nand U9380 (N_9380,N_515,N_2885);
nor U9381 (N_9381,N_1642,N_3702);
nor U9382 (N_9382,N_1918,N_199);
nand U9383 (N_9383,N_951,N_4736);
or U9384 (N_9384,N_4316,N_3981);
or U9385 (N_9385,N_4719,N_3116);
nor U9386 (N_9386,N_294,N_4103);
xnor U9387 (N_9387,N_1114,N_865);
nor U9388 (N_9388,N_4825,N_3602);
nor U9389 (N_9389,N_2195,N_632);
nand U9390 (N_9390,N_3940,N_1248);
nand U9391 (N_9391,N_194,N_4309);
and U9392 (N_9392,N_3922,N_4773);
or U9393 (N_9393,N_4564,N_2941);
and U9394 (N_9394,N_2203,N_3743);
nor U9395 (N_9395,N_1323,N_404);
nor U9396 (N_9396,N_4952,N_849);
and U9397 (N_9397,N_2380,N_2083);
nand U9398 (N_9398,N_2185,N_1705);
or U9399 (N_9399,N_2252,N_3964);
and U9400 (N_9400,N_1125,N_2672);
or U9401 (N_9401,N_4380,N_4195);
nand U9402 (N_9402,N_1228,N_3091);
nor U9403 (N_9403,N_1715,N_84);
and U9404 (N_9404,N_2609,N_4051);
nand U9405 (N_9405,N_1584,N_105);
or U9406 (N_9406,N_4555,N_3871);
or U9407 (N_9407,N_1582,N_3134);
nand U9408 (N_9408,N_3751,N_1876);
nand U9409 (N_9409,N_2164,N_3301);
and U9410 (N_9410,N_1759,N_3863);
or U9411 (N_9411,N_1094,N_664);
and U9412 (N_9412,N_4674,N_2509);
nand U9413 (N_9413,N_2629,N_2141);
nand U9414 (N_9414,N_3673,N_3247);
nor U9415 (N_9415,N_4965,N_3365);
nand U9416 (N_9416,N_893,N_1562);
and U9417 (N_9417,N_930,N_1415);
nor U9418 (N_9418,N_2293,N_1541);
or U9419 (N_9419,N_1486,N_4114);
nor U9420 (N_9420,N_4311,N_127);
nor U9421 (N_9421,N_155,N_3270);
nor U9422 (N_9422,N_4871,N_3996);
and U9423 (N_9423,N_1663,N_2500);
nand U9424 (N_9424,N_3478,N_2407);
nand U9425 (N_9425,N_3605,N_4963);
and U9426 (N_9426,N_1176,N_1845);
and U9427 (N_9427,N_1556,N_2495);
and U9428 (N_9428,N_437,N_3851);
nand U9429 (N_9429,N_31,N_1331);
or U9430 (N_9430,N_876,N_2797);
or U9431 (N_9431,N_4792,N_4793);
xnor U9432 (N_9432,N_3234,N_769);
and U9433 (N_9433,N_2348,N_4702);
and U9434 (N_9434,N_2285,N_2489);
and U9435 (N_9435,N_756,N_1056);
and U9436 (N_9436,N_69,N_3211);
or U9437 (N_9437,N_326,N_3526);
nor U9438 (N_9438,N_652,N_4826);
or U9439 (N_9439,N_1702,N_720);
xnor U9440 (N_9440,N_2118,N_470);
nor U9441 (N_9441,N_566,N_4044);
or U9442 (N_9442,N_2664,N_2631);
or U9443 (N_9443,N_746,N_4427);
or U9444 (N_9444,N_1811,N_4716);
and U9445 (N_9445,N_196,N_1048);
nand U9446 (N_9446,N_3568,N_1889);
xnor U9447 (N_9447,N_2562,N_1972);
xnor U9448 (N_9448,N_1805,N_1888);
nor U9449 (N_9449,N_2821,N_3436);
and U9450 (N_9450,N_3320,N_19);
nand U9451 (N_9451,N_2627,N_581);
nand U9452 (N_9452,N_2143,N_255);
and U9453 (N_9453,N_1763,N_1901);
nand U9454 (N_9454,N_526,N_2567);
or U9455 (N_9455,N_1224,N_4162);
or U9456 (N_9456,N_3970,N_243);
and U9457 (N_9457,N_493,N_3359);
and U9458 (N_9458,N_3126,N_2237);
or U9459 (N_9459,N_4365,N_2348);
nand U9460 (N_9460,N_2887,N_4487);
or U9461 (N_9461,N_190,N_4523);
and U9462 (N_9462,N_3461,N_543);
and U9463 (N_9463,N_4566,N_2497);
and U9464 (N_9464,N_3697,N_1213);
nor U9465 (N_9465,N_4901,N_4960);
and U9466 (N_9466,N_3434,N_2028);
nor U9467 (N_9467,N_4480,N_3482);
nor U9468 (N_9468,N_4128,N_2362);
or U9469 (N_9469,N_199,N_4441);
nor U9470 (N_9470,N_1559,N_4036);
and U9471 (N_9471,N_666,N_2293);
nand U9472 (N_9472,N_4898,N_3008);
and U9473 (N_9473,N_1026,N_255);
nor U9474 (N_9474,N_1136,N_3076);
or U9475 (N_9475,N_4307,N_3099);
or U9476 (N_9476,N_2970,N_848);
xnor U9477 (N_9477,N_4478,N_2681);
nand U9478 (N_9478,N_4367,N_817);
or U9479 (N_9479,N_4747,N_4649);
and U9480 (N_9480,N_2840,N_4972);
and U9481 (N_9481,N_2902,N_3908);
or U9482 (N_9482,N_4298,N_4304);
nand U9483 (N_9483,N_3254,N_2166);
nor U9484 (N_9484,N_2580,N_2866);
or U9485 (N_9485,N_2206,N_2636);
and U9486 (N_9486,N_754,N_1698);
and U9487 (N_9487,N_4393,N_4408);
nor U9488 (N_9488,N_680,N_3647);
nor U9489 (N_9489,N_1893,N_3480);
nand U9490 (N_9490,N_4409,N_1662);
nor U9491 (N_9491,N_4045,N_2166);
or U9492 (N_9492,N_3770,N_1349);
and U9493 (N_9493,N_250,N_1362);
nor U9494 (N_9494,N_651,N_75);
nand U9495 (N_9495,N_1961,N_1746);
nor U9496 (N_9496,N_58,N_274);
or U9497 (N_9497,N_1846,N_2580);
and U9498 (N_9498,N_1168,N_3926);
nor U9499 (N_9499,N_2116,N_4506);
nand U9500 (N_9500,N_123,N_4337);
nor U9501 (N_9501,N_4052,N_3305);
nor U9502 (N_9502,N_3374,N_785);
nor U9503 (N_9503,N_176,N_183);
or U9504 (N_9504,N_3851,N_2226);
and U9505 (N_9505,N_1490,N_2678);
nand U9506 (N_9506,N_2685,N_2854);
nor U9507 (N_9507,N_9,N_4809);
nor U9508 (N_9508,N_2004,N_3972);
or U9509 (N_9509,N_3889,N_1172);
or U9510 (N_9510,N_2503,N_4506);
nor U9511 (N_9511,N_4281,N_4636);
nor U9512 (N_9512,N_4265,N_353);
nand U9513 (N_9513,N_865,N_4596);
or U9514 (N_9514,N_695,N_1259);
and U9515 (N_9515,N_25,N_4005);
and U9516 (N_9516,N_2632,N_3075);
and U9517 (N_9517,N_4475,N_4080);
xor U9518 (N_9518,N_1171,N_486);
or U9519 (N_9519,N_4310,N_4464);
or U9520 (N_9520,N_2666,N_3998);
nor U9521 (N_9521,N_2454,N_2721);
xnor U9522 (N_9522,N_4549,N_1965);
or U9523 (N_9523,N_2867,N_3139);
or U9524 (N_9524,N_3855,N_2988);
xnor U9525 (N_9525,N_2332,N_1935);
nand U9526 (N_9526,N_3441,N_2895);
and U9527 (N_9527,N_593,N_1925);
and U9528 (N_9528,N_4884,N_11);
or U9529 (N_9529,N_4155,N_2688);
nand U9530 (N_9530,N_2166,N_1206);
or U9531 (N_9531,N_3589,N_47);
or U9532 (N_9532,N_1157,N_3285);
or U9533 (N_9533,N_1141,N_3482);
nand U9534 (N_9534,N_58,N_4408);
nand U9535 (N_9535,N_4719,N_2054);
xor U9536 (N_9536,N_3620,N_3749);
nor U9537 (N_9537,N_3102,N_1671);
or U9538 (N_9538,N_4915,N_3336);
nor U9539 (N_9539,N_4983,N_1630);
and U9540 (N_9540,N_4242,N_2279);
nand U9541 (N_9541,N_1737,N_434);
or U9542 (N_9542,N_3257,N_2771);
nand U9543 (N_9543,N_4027,N_362);
nand U9544 (N_9544,N_1017,N_910);
and U9545 (N_9545,N_3235,N_2421);
nand U9546 (N_9546,N_2826,N_1272);
or U9547 (N_9547,N_2609,N_2015);
nor U9548 (N_9548,N_1151,N_2910);
nand U9549 (N_9549,N_3271,N_3162);
and U9550 (N_9550,N_2309,N_4944);
or U9551 (N_9551,N_3253,N_2317);
xnor U9552 (N_9552,N_3916,N_3546);
nor U9553 (N_9553,N_2442,N_3378);
nand U9554 (N_9554,N_2471,N_837);
nor U9555 (N_9555,N_3348,N_1439);
nor U9556 (N_9556,N_932,N_3313);
or U9557 (N_9557,N_3396,N_1360);
and U9558 (N_9558,N_2612,N_1030);
nor U9559 (N_9559,N_3330,N_2499);
or U9560 (N_9560,N_3085,N_3616);
nand U9561 (N_9561,N_3740,N_709);
nor U9562 (N_9562,N_3862,N_4998);
xor U9563 (N_9563,N_3189,N_605);
nor U9564 (N_9564,N_467,N_4399);
and U9565 (N_9565,N_1656,N_3541);
or U9566 (N_9566,N_4549,N_581);
nor U9567 (N_9567,N_2903,N_1973);
nand U9568 (N_9568,N_1210,N_4106);
or U9569 (N_9569,N_56,N_440);
nor U9570 (N_9570,N_48,N_2185);
or U9571 (N_9571,N_79,N_4000);
xnor U9572 (N_9572,N_442,N_3331);
nand U9573 (N_9573,N_577,N_1138);
nand U9574 (N_9574,N_3846,N_679);
nand U9575 (N_9575,N_4796,N_3491);
nor U9576 (N_9576,N_3828,N_3083);
and U9577 (N_9577,N_4320,N_274);
nand U9578 (N_9578,N_4808,N_2039);
nand U9579 (N_9579,N_3450,N_866);
and U9580 (N_9580,N_2007,N_1539);
nand U9581 (N_9581,N_1232,N_423);
nor U9582 (N_9582,N_3502,N_3079);
and U9583 (N_9583,N_865,N_4879);
xor U9584 (N_9584,N_1679,N_3005);
or U9585 (N_9585,N_206,N_1457);
nor U9586 (N_9586,N_3182,N_2886);
and U9587 (N_9587,N_3628,N_3853);
and U9588 (N_9588,N_3424,N_2246);
nor U9589 (N_9589,N_3726,N_4891);
nor U9590 (N_9590,N_911,N_3510);
nor U9591 (N_9591,N_659,N_4373);
and U9592 (N_9592,N_1339,N_723);
xnor U9593 (N_9593,N_4891,N_297);
nor U9594 (N_9594,N_4004,N_601);
nor U9595 (N_9595,N_2373,N_3076);
nand U9596 (N_9596,N_1566,N_2733);
or U9597 (N_9597,N_923,N_3481);
or U9598 (N_9598,N_1,N_3772);
nor U9599 (N_9599,N_633,N_1198);
and U9600 (N_9600,N_2634,N_850);
and U9601 (N_9601,N_2542,N_1360);
nand U9602 (N_9602,N_2860,N_2201);
nor U9603 (N_9603,N_463,N_2307);
nand U9604 (N_9604,N_3976,N_2084);
nor U9605 (N_9605,N_441,N_336);
nor U9606 (N_9606,N_4812,N_1776);
nor U9607 (N_9607,N_4189,N_4476);
or U9608 (N_9608,N_3779,N_2163);
nor U9609 (N_9609,N_824,N_3586);
and U9610 (N_9610,N_19,N_302);
xor U9611 (N_9611,N_2979,N_2239);
or U9612 (N_9612,N_2413,N_3638);
nand U9613 (N_9613,N_122,N_2581);
nand U9614 (N_9614,N_2299,N_4460);
and U9615 (N_9615,N_72,N_2369);
or U9616 (N_9616,N_2745,N_1003);
or U9617 (N_9617,N_3680,N_857);
or U9618 (N_9618,N_1928,N_3240);
or U9619 (N_9619,N_4481,N_4556);
nor U9620 (N_9620,N_2256,N_3039);
nand U9621 (N_9621,N_4863,N_1715);
or U9622 (N_9622,N_4339,N_2959);
or U9623 (N_9623,N_4632,N_3609);
nand U9624 (N_9624,N_2820,N_2536);
nand U9625 (N_9625,N_3114,N_3330);
or U9626 (N_9626,N_1241,N_1743);
nand U9627 (N_9627,N_2971,N_1912);
and U9628 (N_9628,N_2192,N_2259);
or U9629 (N_9629,N_4713,N_2310);
and U9630 (N_9630,N_3345,N_1495);
nor U9631 (N_9631,N_1496,N_4807);
nor U9632 (N_9632,N_76,N_2521);
or U9633 (N_9633,N_2826,N_4036);
or U9634 (N_9634,N_432,N_441);
or U9635 (N_9635,N_4983,N_4533);
or U9636 (N_9636,N_2670,N_3488);
or U9637 (N_9637,N_899,N_862);
and U9638 (N_9638,N_3243,N_1089);
nand U9639 (N_9639,N_3827,N_4530);
and U9640 (N_9640,N_4436,N_619);
nand U9641 (N_9641,N_380,N_1572);
nor U9642 (N_9642,N_3243,N_2988);
and U9643 (N_9643,N_2129,N_2925);
nor U9644 (N_9644,N_3397,N_3076);
and U9645 (N_9645,N_3735,N_1926);
nand U9646 (N_9646,N_1371,N_36);
or U9647 (N_9647,N_4594,N_1245);
nor U9648 (N_9648,N_4425,N_4215);
and U9649 (N_9649,N_2085,N_748);
nor U9650 (N_9650,N_4929,N_1500);
nor U9651 (N_9651,N_1276,N_2716);
nor U9652 (N_9652,N_3421,N_431);
and U9653 (N_9653,N_4503,N_4965);
nor U9654 (N_9654,N_2877,N_4480);
nand U9655 (N_9655,N_4004,N_2493);
nand U9656 (N_9656,N_3909,N_4745);
and U9657 (N_9657,N_2987,N_2890);
and U9658 (N_9658,N_4417,N_2650);
or U9659 (N_9659,N_1928,N_1555);
or U9660 (N_9660,N_3161,N_3388);
or U9661 (N_9661,N_4674,N_4355);
or U9662 (N_9662,N_4654,N_2150);
nand U9663 (N_9663,N_2718,N_1282);
and U9664 (N_9664,N_1897,N_2067);
nand U9665 (N_9665,N_1791,N_144);
and U9666 (N_9666,N_939,N_4089);
nand U9667 (N_9667,N_3893,N_1074);
and U9668 (N_9668,N_2052,N_3397);
nand U9669 (N_9669,N_4915,N_3800);
or U9670 (N_9670,N_1890,N_2353);
or U9671 (N_9671,N_2965,N_3302);
nand U9672 (N_9672,N_2090,N_2641);
nand U9673 (N_9673,N_3846,N_1766);
xor U9674 (N_9674,N_3591,N_4343);
or U9675 (N_9675,N_1070,N_996);
xor U9676 (N_9676,N_3851,N_817);
or U9677 (N_9677,N_3089,N_1935);
nand U9678 (N_9678,N_1199,N_3834);
nand U9679 (N_9679,N_4995,N_345);
nand U9680 (N_9680,N_4953,N_4966);
and U9681 (N_9681,N_1715,N_4102);
nand U9682 (N_9682,N_671,N_425);
nor U9683 (N_9683,N_2737,N_2518);
or U9684 (N_9684,N_3036,N_3285);
and U9685 (N_9685,N_2958,N_1636);
nor U9686 (N_9686,N_976,N_2328);
nand U9687 (N_9687,N_1722,N_4663);
or U9688 (N_9688,N_2069,N_1882);
nand U9689 (N_9689,N_4659,N_3998);
nand U9690 (N_9690,N_4801,N_2151);
or U9691 (N_9691,N_30,N_4118);
nor U9692 (N_9692,N_244,N_1709);
and U9693 (N_9693,N_4597,N_1080);
nor U9694 (N_9694,N_2809,N_1412);
or U9695 (N_9695,N_4002,N_1329);
or U9696 (N_9696,N_4760,N_1661);
or U9697 (N_9697,N_1636,N_4795);
nand U9698 (N_9698,N_2889,N_1102);
or U9699 (N_9699,N_1984,N_2503);
nand U9700 (N_9700,N_2395,N_253);
and U9701 (N_9701,N_3220,N_4065);
nand U9702 (N_9702,N_4633,N_890);
nand U9703 (N_9703,N_2075,N_4701);
and U9704 (N_9704,N_3612,N_1109);
nor U9705 (N_9705,N_2577,N_1384);
or U9706 (N_9706,N_2456,N_136);
nor U9707 (N_9707,N_1961,N_3707);
nand U9708 (N_9708,N_4515,N_3184);
xnor U9709 (N_9709,N_75,N_4999);
or U9710 (N_9710,N_4105,N_2489);
and U9711 (N_9711,N_1602,N_1944);
or U9712 (N_9712,N_4596,N_1952);
or U9713 (N_9713,N_2372,N_3456);
nor U9714 (N_9714,N_2715,N_2);
or U9715 (N_9715,N_2891,N_4361);
and U9716 (N_9716,N_4461,N_1169);
nor U9717 (N_9717,N_170,N_1044);
nand U9718 (N_9718,N_1897,N_2454);
nand U9719 (N_9719,N_660,N_1948);
and U9720 (N_9720,N_3453,N_4837);
nor U9721 (N_9721,N_1799,N_3889);
nor U9722 (N_9722,N_3626,N_1906);
nand U9723 (N_9723,N_3400,N_2568);
or U9724 (N_9724,N_1111,N_3817);
nor U9725 (N_9725,N_4454,N_1479);
nor U9726 (N_9726,N_2365,N_1967);
and U9727 (N_9727,N_3287,N_2505);
or U9728 (N_9728,N_1581,N_1563);
and U9729 (N_9729,N_2986,N_296);
or U9730 (N_9730,N_3516,N_3076);
nor U9731 (N_9731,N_1514,N_3694);
and U9732 (N_9732,N_2980,N_2897);
or U9733 (N_9733,N_555,N_1150);
nand U9734 (N_9734,N_2115,N_2848);
nor U9735 (N_9735,N_547,N_3228);
nand U9736 (N_9736,N_533,N_4568);
or U9737 (N_9737,N_1891,N_4644);
nand U9738 (N_9738,N_2055,N_2145);
nand U9739 (N_9739,N_3427,N_49);
nor U9740 (N_9740,N_4799,N_3273);
and U9741 (N_9741,N_2544,N_2725);
nor U9742 (N_9742,N_3863,N_251);
and U9743 (N_9743,N_1672,N_4654);
and U9744 (N_9744,N_3386,N_4080);
nor U9745 (N_9745,N_3609,N_1908);
nor U9746 (N_9746,N_3686,N_2502);
or U9747 (N_9747,N_2724,N_9);
or U9748 (N_9748,N_3874,N_1211);
or U9749 (N_9749,N_3704,N_1187);
nand U9750 (N_9750,N_2528,N_2141);
or U9751 (N_9751,N_4416,N_3602);
nor U9752 (N_9752,N_3552,N_2929);
nand U9753 (N_9753,N_2166,N_687);
or U9754 (N_9754,N_2135,N_2748);
nand U9755 (N_9755,N_3890,N_790);
or U9756 (N_9756,N_2235,N_4100);
or U9757 (N_9757,N_2720,N_3992);
or U9758 (N_9758,N_86,N_3561);
nor U9759 (N_9759,N_1984,N_2065);
and U9760 (N_9760,N_1974,N_417);
and U9761 (N_9761,N_3708,N_1495);
and U9762 (N_9762,N_2041,N_232);
xor U9763 (N_9763,N_4474,N_853);
nand U9764 (N_9764,N_4118,N_3950);
and U9765 (N_9765,N_3457,N_1157);
nor U9766 (N_9766,N_4348,N_4653);
and U9767 (N_9767,N_4788,N_3216);
and U9768 (N_9768,N_1339,N_579);
nand U9769 (N_9769,N_659,N_4632);
or U9770 (N_9770,N_3012,N_3617);
nor U9771 (N_9771,N_3572,N_354);
nand U9772 (N_9772,N_1107,N_2170);
nand U9773 (N_9773,N_2004,N_2015);
nor U9774 (N_9774,N_2229,N_3729);
or U9775 (N_9775,N_3482,N_3876);
or U9776 (N_9776,N_758,N_2298);
and U9777 (N_9777,N_4488,N_4949);
or U9778 (N_9778,N_3018,N_295);
or U9779 (N_9779,N_2923,N_4728);
and U9780 (N_9780,N_4653,N_4648);
and U9781 (N_9781,N_3537,N_1270);
and U9782 (N_9782,N_3745,N_2037);
or U9783 (N_9783,N_4650,N_4086);
nor U9784 (N_9784,N_3790,N_2106);
nand U9785 (N_9785,N_3142,N_3117);
nand U9786 (N_9786,N_2001,N_2858);
or U9787 (N_9787,N_2576,N_3543);
nor U9788 (N_9788,N_388,N_3486);
or U9789 (N_9789,N_1222,N_383);
and U9790 (N_9790,N_25,N_4254);
and U9791 (N_9791,N_4543,N_4890);
or U9792 (N_9792,N_1709,N_2718);
nor U9793 (N_9793,N_978,N_560);
nor U9794 (N_9794,N_1719,N_2340);
and U9795 (N_9795,N_2272,N_1678);
nand U9796 (N_9796,N_2430,N_400);
nand U9797 (N_9797,N_3265,N_2410);
and U9798 (N_9798,N_883,N_1759);
and U9799 (N_9799,N_2063,N_4098);
and U9800 (N_9800,N_1590,N_1699);
or U9801 (N_9801,N_2315,N_1531);
nor U9802 (N_9802,N_2330,N_688);
or U9803 (N_9803,N_4641,N_1816);
and U9804 (N_9804,N_13,N_4706);
and U9805 (N_9805,N_1414,N_307);
or U9806 (N_9806,N_4247,N_550);
and U9807 (N_9807,N_4995,N_772);
and U9808 (N_9808,N_4689,N_742);
or U9809 (N_9809,N_2589,N_2620);
or U9810 (N_9810,N_2133,N_3542);
or U9811 (N_9811,N_916,N_4302);
nand U9812 (N_9812,N_2957,N_1183);
nor U9813 (N_9813,N_875,N_4967);
or U9814 (N_9814,N_1528,N_389);
or U9815 (N_9815,N_3377,N_591);
nor U9816 (N_9816,N_3948,N_2649);
nand U9817 (N_9817,N_1853,N_4291);
or U9818 (N_9818,N_3190,N_3583);
nand U9819 (N_9819,N_3938,N_1851);
and U9820 (N_9820,N_881,N_2780);
or U9821 (N_9821,N_4108,N_2529);
or U9822 (N_9822,N_4831,N_1788);
nand U9823 (N_9823,N_2228,N_3985);
and U9824 (N_9824,N_1079,N_1274);
nor U9825 (N_9825,N_3594,N_476);
and U9826 (N_9826,N_2774,N_3358);
or U9827 (N_9827,N_4731,N_3032);
and U9828 (N_9828,N_3245,N_975);
and U9829 (N_9829,N_4358,N_1985);
nor U9830 (N_9830,N_3532,N_4906);
nor U9831 (N_9831,N_4209,N_777);
or U9832 (N_9832,N_4878,N_539);
nor U9833 (N_9833,N_3195,N_1051);
and U9834 (N_9834,N_4361,N_1621);
nor U9835 (N_9835,N_3967,N_4644);
nand U9836 (N_9836,N_3999,N_1598);
xnor U9837 (N_9837,N_1787,N_3641);
or U9838 (N_9838,N_4381,N_3958);
or U9839 (N_9839,N_4467,N_2990);
and U9840 (N_9840,N_2400,N_107);
and U9841 (N_9841,N_938,N_1701);
nor U9842 (N_9842,N_4377,N_998);
and U9843 (N_9843,N_2106,N_3906);
nand U9844 (N_9844,N_2231,N_3939);
xor U9845 (N_9845,N_2327,N_1336);
nand U9846 (N_9846,N_4148,N_2609);
nor U9847 (N_9847,N_2665,N_3355);
xnor U9848 (N_9848,N_816,N_4163);
nor U9849 (N_9849,N_3846,N_4804);
and U9850 (N_9850,N_3709,N_848);
or U9851 (N_9851,N_421,N_2686);
nor U9852 (N_9852,N_2063,N_4441);
or U9853 (N_9853,N_2842,N_1976);
nor U9854 (N_9854,N_2540,N_3984);
and U9855 (N_9855,N_4481,N_1159);
nand U9856 (N_9856,N_3019,N_4073);
nand U9857 (N_9857,N_418,N_840);
and U9858 (N_9858,N_2910,N_2891);
and U9859 (N_9859,N_4185,N_1191);
or U9860 (N_9860,N_3688,N_1325);
nor U9861 (N_9861,N_3217,N_4907);
or U9862 (N_9862,N_4417,N_4872);
and U9863 (N_9863,N_1594,N_2977);
xor U9864 (N_9864,N_140,N_1876);
nor U9865 (N_9865,N_245,N_501);
and U9866 (N_9866,N_4810,N_924);
or U9867 (N_9867,N_4322,N_2136);
nand U9868 (N_9868,N_941,N_2076);
nor U9869 (N_9869,N_952,N_4493);
nor U9870 (N_9870,N_2464,N_4145);
nand U9871 (N_9871,N_4320,N_312);
and U9872 (N_9872,N_255,N_4441);
or U9873 (N_9873,N_2117,N_3254);
and U9874 (N_9874,N_2860,N_4353);
or U9875 (N_9875,N_4855,N_2659);
nand U9876 (N_9876,N_233,N_944);
nand U9877 (N_9877,N_2092,N_184);
and U9878 (N_9878,N_556,N_1562);
and U9879 (N_9879,N_2649,N_509);
nand U9880 (N_9880,N_3286,N_3119);
or U9881 (N_9881,N_4836,N_3344);
nand U9882 (N_9882,N_3688,N_1486);
nand U9883 (N_9883,N_1323,N_415);
nand U9884 (N_9884,N_2200,N_4364);
nand U9885 (N_9885,N_4920,N_4230);
nand U9886 (N_9886,N_3521,N_4298);
or U9887 (N_9887,N_3505,N_3208);
nor U9888 (N_9888,N_2414,N_2652);
nor U9889 (N_9889,N_3170,N_814);
nor U9890 (N_9890,N_2780,N_719);
nor U9891 (N_9891,N_4884,N_2210);
or U9892 (N_9892,N_2090,N_1018);
nand U9893 (N_9893,N_959,N_4102);
and U9894 (N_9894,N_4363,N_4343);
and U9895 (N_9895,N_176,N_3770);
nand U9896 (N_9896,N_561,N_4053);
nand U9897 (N_9897,N_1820,N_632);
xnor U9898 (N_9898,N_3425,N_4801);
or U9899 (N_9899,N_3078,N_4180);
nor U9900 (N_9900,N_3410,N_510);
xor U9901 (N_9901,N_649,N_2914);
and U9902 (N_9902,N_3701,N_4696);
nand U9903 (N_9903,N_3243,N_3961);
and U9904 (N_9904,N_486,N_171);
and U9905 (N_9905,N_26,N_694);
and U9906 (N_9906,N_360,N_953);
nand U9907 (N_9907,N_4089,N_2223);
and U9908 (N_9908,N_2747,N_4800);
nand U9909 (N_9909,N_4487,N_7);
and U9910 (N_9910,N_2236,N_3525);
nor U9911 (N_9911,N_1141,N_2714);
nand U9912 (N_9912,N_82,N_3030);
or U9913 (N_9913,N_1555,N_1451);
nor U9914 (N_9914,N_982,N_2188);
nor U9915 (N_9915,N_4814,N_2112);
nand U9916 (N_9916,N_4822,N_3423);
nor U9917 (N_9917,N_4937,N_1609);
and U9918 (N_9918,N_2971,N_1835);
nor U9919 (N_9919,N_1455,N_4554);
or U9920 (N_9920,N_4050,N_2334);
and U9921 (N_9921,N_176,N_1010);
or U9922 (N_9922,N_2513,N_601);
or U9923 (N_9923,N_4034,N_3512);
or U9924 (N_9924,N_4582,N_446);
or U9925 (N_9925,N_246,N_3866);
nor U9926 (N_9926,N_2133,N_3920);
or U9927 (N_9927,N_4518,N_377);
nand U9928 (N_9928,N_2563,N_867);
or U9929 (N_9929,N_475,N_4579);
nor U9930 (N_9930,N_1414,N_2091);
nand U9931 (N_9931,N_1261,N_3117);
nor U9932 (N_9932,N_3394,N_4866);
or U9933 (N_9933,N_2961,N_3886);
nor U9934 (N_9934,N_3763,N_2920);
or U9935 (N_9935,N_906,N_2981);
nand U9936 (N_9936,N_2618,N_4297);
xnor U9937 (N_9937,N_4260,N_3212);
or U9938 (N_9938,N_319,N_2860);
nand U9939 (N_9939,N_1515,N_4104);
xnor U9940 (N_9940,N_479,N_3341);
nor U9941 (N_9941,N_4228,N_87);
or U9942 (N_9942,N_2359,N_3950);
nand U9943 (N_9943,N_571,N_3108);
nand U9944 (N_9944,N_2943,N_1604);
nor U9945 (N_9945,N_1875,N_1208);
nand U9946 (N_9946,N_259,N_2490);
and U9947 (N_9947,N_1165,N_4636);
and U9948 (N_9948,N_1546,N_1740);
and U9949 (N_9949,N_272,N_1338);
nor U9950 (N_9950,N_3385,N_3258);
nand U9951 (N_9951,N_483,N_2940);
nor U9952 (N_9952,N_4081,N_1816);
and U9953 (N_9953,N_4534,N_4834);
nand U9954 (N_9954,N_4373,N_820);
nor U9955 (N_9955,N_649,N_267);
nand U9956 (N_9956,N_619,N_2424);
and U9957 (N_9957,N_1289,N_258);
or U9958 (N_9958,N_1227,N_3115);
or U9959 (N_9959,N_116,N_3184);
xnor U9960 (N_9960,N_867,N_4890);
nand U9961 (N_9961,N_3266,N_4888);
or U9962 (N_9962,N_2769,N_3371);
and U9963 (N_9963,N_3658,N_107);
nand U9964 (N_9964,N_172,N_4672);
and U9965 (N_9965,N_4528,N_1031);
nor U9966 (N_9966,N_4363,N_3174);
or U9967 (N_9967,N_949,N_3376);
nor U9968 (N_9968,N_1409,N_2580);
nor U9969 (N_9969,N_2179,N_20);
nand U9970 (N_9970,N_4562,N_599);
and U9971 (N_9971,N_4084,N_4759);
nor U9972 (N_9972,N_2352,N_707);
nand U9973 (N_9973,N_4488,N_896);
and U9974 (N_9974,N_4606,N_2261);
nand U9975 (N_9975,N_3401,N_2771);
and U9976 (N_9976,N_4309,N_3336);
nor U9977 (N_9977,N_394,N_4553);
and U9978 (N_9978,N_2884,N_3601);
nor U9979 (N_9979,N_4351,N_4583);
nor U9980 (N_9980,N_2645,N_1327);
nor U9981 (N_9981,N_2419,N_187);
or U9982 (N_9982,N_4295,N_1934);
and U9983 (N_9983,N_112,N_1719);
nand U9984 (N_9984,N_3395,N_4168);
nand U9985 (N_9985,N_2108,N_203);
nand U9986 (N_9986,N_1803,N_1043);
nor U9987 (N_9987,N_1921,N_520);
and U9988 (N_9988,N_4032,N_1475);
nor U9989 (N_9989,N_3070,N_168);
and U9990 (N_9990,N_4781,N_1922);
nand U9991 (N_9991,N_2290,N_3206);
and U9992 (N_9992,N_2001,N_2012);
nor U9993 (N_9993,N_3425,N_2931);
or U9994 (N_9994,N_2529,N_4835);
and U9995 (N_9995,N_1845,N_904);
or U9996 (N_9996,N_1932,N_3555);
xnor U9997 (N_9997,N_2293,N_437);
and U9998 (N_9998,N_835,N_4373);
nand U9999 (N_9999,N_4134,N_4124);
and UO_0 (O_0,N_8598,N_6189);
nor UO_1 (O_1,N_5134,N_5334);
nor UO_2 (O_2,N_5386,N_8110);
nand UO_3 (O_3,N_9915,N_9771);
nand UO_4 (O_4,N_9738,N_9066);
or UO_5 (O_5,N_5478,N_7421);
xor UO_6 (O_6,N_6211,N_5355);
nand UO_7 (O_7,N_5728,N_5544);
nand UO_8 (O_8,N_7458,N_7583);
nand UO_9 (O_9,N_9489,N_5221);
nand UO_10 (O_10,N_9136,N_5705);
nand UO_11 (O_11,N_8434,N_6218);
nor UO_12 (O_12,N_7716,N_5503);
nand UO_13 (O_13,N_5155,N_8328);
or UO_14 (O_14,N_7637,N_9355);
or UO_15 (O_15,N_9339,N_6098);
or UO_16 (O_16,N_5859,N_6061);
nor UO_17 (O_17,N_7236,N_5771);
nand UO_18 (O_18,N_6675,N_5640);
or UO_19 (O_19,N_8073,N_5548);
nand UO_20 (O_20,N_7175,N_7357);
nor UO_21 (O_21,N_7747,N_8829);
or UO_22 (O_22,N_9457,N_9217);
nand UO_23 (O_23,N_5876,N_9475);
nand UO_24 (O_24,N_5766,N_6854);
or UO_25 (O_25,N_7755,N_5989);
and UO_26 (O_26,N_5020,N_9684);
nand UO_27 (O_27,N_6213,N_7883);
or UO_28 (O_28,N_9545,N_8317);
nand UO_29 (O_29,N_5136,N_7996);
and UO_30 (O_30,N_7569,N_9060);
nor UO_31 (O_31,N_6307,N_8902);
and UO_32 (O_32,N_9958,N_9076);
nand UO_33 (O_33,N_5521,N_8891);
nor UO_34 (O_34,N_9458,N_7290);
or UO_35 (O_35,N_8002,N_7628);
or UO_36 (O_36,N_9605,N_5925);
and UO_37 (O_37,N_8831,N_7442);
nand UO_38 (O_38,N_9970,N_5070);
nand UO_39 (O_39,N_5870,N_6379);
or UO_40 (O_40,N_8363,N_7949);
or UO_41 (O_41,N_8089,N_7035);
nand UO_42 (O_42,N_9146,N_7578);
and UO_43 (O_43,N_9990,N_8368);
and UO_44 (O_44,N_7938,N_6339);
xnor UO_45 (O_45,N_7582,N_9147);
and UO_46 (O_46,N_8796,N_6475);
nor UO_47 (O_47,N_8481,N_8597);
or UO_48 (O_48,N_9371,N_5873);
and UO_49 (O_49,N_6177,N_5200);
or UO_50 (O_50,N_8780,N_5270);
and UO_51 (O_51,N_5737,N_9503);
nor UO_52 (O_52,N_6783,N_6318);
nor UO_53 (O_53,N_9737,N_8250);
xor UO_54 (O_54,N_7049,N_8124);
nand UO_55 (O_55,N_9379,N_9947);
nand UO_56 (O_56,N_9277,N_6624);
nor UO_57 (O_57,N_9143,N_9312);
xor UO_58 (O_58,N_7071,N_9908);
nand UO_59 (O_59,N_7686,N_6420);
nand UO_60 (O_60,N_8261,N_5955);
nor UO_61 (O_61,N_5231,N_8390);
nor UO_62 (O_62,N_7550,N_5186);
nand UO_63 (O_63,N_7102,N_5865);
nand UO_64 (O_64,N_7679,N_8427);
or UO_65 (O_65,N_8857,N_9207);
nor UO_66 (O_66,N_8942,N_8437);
nor UO_67 (O_67,N_9837,N_8495);
or UO_68 (O_68,N_8890,N_8330);
nor UO_69 (O_69,N_9902,N_5677);
or UO_70 (O_70,N_8341,N_7935);
nand UO_71 (O_71,N_7137,N_6136);
nor UO_72 (O_72,N_9216,N_7203);
nand UO_73 (O_73,N_5847,N_7767);
and UO_74 (O_74,N_8405,N_7200);
or UO_75 (O_75,N_6151,N_8357);
or UO_76 (O_76,N_9986,N_9331);
nand UO_77 (O_77,N_9675,N_5042);
and UO_78 (O_78,N_8067,N_5214);
nor UO_79 (O_79,N_5276,N_8070);
nor UO_80 (O_80,N_8229,N_8923);
and UO_81 (O_81,N_6202,N_6469);
or UO_82 (O_82,N_6694,N_7879);
nor UO_83 (O_83,N_7307,N_8924);
nor UO_84 (O_84,N_5985,N_7094);
nand UO_85 (O_85,N_9100,N_7511);
or UO_86 (O_86,N_6735,N_9852);
nand UO_87 (O_87,N_8309,N_6220);
or UO_88 (O_88,N_5153,N_7598);
xnor UO_89 (O_89,N_6705,N_5391);
nor UO_90 (O_90,N_7590,N_8322);
nand UO_91 (O_91,N_9424,N_8922);
nor UO_92 (O_92,N_9607,N_6827);
xnor UO_93 (O_93,N_9812,N_5067);
and UO_94 (O_94,N_5370,N_6560);
and UO_95 (O_95,N_5307,N_5822);
and UO_96 (O_96,N_9614,N_9383);
nand UO_97 (O_97,N_6041,N_8763);
and UO_98 (O_98,N_5255,N_8315);
xor UO_99 (O_99,N_6270,N_8337);
or UO_100 (O_100,N_6463,N_7532);
nor UO_101 (O_101,N_6761,N_7995);
nand UO_102 (O_102,N_5192,N_6107);
and UO_103 (O_103,N_7677,N_9090);
nor UO_104 (O_104,N_9558,N_5234);
and UO_105 (O_105,N_7557,N_6702);
or UO_106 (O_106,N_5271,N_6736);
nor UO_107 (O_107,N_8214,N_9944);
nand UO_108 (O_108,N_9745,N_6908);
nand UO_109 (O_109,N_8870,N_8079);
or UO_110 (O_110,N_7846,N_5852);
or UO_111 (O_111,N_8592,N_5013);
nor UO_112 (O_112,N_8954,N_9418);
or UO_113 (O_113,N_9401,N_8200);
nand UO_114 (O_114,N_5601,N_5762);
and UO_115 (O_115,N_9604,N_5621);
or UO_116 (O_116,N_7393,N_8058);
nor UO_117 (O_117,N_5862,N_7843);
and UO_118 (O_118,N_5169,N_5472);
nand UO_119 (O_119,N_7813,N_9730);
or UO_120 (O_120,N_6371,N_6424);
and UO_121 (O_121,N_7856,N_7558);
nor UO_122 (O_122,N_5977,N_7069);
nor UO_123 (O_123,N_8952,N_8103);
or UO_124 (O_124,N_8137,N_5899);
and UO_125 (O_125,N_9054,N_8411);
and UO_126 (O_126,N_8100,N_7096);
nor UO_127 (O_127,N_6498,N_9250);
nor UO_128 (O_128,N_8052,N_8059);
nor UO_129 (O_129,N_6242,N_7509);
xnor UO_130 (O_130,N_9116,N_6855);
or UO_131 (O_131,N_5981,N_5321);
or UO_132 (O_132,N_8822,N_7176);
nand UO_133 (O_133,N_9195,N_5225);
and UO_134 (O_134,N_8778,N_6103);
or UO_135 (O_135,N_8758,N_9713);
or UO_136 (O_136,N_6750,N_8507);
nand UO_137 (O_137,N_6353,N_9827);
nand UO_138 (O_138,N_9751,N_7770);
or UO_139 (O_139,N_7559,N_7202);
and UO_140 (O_140,N_7502,N_6078);
or UO_141 (O_141,N_9756,N_9749);
nand UO_142 (O_142,N_5597,N_9861);
or UO_143 (O_143,N_7450,N_6873);
xor UO_144 (O_144,N_7121,N_7903);
or UO_145 (O_145,N_5662,N_5128);
or UO_146 (O_146,N_5571,N_9050);
nand UO_147 (O_147,N_6868,N_6237);
nor UO_148 (O_148,N_6878,N_6143);
nand UO_149 (O_149,N_9234,N_9820);
nor UO_150 (O_150,N_7118,N_5213);
nor UO_151 (O_151,N_9942,N_6661);
and UO_152 (O_152,N_5209,N_5806);
nand UO_153 (O_153,N_6127,N_7024);
nand UO_154 (O_154,N_7966,N_7242);
nor UO_155 (O_155,N_7310,N_8130);
or UO_156 (O_156,N_7065,N_6239);
and UO_157 (O_157,N_6315,N_7427);
or UO_158 (O_158,N_6505,N_8948);
or UO_159 (O_159,N_8361,N_6481);
nor UO_160 (O_160,N_8339,N_5826);
and UO_161 (O_161,N_6611,N_7623);
or UO_162 (O_162,N_5693,N_8134);
or UO_163 (O_163,N_7705,N_9222);
or UO_164 (O_164,N_7144,N_5863);
nor UO_165 (O_165,N_8715,N_8340);
or UO_166 (O_166,N_8677,N_9473);
and UO_167 (O_167,N_7886,N_5126);
nand UO_168 (O_168,N_5181,N_7457);
or UO_169 (O_169,N_9522,N_8521);
nand UO_170 (O_170,N_5482,N_9415);
nor UO_171 (O_171,N_6634,N_9982);
nor UO_172 (O_172,N_9498,N_5379);
nand UO_173 (O_173,N_5253,N_5403);
nand UO_174 (O_174,N_7685,N_8231);
nand UO_175 (O_175,N_9440,N_9588);
and UO_176 (O_176,N_8502,N_8406);
and UO_177 (O_177,N_6393,N_7530);
and UO_178 (O_178,N_9348,N_6225);
nor UO_179 (O_179,N_7790,N_7189);
nand UO_180 (O_180,N_5577,N_8743);
xnor UO_181 (O_181,N_9188,N_5112);
and UO_182 (O_182,N_9098,N_6494);
nand UO_183 (O_183,N_5460,N_8319);
nor UO_184 (O_184,N_7420,N_8996);
nand UO_185 (O_185,N_8702,N_9665);
or UO_186 (O_186,N_9907,N_8577);
nand UO_187 (O_187,N_9139,N_9006);
nand UO_188 (O_188,N_9936,N_7085);
nor UO_189 (O_189,N_9454,N_7003);
nand UO_190 (O_190,N_6576,N_9764);
nor UO_191 (O_191,N_7356,N_7104);
nand UO_192 (O_192,N_5110,N_7297);
and UO_193 (O_193,N_5080,N_5339);
nor UO_194 (O_194,N_5696,N_7862);
nand UO_195 (O_195,N_5467,N_8804);
nand UO_196 (O_196,N_7109,N_7806);
and UO_197 (O_197,N_7403,N_6453);
nand UO_198 (O_198,N_6106,N_5637);
nor UO_199 (O_199,N_8213,N_6024);
and UO_200 (O_200,N_8910,N_5437);
or UO_201 (O_201,N_8639,N_6745);
nor UO_202 (O_202,N_6122,N_8460);
nand UO_203 (O_203,N_8737,N_6445);
and UO_204 (O_204,N_5280,N_7327);
nand UO_205 (O_205,N_7162,N_7306);
nor UO_206 (O_206,N_5631,N_6996);
nand UO_207 (O_207,N_6960,N_6703);
and UO_208 (O_208,N_7480,N_9297);
nor UO_209 (O_209,N_5517,N_9600);
nand UO_210 (O_210,N_7371,N_9435);
and UO_211 (O_211,N_6171,N_8634);
and UO_212 (O_212,N_6536,N_6080);
and UO_213 (O_213,N_8935,N_6981);
nor UO_214 (O_214,N_5596,N_5362);
nor UO_215 (O_215,N_7842,N_5513);
nor UO_216 (O_216,N_6622,N_5257);
nand UO_217 (O_217,N_6713,N_9377);
nand UO_218 (O_218,N_5167,N_6336);
and UO_219 (O_219,N_7149,N_9563);
nor UO_220 (O_220,N_5432,N_7596);
nand UO_221 (O_221,N_5609,N_7508);
or UO_222 (O_222,N_5419,N_6815);
and UO_223 (O_223,N_9243,N_7962);
nand UO_224 (O_224,N_8268,N_9621);
and UO_225 (O_225,N_7880,N_6541);
and UO_226 (O_226,N_6386,N_8273);
or UO_227 (O_227,N_5625,N_5821);
nand UO_228 (O_228,N_6825,N_7436);
nor UO_229 (O_229,N_8299,N_9004);
and UO_230 (O_230,N_7984,N_6973);
nand UO_231 (O_231,N_5014,N_9064);
and UO_232 (O_232,N_7401,N_8065);
nor UO_233 (O_233,N_6490,N_9030);
and UO_234 (O_234,N_6645,N_5587);
xor UO_235 (O_235,N_6626,N_9308);
nor UO_236 (O_236,N_9893,N_6488);
nor UO_237 (O_237,N_8108,N_7057);
nand UO_238 (O_238,N_7915,N_7142);
or UO_239 (O_239,N_7045,N_7285);
nor UO_240 (O_240,N_7979,N_7370);
or UO_241 (O_241,N_5927,N_7753);
or UO_242 (O_242,N_9258,N_9559);
nand UO_243 (O_243,N_9570,N_6967);
nor UO_244 (O_244,N_9267,N_8176);
or UO_245 (O_245,N_9875,N_5172);
and UO_246 (O_246,N_6092,N_5756);
nor UO_247 (O_247,N_5100,N_5942);
and UO_248 (O_248,N_5782,N_9229);
or UO_249 (O_249,N_6752,N_7851);
nand UO_250 (O_250,N_7037,N_6053);
and UO_251 (O_251,N_6313,N_5506);
or UO_252 (O_252,N_8062,N_5289);
nor UO_253 (O_253,N_5951,N_9387);
or UO_254 (O_254,N_7028,N_6502);
nand UO_255 (O_255,N_9316,N_9187);
and UO_256 (O_256,N_5018,N_9298);
or UO_257 (O_257,N_5036,N_6905);
or UO_258 (O_258,N_5626,N_9985);
nor UO_259 (O_259,N_6864,N_9142);
or UO_260 (O_260,N_5986,N_5554);
nand UO_261 (O_261,N_7900,N_7207);
or UO_262 (O_262,N_7261,N_5351);
or UO_263 (O_263,N_5141,N_5984);
or UO_264 (O_264,N_9131,N_6497);
or UO_265 (O_265,N_7882,N_6314);
nand UO_266 (O_266,N_7342,N_5353);
nand UO_267 (O_267,N_9869,N_9808);
or UO_268 (O_268,N_8294,N_8833);
nand UO_269 (O_269,N_6008,N_5058);
or UO_270 (O_270,N_6749,N_9357);
nor UO_271 (O_271,N_7603,N_9138);
nor UO_272 (O_272,N_5190,N_8295);
nor UO_273 (O_273,N_7731,N_9903);
nor UO_274 (O_274,N_9775,N_8043);
and UO_275 (O_275,N_7488,N_7772);
or UO_276 (O_276,N_6384,N_5468);
or UO_277 (O_277,N_7981,N_8487);
or UO_278 (O_278,N_6887,N_5962);
nand UO_279 (O_279,N_6030,N_8203);
and UO_280 (O_280,N_9799,N_8346);
or UO_281 (O_281,N_9329,N_8312);
nor UO_282 (O_282,N_9324,N_6426);
nor UO_283 (O_283,N_5458,N_6742);
nand UO_284 (O_284,N_9422,N_6663);
nor UO_285 (O_285,N_9159,N_6780);
and UO_286 (O_286,N_8125,N_6456);
nand UO_287 (O_287,N_5064,N_7040);
and UO_288 (O_288,N_6205,N_6025);
nor UO_289 (O_289,N_8478,N_8704);
nor UO_290 (O_290,N_5407,N_6737);
nor UO_291 (O_291,N_6826,N_7079);
or UO_292 (O_292,N_9996,N_7850);
nor UO_293 (O_293,N_8520,N_8090);
nand UO_294 (O_294,N_5538,N_6467);
nand UO_295 (O_295,N_5005,N_6184);
and UO_296 (O_296,N_8366,N_8398);
nor UO_297 (O_297,N_7288,N_7857);
or UO_298 (O_298,N_6948,N_8423);
nand UO_299 (O_299,N_5645,N_7074);
or UO_300 (O_300,N_7902,N_7061);
nand UO_301 (O_301,N_8265,N_8466);
and UO_302 (O_302,N_8054,N_8574);
nand UO_303 (O_303,N_5254,N_8854);
and UO_304 (O_304,N_6448,N_8937);
and UO_305 (O_305,N_9956,N_6309);
or UO_306 (O_306,N_9537,N_5476);
nor UO_307 (O_307,N_8852,N_8516);
or UO_308 (O_308,N_7812,N_8329);
nand UO_309 (O_309,N_5834,N_5043);
or UO_310 (O_310,N_7525,N_6599);
and UO_311 (O_311,N_7796,N_7631);
or UO_312 (O_312,N_5120,N_6332);
nand UO_313 (O_313,N_8496,N_7968);
or UO_314 (O_314,N_9606,N_9719);
or UO_315 (O_315,N_8246,N_8094);
or UO_316 (O_316,N_8228,N_6414);
and UO_317 (O_317,N_6770,N_5227);
nand UO_318 (O_318,N_6447,N_6470);
and UO_319 (O_319,N_5878,N_6292);
nand UO_320 (O_320,N_5305,N_6405);
nor UO_321 (O_321,N_9926,N_9830);
or UO_322 (O_322,N_5971,N_9581);
nand UO_323 (O_323,N_7013,N_6056);
nor UO_324 (O_324,N_8575,N_5035);
and UO_325 (O_325,N_5273,N_9727);
nand UO_326 (O_326,N_6176,N_5777);
and UO_327 (O_327,N_8662,N_9672);
nor UO_328 (O_328,N_6436,N_7785);
nor UO_329 (O_329,N_5099,N_5267);
nand UO_330 (O_330,N_6831,N_6817);
or UO_331 (O_331,N_5290,N_6533);
or UO_332 (O_332,N_9214,N_6229);
and UO_333 (O_333,N_7269,N_5930);
and UO_334 (O_334,N_9041,N_7978);
nand UO_335 (O_335,N_9128,N_7787);
or UO_336 (O_336,N_9747,N_5081);
and UO_337 (O_337,N_7866,N_5868);
nand UO_338 (O_338,N_5886,N_8126);
and UO_339 (O_339,N_7352,N_9381);
or UO_340 (O_340,N_6289,N_7173);
nor UO_341 (O_341,N_5363,N_8671);
nand UO_342 (O_342,N_7728,N_5183);
and UO_343 (O_343,N_6789,N_7808);
or UO_344 (O_344,N_5512,N_6580);
or UO_345 (O_345,N_6643,N_9448);
and UO_346 (O_346,N_7194,N_6363);
or UO_347 (O_347,N_7097,N_6804);
and UO_348 (O_348,N_8619,N_9923);
xnor UO_349 (O_349,N_5956,N_8400);
nor UO_350 (O_350,N_5522,N_6846);
xnor UO_351 (O_351,N_5883,N_7046);
or UO_352 (O_352,N_8624,N_9599);
or UO_353 (O_353,N_5987,N_6692);
nor UO_354 (O_354,N_5384,N_5057);
nand UO_355 (O_355,N_7892,N_5681);
or UO_356 (O_356,N_8506,N_8732);
nor UO_357 (O_357,N_5433,N_8031);
and UO_358 (O_358,N_9698,N_6959);
nand UO_359 (O_359,N_7470,N_6347);
nor UO_360 (O_360,N_8561,N_6458);
nand UO_361 (O_361,N_8413,N_7122);
or UO_362 (O_362,N_8015,N_9446);
nand UO_363 (O_363,N_7552,N_5297);
and UO_364 (O_364,N_9168,N_5083);
nor UO_365 (O_365,N_7295,N_8553);
nor UO_366 (O_366,N_5795,N_5223);
and UO_367 (O_367,N_6682,N_5959);
nor UO_368 (O_368,N_6975,N_5980);
or UO_369 (O_369,N_7896,N_7561);
or UO_370 (O_370,N_7641,N_6767);
nand UO_371 (O_371,N_5357,N_9882);
nor UO_372 (O_372,N_6268,N_5119);
nand UO_373 (O_373,N_5203,N_5770);
or UO_374 (O_374,N_6259,N_6422);
nand UO_375 (O_375,N_6719,N_9282);
nand UO_376 (O_376,N_5196,N_5579);
and UO_377 (O_377,N_8071,N_6330);
and UO_378 (O_378,N_7958,N_9426);
nor UO_379 (O_379,N_5837,N_8940);
and UO_380 (O_380,N_6057,N_6357);
nor UO_381 (O_381,N_7026,N_8904);
and UO_382 (O_382,N_5111,N_7693);
and UO_383 (O_383,N_6796,N_9202);
nand UO_384 (O_384,N_7032,N_6740);
nor UO_385 (O_385,N_7008,N_7651);
or UO_386 (O_386,N_5532,N_7246);
nand UO_387 (O_387,N_5037,N_5844);
nor UO_388 (O_388,N_9080,N_6069);
nand UO_389 (O_389,N_5101,N_5519);
or UO_390 (O_390,N_6808,N_9326);
nand UO_391 (O_391,N_8030,N_8119);
or UO_392 (O_392,N_8422,N_7726);
nor UO_393 (O_393,N_6305,N_5804);
nor UO_394 (O_394,N_8482,N_5368);
nor UO_395 (O_395,N_8061,N_6508);
nand UO_396 (O_396,N_8788,N_8826);
or UO_397 (O_397,N_5185,N_7405);
and UO_398 (O_398,N_8714,N_6923);
and UO_399 (O_399,N_8115,N_6655);
or UO_400 (O_400,N_6418,N_9507);
nand UO_401 (O_401,N_6528,N_5616);
and UO_402 (O_402,N_5440,N_7840);
nor UO_403 (O_403,N_6793,N_6914);
or UO_404 (O_404,N_9190,N_5842);
or UO_405 (O_405,N_5508,N_5354);
nand UO_406 (O_406,N_9710,N_7634);
nand UO_407 (O_407,N_6672,N_9285);
nand UO_408 (O_408,N_7604,N_6810);
nand UO_409 (O_409,N_7937,N_8032);
xor UO_410 (O_410,N_8451,N_8622);
and UO_411 (O_411,N_6193,N_5139);
or UO_412 (O_412,N_7639,N_6899);
or UO_413 (O_413,N_7522,N_9833);
or UO_414 (O_414,N_8118,N_9042);
nand UO_415 (O_415,N_5734,N_7536);
nor UO_416 (O_416,N_7099,N_5471);
and UO_417 (O_417,N_6697,N_7798);
and UO_418 (O_418,N_6530,N_7626);
or UO_419 (O_419,N_8899,N_9575);
nor UO_420 (O_420,N_9449,N_8627);
or UO_421 (O_421,N_9465,N_9850);
or UO_422 (O_422,N_8892,N_6799);
nor UO_423 (O_423,N_9427,N_8961);
or UO_424 (O_424,N_8132,N_8323);
or UO_425 (O_425,N_5992,N_8230);
and UO_426 (O_426,N_8260,N_8873);
nand UO_427 (O_427,N_9912,N_7397);
or UO_428 (O_428,N_5275,N_8686);
and UO_429 (O_429,N_8519,N_8350);
nand UO_430 (O_430,N_5885,N_6577);
nor UO_431 (O_431,N_6895,N_5960);
nand UO_432 (O_432,N_6192,N_9074);
and UO_433 (O_433,N_8977,N_7983);
nor UO_434 (O_434,N_9802,N_7618);
nor UO_435 (O_435,N_5539,N_6801);
and UO_436 (O_436,N_6939,N_7800);
and UO_437 (O_437,N_7826,N_5816);
and UO_438 (O_438,N_8705,N_7302);
or UO_439 (O_439,N_6302,N_6255);
nand UO_440 (O_440,N_5121,N_6464);
or UO_441 (O_441,N_5342,N_6381);
and UO_442 (O_442,N_7438,N_6049);
nand UO_443 (O_443,N_8453,N_6394);
or UO_444 (O_444,N_7518,N_5452);
and UO_445 (O_445,N_5011,N_6961);
nand UO_446 (O_446,N_5288,N_5772);
or UO_447 (O_447,N_9792,N_6310);
or UO_448 (O_448,N_9924,N_5751);
and UO_449 (O_449,N_6773,N_9686);
nor UO_450 (O_450,N_9151,N_7341);
nand UO_451 (O_451,N_8147,N_7055);
and UO_452 (O_452,N_9735,N_6532);
nand UO_453 (O_453,N_9351,N_8544);
and UO_454 (O_454,N_7757,N_6409);
nand UO_455 (O_455,N_7853,N_9275);
and UO_456 (O_456,N_6130,N_8187);
nor UO_457 (O_457,N_5910,N_9091);
nand UO_458 (O_458,N_5877,N_7919);
nand UO_459 (O_459,N_8475,N_7745);
nor UO_460 (O_460,N_9846,N_7537);
nand UO_461 (O_461,N_6641,N_9549);
and UO_462 (O_462,N_8604,N_7116);
and UO_463 (O_463,N_6304,N_7400);
nand UO_464 (O_464,N_9325,N_8184);
and UO_465 (O_465,N_5610,N_6687);
or UO_466 (O_466,N_8643,N_6235);
xor UO_467 (O_467,N_6988,N_6281);
xnor UO_468 (O_468,N_9266,N_7971);
nand UO_469 (O_469,N_8790,N_9911);
xnor UO_470 (O_470,N_5608,N_5168);
and UO_471 (O_471,N_6830,N_7712);
nor UO_472 (O_472,N_6906,N_7895);
and UO_473 (O_473,N_7131,N_7969);
xnor UO_474 (O_474,N_7492,N_7072);
nor UO_475 (O_475,N_8056,N_7058);
nand UO_476 (O_476,N_5446,N_7760);
nand UO_477 (O_477,N_5599,N_8797);
nor UO_478 (O_478,N_9673,N_8293);
and UO_479 (O_479,N_8166,N_5041);
nand UO_480 (O_480,N_9744,N_8959);
nor UO_481 (O_481,N_9796,N_6935);
or UO_482 (O_482,N_9533,N_8847);
nor UO_483 (O_483,N_8074,N_8352);
and UO_484 (O_484,N_5917,N_8226);
nand UO_485 (O_485,N_9482,N_6060);
nand UO_486 (O_486,N_5406,N_8020);
or UO_487 (O_487,N_5248,N_9643);
or UO_488 (O_488,N_6093,N_5118);
nor UO_489 (O_489,N_5828,N_7444);
and UO_490 (O_490,N_7733,N_7923);
or UO_491 (O_491,N_7305,N_9920);
and UO_492 (O_492,N_7062,N_8017);
nor UO_493 (O_493,N_8936,N_8105);
nor UO_494 (O_494,N_6167,N_9340);
and UO_495 (O_495,N_6872,N_8649);
or UO_496 (O_496,N_5469,N_8582);
nor UO_497 (O_497,N_9194,N_7208);
nand UO_498 (O_498,N_7320,N_8036);
xnor UO_499 (O_499,N_6044,N_7916);
or UO_500 (O_500,N_8397,N_6356);
nor UO_501 (O_501,N_8990,N_5997);
and UO_502 (O_502,N_8562,N_7174);
nand UO_503 (O_503,N_6602,N_6311);
or UO_504 (O_504,N_9126,N_6954);
nand UO_505 (O_505,N_8876,N_7524);
nand UO_506 (O_506,N_5536,N_9252);
or UO_507 (O_507,N_6161,N_9445);
and UO_508 (O_508,N_6390,N_8573);
and UO_509 (O_509,N_9781,N_5820);
nand UO_510 (O_510,N_5802,N_5375);
and UO_511 (O_511,N_5263,N_8389);
and UO_512 (O_512,N_9556,N_6708);
nand UO_513 (O_513,N_9213,N_5068);
nor UO_514 (O_514,N_8967,N_7257);
or UO_515 (O_515,N_5749,N_9467);
nand UO_516 (O_516,N_5628,N_7528);
nand UO_517 (O_517,N_8048,N_7933);
nand UO_518 (O_518,N_7725,N_9813);
nand UO_519 (O_519,N_5524,N_8655);
and UO_520 (O_520,N_8896,N_9205);
or UO_521 (O_521,N_8995,N_6834);
nor UO_522 (O_522,N_9253,N_7735);
nand UO_523 (O_523,N_9725,N_5796);
and UO_524 (O_524,N_6527,N_7844);
nor UO_525 (O_525,N_5869,N_7573);
or UO_526 (O_526,N_8808,N_7545);
nand UO_527 (O_527,N_8844,N_9582);
and UO_528 (O_528,N_9815,N_8414);
nand UO_529 (O_529,N_8943,N_6738);
nor UO_530 (O_530,N_7988,N_9822);
or UO_531 (O_531,N_7413,N_5708);
and UO_532 (O_532,N_7974,N_6100);
nand UO_533 (O_533,N_6099,N_6465);
or UO_534 (O_534,N_8376,N_8149);
or UO_535 (O_535,N_7009,N_9626);
or UO_536 (O_536,N_7673,N_7908);
xor UO_537 (O_537,N_6133,N_8616);
nand UO_538 (O_538,N_9690,N_5398);
nand UO_539 (O_539,N_5694,N_9951);
nor UO_540 (O_540,N_9670,N_8975);
or UO_541 (O_541,N_9263,N_5813);
xor UO_542 (O_542,N_5151,N_5660);
xnor UO_543 (O_543,N_5466,N_7332);
and UO_544 (O_544,N_9400,N_5441);
nor UO_545 (O_545,N_8949,N_7911);
nor UO_546 (O_546,N_7945,N_7534);
nor UO_547 (O_547,N_6859,N_8884);
and UO_548 (O_548,N_5994,N_6250);
and UO_549 (O_549,N_9358,N_5028);
nor UO_550 (O_550,N_9906,N_8840);
and UO_551 (O_551,N_5303,N_6896);
nor UO_552 (O_552,N_9651,N_9900);
or UO_553 (O_553,N_7620,N_9341);
or UO_554 (O_554,N_8469,N_9757);
nor UO_555 (O_555,N_5801,N_9478);
nor UO_556 (O_556,N_7318,N_8965);
or UO_557 (O_557,N_9497,N_8614);
nand UO_558 (O_558,N_8631,N_5238);
and UO_559 (O_559,N_7493,N_7133);
or UO_560 (O_560,N_7678,N_5264);
or UO_561 (O_561,N_9644,N_9639);
and UO_562 (O_562,N_6459,N_5779);
nand UO_563 (O_563,N_9012,N_6786);
or UO_564 (O_564,N_5604,N_7498);
nand UO_565 (O_565,N_8689,N_6271);
nor UO_566 (O_566,N_7303,N_8278);
xor UO_567 (O_567,N_6163,N_6217);
nor UO_568 (O_568,N_5655,N_9697);
or UO_569 (O_569,N_8531,N_7237);
nand UO_570 (O_570,N_8359,N_9722);
nand UO_571 (O_571,N_7479,N_9079);
nor UO_572 (O_572,N_5814,N_5691);
nor UO_573 (O_573,N_9070,N_5024);
nor UO_574 (O_574,N_7586,N_5600);
nand UO_575 (O_575,N_7019,N_8204);
nand UO_576 (O_576,N_7343,N_6263);
nand UO_577 (O_577,N_7240,N_9488);
nor UO_578 (O_578,N_7717,N_7991);
nand UO_579 (O_579,N_8645,N_6877);
nand UO_580 (O_580,N_5664,N_9904);
or UO_581 (O_581,N_6681,N_8318);
nand UO_582 (O_582,N_5652,N_7084);
nor UO_583 (O_583,N_8979,N_5651);
nand UO_584 (O_584,N_8779,N_6617);
nand UO_585 (O_585,N_8980,N_6196);
and UO_586 (O_586,N_8374,N_7279);
nand UO_587 (O_587,N_6774,N_7683);
and UO_588 (O_588,N_8933,N_5158);
and UO_589 (O_589,N_7887,N_5090);
nand UO_590 (O_590,N_6408,N_8165);
or UO_591 (O_591,N_5946,N_5445);
and UO_592 (O_592,N_7163,N_9666);
or UO_593 (O_593,N_8872,N_6565);
nand UO_594 (O_594,N_8770,N_7765);
nand UO_595 (O_595,N_7186,N_6698);
or UO_596 (O_596,N_5653,N_7463);
nor UO_597 (O_597,N_7827,N_6254);
nor UO_598 (O_598,N_9442,N_6327);
nor UO_599 (O_599,N_9046,N_7425);
or UO_600 (O_600,N_7266,N_5632);
and UO_601 (O_601,N_6922,N_9492);
and UO_602 (O_602,N_5630,N_5348);
nand UO_603 (O_603,N_8569,N_8670);
and UO_604 (O_604,N_9878,N_8308);
nor UO_605 (O_605,N_8775,N_6998);
nor UO_606 (O_606,N_8838,N_8659);
nand UO_607 (O_607,N_7276,N_6433);
nor UO_608 (O_608,N_6871,N_8971);
or UO_609 (O_609,N_9338,N_6260);
xnor UO_610 (O_610,N_9078,N_9270);
nand UO_611 (O_611,N_9224,N_6632);
and UO_612 (O_612,N_8360,N_6400);
and UO_613 (O_613,N_8491,N_8356);
and UO_614 (O_614,N_6275,N_5097);
nor UO_615 (O_615,N_7749,N_5247);
or UO_616 (O_616,N_8183,N_6563);
nand UO_617 (O_617,N_9832,N_6264);
nand UO_618 (O_618,N_7471,N_9825);
and UO_619 (O_619,N_8730,N_9546);
nand UO_620 (O_620,N_8143,N_7932);
nor UO_621 (O_621,N_5717,N_5333);
nand UO_622 (O_622,N_9230,N_6385);
nand UO_623 (O_623,N_7574,N_9220);
or UO_624 (O_624,N_9980,N_9841);
and UO_625 (O_625,N_9810,N_6757);
nand UO_626 (O_626,N_5125,N_5062);
nand UO_627 (O_627,N_6512,N_6373);
nor UO_628 (O_628,N_9019,N_5936);
and UO_629 (O_629,N_6633,N_6779);
nor UO_630 (O_630,N_8430,N_7675);
nor UO_631 (O_631,N_8757,N_8522);
nor UO_632 (O_632,N_5332,N_5377);
nor UO_633 (O_633,N_8957,N_8976);
or UO_634 (O_634,N_9680,N_5975);
and UO_635 (O_635,N_7655,N_5619);
nor UO_636 (O_636,N_7501,N_5054);
and UO_637 (O_637,N_9288,N_6969);
nand UO_638 (O_638,N_5022,N_7539);
or UO_639 (O_639,N_6296,N_9172);
nor UO_640 (O_640,N_5726,N_6345);
or UO_641 (O_641,N_5415,N_7544);
nand UO_642 (O_642,N_7873,N_5784);
or UO_643 (O_643,N_8155,N_5665);
nand UO_644 (O_644,N_6568,N_7961);
nand UO_645 (O_645,N_6853,N_6838);
or UO_646 (O_646,N_7994,N_7483);
nand UO_647 (O_647,N_7848,N_6968);
or UO_648 (O_648,N_6819,N_7630);
or UO_649 (O_649,N_5338,N_6081);
and UO_650 (O_650,N_6321,N_9597);
nand UO_651 (O_651,N_9838,N_5256);
or UO_652 (O_652,N_6197,N_8490);
nand UO_653 (O_653,N_9048,N_7758);
nor UO_654 (O_654,N_8603,N_6542);
nor UO_655 (O_655,N_6942,N_8620);
and UO_656 (O_656,N_8331,N_9791);
nor UO_657 (O_657,N_5598,N_9286);
nand UO_658 (O_658,N_9591,N_6526);
nor UO_659 (O_659,N_6168,N_6715);
or UO_660 (O_660,N_5891,N_9496);
and UO_661 (O_661,N_9122,N_6913);
and UO_662 (O_662,N_7825,N_9113);
xor UO_663 (O_663,N_6155,N_8684);
or UO_664 (O_664,N_7526,N_9623);
nand UO_665 (O_665,N_8885,N_5765);
or UO_666 (O_666,N_7831,N_8212);
or UO_667 (O_667,N_6104,N_6581);
nand UO_668 (O_668,N_6656,N_5344);
nand UO_669 (O_669,N_6166,N_6972);
nand UO_670 (O_670,N_8698,N_5052);
and UO_671 (O_671,N_8589,N_7653);
or UO_672 (O_672,N_6564,N_6297);
nand UO_673 (O_673,N_5947,N_9768);
nand UO_674 (O_674,N_8313,N_9585);
nor UO_675 (O_675,N_8338,N_9027);
and UO_676 (O_676,N_8966,N_7993);
and UO_677 (O_677,N_9922,N_7296);
nor UO_678 (O_678,N_9118,N_5304);
and UO_679 (O_679,N_6559,N_6951);
xor UO_680 (O_680,N_6829,N_9404);
or UO_681 (O_681,N_7051,N_7907);
or UO_682 (O_682,N_7531,N_7367);
xor UO_683 (O_683,N_8162,N_7689);
nor UO_684 (O_684,N_9595,N_9578);
or UO_685 (O_685,N_8532,N_8505);
nor UO_686 (O_686,N_6837,N_5659);
nand UO_687 (O_687,N_6665,N_9840);
nand UO_688 (O_688,N_9092,N_9317);
nor UO_689 (O_689,N_7225,N_7277);
nand UO_690 (O_690,N_8930,N_5793);
xor UO_691 (O_691,N_6474,N_8501);
nor UO_692 (O_692,N_9762,N_9119);
and UO_693 (O_693,N_5594,N_8419);
and UO_694 (O_694,N_7105,N_9043);
nand UO_695 (O_695,N_8735,N_7495);
nor UO_696 (O_696,N_7967,N_5686);
nand UO_697 (O_697,N_9425,N_6028);
and UO_698 (O_698,N_8001,N_6875);
and UO_699 (O_699,N_8171,N_9629);
or UO_700 (O_700,N_5781,N_5500);
nand UO_701 (O_701,N_9443,N_5487);
nand UO_702 (O_702,N_6503,N_6690);
and UO_703 (O_703,N_9603,N_8635);
nand UO_704 (O_704,N_5939,N_6891);
and UO_705 (O_705,N_6188,N_9501);
and UO_706 (O_706,N_6716,N_8632);
or UO_707 (O_707,N_6210,N_6584);
nor UO_708 (O_708,N_8034,N_8534);
nand UO_709 (O_709,N_5838,N_5218);
and UO_710 (O_710,N_6017,N_9806);
nand UO_711 (O_711,N_6962,N_9315);
nand UO_712 (O_712,N_5970,N_6573);
nand UO_713 (O_713,N_6765,N_8220);
nand UO_714 (O_714,N_7836,N_8354);
and UO_715 (O_715,N_9919,N_5165);
and UO_716 (O_716,N_9067,N_8865);
nor UO_717 (O_717,N_8740,N_7211);
and UO_718 (O_718,N_7838,N_5514);
nand UO_719 (O_719,N_7106,N_6523);
and UO_720 (O_720,N_5427,N_7117);
nor UO_721 (O_721,N_8272,N_6734);
nand UO_722 (O_722,N_6063,N_7369);
and UO_723 (O_723,N_7670,N_9433);
nand UO_724 (O_724,N_5582,N_5996);
and UO_725 (O_725,N_8461,N_9441);
nor UO_726 (O_726,N_7833,N_8136);
or UO_727 (O_727,N_7212,N_7845);
or UO_728 (O_728,N_7179,N_8279);
and UO_729 (O_729,N_5888,N_5545);
and UO_730 (O_730,N_7092,N_6190);
nor UO_731 (O_731,N_6340,N_8650);
or UO_732 (O_732,N_8160,N_7871);
xor UO_733 (O_733,N_8787,N_5301);
and UO_734 (O_734,N_9160,N_9167);
nand UO_735 (O_735,N_6120,N_9618);
and UO_736 (O_736,N_9051,N_7987);
nand UO_737 (O_737,N_9865,N_7054);
nand UO_738 (O_738,N_5093,N_9024);
or UO_739 (O_739,N_6768,N_5807);
or UO_740 (O_740,N_9569,N_5505);
and UO_741 (O_741,N_9010,N_7233);
nand UO_742 (O_742,N_5527,N_5222);
and UO_743 (O_743,N_6164,N_8111);
or UO_744 (O_744,N_9760,N_9772);
and UO_745 (O_745,N_8742,N_7519);
nand UO_746 (O_746,N_9784,N_5450);
and UO_747 (O_747,N_8385,N_9097);
nand UO_748 (O_748,N_8676,N_8938);
nor UO_749 (O_749,N_7298,N_8087);
or UO_750 (O_750,N_8736,N_9876);
and UO_751 (O_751,N_6088,N_5680);
nor UO_752 (O_752,N_9141,N_8098);
or UO_753 (O_753,N_6607,N_8424);
nand UO_754 (O_754,N_9293,N_8889);
nand UO_755 (O_755,N_6521,N_7794);
or UO_756 (O_756,N_9929,N_6156);
or UO_757 (O_757,N_8066,N_8114);
nand UO_758 (O_758,N_6771,N_8618);
or UO_759 (O_759,N_6269,N_7111);
nor UO_760 (O_760,N_6415,N_6109);
or UO_761 (O_761,N_6549,N_7168);
nor UO_762 (O_762,N_9349,N_8968);
or UO_763 (O_763,N_7317,N_9000);
or UO_764 (O_764,N_9455,N_5274);
nor UO_765 (O_765,N_8144,N_6034);
or UO_766 (O_766,N_8628,N_8637);
xnor UO_767 (O_767,N_5924,N_9278);
nor UO_768 (O_768,N_8570,N_6303);
nand UO_769 (O_769,N_7778,N_8382);
nand UO_770 (O_770,N_7464,N_6288);
nand UO_771 (O_771,N_6361,N_9562);
and UO_772 (O_772,N_7152,N_7059);
nor UO_773 (O_773,N_7952,N_8131);
and UO_774 (O_774,N_8392,N_6185);
nor UO_775 (O_775,N_8488,N_9968);
and UO_776 (O_776,N_8718,N_6955);
and UO_777 (O_777,N_7360,N_8759);
nor UO_778 (O_778,N_6699,N_5976);
and UO_779 (O_779,N_7560,N_9257);
nand UO_780 (O_780,N_5135,N_8086);
nor UO_781 (O_781,N_6293,N_6650);
and UO_782 (O_782,N_6696,N_6707);
nor UO_783 (O_783,N_6095,N_6791);
nand UO_784 (O_784,N_5228,N_8431);
nand UO_785 (O_785,N_8191,N_8665);
nor UO_786 (O_786,N_8610,N_9161);
or UO_787 (O_787,N_5941,N_8407);
nor UO_788 (O_788,N_9972,N_7549);
nand UO_789 (O_789,N_7461,N_9758);
or UO_790 (O_790,N_9694,N_6431);
or UO_791 (O_791,N_6865,N_7823);
and UO_792 (O_792,N_6147,N_8508);
and UO_793 (O_793,N_5607,N_5736);
and UO_794 (O_794,N_7336,N_6153);
nand UO_795 (O_795,N_6139,N_6320);
or UO_796 (O_796,N_9251,N_6806);
nor UO_797 (O_797,N_9026,N_9398);
and UO_798 (O_798,N_9828,N_6720);
or UO_799 (O_799,N_9095,N_7874);
and UO_800 (O_800,N_7112,N_7432);
nor UO_801 (O_801,N_8941,N_5864);
and UO_802 (O_802,N_8560,N_7351);
nor UO_803 (O_803,N_6026,N_5810);
nor UO_804 (O_804,N_8800,N_8626);
nor UO_805 (O_805,N_9233,N_7132);
or UO_806 (O_806,N_5573,N_6284);
nand UO_807 (O_807,N_9346,N_9598);
and UO_808 (O_808,N_9765,N_6131);
or UO_809 (O_809,N_8444,N_9111);
nand UO_810 (O_810,N_8669,N_5138);
nor UO_811 (O_811,N_9487,N_6818);
or UO_812 (O_812,N_9959,N_5109);
and UO_813 (O_813,N_5715,N_7629);
nand UO_814 (O_814,N_8934,N_5161);
nor UO_815 (O_815,N_8906,N_8994);
and UO_816 (O_816,N_9682,N_5998);
and UO_817 (O_817,N_7156,N_7482);
and UO_818 (O_818,N_6930,N_9659);
and UO_819 (O_819,N_6403,N_9883);
or UO_820 (O_820,N_7801,N_7682);
nand UO_821 (O_821,N_6322,N_6477);
and UO_822 (O_822,N_9154,N_7243);
nor UO_823 (O_823,N_7898,N_7182);
nand UO_824 (O_824,N_9343,N_8638);
and UO_825 (O_825,N_7665,N_6035);
nor UO_826 (O_826,N_7643,N_5758);
nand UO_827 (O_827,N_7067,N_5116);
or UO_828 (O_828,N_5739,N_8551);
and UO_829 (O_829,N_5954,N_7698);
nor UO_830 (O_830,N_7736,N_8761);
or UO_831 (O_831,N_7893,N_6539);
nor UO_832 (O_832,N_8386,N_5938);
and UO_833 (O_833,N_9509,N_5473);
or UO_834 (O_834,N_5892,N_5968);
nand UO_835 (O_835,N_5874,N_8660);
nand UO_836 (O_836,N_6073,N_9683);
nand UO_837 (O_837,N_7542,N_8509);
nand UO_838 (O_838,N_6267,N_5848);
nor UO_839 (O_839,N_5345,N_7366);
nor UO_840 (O_840,N_9889,N_8984);
or UO_841 (O_841,N_7478,N_8450);
and UO_842 (O_842,N_5311,N_7910);
nor UO_843 (O_843,N_8477,N_7280);
nor UO_844 (O_844,N_9268,N_7139);
nor UO_845 (O_845,N_9388,N_8050);
or UO_846 (O_846,N_9292,N_9879);
and UO_847 (O_847,N_7252,N_7870);
and UO_848 (O_848,N_5008,N_5242);
or UO_849 (O_849,N_7607,N_9705);
or UO_850 (O_850,N_9524,N_7023);
nand UO_851 (O_851,N_8712,N_5791);
or UO_852 (O_852,N_7533,N_7672);
or UO_853 (O_853,N_9206,N_7220);
and UO_854 (O_854,N_8138,N_8245);
nor UO_855 (O_855,N_7849,N_7021);
nand UO_856 (O_856,N_6338,N_6583);
nand UO_857 (O_857,N_7330,N_7816);
nor UO_858 (O_858,N_7783,N_7547);
nand UO_859 (O_859,N_9880,N_6300);
nand UO_860 (O_860,N_9307,N_9998);
and UO_861 (O_861,N_7829,N_6840);
nor UO_862 (O_862,N_6134,N_9824);
or UO_863 (O_863,N_5673,N_7503);
nand UO_864 (O_864,N_5217,N_7741);
nand UO_865 (O_865,N_7235,N_9976);
or UO_866 (O_866,N_7711,N_9246);
or UO_867 (O_867,N_5644,N_7344);
or UO_868 (O_868,N_9851,N_5150);
nand UO_869 (O_869,N_8355,N_5034);
nand UO_870 (O_870,N_5916,N_8037);
nand UO_871 (O_871,N_8903,N_5943);
nor UO_872 (O_872,N_6884,N_5572);
nor UO_873 (O_873,N_7222,N_7083);
or UO_874 (O_874,N_9941,N_9459);
or UO_875 (O_875,N_8690,N_7391);
or UO_876 (O_876,N_7805,N_5858);
nor UO_877 (O_877,N_8076,N_9527);
or UO_878 (O_878,N_9635,N_7597);
and UO_879 (O_879,N_6516,N_7647);
or UO_880 (O_880,N_5509,N_8394);
and UO_881 (O_881,N_9320,N_6222);
and UO_882 (O_882,N_7018,N_7710);
or UO_883 (O_883,N_7375,N_7752);
and UO_884 (O_884,N_8850,N_6727);
and UO_885 (O_885,N_8549,N_8327);
nand UO_886 (O_886,N_9676,N_7196);
nand UO_887 (O_887,N_6937,N_5031);
and UO_888 (O_888,N_9513,N_8492);
nor UO_889 (O_889,N_8749,N_6387);
and UO_890 (O_890,N_7918,N_7746);
nand UO_891 (O_891,N_7602,N_7797);
or UO_892 (O_892,N_9695,N_8525);
nand UO_893 (O_893,N_9661,N_5173);
or UO_894 (O_894,N_6653,N_6441);
and UO_895 (O_895,N_5763,N_9269);
and UO_896 (O_896,N_9380,N_9729);
nor UO_897 (O_897,N_6172,N_8606);
and UO_898 (O_898,N_9290,N_8674);
nor UO_899 (O_899,N_9402,N_7080);
and UO_900 (O_900,N_7761,N_6111);
and UO_901 (O_901,N_6613,N_9181);
nor UO_902 (O_902,N_8880,N_7500);
nand UO_903 (O_903,N_7414,N_5201);
and UO_904 (O_904,N_5488,N_7591);
nor UO_905 (O_905,N_7229,N_5258);
or UO_906 (O_906,N_9786,N_9306);
nand UO_907 (O_907,N_8498,N_5692);
or UO_908 (O_908,N_8276,N_6256);
and UO_909 (O_909,N_7964,N_9521);
or UO_910 (O_910,N_8500,N_6811);
and UO_911 (O_911,N_9891,N_9712);
or UO_912 (O_912,N_7609,N_9238);
and UO_913 (O_913,N_9184,N_7025);
or UO_914 (O_914,N_9460,N_6232);
nor UO_915 (O_915,N_5563,N_5965);
nand UO_916 (O_916,N_6160,N_6212);
nor UO_917 (O_917,N_7068,N_9536);
nand UO_918 (O_918,N_7205,N_8504);
nand UO_919 (O_919,N_5292,N_7204);
nor UO_920 (O_920,N_8821,N_5343);
nand UO_921 (O_921,N_6636,N_7906);
and UO_922 (O_922,N_8241,N_8540);
xnor UO_923 (O_923,N_6325,N_8343);
nor UO_924 (O_924,N_5683,N_7451);
and UO_925 (O_925,N_5709,N_9755);
and UO_926 (O_926,N_7433,N_6116);
or UO_927 (O_927,N_5170,N_6186);
nor UO_928 (O_928,N_7600,N_6755);
or UO_929 (O_929,N_6620,N_9189);
or UO_930 (O_930,N_9087,N_5486);
nor UO_931 (O_931,N_5900,N_5603);
or UO_932 (O_932,N_6732,N_8981);
and UO_933 (O_933,N_5088,N_8564);
nor UO_934 (O_934,N_9646,N_9872);
nor UO_935 (O_935,N_8378,N_9210);
or UO_936 (O_936,N_8652,N_5329);
or UO_937 (O_937,N_8530,N_7048);
or UO_938 (O_938,N_6949,N_6522);
nand UO_939 (O_939,N_9471,N_5340);
nand UO_940 (O_940,N_9372,N_5746);
nor UO_941 (O_941,N_9280,N_9518);
nand UO_942 (O_942,N_7348,N_7638);
nor UO_943 (O_943,N_5764,N_6711);
and UO_944 (O_944,N_7262,N_5672);
xnor UO_945 (O_945,N_8240,N_7066);
and UO_946 (O_946,N_9688,N_7361);
nand UO_947 (O_947,N_9589,N_9374);
or UO_948 (O_948,N_9135,N_8843);
and UO_949 (O_949,N_6615,N_8219);
nor UO_950 (O_950,N_9215,N_8898);
and UO_951 (O_951,N_6455,N_7663);
or UO_952 (O_952,N_6710,N_9818);
xnor UO_953 (O_953,N_8862,N_6987);
nand UO_954 (O_954,N_8657,N_5757);
nand UO_955 (O_955,N_8777,N_7739);
nor UO_956 (O_956,N_5009,N_8210);
and UO_957 (O_957,N_7210,N_9032);
xor UO_958 (O_958,N_7217,N_9271);
nand UO_959 (O_959,N_7818,N_6039);
nor UO_960 (O_960,N_9669,N_8887);
xor UO_961 (O_961,N_8471,N_7115);
nor UO_962 (O_962,N_9287,N_9742);
nand UO_963 (O_963,N_6798,N_9774);
and UO_964 (O_964,N_7636,N_8612);
and UO_965 (O_965,N_6117,N_5380);
nor UO_966 (O_966,N_5658,N_8728);
or UO_967 (O_967,N_9842,N_8909);
and UO_968 (O_968,N_6496,N_7562);
or UO_969 (O_969,N_5895,N_8455);
or UO_970 (O_970,N_9208,N_5039);
nor UO_971 (O_971,N_7250,N_7384);
nor UO_972 (O_972,N_9177,N_7044);
nor UO_973 (O_973,N_8257,N_8102);
and UO_974 (O_974,N_9974,N_8449);
and UO_975 (O_975,N_8215,N_5591);
xnor UO_976 (O_976,N_6971,N_5360);
and UO_977 (O_977,N_8701,N_8145);
nor UO_978 (O_978,N_9130,N_8112);
nand UO_979 (O_979,N_6612,N_7124);
nor UO_980 (O_980,N_8914,N_5786);
nor UO_981 (O_981,N_7155,N_6919);
nand UO_982 (O_982,N_7720,N_5620);
or UO_983 (O_983,N_9962,N_7416);
and UO_984 (O_984,N_7095,N_8550);
and UO_985 (O_985,N_8584,N_5382);
nand UO_986 (O_986,N_6501,N_5207);
or UO_987 (O_987,N_7402,N_7270);
or UO_988 (O_988,N_6870,N_5533);
nor UO_989 (O_989,N_9318,N_7056);
and UO_990 (O_990,N_6010,N_6912);
nor UO_991 (O_991,N_7082,N_7516);
nand UO_992 (O_992,N_7338,N_9835);
nand UO_993 (O_993,N_9453,N_9740);
nand UO_994 (O_994,N_7325,N_8193);
and UO_995 (O_995,N_6561,N_8699);
and UO_996 (O_996,N_9337,N_5701);
xnor UO_997 (O_997,N_5326,N_5318);
or UO_998 (O_998,N_5730,N_8412);
and UO_999 (O_999,N_9276,N_6344);
nand UO_1000 (O_1000,N_5281,N_8806);
nor UO_1001 (O_1001,N_5178,N_6372);
and UO_1002 (O_1002,N_6005,N_9444);
or UO_1003 (O_1003,N_5646,N_6892);
or UO_1004 (O_1004,N_9711,N_5972);
or UO_1005 (O_1005,N_9432,N_5239);
and UO_1006 (O_1006,N_8988,N_8045);
and UO_1007 (O_1007,N_7588,N_7697);
xnor UO_1008 (O_1008,N_6097,N_8672);
nand UO_1009 (O_1009,N_8253,N_8303);
or UO_1010 (O_1010,N_5078,N_9245);
nand UO_1011 (O_1011,N_7506,N_7128);
nand UO_1012 (O_1012,N_9573,N_6351);
or UO_1013 (O_1013,N_5220,N_6587);
nor UO_1014 (O_1014,N_5277,N_5226);
and UO_1015 (O_1015,N_9662,N_5470);
xor UO_1016 (O_1016,N_7570,N_9035);
nand UO_1017 (O_1017,N_9530,N_9510);
nor UO_1018 (O_1018,N_8837,N_9369);
and UO_1019 (O_1019,N_5497,N_9763);
or UO_1020 (O_1020,N_5265,N_5046);
or UO_1021 (O_1021,N_9093,N_8028);
and UO_1022 (O_1022,N_8766,N_8703);
or UO_1023 (O_1023,N_8602,N_9811);
and UO_1024 (O_1024,N_9704,N_6883);
and UO_1025 (O_1025,N_6880,N_5835);
and UO_1026 (O_1026,N_8836,N_9845);
xor UO_1027 (O_1027,N_7732,N_5839);
xor UO_1028 (O_1028,N_9472,N_9905);
and UO_1029 (O_1029,N_6023,N_8950);
nor UO_1030 (O_1030,N_8986,N_9466);
nor UO_1031 (O_1031,N_6683,N_7865);
and UO_1032 (O_1032,N_5833,N_8794);
or UO_1033 (O_1033,N_7226,N_5202);
nand UO_1034 (O_1034,N_9386,N_7388);
or UO_1035 (O_1035,N_8387,N_6894);
nand UO_1036 (O_1036,N_6813,N_5224);
and UO_1037 (O_1037,N_7936,N_6421);
nor UO_1038 (O_1038,N_6667,N_9470);
and UO_1039 (O_1039,N_7170,N_9073);
and UO_1040 (O_1040,N_7889,N_5283);
nand UO_1041 (O_1041,N_5944,N_5707);
and UO_1042 (O_1042,N_7101,N_8003);
nor UO_1043 (O_1043,N_8881,N_5381);
nand UO_1044 (O_1044,N_7439,N_8280);
nand UO_1045 (O_1045,N_6616,N_5372);
xor UO_1046 (O_1046,N_9925,N_7815);
nor UO_1047 (O_1047,N_6110,N_8194);
or UO_1048 (O_1048,N_8016,N_6157);
nor UO_1049 (O_1049,N_6001,N_5932);
nand UO_1050 (O_1050,N_7657,N_7497);
nand UO_1051 (O_1051,N_8815,N_8554);
and UO_1052 (O_1052,N_9008,N_5105);
nand UO_1053 (O_1053,N_5564,N_7704);
or UO_1054 (O_1054,N_5142,N_8809);
nand UO_1055 (O_1055,N_8064,N_9913);
nand UO_1056 (O_1056,N_6893,N_9770);
nand UO_1057 (O_1057,N_6795,N_9103);
nor UO_1058 (O_1058,N_5811,N_5038);
nand UO_1059 (O_1059,N_6146,N_8696);
and UO_1060 (O_1060,N_5993,N_8900);
nand UO_1061 (O_1061,N_5518,N_9935);
nand UO_1062 (O_1062,N_7819,N_9173);
nand UO_1063 (O_1063,N_9612,N_5492);
nor UO_1064 (O_1064,N_6223,N_8234);
nand UO_1065 (O_1065,N_5634,N_8636);
nor UO_1066 (O_1066,N_8109,N_9899);
and UO_1067 (O_1067,N_5087,N_8420);
nor UO_1068 (O_1068,N_5738,N_5583);
nand UO_1069 (O_1069,N_9107,N_6700);
and UO_1070 (O_1070,N_6601,N_8345);
nand UO_1071 (O_1071,N_6927,N_9885);
nor UO_1072 (O_1072,N_6823,N_6614);
and UO_1073 (O_1073,N_9330,N_8348);
nor UO_1074 (O_1074,N_8306,N_6369);
or UO_1075 (O_1075,N_7939,N_5732);
nand UO_1076 (O_1076,N_7690,N_5180);
or UO_1077 (O_1077,N_7090,N_8188);
and UO_1078 (O_1078,N_6295,N_5531);
nand UO_1079 (O_1079,N_8926,N_8404);
nand UO_1080 (O_1080,N_8128,N_8524);
nor UO_1081 (O_1081,N_9715,N_6965);
nor UO_1082 (O_1082,N_7820,N_8106);
or UO_1083 (O_1083,N_6659,N_8956);
and UO_1084 (O_1084,N_9809,N_7992);
or UO_1085 (O_1085,N_7773,N_7195);
or UO_1086 (O_1086,N_6807,N_9493);
nor UO_1087 (O_1087,N_9608,N_5188);
nand UO_1088 (O_1088,N_6493,N_9724);
nand UO_1089 (O_1089,N_8535,N_7038);
or UO_1090 (O_1090,N_5327,N_6729);
nand UO_1091 (O_1091,N_8290,N_8722);
nor UO_1092 (O_1092,N_7373,N_8334);
nor UO_1093 (O_1093,N_8731,N_7022);
nor UO_1094 (O_1094,N_7466,N_8653);
nor UO_1095 (O_1095,N_5767,N_9014);
nand UO_1096 (O_1096,N_8772,N_8982);
nor UO_1097 (O_1097,N_8538,N_8452);
nor UO_1098 (O_1098,N_8605,N_6417);
or UO_1099 (O_1099,N_8608,N_8201);
or UO_1100 (O_1100,N_5144,N_8101);
and UO_1101 (O_1101,N_7869,N_6668);
or UO_1102 (O_1102,N_6346,N_7606);
nor UO_1103 (O_1103,N_5047,N_7383);
nand UO_1104 (O_1104,N_9239,N_7180);
nand UO_1105 (O_1105,N_5159,N_6245);
nor UO_1106 (O_1106,N_8739,N_7947);
nand UO_1107 (O_1107,N_9689,N_8206);
nand UO_1108 (O_1108,N_6121,N_9390);
nand UO_1109 (O_1109,N_7517,N_9999);
nor UO_1110 (O_1110,N_6007,N_5324);
nand UO_1111 (O_1111,N_5952,N_5661);
xnor UO_1112 (O_1112,N_6071,N_5021);
nand UO_1113 (O_1113,N_6142,N_7185);
nor UO_1114 (O_1114,N_7627,N_6941);
or UO_1115 (O_1115,N_5723,N_7510);
nor UO_1116 (O_1116,N_5229,N_5654);
xnor UO_1117 (O_1117,N_6596,N_5102);
nand UO_1118 (O_1118,N_9897,N_8078);
or UO_1119 (O_1119,N_9144,N_6413);
nand UO_1120 (O_1120,N_8768,N_6238);
or UO_1121 (O_1121,N_5568,N_9514);
or UO_1122 (O_1122,N_9706,N_5325);
or UO_1123 (O_1123,N_5560,N_5958);
nand UO_1124 (O_1124,N_5666,N_8039);
or UO_1125 (O_1125,N_7119,N_5671);
or UO_1126 (O_1126,N_9156,N_8099);
or UO_1127 (O_1127,N_5016,N_9650);
nand UO_1128 (O_1128,N_9708,N_9481);
and UO_1129 (O_1129,N_6228,N_6860);
nor UO_1130 (O_1130,N_5576,N_9058);
nor UO_1131 (O_1131,N_9619,N_9641);
and UO_1132 (O_1132,N_9461,N_5435);
or UO_1133 (O_1133,N_9104,N_6982);
and UO_1134 (O_1134,N_6651,N_8515);
nand UO_1135 (O_1135,N_6680,N_5722);
nor UO_1136 (O_1136,N_6515,N_8513);
or UO_1137 (O_1137,N_5846,N_5881);
or UO_1138 (O_1138,N_8186,N_8271);
or UO_1139 (O_1139,N_6209,N_8545);
or UO_1140 (O_1140,N_5194,N_9785);
nor UO_1141 (O_1141,N_5056,N_8285);
or UO_1142 (O_1142,N_5443,N_6963);
and UO_1143 (O_1143,N_7985,N_8576);
or UO_1144 (O_1144,N_8648,N_5094);
and UO_1145 (O_1145,N_8457,N_6835);
or UO_1146 (O_1146,N_9469,N_7039);
xor UO_1147 (O_1147,N_5480,N_6075);
or UO_1148 (O_1148,N_7454,N_9023);
and UO_1149 (O_1149,N_7263,N_7353);
or UO_1150 (O_1150,N_6316,N_8773);
and UO_1151 (O_1151,N_7580,N_9776);
nand UO_1152 (O_1152,N_7120,N_9003);
and UO_1153 (O_1153,N_8537,N_6301);
nor UO_1154 (O_1154,N_8256,N_7468);
or UO_1155 (O_1155,N_7004,N_5743);
or UO_1156 (O_1156,N_5439,N_7372);
nor UO_1157 (O_1157,N_9709,N_8454);
and UO_1158 (O_1158,N_8752,N_6180);
or UO_1159 (O_1159,N_9731,N_9169);
nor UO_1160 (O_1160,N_8081,N_8262);
nor UO_1161 (O_1161,N_5983,N_8146);
nor UO_1162 (O_1162,N_9702,N_7006);
nor UO_1163 (O_1163,N_7948,N_6903);
nor UO_1164 (O_1164,N_8587,N_7033);
and UO_1165 (O_1165,N_5177,N_8107);
nor UO_1166 (O_1166,N_6328,N_5060);
nand UO_1167 (O_1167,N_7424,N_9367);
nand UO_1168 (O_1168,N_8196,N_6814);
and UO_1169 (O_1169,N_5748,N_5851);
and UO_1170 (O_1170,N_9494,N_5189);
nand UO_1171 (O_1171,N_8823,N_8819);
nor UO_1172 (O_1172,N_6423,N_6395);
nor UO_1173 (O_1173,N_7378,N_8964);
nand UO_1174 (O_1174,N_5949,N_8336);
nand UO_1175 (O_1175,N_7997,N_6944);
or UO_1176 (O_1176,N_5935,N_5233);
nand UO_1177 (O_1177,N_8408,N_9451);
nor UO_1178 (O_1178,N_7934,N_9490);
and UO_1179 (O_1179,N_8987,N_9291);
nor UO_1180 (O_1180,N_6510,N_6635);
nand UO_1181 (O_1181,N_6126,N_7409);
and UO_1182 (O_1182,N_8164,N_7010);
or UO_1183 (O_1183,N_6429,N_9795);
or UO_1184 (O_1184,N_6647,N_5698);
nor UO_1185 (O_1185,N_9655,N_9940);
or UO_1186 (O_1186,N_9028,N_5298);
nor UO_1187 (O_1187,N_8395,N_5725);
or UO_1188 (O_1188,N_5523,N_7091);
xor UO_1189 (O_1189,N_6828,N_6000);
nor UO_1190 (O_1190,N_6547,N_7434);
and UO_1191 (O_1191,N_6112,N_8300);
or UO_1192 (O_1192,N_7292,N_7727);
or UO_1193 (O_1193,N_6525,N_6676);
or UO_1194 (O_1194,N_8782,N_9587);
xor UO_1195 (O_1195,N_9328,N_5800);
nor UO_1196 (O_1196,N_9430,N_9016);
nor UO_1197 (O_1197,N_8929,N_6558);
xor UO_1198 (O_1198,N_9485,N_8180);
nor UO_1199 (O_1199,N_6298,N_9590);
or UO_1200 (O_1200,N_9327,N_8247);
nor UO_1201 (O_1201,N_8292,N_7283);
and UO_1202 (O_1202,N_7659,N_6401);
nand UO_1203 (O_1203,N_8991,N_7514);
nor UO_1204 (O_1204,N_5567,N_9938);
or UO_1205 (O_1205,N_5436,N_5685);
nand UO_1206 (O_1206,N_8617,N_5551);
nand UO_1207 (O_1207,N_6195,N_7548);
nand UO_1208 (O_1208,N_5465,N_5291);
nand UO_1209 (O_1209,N_6040,N_6076);
or UO_1210 (O_1210,N_9347,N_8489);
or UO_1211 (O_1211,N_8673,N_7428);
or UO_1212 (O_1212,N_8027,N_8568);
and UO_1213 (O_1213,N_9805,N_6640);
or UO_1214 (O_1214,N_5920,N_6425);
nand UO_1215 (O_1215,N_8362,N_8820);
nor UO_1216 (O_1216,N_5915,N_8858);
or UO_1217 (O_1217,N_8024,N_7718);
and UO_1218 (O_1218,N_9294,N_6047);
nand UO_1219 (O_1219,N_6440,N_5114);
nor UO_1220 (O_1220,N_7209,N_9801);
and UO_1221 (O_1221,N_7191,N_9873);
and UO_1222 (O_1222,N_8511,N_5098);
nand UO_1223 (O_1223,N_9864,N_8783);
nand UO_1224 (O_1224,N_9013,N_9186);
and UO_1225 (O_1225,N_5163,N_8156);
nand UO_1226 (O_1226,N_7148,N_5627);
and UO_1227 (O_1227,N_9534,N_8391);
or UO_1228 (O_1228,N_8548,N_6976);
nand UO_1229 (O_1229,N_5982,N_7652);
and UO_1230 (O_1230,N_6354,N_7917);
or UO_1231 (O_1231,N_9767,N_9299);
nand UO_1232 (O_1232,N_8680,N_7380);
or UO_1233 (O_1233,N_5361,N_9480);
nor UO_1234 (O_1234,N_6484,N_7914);
and UO_1235 (O_1235,N_5507,N_7688);
or UO_1236 (O_1236,N_9544,N_6608);
or UO_1237 (O_1237,N_8908,N_5588);
and UO_1238 (O_1238,N_8022,N_6677);
and UO_1239 (O_1239,N_6115,N_5219);
nand UO_1240 (O_1240,N_6658,N_5879);
nand UO_1241 (O_1241,N_5783,N_6592);
and UO_1242 (O_1242,N_6802,N_7830);
and UO_1243 (O_1243,N_7662,N_6994);
or UO_1244 (O_1244,N_9790,N_8586);
and UO_1245 (O_1245,N_7781,N_6900);
and UO_1246 (O_1246,N_6534,N_7476);
nor UO_1247 (O_1247,N_6609,N_9726);
nand UO_1248 (O_1248,N_9649,N_9056);
or UO_1249 (O_1249,N_7855,N_8281);
and UO_1250 (O_1250,N_9611,N_9406);
nand UO_1251 (O_1251,N_9040,N_7249);
and UO_1252 (O_1252,N_9971,N_7355);
or UO_1253 (O_1253,N_6885,N_7563);
nor UO_1254 (O_1254,N_9505,N_6243);
or UO_1255 (O_1255,N_5373,N_6701);
and UO_1256 (O_1256,N_9105,N_5317);
or UO_1257 (O_1257,N_7779,N_7839);
and UO_1258 (O_1258,N_8566,N_9783);
nand UO_1259 (O_1259,N_9015,N_6428);
nor UO_1260 (O_1260,N_5526,N_5413);
nand UO_1261 (O_1261,N_7624,N_5252);
nand UO_1262 (O_1262,N_5328,N_6391);
nand UO_1263 (O_1263,N_6709,N_6598);
and UO_1264 (O_1264,N_5330,N_7273);
nand UO_1265 (O_1265,N_8853,N_7005);
nor UO_1266 (O_1266,N_9029,N_7184);
nor UO_1267 (O_1267,N_9613,N_8713);
or UO_1268 (O_1268,N_7714,N_8641);
and UO_1269 (O_1269,N_9089,N_5824);
nand UO_1270 (O_1270,N_9360,N_6335);
nor UO_1271 (O_1271,N_9894,N_5000);
nand UO_1272 (O_1272,N_7668,N_8296);
or UO_1273 (O_1273,N_6569,N_7396);
nor UO_1274 (O_1274,N_9385,N_5428);
nor UO_1275 (O_1275,N_9523,N_8266);
and UO_1276 (O_1276,N_5308,N_8150);
nand UO_1277 (O_1277,N_9225,N_6787);
or UO_1278 (O_1278,N_7617,N_7960);
or UO_1279 (O_1279,N_5019,N_9858);
or UO_1280 (O_1280,N_9633,N_7515);
nor UO_1281 (O_1281,N_9918,N_6520);
and UO_1282 (O_1282,N_6038,N_5048);
nand UO_1283 (O_1283,N_7146,N_5369);
nor UO_1284 (O_1284,N_9632,N_9652);
nand UO_1285 (O_1285,N_6621,N_9766);
and UO_1286 (O_1286,N_6132,N_8647);
nor UO_1287 (O_1287,N_6833,N_9975);
xnor UO_1288 (O_1288,N_9289,N_9332);
or UO_1289 (O_1289,N_8518,N_6956);
nor UO_1290 (O_1290,N_7354,N_7709);
and UO_1291 (O_1291,N_9748,N_6135);
nand UO_1292 (O_1292,N_9483,N_8734);
or UO_1293 (O_1293,N_7611,N_6557);
and UO_1294 (O_1294,N_5015,N_5299);
and UO_1295 (O_1295,N_6794,N_7481);
or UO_1296 (O_1296,N_5541,N_9789);
and UO_1297 (O_1297,N_6002,N_7740);
or UO_1298 (O_1298,N_8446,N_6378);
nor UO_1299 (O_1299,N_5401,N_7943);
and UO_1300 (O_1300,N_9703,N_6273);
nand UO_1301 (O_1301,N_6137,N_9231);
and UO_1302 (O_1302,N_8683,N_9631);
nor UO_1303 (O_1303,N_5830,N_8972);
xnor UO_1304 (O_1304,N_8646,N_9241);
nor UO_1305 (O_1305,N_5908,N_5383);
and UO_1306 (O_1306,N_7494,N_8401);
nand UO_1307 (O_1307,N_8697,N_5160);
and UO_1308 (O_1308,N_5245,N_5501);
nor UO_1309 (O_1309,N_8494,N_9987);
or UO_1310 (O_1310,N_8380,N_5129);
nor UO_1311 (O_1311,N_6518,N_5912);
nor UO_1312 (O_1312,N_9397,N_5933);
nand UO_1313 (O_1313,N_9714,N_6866);
nand UO_1314 (O_1314,N_5146,N_6943);
xor UO_1315 (O_1315,N_5832,N_6187);
or UO_1316 (O_1316,N_5418,N_9350);
nor UO_1317 (O_1317,N_9586,N_5829);
and UO_1318 (O_1318,N_8827,N_9196);
nor UO_1319 (O_1319,N_6411,N_5902);
nor UO_1320 (O_1320,N_9814,N_7282);
nand UO_1321 (O_1321,N_9486,N_5461);
and UO_1322 (O_1322,N_6362,N_7154);
nor UO_1323 (O_1323,N_6674,N_8539);
nor UO_1324 (O_1324,N_6619,N_7695);
and UO_1325 (O_1325,N_8583,N_8784);
nor UO_1326 (O_1326,N_6279,N_9431);
nand UO_1327 (O_1327,N_8816,N_6241);
or UO_1328 (O_1328,N_8014,N_5668);
or UO_1329 (O_1329,N_8510,N_6989);
and UO_1330 (O_1330,N_8693,N_7455);
nor UO_1331 (O_1331,N_9491,N_9166);
nand UO_1332 (O_1332,N_9561,N_9856);
or UO_1333 (O_1333,N_6517,N_8578);
or UO_1334 (O_1334,N_6495,N_6036);
nand UO_1335 (O_1335,N_7587,N_8556);
and UO_1336 (O_1336,N_6094,N_7809);
nor UO_1337 (O_1337,N_8916,N_9979);
or UO_1338 (O_1338,N_9995,N_7529);
and UO_1339 (O_1339,N_5371,N_5778);
nand UO_1340 (O_1340,N_5341,N_6777);
or UO_1341 (O_1341,N_9888,N_8223);
and UO_1342 (O_1342,N_7799,N_9520);
and UO_1343 (O_1343,N_7706,N_5385);
nor UO_1344 (O_1344,N_6918,N_9699);
nand UO_1345 (O_1345,N_9528,N_6723);
or UO_1346 (O_1346,N_8688,N_5540);
nand UO_1347 (O_1347,N_9219,N_7440);
and UO_1348 (O_1348,N_9232,N_5741);
nor UO_1349 (O_1349,N_6857,N_6468);
and UO_1350 (O_1350,N_7275,N_7075);
or UO_1351 (O_1351,N_7475,N_5421);
and UO_1352 (O_1352,N_6725,N_7614);
nor UO_1353 (O_1353,N_6631,N_9862);
xor UO_1354 (O_1354,N_8053,N_7272);
or UO_1355 (O_1355,N_5358,N_9474);
nor UO_1356 (O_1356,N_9868,N_6848);
nand UO_1357 (O_1357,N_8985,N_5639);
and UO_1358 (O_1358,N_9005,N_6566);
and UO_1359 (O_1359,N_9384,N_9601);
or UO_1360 (O_1360,N_5797,N_8868);
nor UO_1361 (O_1361,N_5967,N_5199);
or UO_1362 (O_1362,N_9525,N_8579);
or UO_1363 (O_1363,N_7043,N_9022);
or UO_1364 (O_1364,N_6003,N_8667);
nor UO_1365 (O_1365,N_8117,N_9477);
or UO_1366 (O_1366,N_8127,N_8497);
nor UO_1367 (O_1367,N_7847,N_6540);
nor UO_1368 (O_1368,N_8480,N_9218);
nand UO_1369 (O_1369,N_5287,N_8410);
nand UO_1370 (O_1370,N_5918,N_9532);
or UO_1371 (O_1371,N_9197,N_9817);
and UO_1372 (O_1372,N_6578,N_8282);
nor UO_1373 (O_1373,N_5464,N_9011);
nor UO_1374 (O_1374,N_7828,N_7955);
and UO_1375 (O_1375,N_5622,N_5769);
nand UO_1376 (O_1376,N_9937,N_5259);
or UO_1377 (O_1377,N_9741,N_5695);
and UO_1378 (O_1378,N_5866,N_5511);
nor UO_1379 (O_1379,N_9778,N_5074);
and UO_1380 (O_1380,N_7976,N_5774);
and UO_1381 (O_1381,N_6140,N_6852);
nor UO_1382 (O_1382,N_6473,N_7221);
nand UO_1383 (O_1383,N_5313,N_8486);
nand UO_1384 (O_1384,N_7579,N_9099);
and UO_1385 (O_1385,N_7610,N_8088);
xor UO_1386 (O_1386,N_9574,N_6760);
and UO_1387 (O_1387,N_7681,N_7861);
and UO_1388 (O_1388,N_9679,N_6451);
nor UO_1389 (O_1389,N_6443,N_9681);
or UO_1390 (O_1390,N_8875,N_9363);
nor UO_1391 (O_1391,N_5718,N_7692);
nor UO_1392 (O_1392,N_5127,N_8681);
nor UO_1393 (O_1393,N_9226,N_5049);
or UO_1394 (O_1394,N_6678,N_8344);
or UO_1395 (O_1395,N_5408,N_8755);
nor UO_1396 (O_1396,N_8332,N_5714);
nand UO_1397 (O_1397,N_6224,N_6572);
or UO_1398 (O_1398,N_5266,N_9867);
nor UO_1399 (O_1399,N_7832,N_8599);
nand UO_1400 (O_1400,N_5905,N_9953);
and UO_1401 (O_1401,N_5742,N_8314);
and UO_1402 (O_1402,N_6579,N_5143);
or UO_1403 (O_1403,N_7328,N_7293);
or UO_1404 (O_1404,N_8720,N_9580);
nand UO_1405 (O_1405,N_7859,N_8349);
nor UO_1406 (O_1406,N_9950,N_7957);
and UO_1407 (O_1407,N_9302,N_8316);
and UO_1408 (O_1408,N_9157,N_7764);
and UO_1409 (O_1409,N_8753,N_6334);
or UO_1410 (O_1410,N_8429,N_7417);
and UO_1411 (O_1411,N_6776,N_9200);
nand UO_1412 (O_1412,N_7077,N_7931);
nor UO_1413 (O_1413,N_9860,N_5012);
or UO_1414 (O_1414,N_9954,N_8046);
or UO_1415 (O_1415,N_6406,N_6198);
or UO_1416 (O_1416,N_8375,N_7248);
or UO_1417 (O_1417,N_7253,N_5456);
nand UO_1418 (O_1418,N_7793,N_5208);
nand UO_1419 (O_1419,N_9550,N_5780);
and UO_1420 (O_1420,N_9413,N_6331);
nor UO_1421 (O_1421,N_7002,N_8235);
nand UO_1422 (O_1422,N_5606,N_8232);
and UO_1423 (O_1423,N_9692,N_6125);
and UO_1424 (O_1424,N_9021,N_9045);
and UO_1425 (O_1425,N_7742,N_5697);
nand UO_1426 (O_1426,N_5400,N_6485);
and UO_1427 (O_1427,N_7198,N_8005);
nand UO_1428 (O_1428,N_6312,N_8591);
nand UO_1429 (O_1429,N_5845,N_8543);
or UO_1430 (O_1430,N_8305,N_5204);
nor UO_1431 (O_1431,N_5055,N_5366);
nand UO_1432 (O_1432,N_8051,N_7658);
and UO_1433 (O_1433,N_9564,N_8325);
nor UO_1434 (O_1434,N_9567,N_9133);
or UO_1435 (O_1435,N_9700,N_6809);
and UO_1436 (O_1436,N_7999,N_6595);
or UO_1437 (O_1437,N_6398,N_7460);
nor UO_1438 (O_1438,N_6504,N_8793);
and UO_1439 (O_1439,N_6984,N_8254);
and UO_1440 (O_1440,N_5823,N_9638);
nand UO_1441 (O_1441,N_7036,N_8764);
nand UO_1442 (O_1442,N_6766,N_6816);
xnor UO_1443 (O_1443,N_9761,N_5711);
and UO_1444 (O_1444,N_8960,N_6082);
nand UO_1445 (O_1445,N_7289,N_6306);
and UO_1446 (O_1446,N_5269,N_5964);
nor UO_1447 (O_1447,N_7169,N_8754);
or UO_1448 (O_1448,N_7347,N_7431);
or UO_1449 (O_1449,N_8019,N_8075);
xor UO_1450 (O_1450,N_8233,N_9192);
and UO_1451 (O_1451,N_9412,N_5688);
nor UO_1452 (O_1452,N_7029,N_8871);
nand UO_1453 (O_1453,N_8830,N_9642);
and UO_1454 (O_1454,N_8288,N_6995);
or UO_1455 (O_1455,N_5438,N_7523);
nand UO_1456 (O_1456,N_5897,N_7188);
and UO_1457 (O_1457,N_9121,N_6660);
and UO_1458 (O_1458,N_6079,N_6990);
nor UO_1459 (O_1459,N_6037,N_5115);
and UO_1460 (O_1460,N_7265,N_5425);
nor UO_1461 (O_1461,N_8168,N_5123);
or UO_1462 (O_1462,N_8202,N_7490);
nor UO_1463 (O_1463,N_5733,N_8963);
nor UO_1464 (O_1464,N_8425,N_7000);
or UO_1465 (O_1465,N_6781,N_9436);
or UO_1466 (O_1466,N_9353,N_5084);
or UO_1467 (O_1467,N_9516,N_9866);
nor UO_1468 (O_1468,N_9018,N_7041);
or UO_1469 (O_1469,N_7708,N_5735);
or UO_1470 (O_1470,N_9625,N_7650);
or UO_1471 (O_1471,N_8381,N_5030);
nor UO_1472 (O_1472,N_6717,N_8547);
nor UO_1473 (O_1473,N_5294,N_9963);
nor UO_1474 (O_1474,N_5759,N_6249);
and UO_1475 (O_1475,N_7014,N_5010);
nor UO_1476 (O_1476,N_6858,N_5836);
and UO_1477 (O_1477,N_9609,N_7015);
and UO_1478 (O_1478,N_5356,N_5713);
nand UO_1479 (O_1479,N_5335,N_7912);
nor UO_1480 (O_1480,N_5306,N_7362);
xnor UO_1481 (O_1481,N_6714,N_9059);
or UO_1482 (O_1482,N_5481,N_5040);
and UO_1483 (O_1483,N_5493,N_6869);
and UO_1484 (O_1484,N_8694,N_6492);
or UO_1485 (O_1485,N_7313,N_6629);
or UO_1486 (O_1486,N_6782,N_6863);
nand UO_1487 (O_1487,N_5589,N_8565);
and UO_1488 (O_1488,N_6019,N_9244);
nor UO_1489 (O_1489,N_7595,N_7224);
nor UO_1490 (O_1490,N_8707,N_5426);
and UO_1491 (O_1491,N_5430,N_6901);
nand UO_1492 (O_1492,N_9992,N_9624);
and UO_1493 (O_1493,N_9794,N_9780);
nand UO_1494 (O_1494,N_8691,N_7754);
or UO_1495 (O_1495,N_9560,N_8523);
or UO_1496 (O_1496,N_5921,N_9565);
nand UO_1497 (O_1497,N_6764,N_6219);
or UO_1498 (O_1498,N_8781,N_8559);
or UO_1499 (O_1499,N_5147,N_5387);
endmodule