module basic_500_3000_500_60_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_409,In_397);
nand U1 (N_1,In_343,In_160);
nand U2 (N_2,In_337,In_32);
nor U3 (N_3,In_176,In_81);
nor U4 (N_4,In_139,In_499);
nand U5 (N_5,In_171,In_490);
or U6 (N_6,In_292,In_447);
nor U7 (N_7,In_443,In_145);
xor U8 (N_8,In_291,In_430);
or U9 (N_9,In_427,In_98);
nor U10 (N_10,In_393,In_424);
and U11 (N_11,In_129,In_440);
and U12 (N_12,In_357,In_166);
nor U13 (N_13,In_332,In_163);
nor U14 (N_14,In_240,In_419);
nor U15 (N_15,In_186,In_44);
or U16 (N_16,In_191,In_190);
and U17 (N_17,In_152,In_368);
nor U18 (N_18,In_156,In_297);
nand U19 (N_19,In_216,In_132);
and U20 (N_20,In_41,In_298);
nor U21 (N_21,In_210,In_229);
nor U22 (N_22,In_420,In_97);
or U23 (N_23,In_91,In_80);
nand U24 (N_24,In_154,In_261);
nor U25 (N_25,In_50,In_365);
nor U26 (N_26,In_144,In_476);
nor U27 (N_27,In_151,In_199);
nand U28 (N_28,In_62,In_12);
nor U29 (N_29,In_40,In_406);
and U30 (N_30,In_267,In_200);
and U31 (N_31,In_329,In_95);
nor U32 (N_32,In_354,In_286);
nor U33 (N_33,In_173,In_413);
nor U34 (N_34,In_121,In_169);
nand U35 (N_35,In_219,In_319);
and U36 (N_36,In_164,In_101);
nor U37 (N_37,In_260,In_223);
nor U38 (N_38,In_435,In_454);
and U39 (N_39,In_475,In_345);
nor U40 (N_40,In_324,In_19);
and U41 (N_41,In_10,In_271);
nor U42 (N_42,In_64,In_432);
or U43 (N_43,In_110,In_484);
and U44 (N_44,In_63,In_301);
or U45 (N_45,In_134,In_361);
nor U46 (N_46,In_20,In_177);
or U47 (N_47,In_441,In_211);
nor U48 (N_48,In_446,In_133);
and U49 (N_49,In_13,In_493);
nand U50 (N_50,In_308,In_92);
nand U51 (N_51,In_305,In_328);
or U52 (N_52,In_123,In_233);
or U53 (N_53,In_6,In_348);
or U54 (N_54,In_27,In_76);
or U55 (N_55,In_52,In_417);
or U56 (N_56,In_55,In_374);
and U57 (N_57,In_262,N_29);
nor U58 (N_58,In_407,In_53);
nand U59 (N_59,In_1,In_477);
nand U60 (N_60,In_46,In_356);
or U61 (N_61,In_203,In_180);
nor U62 (N_62,In_181,In_71);
nor U63 (N_63,In_347,In_438);
nor U64 (N_64,In_436,In_296);
and U65 (N_65,In_54,In_450);
and U66 (N_66,In_135,In_138);
and U67 (N_67,In_136,In_366);
nand U68 (N_68,In_363,In_483);
or U69 (N_69,N_10,In_14);
or U70 (N_70,In_100,In_353);
nor U71 (N_71,In_220,N_7);
or U72 (N_72,In_57,In_414);
and U73 (N_73,In_187,In_444);
or U74 (N_74,In_4,In_445);
and U75 (N_75,In_464,In_496);
nor U76 (N_76,In_491,In_395);
or U77 (N_77,In_472,In_205);
or U78 (N_78,In_84,In_431);
and U79 (N_79,In_290,In_346);
or U80 (N_80,In_172,In_344);
nor U81 (N_81,In_412,In_273);
nor U82 (N_82,In_388,In_167);
nand U83 (N_83,In_178,N_49);
nor U84 (N_84,In_299,In_94);
nor U85 (N_85,In_396,In_33);
or U86 (N_86,In_195,N_16);
nor U87 (N_87,N_33,In_162);
nand U88 (N_88,In_462,In_140);
or U89 (N_89,In_196,N_20);
nor U90 (N_90,In_482,In_352);
nand U91 (N_91,N_23,In_75);
or U92 (N_92,N_24,In_460);
and U93 (N_93,In_351,In_26);
and U94 (N_94,In_453,In_125);
xor U95 (N_95,In_113,In_340);
nor U96 (N_96,In_36,In_227);
or U97 (N_97,In_147,In_194);
nor U98 (N_98,In_142,N_22);
nor U99 (N_99,In_115,In_465);
or U100 (N_100,In_197,In_120);
nor U101 (N_101,In_108,N_25);
and U102 (N_102,In_48,In_24);
nor U103 (N_103,In_258,N_83);
or U104 (N_104,In_248,In_467);
nor U105 (N_105,In_170,N_12);
and U106 (N_106,In_333,In_96);
and U107 (N_107,In_391,In_21);
and U108 (N_108,N_38,In_479);
and U109 (N_109,In_497,In_266);
nand U110 (N_110,In_425,In_434);
nand U111 (N_111,In_208,N_48);
and U112 (N_112,In_313,In_452);
and U113 (N_113,In_410,N_69);
or U114 (N_114,In_402,In_252);
and U115 (N_115,N_89,N_3);
nor U116 (N_116,In_327,In_43);
nand U117 (N_117,In_183,In_349);
or U118 (N_118,In_433,In_377);
or U119 (N_119,In_283,In_9);
and U120 (N_120,In_274,In_331);
nand U121 (N_121,In_237,In_279);
nand U122 (N_122,In_486,N_39);
and U123 (N_123,N_61,In_179);
or U124 (N_124,N_78,In_380);
nor U125 (N_125,In_82,In_466);
nor U126 (N_126,N_80,In_378);
and U127 (N_127,N_98,N_87);
and U128 (N_128,In_330,In_66);
and U129 (N_129,In_270,In_399);
nor U130 (N_130,In_280,In_241);
or U131 (N_131,In_246,In_107);
nor U132 (N_132,In_16,In_360);
or U133 (N_133,In_214,N_63);
or U134 (N_134,In_238,N_21);
nor U135 (N_135,In_311,In_251);
nor U136 (N_136,N_74,In_65);
or U137 (N_137,In_489,In_358);
and U138 (N_138,N_36,N_31);
nand U139 (N_139,In_458,In_306);
or U140 (N_140,In_15,In_56);
and U141 (N_141,N_32,In_303);
and U142 (N_142,In_369,In_60);
nand U143 (N_143,In_45,In_304);
and U144 (N_144,In_137,In_99);
and U145 (N_145,In_253,In_153);
or U146 (N_146,In_480,N_5);
nand U147 (N_147,In_335,In_7);
or U148 (N_148,N_15,In_422);
or U149 (N_149,N_75,In_429);
xnor U150 (N_150,In_487,In_317);
and U151 (N_151,N_124,In_161);
or U152 (N_152,In_481,In_492);
xor U153 (N_153,In_293,In_403);
nand U154 (N_154,In_459,In_264);
or U155 (N_155,N_139,In_217);
and U156 (N_156,N_141,In_89);
nor U157 (N_157,N_125,In_159);
nand U158 (N_158,In_272,In_103);
and U159 (N_159,In_78,In_404);
and U160 (N_160,In_18,N_137);
nand U161 (N_161,In_127,In_371);
and U162 (N_162,In_468,N_53);
nor U163 (N_163,N_81,N_106);
or U164 (N_164,N_132,In_288);
and U165 (N_165,In_37,In_143);
and U166 (N_166,In_442,In_321);
nor U167 (N_167,In_93,In_392);
nand U168 (N_168,N_44,In_204);
nor U169 (N_169,In_307,In_206);
or U170 (N_170,In_326,In_394);
nand U171 (N_171,In_11,In_281);
and U172 (N_172,In_86,In_38);
nor U173 (N_173,N_148,N_47);
nand U174 (N_174,In_265,N_58);
xnor U175 (N_175,In_373,N_135);
or U176 (N_176,In_116,In_322);
and U177 (N_177,In_385,N_55);
and U178 (N_178,In_259,In_249);
or U179 (N_179,In_174,N_56);
and U180 (N_180,In_209,In_478);
or U181 (N_181,In_59,N_116);
and U182 (N_182,N_127,In_29);
and U183 (N_183,In_287,In_83);
and U184 (N_184,N_149,In_119);
or U185 (N_185,N_73,N_72);
nand U186 (N_186,In_473,In_325);
nand U187 (N_187,In_193,In_106);
nor U188 (N_188,N_57,In_312);
and U189 (N_189,In_185,N_140);
or U190 (N_190,N_27,N_45);
and U191 (N_191,In_168,N_42);
nor U192 (N_192,In_285,N_59);
nand U193 (N_193,In_201,N_79);
nand U194 (N_194,N_30,N_93);
or U195 (N_195,N_147,N_108);
nor U196 (N_196,N_129,N_115);
and U197 (N_197,N_138,In_245);
and U198 (N_198,In_372,N_136);
or U199 (N_199,In_117,In_318);
and U200 (N_200,In_5,In_239);
nand U201 (N_201,In_236,N_190);
nor U202 (N_202,N_194,N_197);
or U203 (N_203,In_350,In_231);
nand U204 (N_204,N_4,N_40);
nand U205 (N_205,In_213,N_37);
or U206 (N_206,In_457,In_122);
nor U207 (N_207,In_471,In_426);
nand U208 (N_208,In_254,N_9);
or U209 (N_209,In_275,In_367);
nor U210 (N_210,In_221,In_87);
or U211 (N_211,In_49,In_418);
nand U212 (N_212,In_470,N_186);
nor U213 (N_213,N_107,N_65);
and U214 (N_214,N_122,N_185);
nand U215 (N_215,N_94,N_182);
nor U216 (N_216,In_131,In_28);
nor U217 (N_217,In_302,N_1);
and U218 (N_218,In_314,N_99);
or U219 (N_219,N_153,In_423);
nor U220 (N_220,In_0,N_134);
and U221 (N_221,N_174,N_14);
and U222 (N_222,N_118,In_39);
nor U223 (N_223,N_170,In_461);
nand U224 (N_224,In_411,In_155);
or U225 (N_225,In_35,In_455);
nand U226 (N_226,In_376,N_144);
or U227 (N_227,N_95,In_73);
nor U228 (N_228,N_111,In_428);
and U229 (N_229,In_188,N_198);
or U230 (N_230,In_198,In_146);
and U231 (N_231,In_189,N_121);
or U232 (N_232,N_100,N_151);
nand U233 (N_233,In_141,In_289);
nor U234 (N_234,N_187,N_178);
nor U235 (N_235,N_119,In_109);
nor U236 (N_236,In_370,In_495);
nor U237 (N_237,In_255,N_133);
nor U238 (N_238,N_166,In_456);
or U239 (N_239,In_243,In_157);
and U240 (N_240,N_90,In_309);
nand U241 (N_241,N_82,In_118);
nand U242 (N_242,N_171,In_320);
nor U243 (N_243,In_338,In_23);
or U244 (N_244,In_105,In_226);
or U245 (N_245,In_421,In_112);
xor U246 (N_246,In_439,N_143);
nor U247 (N_247,In_384,N_103);
or U248 (N_248,In_310,In_400);
and U249 (N_249,N_71,N_46);
nand U250 (N_250,In_250,In_224);
nand U251 (N_251,N_110,N_245);
nand U252 (N_252,N_101,In_295);
or U253 (N_253,In_128,N_203);
nor U254 (N_254,N_215,In_362);
or U255 (N_255,N_11,N_50);
or U256 (N_256,In_31,N_246);
nand U257 (N_257,N_244,In_85);
nor U258 (N_258,N_13,In_375);
and U259 (N_259,N_70,N_224);
or U260 (N_260,N_211,N_2);
nand U261 (N_261,N_155,In_339);
xor U262 (N_262,N_192,N_172);
nand U263 (N_263,N_207,N_8);
and U264 (N_264,In_42,In_67);
nor U265 (N_265,N_102,In_382);
nand U266 (N_266,In_90,In_276);
nor U267 (N_267,N_231,N_206);
nor U268 (N_268,N_34,N_154);
or U269 (N_269,In_104,N_67);
and U270 (N_270,N_26,In_222);
and U271 (N_271,N_130,N_201);
nor U272 (N_272,N_180,In_149);
or U273 (N_273,N_223,N_86);
or U274 (N_274,N_84,In_114);
and U275 (N_275,In_256,N_236);
nor U276 (N_276,N_64,In_415);
nand U277 (N_277,N_62,In_202);
or U278 (N_278,In_74,In_448);
nor U279 (N_279,N_169,In_488);
or U280 (N_280,N_54,In_234);
nand U281 (N_281,In_405,In_364);
and U282 (N_282,In_17,N_104);
nand U283 (N_283,In_58,N_168);
nor U284 (N_284,In_336,In_102);
nand U285 (N_285,N_77,N_195);
nor U286 (N_286,N_239,N_183);
nor U287 (N_287,In_3,In_387);
nor U288 (N_288,N_152,N_230);
nor U289 (N_289,In_494,N_60);
nand U290 (N_290,N_237,N_68);
nand U291 (N_291,In_158,In_242);
nor U292 (N_292,N_229,N_196);
nor U293 (N_293,In_257,In_315);
or U294 (N_294,In_449,N_204);
or U295 (N_295,N_96,N_221);
nand U296 (N_296,In_383,In_294);
nand U297 (N_297,In_284,In_22);
and U298 (N_298,In_408,N_43);
nand U299 (N_299,N_205,N_76);
nand U300 (N_300,N_128,N_232);
and U301 (N_301,N_91,In_247);
and U302 (N_302,N_252,N_199);
and U303 (N_303,In_300,In_437);
or U304 (N_304,N_209,N_290);
nand U305 (N_305,N_287,N_216);
or U306 (N_306,In_390,In_232);
nand U307 (N_307,N_255,In_126);
nand U308 (N_308,N_226,N_247);
nand U309 (N_309,In_381,N_288);
and U310 (N_310,In_182,N_175);
nor U311 (N_311,In_72,N_283);
xnor U312 (N_312,N_272,N_238);
nand U313 (N_313,In_124,N_286);
nand U314 (N_314,N_243,N_274);
and U315 (N_315,N_193,N_117);
and U316 (N_316,N_173,N_163);
nor U317 (N_317,N_113,N_235);
xor U318 (N_318,In_463,N_279);
or U319 (N_319,In_34,N_251);
nor U320 (N_320,N_145,In_263);
nor U321 (N_321,N_51,N_263);
or U322 (N_322,N_297,N_167);
nand U323 (N_323,N_292,N_164);
and U324 (N_324,N_261,In_235);
nor U325 (N_325,N_284,N_242);
nand U326 (N_326,N_264,N_92);
and U327 (N_327,In_474,In_88);
and U328 (N_328,N_28,N_281);
and U329 (N_329,N_97,N_259);
nor U330 (N_330,In_148,N_228);
or U331 (N_331,N_217,N_218);
or U332 (N_332,N_250,In_341);
nand U333 (N_333,N_241,N_179);
nand U334 (N_334,N_159,In_68);
nor U335 (N_335,N_17,N_184);
and U336 (N_336,N_156,N_213);
nand U337 (N_337,In_228,N_131);
and U338 (N_338,N_269,In_244);
or U339 (N_339,N_296,N_162);
nand U340 (N_340,In_342,N_262);
and U341 (N_341,N_150,N_160);
xnor U342 (N_342,N_227,In_218);
nor U343 (N_343,In_278,N_299);
xor U344 (N_344,N_298,N_200);
or U345 (N_345,In_77,In_451);
or U346 (N_346,N_293,In_70);
and U347 (N_347,N_289,In_469);
or U348 (N_348,In_130,In_225);
or U349 (N_349,N_158,N_257);
xor U350 (N_350,N_294,N_343);
nand U351 (N_351,N_345,N_220);
nand U352 (N_352,N_258,N_6);
and U353 (N_353,N_234,N_181);
or U354 (N_354,In_277,In_230);
xnor U355 (N_355,In_61,N_321);
and U356 (N_356,In_175,N_280);
nor U357 (N_357,In_212,N_225);
and U358 (N_358,N_325,N_328);
and U359 (N_359,N_314,N_332);
and U360 (N_360,N_311,N_189);
or U361 (N_361,N_277,N_0);
and U362 (N_362,N_214,N_329);
or U363 (N_363,N_210,In_150);
nor U364 (N_364,In_268,N_337);
xor U365 (N_365,N_318,N_157);
nor U366 (N_366,N_268,N_253);
nand U367 (N_367,N_256,N_320);
xnor U368 (N_368,N_300,In_359);
nor U369 (N_369,N_344,N_282);
and U370 (N_370,N_306,N_120);
nor U371 (N_371,N_342,N_35);
and U372 (N_372,N_260,In_355);
and U373 (N_373,N_18,In_379);
or U374 (N_374,In_389,N_349);
nand U375 (N_375,N_85,N_276);
or U376 (N_376,N_19,In_79);
or U377 (N_377,N_315,N_348);
or U378 (N_378,N_266,N_275);
or U379 (N_379,N_302,In_47);
and U380 (N_380,N_177,N_346);
or U381 (N_381,N_270,N_126);
and U382 (N_382,N_326,N_327);
and U383 (N_383,N_233,In_51);
or U384 (N_384,N_105,In_316);
or U385 (N_385,N_267,N_347);
and U386 (N_386,N_41,N_254);
or U387 (N_387,N_271,N_265);
nor U388 (N_388,N_222,N_165);
and U389 (N_389,N_123,N_219);
and U390 (N_390,N_339,N_313);
or U391 (N_391,N_333,N_176);
nand U392 (N_392,N_202,N_212);
or U393 (N_393,N_66,N_323);
or U394 (N_394,N_109,N_278);
or U395 (N_395,In_323,N_161);
or U396 (N_396,N_322,N_295);
and U397 (N_397,N_334,N_285);
nor U398 (N_398,In_165,N_308);
nand U399 (N_399,In_69,In_269);
xnor U400 (N_400,N_366,N_303);
and U401 (N_401,N_304,In_282);
and U402 (N_402,N_240,N_380);
and U403 (N_403,N_358,N_375);
nand U404 (N_404,N_381,In_111);
nand U405 (N_405,In_192,In_2);
or U406 (N_406,N_336,N_354);
and U407 (N_407,N_384,In_334);
and U408 (N_408,N_340,N_390);
or U409 (N_409,N_316,N_273);
and U410 (N_410,N_291,In_25);
or U411 (N_411,N_382,In_398);
or U412 (N_412,N_363,N_331);
nand U413 (N_413,N_335,N_377);
nor U414 (N_414,In_416,N_310);
and U415 (N_415,N_317,N_386);
nand U416 (N_416,N_374,N_394);
and U417 (N_417,N_367,N_357);
nand U418 (N_418,N_396,N_362);
nand U419 (N_419,N_350,N_356);
nand U420 (N_420,N_112,N_393);
and U421 (N_421,N_249,N_191);
nor U422 (N_422,N_365,N_307);
nand U423 (N_423,N_188,In_401);
or U424 (N_424,N_389,N_369);
nand U425 (N_425,N_309,N_52);
nor U426 (N_426,N_324,In_485);
or U427 (N_427,N_330,In_215);
or U428 (N_428,N_88,N_385);
nor U429 (N_429,N_319,In_30);
or U430 (N_430,N_378,N_146);
nor U431 (N_431,N_383,N_395);
nor U432 (N_432,N_376,N_398);
nand U433 (N_433,N_248,N_371);
nor U434 (N_434,In_184,In_498);
nand U435 (N_435,N_364,N_379);
and U436 (N_436,N_305,N_360);
nor U437 (N_437,N_397,N_341);
nor U438 (N_438,N_142,In_386);
nand U439 (N_439,N_370,N_372);
nor U440 (N_440,N_352,N_351);
nand U441 (N_441,N_208,N_388);
and U442 (N_442,N_359,In_207);
nand U443 (N_443,N_399,N_114);
or U444 (N_444,N_338,N_312);
nand U445 (N_445,N_368,N_391);
or U446 (N_446,N_392,N_353);
and U447 (N_447,N_387,N_361);
nor U448 (N_448,N_373,N_301);
nand U449 (N_449,N_355,In_8);
and U450 (N_450,N_424,N_431);
and U451 (N_451,N_428,N_447);
and U452 (N_452,N_435,N_423);
nor U453 (N_453,N_427,N_412);
and U454 (N_454,N_432,N_410);
or U455 (N_455,N_439,N_433);
nor U456 (N_456,N_445,N_430);
or U457 (N_457,N_438,N_448);
nor U458 (N_458,N_413,N_443);
and U459 (N_459,N_434,N_444);
nand U460 (N_460,N_442,N_405);
nor U461 (N_461,N_446,N_400);
nand U462 (N_462,N_440,N_414);
or U463 (N_463,N_401,N_416);
nor U464 (N_464,N_408,N_422);
and U465 (N_465,N_419,N_411);
or U466 (N_466,N_421,N_426);
xnor U467 (N_467,N_403,N_425);
nand U468 (N_468,N_415,N_420);
and U469 (N_469,N_402,N_449);
nand U470 (N_470,N_441,N_436);
nor U471 (N_471,N_406,N_417);
nor U472 (N_472,N_429,N_404);
and U473 (N_473,N_409,N_437);
nor U474 (N_474,N_407,N_418);
and U475 (N_475,N_437,N_401);
xor U476 (N_476,N_437,N_417);
and U477 (N_477,N_436,N_448);
nand U478 (N_478,N_400,N_414);
nor U479 (N_479,N_442,N_427);
and U480 (N_480,N_418,N_439);
and U481 (N_481,N_414,N_410);
nand U482 (N_482,N_447,N_441);
nand U483 (N_483,N_445,N_420);
or U484 (N_484,N_443,N_402);
nand U485 (N_485,N_446,N_423);
and U486 (N_486,N_427,N_440);
nor U487 (N_487,N_415,N_423);
nand U488 (N_488,N_437,N_449);
and U489 (N_489,N_441,N_445);
or U490 (N_490,N_449,N_414);
or U491 (N_491,N_436,N_411);
and U492 (N_492,N_412,N_434);
nor U493 (N_493,N_415,N_406);
nand U494 (N_494,N_400,N_440);
and U495 (N_495,N_403,N_415);
nand U496 (N_496,N_445,N_443);
or U497 (N_497,N_438,N_415);
or U498 (N_498,N_412,N_430);
nand U499 (N_499,N_405,N_417);
or U500 (N_500,N_461,N_491);
nand U501 (N_501,N_497,N_469);
and U502 (N_502,N_479,N_465);
and U503 (N_503,N_481,N_490);
or U504 (N_504,N_489,N_474);
or U505 (N_505,N_462,N_482);
and U506 (N_506,N_470,N_455);
nand U507 (N_507,N_476,N_483);
and U508 (N_508,N_463,N_464);
and U509 (N_509,N_475,N_468);
nor U510 (N_510,N_493,N_450);
or U511 (N_511,N_453,N_471);
nor U512 (N_512,N_487,N_494);
nand U513 (N_513,N_486,N_478);
nor U514 (N_514,N_466,N_460);
nand U515 (N_515,N_492,N_477);
nand U516 (N_516,N_485,N_451);
nand U517 (N_517,N_473,N_456);
nor U518 (N_518,N_458,N_459);
and U519 (N_519,N_452,N_498);
and U520 (N_520,N_467,N_488);
nand U521 (N_521,N_472,N_457);
or U522 (N_522,N_454,N_484);
or U523 (N_523,N_480,N_495);
nand U524 (N_524,N_499,N_496);
or U525 (N_525,N_458,N_473);
or U526 (N_526,N_491,N_451);
or U527 (N_527,N_492,N_455);
nand U528 (N_528,N_464,N_492);
and U529 (N_529,N_483,N_451);
nor U530 (N_530,N_452,N_479);
nand U531 (N_531,N_489,N_492);
and U532 (N_532,N_464,N_457);
and U533 (N_533,N_498,N_465);
and U534 (N_534,N_459,N_473);
nand U535 (N_535,N_481,N_450);
and U536 (N_536,N_485,N_476);
xnor U537 (N_537,N_478,N_488);
nor U538 (N_538,N_465,N_488);
or U539 (N_539,N_477,N_482);
nand U540 (N_540,N_457,N_459);
nor U541 (N_541,N_481,N_499);
or U542 (N_542,N_474,N_454);
xnor U543 (N_543,N_461,N_490);
or U544 (N_544,N_463,N_453);
or U545 (N_545,N_472,N_499);
and U546 (N_546,N_497,N_479);
or U547 (N_547,N_470,N_464);
nor U548 (N_548,N_486,N_490);
nor U549 (N_549,N_482,N_453);
and U550 (N_550,N_501,N_518);
or U551 (N_551,N_522,N_535);
or U552 (N_552,N_526,N_539);
nor U553 (N_553,N_546,N_502);
nand U554 (N_554,N_547,N_505);
nand U555 (N_555,N_511,N_527);
and U556 (N_556,N_512,N_538);
and U557 (N_557,N_524,N_517);
nand U558 (N_558,N_500,N_504);
and U559 (N_559,N_542,N_548);
and U560 (N_560,N_515,N_510);
or U561 (N_561,N_534,N_520);
and U562 (N_562,N_503,N_516);
nand U563 (N_563,N_514,N_531);
nand U564 (N_564,N_523,N_528);
or U565 (N_565,N_541,N_537);
or U566 (N_566,N_536,N_521);
and U567 (N_567,N_519,N_507);
nor U568 (N_568,N_532,N_513);
nor U569 (N_569,N_549,N_545);
or U570 (N_570,N_506,N_508);
and U571 (N_571,N_540,N_533);
nand U572 (N_572,N_525,N_543);
and U573 (N_573,N_509,N_544);
nand U574 (N_574,N_530,N_529);
and U575 (N_575,N_544,N_542);
or U576 (N_576,N_507,N_539);
or U577 (N_577,N_536,N_516);
or U578 (N_578,N_503,N_537);
nand U579 (N_579,N_519,N_539);
or U580 (N_580,N_522,N_531);
nand U581 (N_581,N_515,N_512);
nor U582 (N_582,N_512,N_521);
nor U583 (N_583,N_514,N_522);
nor U584 (N_584,N_527,N_517);
nor U585 (N_585,N_542,N_549);
nand U586 (N_586,N_529,N_515);
nand U587 (N_587,N_508,N_542);
nand U588 (N_588,N_527,N_541);
nand U589 (N_589,N_506,N_503);
and U590 (N_590,N_524,N_521);
and U591 (N_591,N_539,N_504);
nand U592 (N_592,N_513,N_549);
nor U593 (N_593,N_521,N_533);
xnor U594 (N_594,N_518,N_544);
or U595 (N_595,N_507,N_501);
and U596 (N_596,N_510,N_540);
nor U597 (N_597,N_531,N_549);
nor U598 (N_598,N_523,N_511);
and U599 (N_599,N_521,N_523);
nor U600 (N_600,N_598,N_589);
nand U601 (N_601,N_574,N_580);
xor U602 (N_602,N_582,N_578);
and U603 (N_603,N_555,N_559);
and U604 (N_604,N_561,N_575);
nand U605 (N_605,N_556,N_553);
or U606 (N_606,N_597,N_587);
nor U607 (N_607,N_584,N_579);
nor U608 (N_608,N_576,N_591);
nor U609 (N_609,N_566,N_592);
and U610 (N_610,N_562,N_581);
nand U611 (N_611,N_565,N_560);
nor U612 (N_612,N_551,N_583);
and U613 (N_613,N_552,N_564);
or U614 (N_614,N_593,N_573);
or U615 (N_615,N_590,N_557);
and U616 (N_616,N_586,N_569);
or U617 (N_617,N_585,N_558);
nor U618 (N_618,N_596,N_563);
or U619 (N_619,N_568,N_595);
or U620 (N_620,N_572,N_554);
and U621 (N_621,N_567,N_588);
nand U622 (N_622,N_550,N_594);
nor U623 (N_623,N_571,N_577);
nor U624 (N_624,N_570,N_599);
nor U625 (N_625,N_561,N_593);
nand U626 (N_626,N_564,N_582);
or U627 (N_627,N_572,N_598);
nor U628 (N_628,N_577,N_583);
and U629 (N_629,N_555,N_569);
or U630 (N_630,N_586,N_588);
or U631 (N_631,N_562,N_591);
nand U632 (N_632,N_575,N_563);
nand U633 (N_633,N_591,N_579);
nor U634 (N_634,N_552,N_560);
nor U635 (N_635,N_568,N_556);
xnor U636 (N_636,N_552,N_550);
and U637 (N_637,N_559,N_551);
or U638 (N_638,N_592,N_553);
nand U639 (N_639,N_571,N_550);
nor U640 (N_640,N_597,N_562);
nand U641 (N_641,N_565,N_569);
and U642 (N_642,N_553,N_581);
or U643 (N_643,N_563,N_577);
xor U644 (N_644,N_597,N_594);
nor U645 (N_645,N_591,N_598);
xnor U646 (N_646,N_574,N_595);
and U647 (N_647,N_559,N_563);
xnor U648 (N_648,N_596,N_591);
and U649 (N_649,N_556,N_578);
or U650 (N_650,N_631,N_637);
nor U651 (N_651,N_610,N_617);
or U652 (N_652,N_648,N_616);
and U653 (N_653,N_640,N_613);
or U654 (N_654,N_619,N_620);
nand U655 (N_655,N_639,N_603);
and U656 (N_656,N_604,N_646);
nor U657 (N_657,N_624,N_644);
nor U658 (N_658,N_611,N_605);
nor U659 (N_659,N_629,N_614);
nand U660 (N_660,N_626,N_632);
and U661 (N_661,N_645,N_630);
and U662 (N_662,N_609,N_636);
nor U663 (N_663,N_600,N_643);
and U664 (N_664,N_607,N_608);
or U665 (N_665,N_634,N_638);
or U666 (N_666,N_642,N_601);
nor U667 (N_667,N_633,N_627);
nand U668 (N_668,N_647,N_641);
xor U669 (N_669,N_628,N_635);
and U670 (N_670,N_612,N_618);
and U671 (N_671,N_625,N_649);
and U672 (N_672,N_623,N_615);
nand U673 (N_673,N_622,N_606);
nand U674 (N_674,N_602,N_621);
or U675 (N_675,N_602,N_606);
or U676 (N_676,N_615,N_611);
nor U677 (N_677,N_636,N_645);
or U678 (N_678,N_613,N_617);
and U679 (N_679,N_617,N_621);
xnor U680 (N_680,N_620,N_609);
nor U681 (N_681,N_640,N_644);
or U682 (N_682,N_632,N_609);
or U683 (N_683,N_621,N_629);
or U684 (N_684,N_647,N_605);
nor U685 (N_685,N_641,N_615);
nor U686 (N_686,N_611,N_622);
nor U687 (N_687,N_632,N_612);
nor U688 (N_688,N_634,N_626);
and U689 (N_689,N_622,N_639);
nand U690 (N_690,N_625,N_614);
or U691 (N_691,N_606,N_649);
nor U692 (N_692,N_638,N_643);
nor U693 (N_693,N_639,N_614);
and U694 (N_694,N_632,N_648);
or U695 (N_695,N_615,N_626);
and U696 (N_696,N_603,N_609);
nor U697 (N_697,N_622,N_620);
nand U698 (N_698,N_602,N_642);
nand U699 (N_699,N_628,N_601);
and U700 (N_700,N_677,N_684);
nand U701 (N_701,N_652,N_665);
and U702 (N_702,N_681,N_668);
nor U703 (N_703,N_691,N_661);
nor U704 (N_704,N_693,N_674);
and U705 (N_705,N_679,N_683);
nor U706 (N_706,N_682,N_662);
or U707 (N_707,N_672,N_667);
nor U708 (N_708,N_654,N_678);
or U709 (N_709,N_659,N_676);
nand U710 (N_710,N_687,N_690);
nand U711 (N_711,N_666,N_658);
and U712 (N_712,N_651,N_680);
nor U713 (N_713,N_670,N_698);
and U714 (N_714,N_660,N_675);
and U715 (N_715,N_699,N_689);
or U716 (N_716,N_673,N_655);
and U717 (N_717,N_653,N_686);
nand U718 (N_718,N_695,N_692);
and U719 (N_719,N_694,N_664);
or U720 (N_720,N_685,N_657);
xor U721 (N_721,N_696,N_688);
or U722 (N_722,N_650,N_656);
or U723 (N_723,N_669,N_671);
nor U724 (N_724,N_697,N_663);
or U725 (N_725,N_660,N_674);
nor U726 (N_726,N_664,N_660);
and U727 (N_727,N_691,N_680);
nand U728 (N_728,N_659,N_661);
and U729 (N_729,N_690,N_676);
and U730 (N_730,N_682,N_697);
xor U731 (N_731,N_688,N_684);
nand U732 (N_732,N_681,N_688);
nand U733 (N_733,N_654,N_664);
nor U734 (N_734,N_693,N_692);
nand U735 (N_735,N_699,N_698);
xor U736 (N_736,N_652,N_656);
or U737 (N_737,N_698,N_664);
and U738 (N_738,N_680,N_666);
nand U739 (N_739,N_662,N_671);
nor U740 (N_740,N_697,N_698);
nand U741 (N_741,N_673,N_699);
and U742 (N_742,N_680,N_687);
nor U743 (N_743,N_697,N_687);
nor U744 (N_744,N_694,N_662);
or U745 (N_745,N_698,N_669);
nor U746 (N_746,N_668,N_672);
and U747 (N_747,N_690,N_681);
nand U748 (N_748,N_654,N_670);
nand U749 (N_749,N_691,N_650);
nand U750 (N_750,N_713,N_737);
or U751 (N_751,N_708,N_745);
and U752 (N_752,N_735,N_743);
nor U753 (N_753,N_709,N_718);
or U754 (N_754,N_726,N_724);
nor U755 (N_755,N_725,N_707);
and U756 (N_756,N_704,N_727);
nor U757 (N_757,N_748,N_738);
or U758 (N_758,N_716,N_729);
and U759 (N_759,N_741,N_723);
nand U760 (N_760,N_701,N_744);
nand U761 (N_761,N_739,N_740);
or U762 (N_762,N_710,N_736);
nand U763 (N_763,N_719,N_732);
nand U764 (N_764,N_715,N_734);
and U765 (N_765,N_712,N_730);
and U766 (N_766,N_742,N_746);
nor U767 (N_767,N_728,N_705);
or U768 (N_768,N_700,N_722);
and U769 (N_769,N_749,N_747);
and U770 (N_770,N_706,N_721);
nor U771 (N_771,N_720,N_733);
or U772 (N_772,N_714,N_702);
or U773 (N_773,N_717,N_711);
nor U774 (N_774,N_731,N_703);
or U775 (N_775,N_721,N_745);
nand U776 (N_776,N_726,N_747);
or U777 (N_777,N_749,N_713);
nand U778 (N_778,N_730,N_738);
nor U779 (N_779,N_715,N_731);
and U780 (N_780,N_728,N_742);
and U781 (N_781,N_718,N_712);
or U782 (N_782,N_748,N_732);
nor U783 (N_783,N_742,N_735);
nand U784 (N_784,N_722,N_716);
and U785 (N_785,N_716,N_706);
or U786 (N_786,N_730,N_713);
nor U787 (N_787,N_700,N_726);
nand U788 (N_788,N_749,N_705);
nor U789 (N_789,N_738,N_734);
or U790 (N_790,N_713,N_705);
or U791 (N_791,N_747,N_710);
nand U792 (N_792,N_746,N_722);
or U793 (N_793,N_703,N_748);
nor U794 (N_794,N_725,N_729);
and U795 (N_795,N_735,N_736);
nor U796 (N_796,N_736,N_731);
and U797 (N_797,N_711,N_745);
or U798 (N_798,N_714,N_718);
and U799 (N_799,N_733,N_731);
nand U800 (N_800,N_756,N_754);
nand U801 (N_801,N_751,N_759);
nor U802 (N_802,N_788,N_767);
nand U803 (N_803,N_785,N_752);
and U804 (N_804,N_789,N_772);
xnor U805 (N_805,N_784,N_755);
or U806 (N_806,N_760,N_774);
or U807 (N_807,N_761,N_753);
and U808 (N_808,N_782,N_790);
nor U809 (N_809,N_793,N_791);
nor U810 (N_810,N_769,N_795);
nand U811 (N_811,N_781,N_783);
or U812 (N_812,N_771,N_787);
nor U813 (N_813,N_780,N_768);
nand U814 (N_814,N_758,N_799);
nor U815 (N_815,N_762,N_750);
nand U816 (N_816,N_778,N_765);
and U817 (N_817,N_757,N_770);
or U818 (N_818,N_797,N_786);
and U819 (N_819,N_796,N_776);
or U820 (N_820,N_779,N_766);
or U821 (N_821,N_777,N_775);
and U822 (N_822,N_798,N_763);
and U823 (N_823,N_794,N_792);
and U824 (N_824,N_764,N_773);
nand U825 (N_825,N_786,N_767);
and U826 (N_826,N_777,N_761);
or U827 (N_827,N_799,N_793);
nor U828 (N_828,N_758,N_791);
or U829 (N_829,N_768,N_795);
nor U830 (N_830,N_788,N_773);
and U831 (N_831,N_777,N_786);
and U832 (N_832,N_772,N_770);
or U833 (N_833,N_769,N_755);
nor U834 (N_834,N_751,N_797);
and U835 (N_835,N_756,N_765);
nor U836 (N_836,N_784,N_778);
nand U837 (N_837,N_782,N_781);
nor U838 (N_838,N_796,N_793);
nor U839 (N_839,N_783,N_773);
and U840 (N_840,N_752,N_755);
nand U841 (N_841,N_798,N_771);
or U842 (N_842,N_774,N_750);
nor U843 (N_843,N_795,N_757);
and U844 (N_844,N_774,N_754);
or U845 (N_845,N_781,N_766);
nor U846 (N_846,N_776,N_787);
and U847 (N_847,N_758,N_767);
nand U848 (N_848,N_784,N_788);
nor U849 (N_849,N_781,N_779);
or U850 (N_850,N_821,N_838);
nor U851 (N_851,N_834,N_803);
or U852 (N_852,N_830,N_805);
and U853 (N_853,N_810,N_846);
or U854 (N_854,N_843,N_819);
nand U855 (N_855,N_820,N_827);
or U856 (N_856,N_832,N_840);
nand U857 (N_857,N_829,N_815);
nor U858 (N_858,N_817,N_847);
nand U859 (N_859,N_816,N_848);
or U860 (N_860,N_841,N_814);
nor U861 (N_861,N_831,N_812);
and U862 (N_862,N_833,N_800);
nor U863 (N_863,N_842,N_813);
nand U864 (N_864,N_844,N_802);
or U865 (N_865,N_806,N_822);
and U866 (N_866,N_849,N_835);
and U867 (N_867,N_807,N_818);
nor U868 (N_868,N_826,N_836);
nor U869 (N_869,N_828,N_845);
nor U870 (N_870,N_808,N_824);
nor U871 (N_871,N_837,N_809);
or U872 (N_872,N_825,N_823);
nor U873 (N_873,N_839,N_801);
nand U874 (N_874,N_811,N_804);
and U875 (N_875,N_806,N_813);
and U876 (N_876,N_801,N_838);
and U877 (N_877,N_834,N_846);
and U878 (N_878,N_805,N_844);
nand U879 (N_879,N_801,N_830);
nor U880 (N_880,N_845,N_844);
and U881 (N_881,N_844,N_828);
nand U882 (N_882,N_834,N_815);
nand U883 (N_883,N_839,N_814);
nor U884 (N_884,N_820,N_805);
nand U885 (N_885,N_836,N_817);
nand U886 (N_886,N_818,N_845);
or U887 (N_887,N_818,N_814);
nor U888 (N_888,N_832,N_831);
or U889 (N_889,N_814,N_838);
and U890 (N_890,N_845,N_843);
nor U891 (N_891,N_814,N_800);
or U892 (N_892,N_846,N_840);
or U893 (N_893,N_811,N_815);
nand U894 (N_894,N_825,N_841);
and U895 (N_895,N_817,N_834);
or U896 (N_896,N_804,N_807);
and U897 (N_897,N_840,N_842);
xor U898 (N_898,N_838,N_834);
or U899 (N_899,N_837,N_847);
or U900 (N_900,N_897,N_894);
nor U901 (N_901,N_872,N_891);
nand U902 (N_902,N_887,N_874);
or U903 (N_903,N_866,N_881);
nor U904 (N_904,N_889,N_854);
nor U905 (N_905,N_879,N_867);
nor U906 (N_906,N_864,N_865);
nand U907 (N_907,N_893,N_883);
and U908 (N_908,N_857,N_877);
or U909 (N_909,N_850,N_855);
xor U910 (N_910,N_899,N_861);
nor U911 (N_911,N_878,N_896);
or U912 (N_912,N_860,N_873);
and U913 (N_913,N_856,N_859);
nor U914 (N_914,N_852,N_898);
nor U915 (N_915,N_886,N_892);
nand U916 (N_916,N_875,N_888);
or U917 (N_917,N_869,N_858);
nand U918 (N_918,N_882,N_853);
and U919 (N_919,N_870,N_871);
nand U920 (N_920,N_851,N_880);
nor U921 (N_921,N_884,N_885);
xor U922 (N_922,N_890,N_868);
and U923 (N_923,N_895,N_863);
and U924 (N_924,N_876,N_862);
nand U925 (N_925,N_862,N_875);
and U926 (N_926,N_897,N_862);
or U927 (N_927,N_893,N_898);
nor U928 (N_928,N_890,N_850);
and U929 (N_929,N_880,N_858);
nor U930 (N_930,N_893,N_880);
and U931 (N_931,N_880,N_853);
or U932 (N_932,N_853,N_864);
nor U933 (N_933,N_884,N_858);
nand U934 (N_934,N_868,N_892);
nor U935 (N_935,N_855,N_853);
and U936 (N_936,N_857,N_891);
nor U937 (N_937,N_884,N_896);
xnor U938 (N_938,N_865,N_887);
and U939 (N_939,N_868,N_858);
or U940 (N_940,N_864,N_893);
and U941 (N_941,N_867,N_874);
and U942 (N_942,N_884,N_895);
or U943 (N_943,N_863,N_875);
nand U944 (N_944,N_898,N_882);
nor U945 (N_945,N_864,N_851);
and U946 (N_946,N_875,N_887);
and U947 (N_947,N_879,N_886);
and U948 (N_948,N_885,N_896);
nor U949 (N_949,N_890,N_872);
or U950 (N_950,N_911,N_915);
and U951 (N_951,N_920,N_916);
and U952 (N_952,N_928,N_929);
or U953 (N_953,N_924,N_930);
and U954 (N_954,N_918,N_937);
or U955 (N_955,N_944,N_921);
or U956 (N_956,N_936,N_902);
and U957 (N_957,N_913,N_919);
nor U958 (N_958,N_946,N_917);
and U959 (N_959,N_939,N_900);
nor U960 (N_960,N_904,N_908);
nand U961 (N_961,N_932,N_914);
or U962 (N_962,N_912,N_941);
nor U963 (N_963,N_925,N_927);
nor U964 (N_964,N_910,N_934);
and U965 (N_965,N_909,N_907);
and U966 (N_966,N_922,N_903);
or U967 (N_967,N_931,N_933);
nor U968 (N_968,N_947,N_923);
nand U969 (N_969,N_935,N_901);
or U970 (N_970,N_949,N_948);
nor U971 (N_971,N_926,N_945);
and U972 (N_972,N_905,N_942);
xnor U973 (N_973,N_938,N_940);
or U974 (N_974,N_943,N_906);
nand U975 (N_975,N_930,N_920);
and U976 (N_976,N_949,N_946);
and U977 (N_977,N_937,N_946);
or U978 (N_978,N_937,N_907);
or U979 (N_979,N_901,N_920);
nand U980 (N_980,N_919,N_925);
and U981 (N_981,N_914,N_909);
or U982 (N_982,N_926,N_915);
nor U983 (N_983,N_924,N_948);
nand U984 (N_984,N_926,N_900);
or U985 (N_985,N_925,N_917);
and U986 (N_986,N_926,N_916);
and U987 (N_987,N_921,N_923);
and U988 (N_988,N_900,N_908);
nand U989 (N_989,N_918,N_928);
and U990 (N_990,N_917,N_949);
nor U991 (N_991,N_924,N_922);
and U992 (N_992,N_912,N_927);
and U993 (N_993,N_931,N_935);
and U994 (N_994,N_901,N_944);
or U995 (N_995,N_946,N_945);
and U996 (N_996,N_921,N_905);
nand U997 (N_997,N_947,N_938);
nor U998 (N_998,N_916,N_930);
nand U999 (N_999,N_936,N_946);
nor U1000 (N_1000,N_960,N_987);
and U1001 (N_1001,N_974,N_970);
or U1002 (N_1002,N_986,N_982);
nor U1003 (N_1003,N_989,N_966);
or U1004 (N_1004,N_979,N_988);
nand U1005 (N_1005,N_995,N_993);
nand U1006 (N_1006,N_991,N_997);
nor U1007 (N_1007,N_998,N_975);
nor U1008 (N_1008,N_972,N_965);
or U1009 (N_1009,N_955,N_990);
nand U1010 (N_1010,N_967,N_992);
and U1011 (N_1011,N_951,N_956);
and U1012 (N_1012,N_999,N_964);
and U1013 (N_1013,N_950,N_980);
nand U1014 (N_1014,N_968,N_983);
nor U1015 (N_1015,N_984,N_954);
nor U1016 (N_1016,N_963,N_969);
and U1017 (N_1017,N_976,N_957);
nor U1018 (N_1018,N_977,N_973);
or U1019 (N_1019,N_962,N_952);
nand U1020 (N_1020,N_978,N_961);
nand U1021 (N_1021,N_971,N_996);
or U1022 (N_1022,N_959,N_958);
nand U1023 (N_1023,N_994,N_985);
and U1024 (N_1024,N_981,N_953);
nand U1025 (N_1025,N_950,N_987);
nand U1026 (N_1026,N_969,N_952);
nand U1027 (N_1027,N_986,N_965);
nand U1028 (N_1028,N_952,N_983);
nor U1029 (N_1029,N_963,N_955);
and U1030 (N_1030,N_981,N_971);
nor U1031 (N_1031,N_997,N_970);
nand U1032 (N_1032,N_971,N_964);
and U1033 (N_1033,N_971,N_999);
nor U1034 (N_1034,N_982,N_973);
nor U1035 (N_1035,N_974,N_988);
nor U1036 (N_1036,N_998,N_983);
nor U1037 (N_1037,N_970,N_959);
or U1038 (N_1038,N_990,N_959);
nand U1039 (N_1039,N_955,N_975);
or U1040 (N_1040,N_989,N_986);
and U1041 (N_1041,N_974,N_973);
nand U1042 (N_1042,N_970,N_995);
and U1043 (N_1043,N_954,N_980);
or U1044 (N_1044,N_985,N_997);
and U1045 (N_1045,N_983,N_971);
nor U1046 (N_1046,N_962,N_991);
nor U1047 (N_1047,N_959,N_978);
nand U1048 (N_1048,N_952,N_978);
or U1049 (N_1049,N_999,N_976);
or U1050 (N_1050,N_1014,N_1038);
and U1051 (N_1051,N_1013,N_1031);
or U1052 (N_1052,N_1020,N_1000);
or U1053 (N_1053,N_1027,N_1007);
nand U1054 (N_1054,N_1015,N_1023);
or U1055 (N_1055,N_1035,N_1024);
nor U1056 (N_1056,N_1026,N_1036);
or U1057 (N_1057,N_1029,N_1003);
nor U1058 (N_1058,N_1016,N_1022);
nand U1059 (N_1059,N_1017,N_1009);
nand U1060 (N_1060,N_1010,N_1032);
nand U1061 (N_1061,N_1019,N_1028);
or U1062 (N_1062,N_1034,N_1048);
nand U1063 (N_1063,N_1044,N_1008);
nand U1064 (N_1064,N_1006,N_1001);
xnor U1065 (N_1065,N_1042,N_1049);
nor U1066 (N_1066,N_1012,N_1011);
nand U1067 (N_1067,N_1018,N_1043);
nand U1068 (N_1068,N_1040,N_1025);
nand U1069 (N_1069,N_1033,N_1037);
and U1070 (N_1070,N_1021,N_1002);
nand U1071 (N_1071,N_1041,N_1047);
and U1072 (N_1072,N_1005,N_1045);
nor U1073 (N_1073,N_1004,N_1030);
nor U1074 (N_1074,N_1046,N_1039);
nand U1075 (N_1075,N_1044,N_1010);
or U1076 (N_1076,N_1025,N_1020);
and U1077 (N_1077,N_1010,N_1027);
and U1078 (N_1078,N_1023,N_1005);
nor U1079 (N_1079,N_1024,N_1013);
and U1080 (N_1080,N_1017,N_1043);
nor U1081 (N_1081,N_1012,N_1022);
or U1082 (N_1082,N_1037,N_1043);
nand U1083 (N_1083,N_1021,N_1008);
or U1084 (N_1084,N_1032,N_1049);
nor U1085 (N_1085,N_1049,N_1015);
or U1086 (N_1086,N_1014,N_1005);
nand U1087 (N_1087,N_1043,N_1048);
and U1088 (N_1088,N_1024,N_1018);
and U1089 (N_1089,N_1030,N_1042);
nor U1090 (N_1090,N_1019,N_1043);
nand U1091 (N_1091,N_1004,N_1041);
nand U1092 (N_1092,N_1035,N_1049);
nand U1093 (N_1093,N_1045,N_1016);
xnor U1094 (N_1094,N_1019,N_1000);
nor U1095 (N_1095,N_1034,N_1044);
and U1096 (N_1096,N_1042,N_1032);
nand U1097 (N_1097,N_1036,N_1039);
and U1098 (N_1098,N_1044,N_1015);
or U1099 (N_1099,N_1035,N_1019);
or U1100 (N_1100,N_1085,N_1074);
nor U1101 (N_1101,N_1090,N_1063);
and U1102 (N_1102,N_1093,N_1088);
xnor U1103 (N_1103,N_1064,N_1059);
nand U1104 (N_1104,N_1080,N_1081);
xnor U1105 (N_1105,N_1052,N_1065);
nand U1106 (N_1106,N_1062,N_1071);
and U1107 (N_1107,N_1099,N_1075);
or U1108 (N_1108,N_1061,N_1072);
and U1109 (N_1109,N_1087,N_1069);
nand U1110 (N_1110,N_1051,N_1060);
nor U1111 (N_1111,N_1054,N_1097);
nand U1112 (N_1112,N_1053,N_1098);
nand U1113 (N_1113,N_1055,N_1091);
nand U1114 (N_1114,N_1094,N_1067);
nor U1115 (N_1115,N_1056,N_1057);
or U1116 (N_1116,N_1066,N_1073);
nand U1117 (N_1117,N_1089,N_1083);
nor U1118 (N_1118,N_1086,N_1079);
xor U1119 (N_1119,N_1096,N_1095);
or U1120 (N_1120,N_1050,N_1092);
and U1121 (N_1121,N_1084,N_1078);
nor U1122 (N_1122,N_1082,N_1058);
nor U1123 (N_1123,N_1068,N_1076);
and U1124 (N_1124,N_1077,N_1070);
and U1125 (N_1125,N_1081,N_1059);
nor U1126 (N_1126,N_1079,N_1076);
and U1127 (N_1127,N_1058,N_1065);
nand U1128 (N_1128,N_1067,N_1069);
nand U1129 (N_1129,N_1072,N_1094);
or U1130 (N_1130,N_1058,N_1087);
nor U1131 (N_1131,N_1088,N_1054);
and U1132 (N_1132,N_1098,N_1095);
or U1133 (N_1133,N_1085,N_1099);
nand U1134 (N_1134,N_1093,N_1053);
nor U1135 (N_1135,N_1087,N_1090);
nor U1136 (N_1136,N_1054,N_1066);
nand U1137 (N_1137,N_1081,N_1093);
and U1138 (N_1138,N_1081,N_1054);
nor U1139 (N_1139,N_1099,N_1072);
nand U1140 (N_1140,N_1056,N_1092);
nor U1141 (N_1141,N_1058,N_1056);
nor U1142 (N_1142,N_1059,N_1062);
nand U1143 (N_1143,N_1070,N_1057);
and U1144 (N_1144,N_1079,N_1050);
and U1145 (N_1145,N_1056,N_1065);
nor U1146 (N_1146,N_1066,N_1080);
nor U1147 (N_1147,N_1068,N_1060);
and U1148 (N_1148,N_1077,N_1058);
nor U1149 (N_1149,N_1096,N_1084);
or U1150 (N_1150,N_1116,N_1140);
and U1151 (N_1151,N_1123,N_1104);
or U1152 (N_1152,N_1106,N_1139);
nand U1153 (N_1153,N_1125,N_1114);
or U1154 (N_1154,N_1110,N_1132);
or U1155 (N_1155,N_1128,N_1105);
nor U1156 (N_1156,N_1109,N_1149);
xnor U1157 (N_1157,N_1112,N_1100);
or U1158 (N_1158,N_1145,N_1148);
nand U1159 (N_1159,N_1130,N_1102);
and U1160 (N_1160,N_1103,N_1134);
nand U1161 (N_1161,N_1141,N_1124);
or U1162 (N_1162,N_1138,N_1146);
and U1163 (N_1163,N_1142,N_1101);
nor U1164 (N_1164,N_1147,N_1120);
nor U1165 (N_1165,N_1136,N_1121);
or U1166 (N_1166,N_1144,N_1108);
nand U1167 (N_1167,N_1111,N_1115);
or U1168 (N_1168,N_1133,N_1122);
or U1169 (N_1169,N_1135,N_1131);
or U1170 (N_1170,N_1126,N_1118);
or U1171 (N_1171,N_1143,N_1127);
nand U1172 (N_1172,N_1119,N_1137);
or U1173 (N_1173,N_1107,N_1129);
or U1174 (N_1174,N_1113,N_1117);
and U1175 (N_1175,N_1140,N_1104);
or U1176 (N_1176,N_1126,N_1107);
nor U1177 (N_1177,N_1109,N_1128);
and U1178 (N_1178,N_1106,N_1137);
nor U1179 (N_1179,N_1130,N_1149);
and U1180 (N_1180,N_1114,N_1112);
nor U1181 (N_1181,N_1106,N_1109);
or U1182 (N_1182,N_1102,N_1144);
or U1183 (N_1183,N_1110,N_1139);
nor U1184 (N_1184,N_1134,N_1125);
or U1185 (N_1185,N_1140,N_1128);
or U1186 (N_1186,N_1122,N_1141);
nand U1187 (N_1187,N_1133,N_1147);
nand U1188 (N_1188,N_1135,N_1146);
nand U1189 (N_1189,N_1114,N_1119);
and U1190 (N_1190,N_1126,N_1108);
xor U1191 (N_1191,N_1136,N_1106);
nand U1192 (N_1192,N_1120,N_1128);
or U1193 (N_1193,N_1105,N_1119);
nand U1194 (N_1194,N_1138,N_1119);
nand U1195 (N_1195,N_1111,N_1131);
nor U1196 (N_1196,N_1104,N_1113);
or U1197 (N_1197,N_1130,N_1121);
and U1198 (N_1198,N_1100,N_1102);
or U1199 (N_1199,N_1118,N_1103);
nor U1200 (N_1200,N_1198,N_1169);
nor U1201 (N_1201,N_1183,N_1177);
nand U1202 (N_1202,N_1189,N_1172);
or U1203 (N_1203,N_1196,N_1178);
nand U1204 (N_1204,N_1166,N_1186);
nor U1205 (N_1205,N_1191,N_1175);
nor U1206 (N_1206,N_1182,N_1192);
and U1207 (N_1207,N_1184,N_1168);
xor U1208 (N_1208,N_1150,N_1194);
and U1209 (N_1209,N_1188,N_1187);
and U1210 (N_1210,N_1153,N_1158);
nand U1211 (N_1211,N_1179,N_1159);
or U1212 (N_1212,N_1165,N_1163);
and U1213 (N_1213,N_1157,N_1195);
nor U1214 (N_1214,N_1173,N_1170);
nand U1215 (N_1215,N_1176,N_1164);
nor U1216 (N_1216,N_1199,N_1181);
nor U1217 (N_1217,N_1160,N_1174);
or U1218 (N_1218,N_1167,N_1193);
or U1219 (N_1219,N_1156,N_1180);
and U1220 (N_1220,N_1162,N_1185);
and U1221 (N_1221,N_1197,N_1151);
and U1222 (N_1222,N_1154,N_1161);
and U1223 (N_1223,N_1190,N_1155);
or U1224 (N_1224,N_1152,N_1171);
or U1225 (N_1225,N_1156,N_1174);
or U1226 (N_1226,N_1187,N_1195);
or U1227 (N_1227,N_1155,N_1162);
and U1228 (N_1228,N_1162,N_1178);
nand U1229 (N_1229,N_1195,N_1154);
nand U1230 (N_1230,N_1182,N_1197);
nor U1231 (N_1231,N_1170,N_1172);
nand U1232 (N_1232,N_1191,N_1190);
and U1233 (N_1233,N_1157,N_1150);
nand U1234 (N_1234,N_1167,N_1166);
and U1235 (N_1235,N_1155,N_1164);
nor U1236 (N_1236,N_1171,N_1159);
nor U1237 (N_1237,N_1178,N_1199);
nor U1238 (N_1238,N_1189,N_1184);
or U1239 (N_1239,N_1170,N_1158);
nand U1240 (N_1240,N_1172,N_1171);
nand U1241 (N_1241,N_1190,N_1181);
nor U1242 (N_1242,N_1187,N_1168);
xor U1243 (N_1243,N_1193,N_1198);
and U1244 (N_1244,N_1159,N_1176);
nor U1245 (N_1245,N_1197,N_1155);
nor U1246 (N_1246,N_1175,N_1165);
nor U1247 (N_1247,N_1170,N_1161);
xor U1248 (N_1248,N_1164,N_1152);
nor U1249 (N_1249,N_1154,N_1188);
and U1250 (N_1250,N_1230,N_1214);
or U1251 (N_1251,N_1238,N_1232);
and U1252 (N_1252,N_1206,N_1201);
and U1253 (N_1253,N_1242,N_1215);
nand U1254 (N_1254,N_1234,N_1200);
or U1255 (N_1255,N_1227,N_1244);
and U1256 (N_1256,N_1237,N_1207);
nand U1257 (N_1257,N_1220,N_1225);
and U1258 (N_1258,N_1239,N_1241);
nand U1259 (N_1259,N_1209,N_1208);
or U1260 (N_1260,N_1243,N_1216);
and U1261 (N_1261,N_1247,N_1231);
and U1262 (N_1262,N_1222,N_1226);
nor U1263 (N_1263,N_1246,N_1211);
and U1264 (N_1264,N_1240,N_1228);
nand U1265 (N_1265,N_1212,N_1203);
nor U1266 (N_1266,N_1205,N_1213);
nor U1267 (N_1267,N_1248,N_1245);
nor U1268 (N_1268,N_1221,N_1202);
nor U1269 (N_1269,N_1223,N_1233);
or U1270 (N_1270,N_1229,N_1219);
nand U1271 (N_1271,N_1224,N_1218);
and U1272 (N_1272,N_1210,N_1217);
and U1273 (N_1273,N_1204,N_1235);
and U1274 (N_1274,N_1236,N_1249);
and U1275 (N_1275,N_1217,N_1225);
and U1276 (N_1276,N_1239,N_1225);
nand U1277 (N_1277,N_1225,N_1243);
nor U1278 (N_1278,N_1237,N_1239);
and U1279 (N_1279,N_1214,N_1215);
or U1280 (N_1280,N_1230,N_1206);
nand U1281 (N_1281,N_1216,N_1231);
and U1282 (N_1282,N_1234,N_1235);
xnor U1283 (N_1283,N_1243,N_1203);
nand U1284 (N_1284,N_1231,N_1230);
nor U1285 (N_1285,N_1228,N_1224);
nor U1286 (N_1286,N_1201,N_1228);
nor U1287 (N_1287,N_1244,N_1223);
nor U1288 (N_1288,N_1223,N_1201);
nand U1289 (N_1289,N_1228,N_1248);
nor U1290 (N_1290,N_1227,N_1204);
nand U1291 (N_1291,N_1203,N_1225);
nor U1292 (N_1292,N_1223,N_1245);
nand U1293 (N_1293,N_1227,N_1246);
or U1294 (N_1294,N_1218,N_1217);
nand U1295 (N_1295,N_1244,N_1205);
and U1296 (N_1296,N_1215,N_1230);
nand U1297 (N_1297,N_1246,N_1225);
nand U1298 (N_1298,N_1215,N_1239);
or U1299 (N_1299,N_1208,N_1237);
and U1300 (N_1300,N_1298,N_1272);
or U1301 (N_1301,N_1284,N_1293);
nand U1302 (N_1302,N_1288,N_1269);
and U1303 (N_1303,N_1291,N_1285);
or U1304 (N_1304,N_1264,N_1265);
nor U1305 (N_1305,N_1297,N_1254);
or U1306 (N_1306,N_1250,N_1286);
nand U1307 (N_1307,N_1276,N_1267);
or U1308 (N_1308,N_1252,N_1273);
nor U1309 (N_1309,N_1257,N_1294);
nand U1310 (N_1310,N_1292,N_1253);
nor U1311 (N_1311,N_1299,N_1290);
nand U1312 (N_1312,N_1289,N_1277);
or U1313 (N_1313,N_1260,N_1251);
nand U1314 (N_1314,N_1283,N_1261);
and U1315 (N_1315,N_1259,N_1287);
nand U1316 (N_1316,N_1268,N_1270);
nor U1317 (N_1317,N_1256,N_1271);
or U1318 (N_1318,N_1282,N_1255);
nand U1319 (N_1319,N_1263,N_1275);
or U1320 (N_1320,N_1279,N_1262);
or U1321 (N_1321,N_1281,N_1258);
or U1322 (N_1322,N_1280,N_1274);
nor U1323 (N_1323,N_1296,N_1278);
or U1324 (N_1324,N_1266,N_1295);
nor U1325 (N_1325,N_1264,N_1286);
or U1326 (N_1326,N_1287,N_1276);
nand U1327 (N_1327,N_1257,N_1264);
or U1328 (N_1328,N_1283,N_1282);
and U1329 (N_1329,N_1269,N_1259);
or U1330 (N_1330,N_1288,N_1257);
nor U1331 (N_1331,N_1264,N_1267);
nor U1332 (N_1332,N_1298,N_1283);
nand U1333 (N_1333,N_1279,N_1298);
or U1334 (N_1334,N_1250,N_1273);
or U1335 (N_1335,N_1288,N_1289);
xor U1336 (N_1336,N_1291,N_1275);
nand U1337 (N_1337,N_1270,N_1258);
nor U1338 (N_1338,N_1282,N_1294);
nand U1339 (N_1339,N_1252,N_1263);
nor U1340 (N_1340,N_1277,N_1270);
and U1341 (N_1341,N_1276,N_1292);
or U1342 (N_1342,N_1250,N_1299);
nand U1343 (N_1343,N_1269,N_1262);
nor U1344 (N_1344,N_1265,N_1276);
and U1345 (N_1345,N_1272,N_1289);
nor U1346 (N_1346,N_1292,N_1285);
nor U1347 (N_1347,N_1290,N_1252);
and U1348 (N_1348,N_1264,N_1275);
and U1349 (N_1349,N_1270,N_1296);
or U1350 (N_1350,N_1337,N_1346);
nand U1351 (N_1351,N_1348,N_1329);
or U1352 (N_1352,N_1338,N_1301);
nand U1353 (N_1353,N_1332,N_1327);
nand U1354 (N_1354,N_1323,N_1305);
nor U1355 (N_1355,N_1304,N_1311);
and U1356 (N_1356,N_1321,N_1300);
nand U1357 (N_1357,N_1342,N_1307);
nand U1358 (N_1358,N_1339,N_1345);
nor U1359 (N_1359,N_1316,N_1306);
nand U1360 (N_1360,N_1335,N_1349);
or U1361 (N_1361,N_1318,N_1330);
nand U1362 (N_1362,N_1317,N_1331);
nand U1363 (N_1363,N_1324,N_1309);
nor U1364 (N_1364,N_1344,N_1333);
nor U1365 (N_1365,N_1319,N_1340);
and U1366 (N_1366,N_1313,N_1322);
nand U1367 (N_1367,N_1308,N_1320);
nor U1368 (N_1368,N_1341,N_1343);
nor U1369 (N_1369,N_1325,N_1303);
nor U1370 (N_1370,N_1336,N_1315);
and U1371 (N_1371,N_1334,N_1310);
nand U1372 (N_1372,N_1312,N_1326);
nand U1373 (N_1373,N_1314,N_1302);
and U1374 (N_1374,N_1347,N_1328);
nor U1375 (N_1375,N_1328,N_1321);
nand U1376 (N_1376,N_1325,N_1302);
nor U1377 (N_1377,N_1333,N_1338);
or U1378 (N_1378,N_1333,N_1320);
and U1379 (N_1379,N_1315,N_1323);
nand U1380 (N_1380,N_1336,N_1340);
or U1381 (N_1381,N_1318,N_1335);
nor U1382 (N_1382,N_1342,N_1336);
and U1383 (N_1383,N_1303,N_1343);
or U1384 (N_1384,N_1319,N_1310);
nor U1385 (N_1385,N_1319,N_1324);
and U1386 (N_1386,N_1333,N_1340);
nor U1387 (N_1387,N_1312,N_1348);
or U1388 (N_1388,N_1339,N_1331);
or U1389 (N_1389,N_1329,N_1314);
nand U1390 (N_1390,N_1307,N_1343);
and U1391 (N_1391,N_1335,N_1344);
nand U1392 (N_1392,N_1337,N_1301);
or U1393 (N_1393,N_1310,N_1333);
and U1394 (N_1394,N_1306,N_1315);
and U1395 (N_1395,N_1334,N_1309);
nor U1396 (N_1396,N_1310,N_1307);
and U1397 (N_1397,N_1307,N_1345);
and U1398 (N_1398,N_1305,N_1337);
and U1399 (N_1399,N_1306,N_1323);
nor U1400 (N_1400,N_1386,N_1355);
nor U1401 (N_1401,N_1384,N_1377);
and U1402 (N_1402,N_1391,N_1354);
or U1403 (N_1403,N_1379,N_1387);
and U1404 (N_1404,N_1352,N_1365);
nand U1405 (N_1405,N_1374,N_1364);
nand U1406 (N_1406,N_1388,N_1373);
nand U1407 (N_1407,N_1389,N_1398);
and U1408 (N_1408,N_1359,N_1394);
xnor U1409 (N_1409,N_1353,N_1372);
nand U1410 (N_1410,N_1375,N_1360);
and U1411 (N_1411,N_1362,N_1357);
nand U1412 (N_1412,N_1390,N_1350);
nand U1413 (N_1413,N_1395,N_1399);
nand U1414 (N_1414,N_1383,N_1367);
nand U1415 (N_1415,N_1385,N_1382);
or U1416 (N_1416,N_1366,N_1356);
or U1417 (N_1417,N_1351,N_1361);
and U1418 (N_1418,N_1371,N_1393);
nor U1419 (N_1419,N_1392,N_1358);
and U1420 (N_1420,N_1363,N_1381);
or U1421 (N_1421,N_1380,N_1396);
nor U1422 (N_1422,N_1368,N_1378);
nand U1423 (N_1423,N_1369,N_1370);
xnor U1424 (N_1424,N_1397,N_1376);
nor U1425 (N_1425,N_1382,N_1389);
or U1426 (N_1426,N_1352,N_1399);
or U1427 (N_1427,N_1390,N_1397);
nor U1428 (N_1428,N_1384,N_1393);
or U1429 (N_1429,N_1387,N_1361);
nor U1430 (N_1430,N_1388,N_1358);
or U1431 (N_1431,N_1382,N_1399);
nand U1432 (N_1432,N_1365,N_1358);
nor U1433 (N_1433,N_1385,N_1363);
nand U1434 (N_1434,N_1391,N_1386);
nand U1435 (N_1435,N_1358,N_1359);
nand U1436 (N_1436,N_1366,N_1372);
or U1437 (N_1437,N_1398,N_1360);
xnor U1438 (N_1438,N_1355,N_1389);
nand U1439 (N_1439,N_1360,N_1386);
or U1440 (N_1440,N_1351,N_1367);
and U1441 (N_1441,N_1361,N_1365);
nor U1442 (N_1442,N_1360,N_1354);
nor U1443 (N_1443,N_1375,N_1356);
nor U1444 (N_1444,N_1359,N_1353);
or U1445 (N_1445,N_1377,N_1389);
or U1446 (N_1446,N_1366,N_1367);
or U1447 (N_1447,N_1351,N_1362);
or U1448 (N_1448,N_1365,N_1359);
or U1449 (N_1449,N_1385,N_1397);
or U1450 (N_1450,N_1415,N_1429);
and U1451 (N_1451,N_1438,N_1442);
nand U1452 (N_1452,N_1426,N_1449);
or U1453 (N_1453,N_1440,N_1414);
or U1454 (N_1454,N_1444,N_1420);
nor U1455 (N_1455,N_1407,N_1443);
and U1456 (N_1456,N_1405,N_1412);
nand U1457 (N_1457,N_1427,N_1428);
and U1458 (N_1458,N_1418,N_1421);
and U1459 (N_1459,N_1431,N_1437);
nand U1460 (N_1460,N_1406,N_1441);
nand U1461 (N_1461,N_1417,N_1409);
and U1462 (N_1462,N_1402,N_1425);
or U1463 (N_1463,N_1439,N_1447);
or U1464 (N_1464,N_1413,N_1403);
or U1465 (N_1465,N_1423,N_1445);
nor U1466 (N_1466,N_1424,N_1404);
nor U1467 (N_1467,N_1408,N_1436);
or U1468 (N_1468,N_1434,N_1411);
or U1469 (N_1469,N_1401,N_1416);
xnor U1470 (N_1470,N_1422,N_1410);
or U1471 (N_1471,N_1432,N_1430);
or U1472 (N_1472,N_1433,N_1419);
nand U1473 (N_1473,N_1435,N_1400);
or U1474 (N_1474,N_1446,N_1448);
and U1475 (N_1475,N_1415,N_1422);
or U1476 (N_1476,N_1428,N_1417);
and U1477 (N_1477,N_1446,N_1443);
nor U1478 (N_1478,N_1419,N_1424);
nor U1479 (N_1479,N_1418,N_1444);
nand U1480 (N_1480,N_1435,N_1407);
or U1481 (N_1481,N_1416,N_1423);
nand U1482 (N_1482,N_1418,N_1425);
xor U1483 (N_1483,N_1444,N_1415);
nand U1484 (N_1484,N_1422,N_1414);
and U1485 (N_1485,N_1422,N_1418);
and U1486 (N_1486,N_1408,N_1406);
and U1487 (N_1487,N_1440,N_1422);
nand U1488 (N_1488,N_1441,N_1430);
nand U1489 (N_1489,N_1427,N_1400);
and U1490 (N_1490,N_1437,N_1449);
and U1491 (N_1491,N_1424,N_1438);
nand U1492 (N_1492,N_1443,N_1415);
or U1493 (N_1493,N_1411,N_1417);
nor U1494 (N_1494,N_1418,N_1431);
nand U1495 (N_1495,N_1427,N_1426);
nor U1496 (N_1496,N_1415,N_1438);
and U1497 (N_1497,N_1417,N_1400);
and U1498 (N_1498,N_1433,N_1438);
or U1499 (N_1499,N_1418,N_1447);
nor U1500 (N_1500,N_1478,N_1460);
nand U1501 (N_1501,N_1497,N_1482);
nor U1502 (N_1502,N_1471,N_1458);
or U1503 (N_1503,N_1459,N_1474);
nor U1504 (N_1504,N_1499,N_1451);
or U1505 (N_1505,N_1455,N_1456);
nor U1506 (N_1506,N_1465,N_1463);
and U1507 (N_1507,N_1485,N_1481);
nand U1508 (N_1508,N_1492,N_1462);
nor U1509 (N_1509,N_1498,N_1452);
nand U1510 (N_1510,N_1494,N_1457);
nor U1511 (N_1511,N_1470,N_1484);
nor U1512 (N_1512,N_1486,N_1489);
and U1513 (N_1513,N_1467,N_1477);
nand U1514 (N_1514,N_1475,N_1488);
or U1515 (N_1515,N_1453,N_1472);
or U1516 (N_1516,N_1450,N_1495);
or U1517 (N_1517,N_1491,N_1487);
or U1518 (N_1518,N_1496,N_1461);
and U1519 (N_1519,N_1464,N_1454);
or U1520 (N_1520,N_1490,N_1473);
nor U1521 (N_1521,N_1466,N_1480);
nor U1522 (N_1522,N_1479,N_1469);
and U1523 (N_1523,N_1483,N_1468);
or U1524 (N_1524,N_1493,N_1476);
nand U1525 (N_1525,N_1469,N_1451);
and U1526 (N_1526,N_1496,N_1483);
nor U1527 (N_1527,N_1476,N_1463);
nand U1528 (N_1528,N_1485,N_1491);
and U1529 (N_1529,N_1461,N_1465);
and U1530 (N_1530,N_1474,N_1475);
and U1531 (N_1531,N_1451,N_1456);
and U1532 (N_1532,N_1492,N_1496);
nor U1533 (N_1533,N_1485,N_1486);
and U1534 (N_1534,N_1479,N_1482);
and U1535 (N_1535,N_1487,N_1481);
or U1536 (N_1536,N_1450,N_1469);
nor U1537 (N_1537,N_1456,N_1462);
nand U1538 (N_1538,N_1464,N_1497);
nor U1539 (N_1539,N_1469,N_1463);
nor U1540 (N_1540,N_1460,N_1470);
or U1541 (N_1541,N_1472,N_1498);
nor U1542 (N_1542,N_1496,N_1498);
nor U1543 (N_1543,N_1457,N_1455);
and U1544 (N_1544,N_1493,N_1491);
nand U1545 (N_1545,N_1462,N_1469);
xor U1546 (N_1546,N_1456,N_1485);
nor U1547 (N_1547,N_1487,N_1460);
and U1548 (N_1548,N_1462,N_1486);
nor U1549 (N_1549,N_1482,N_1498);
nand U1550 (N_1550,N_1501,N_1537);
or U1551 (N_1551,N_1506,N_1527);
or U1552 (N_1552,N_1514,N_1544);
nand U1553 (N_1553,N_1510,N_1534);
nor U1554 (N_1554,N_1531,N_1542);
nand U1555 (N_1555,N_1549,N_1536);
and U1556 (N_1556,N_1508,N_1504);
nor U1557 (N_1557,N_1511,N_1543);
nor U1558 (N_1558,N_1546,N_1532);
or U1559 (N_1559,N_1512,N_1526);
nand U1560 (N_1560,N_1513,N_1545);
xor U1561 (N_1561,N_1541,N_1548);
xnor U1562 (N_1562,N_1516,N_1539);
nand U1563 (N_1563,N_1503,N_1540);
nand U1564 (N_1564,N_1509,N_1529);
or U1565 (N_1565,N_1528,N_1547);
nor U1566 (N_1566,N_1530,N_1507);
nand U1567 (N_1567,N_1533,N_1523);
nand U1568 (N_1568,N_1538,N_1517);
and U1569 (N_1569,N_1518,N_1519);
or U1570 (N_1570,N_1515,N_1524);
nor U1571 (N_1571,N_1525,N_1521);
or U1572 (N_1572,N_1520,N_1502);
nand U1573 (N_1573,N_1505,N_1500);
and U1574 (N_1574,N_1522,N_1535);
and U1575 (N_1575,N_1513,N_1535);
or U1576 (N_1576,N_1523,N_1515);
nor U1577 (N_1577,N_1506,N_1504);
and U1578 (N_1578,N_1542,N_1510);
nor U1579 (N_1579,N_1547,N_1503);
and U1580 (N_1580,N_1501,N_1525);
nor U1581 (N_1581,N_1536,N_1542);
or U1582 (N_1582,N_1516,N_1537);
nand U1583 (N_1583,N_1534,N_1505);
and U1584 (N_1584,N_1506,N_1544);
nand U1585 (N_1585,N_1530,N_1528);
nor U1586 (N_1586,N_1525,N_1536);
nor U1587 (N_1587,N_1544,N_1528);
or U1588 (N_1588,N_1536,N_1500);
and U1589 (N_1589,N_1540,N_1547);
nand U1590 (N_1590,N_1502,N_1522);
or U1591 (N_1591,N_1529,N_1541);
nor U1592 (N_1592,N_1529,N_1543);
nand U1593 (N_1593,N_1528,N_1507);
or U1594 (N_1594,N_1503,N_1509);
nor U1595 (N_1595,N_1540,N_1526);
or U1596 (N_1596,N_1540,N_1536);
nor U1597 (N_1597,N_1536,N_1506);
and U1598 (N_1598,N_1543,N_1525);
xor U1599 (N_1599,N_1546,N_1537);
and U1600 (N_1600,N_1589,N_1584);
or U1601 (N_1601,N_1578,N_1566);
and U1602 (N_1602,N_1590,N_1565);
and U1603 (N_1603,N_1568,N_1594);
and U1604 (N_1604,N_1570,N_1554);
nor U1605 (N_1605,N_1579,N_1551);
nand U1606 (N_1606,N_1599,N_1556);
nand U1607 (N_1607,N_1583,N_1591);
nor U1608 (N_1608,N_1552,N_1564);
nand U1609 (N_1609,N_1575,N_1581);
or U1610 (N_1610,N_1576,N_1595);
or U1611 (N_1611,N_1557,N_1598);
and U1612 (N_1612,N_1593,N_1587);
nor U1613 (N_1613,N_1550,N_1553);
or U1614 (N_1614,N_1592,N_1574);
nor U1615 (N_1615,N_1597,N_1569);
and U1616 (N_1616,N_1559,N_1571);
nor U1617 (N_1617,N_1596,N_1558);
and U1618 (N_1618,N_1573,N_1580);
or U1619 (N_1619,N_1588,N_1586);
and U1620 (N_1620,N_1562,N_1555);
nand U1621 (N_1621,N_1572,N_1567);
nand U1622 (N_1622,N_1585,N_1577);
and U1623 (N_1623,N_1582,N_1563);
and U1624 (N_1624,N_1561,N_1560);
nand U1625 (N_1625,N_1574,N_1564);
or U1626 (N_1626,N_1552,N_1589);
and U1627 (N_1627,N_1594,N_1560);
and U1628 (N_1628,N_1562,N_1579);
nand U1629 (N_1629,N_1578,N_1573);
nor U1630 (N_1630,N_1580,N_1596);
nand U1631 (N_1631,N_1584,N_1583);
or U1632 (N_1632,N_1570,N_1599);
nand U1633 (N_1633,N_1566,N_1586);
or U1634 (N_1634,N_1565,N_1555);
or U1635 (N_1635,N_1597,N_1592);
xor U1636 (N_1636,N_1552,N_1578);
and U1637 (N_1637,N_1563,N_1584);
or U1638 (N_1638,N_1571,N_1582);
or U1639 (N_1639,N_1578,N_1564);
and U1640 (N_1640,N_1577,N_1554);
and U1641 (N_1641,N_1569,N_1572);
nand U1642 (N_1642,N_1569,N_1580);
nand U1643 (N_1643,N_1595,N_1597);
nand U1644 (N_1644,N_1559,N_1573);
nand U1645 (N_1645,N_1562,N_1599);
xnor U1646 (N_1646,N_1593,N_1556);
nand U1647 (N_1647,N_1595,N_1586);
or U1648 (N_1648,N_1595,N_1553);
and U1649 (N_1649,N_1593,N_1597);
nor U1650 (N_1650,N_1618,N_1605);
nand U1651 (N_1651,N_1644,N_1641);
and U1652 (N_1652,N_1602,N_1633);
or U1653 (N_1653,N_1613,N_1627);
and U1654 (N_1654,N_1634,N_1608);
and U1655 (N_1655,N_1604,N_1630);
nor U1656 (N_1656,N_1611,N_1623);
nand U1657 (N_1657,N_1624,N_1635);
nor U1658 (N_1658,N_1615,N_1637);
or U1659 (N_1659,N_1600,N_1648);
or U1660 (N_1660,N_1601,N_1638);
or U1661 (N_1661,N_1629,N_1610);
nor U1662 (N_1662,N_1616,N_1603);
nor U1663 (N_1663,N_1639,N_1646);
nand U1664 (N_1664,N_1621,N_1625);
nor U1665 (N_1665,N_1607,N_1642);
xor U1666 (N_1666,N_1612,N_1626);
or U1667 (N_1667,N_1645,N_1640);
and U1668 (N_1668,N_1606,N_1614);
nor U1669 (N_1669,N_1643,N_1649);
nand U1670 (N_1670,N_1619,N_1636);
nand U1671 (N_1671,N_1631,N_1609);
nor U1672 (N_1672,N_1632,N_1647);
nor U1673 (N_1673,N_1617,N_1628);
or U1674 (N_1674,N_1620,N_1622);
nor U1675 (N_1675,N_1639,N_1645);
and U1676 (N_1676,N_1616,N_1628);
nor U1677 (N_1677,N_1634,N_1630);
and U1678 (N_1678,N_1623,N_1635);
and U1679 (N_1679,N_1633,N_1607);
nand U1680 (N_1680,N_1629,N_1624);
nand U1681 (N_1681,N_1649,N_1636);
and U1682 (N_1682,N_1602,N_1613);
or U1683 (N_1683,N_1633,N_1639);
nand U1684 (N_1684,N_1607,N_1604);
and U1685 (N_1685,N_1638,N_1649);
nor U1686 (N_1686,N_1645,N_1609);
nand U1687 (N_1687,N_1602,N_1639);
nand U1688 (N_1688,N_1615,N_1648);
nand U1689 (N_1689,N_1633,N_1640);
and U1690 (N_1690,N_1610,N_1649);
or U1691 (N_1691,N_1607,N_1608);
nand U1692 (N_1692,N_1618,N_1602);
or U1693 (N_1693,N_1621,N_1631);
or U1694 (N_1694,N_1613,N_1622);
nor U1695 (N_1695,N_1640,N_1605);
and U1696 (N_1696,N_1637,N_1626);
nor U1697 (N_1697,N_1626,N_1620);
nor U1698 (N_1698,N_1601,N_1604);
or U1699 (N_1699,N_1618,N_1604);
nor U1700 (N_1700,N_1663,N_1695);
nor U1701 (N_1701,N_1651,N_1671);
or U1702 (N_1702,N_1686,N_1653);
and U1703 (N_1703,N_1657,N_1658);
and U1704 (N_1704,N_1661,N_1660);
or U1705 (N_1705,N_1685,N_1679);
or U1706 (N_1706,N_1673,N_1662);
nand U1707 (N_1707,N_1693,N_1699);
or U1708 (N_1708,N_1670,N_1692);
nand U1709 (N_1709,N_1681,N_1683);
and U1710 (N_1710,N_1665,N_1694);
nand U1711 (N_1711,N_1652,N_1691);
and U1712 (N_1712,N_1659,N_1678);
nor U1713 (N_1713,N_1677,N_1680);
nand U1714 (N_1714,N_1682,N_1668);
and U1715 (N_1715,N_1689,N_1666);
or U1716 (N_1716,N_1684,N_1697);
or U1717 (N_1717,N_1676,N_1655);
nor U1718 (N_1718,N_1656,N_1690);
nand U1719 (N_1719,N_1698,N_1669);
nand U1720 (N_1720,N_1667,N_1687);
or U1721 (N_1721,N_1696,N_1672);
or U1722 (N_1722,N_1674,N_1664);
and U1723 (N_1723,N_1654,N_1675);
nor U1724 (N_1724,N_1650,N_1688);
or U1725 (N_1725,N_1658,N_1672);
or U1726 (N_1726,N_1653,N_1685);
nor U1727 (N_1727,N_1690,N_1650);
nand U1728 (N_1728,N_1689,N_1672);
or U1729 (N_1729,N_1681,N_1674);
nor U1730 (N_1730,N_1682,N_1693);
and U1731 (N_1731,N_1684,N_1654);
and U1732 (N_1732,N_1693,N_1667);
and U1733 (N_1733,N_1685,N_1668);
and U1734 (N_1734,N_1691,N_1659);
or U1735 (N_1735,N_1697,N_1661);
and U1736 (N_1736,N_1653,N_1684);
nor U1737 (N_1737,N_1653,N_1665);
and U1738 (N_1738,N_1654,N_1662);
or U1739 (N_1739,N_1661,N_1655);
or U1740 (N_1740,N_1688,N_1683);
and U1741 (N_1741,N_1658,N_1666);
xnor U1742 (N_1742,N_1665,N_1697);
and U1743 (N_1743,N_1676,N_1661);
and U1744 (N_1744,N_1662,N_1678);
and U1745 (N_1745,N_1688,N_1694);
or U1746 (N_1746,N_1664,N_1661);
nor U1747 (N_1747,N_1685,N_1659);
nor U1748 (N_1748,N_1660,N_1685);
nor U1749 (N_1749,N_1691,N_1653);
nor U1750 (N_1750,N_1734,N_1708);
or U1751 (N_1751,N_1705,N_1739);
or U1752 (N_1752,N_1730,N_1706);
and U1753 (N_1753,N_1726,N_1745);
and U1754 (N_1754,N_1728,N_1744);
and U1755 (N_1755,N_1723,N_1743);
nand U1756 (N_1756,N_1740,N_1719);
nor U1757 (N_1757,N_1732,N_1749);
and U1758 (N_1758,N_1713,N_1735);
or U1759 (N_1759,N_1701,N_1725);
nor U1760 (N_1760,N_1727,N_1709);
nor U1761 (N_1761,N_1747,N_1733);
and U1762 (N_1762,N_1711,N_1717);
and U1763 (N_1763,N_1738,N_1704);
or U1764 (N_1764,N_1746,N_1721);
nand U1765 (N_1765,N_1714,N_1715);
or U1766 (N_1766,N_1710,N_1748);
or U1767 (N_1767,N_1720,N_1712);
xor U1768 (N_1768,N_1702,N_1722);
nand U1769 (N_1769,N_1700,N_1731);
and U1770 (N_1770,N_1724,N_1729);
nor U1771 (N_1771,N_1707,N_1736);
nor U1772 (N_1772,N_1741,N_1716);
nand U1773 (N_1773,N_1737,N_1718);
xor U1774 (N_1774,N_1742,N_1703);
nor U1775 (N_1775,N_1722,N_1731);
nand U1776 (N_1776,N_1714,N_1731);
nor U1777 (N_1777,N_1716,N_1705);
nor U1778 (N_1778,N_1737,N_1724);
or U1779 (N_1779,N_1714,N_1745);
and U1780 (N_1780,N_1744,N_1707);
or U1781 (N_1781,N_1744,N_1708);
nor U1782 (N_1782,N_1714,N_1718);
and U1783 (N_1783,N_1741,N_1711);
nor U1784 (N_1784,N_1713,N_1748);
nor U1785 (N_1785,N_1748,N_1722);
nand U1786 (N_1786,N_1723,N_1705);
and U1787 (N_1787,N_1724,N_1722);
and U1788 (N_1788,N_1744,N_1703);
nand U1789 (N_1789,N_1745,N_1744);
and U1790 (N_1790,N_1723,N_1706);
and U1791 (N_1791,N_1737,N_1744);
or U1792 (N_1792,N_1741,N_1747);
or U1793 (N_1793,N_1734,N_1722);
or U1794 (N_1794,N_1716,N_1724);
nor U1795 (N_1795,N_1703,N_1722);
nand U1796 (N_1796,N_1746,N_1706);
nor U1797 (N_1797,N_1716,N_1723);
nand U1798 (N_1798,N_1747,N_1714);
and U1799 (N_1799,N_1737,N_1710);
and U1800 (N_1800,N_1760,N_1755);
nor U1801 (N_1801,N_1758,N_1779);
or U1802 (N_1802,N_1790,N_1782);
or U1803 (N_1803,N_1791,N_1781);
and U1804 (N_1804,N_1795,N_1773);
or U1805 (N_1805,N_1759,N_1789);
and U1806 (N_1806,N_1785,N_1769);
nor U1807 (N_1807,N_1761,N_1770);
xor U1808 (N_1808,N_1757,N_1774);
or U1809 (N_1809,N_1772,N_1797);
or U1810 (N_1810,N_1777,N_1762);
nand U1811 (N_1811,N_1756,N_1778);
nand U1812 (N_1812,N_1796,N_1794);
nand U1813 (N_1813,N_1788,N_1799);
and U1814 (N_1814,N_1751,N_1798);
and U1815 (N_1815,N_1771,N_1765);
nor U1816 (N_1816,N_1753,N_1775);
and U1817 (N_1817,N_1786,N_1754);
xnor U1818 (N_1818,N_1780,N_1783);
nand U1819 (N_1819,N_1763,N_1767);
nor U1820 (N_1820,N_1752,N_1793);
and U1821 (N_1821,N_1776,N_1766);
nor U1822 (N_1822,N_1764,N_1750);
nand U1823 (N_1823,N_1784,N_1792);
nor U1824 (N_1824,N_1787,N_1768);
or U1825 (N_1825,N_1753,N_1778);
and U1826 (N_1826,N_1796,N_1774);
nor U1827 (N_1827,N_1763,N_1762);
or U1828 (N_1828,N_1754,N_1777);
and U1829 (N_1829,N_1778,N_1769);
nand U1830 (N_1830,N_1796,N_1791);
and U1831 (N_1831,N_1760,N_1758);
and U1832 (N_1832,N_1751,N_1787);
or U1833 (N_1833,N_1793,N_1753);
nor U1834 (N_1834,N_1751,N_1781);
or U1835 (N_1835,N_1778,N_1788);
nand U1836 (N_1836,N_1787,N_1799);
or U1837 (N_1837,N_1786,N_1782);
nor U1838 (N_1838,N_1759,N_1771);
nand U1839 (N_1839,N_1791,N_1769);
or U1840 (N_1840,N_1798,N_1789);
or U1841 (N_1841,N_1771,N_1790);
nand U1842 (N_1842,N_1781,N_1799);
and U1843 (N_1843,N_1751,N_1791);
nor U1844 (N_1844,N_1782,N_1780);
xor U1845 (N_1845,N_1755,N_1779);
and U1846 (N_1846,N_1772,N_1763);
nand U1847 (N_1847,N_1756,N_1794);
nand U1848 (N_1848,N_1760,N_1761);
nand U1849 (N_1849,N_1763,N_1777);
nor U1850 (N_1850,N_1825,N_1803);
nor U1851 (N_1851,N_1800,N_1831);
nor U1852 (N_1852,N_1812,N_1849);
xor U1853 (N_1853,N_1845,N_1819);
nand U1854 (N_1854,N_1814,N_1817);
nor U1855 (N_1855,N_1844,N_1821);
or U1856 (N_1856,N_1826,N_1805);
or U1857 (N_1857,N_1833,N_1824);
or U1858 (N_1858,N_1811,N_1801);
nor U1859 (N_1859,N_1835,N_1830);
or U1860 (N_1860,N_1807,N_1809);
nand U1861 (N_1861,N_1816,N_1829);
nand U1862 (N_1862,N_1839,N_1823);
nor U1863 (N_1863,N_1843,N_1846);
or U1864 (N_1864,N_1818,N_1827);
nor U1865 (N_1865,N_1841,N_1806);
and U1866 (N_1866,N_1834,N_1832);
nor U1867 (N_1867,N_1804,N_1836);
and U1868 (N_1868,N_1820,N_1822);
or U1869 (N_1869,N_1802,N_1828);
and U1870 (N_1870,N_1815,N_1847);
nand U1871 (N_1871,N_1808,N_1842);
and U1872 (N_1872,N_1837,N_1838);
and U1873 (N_1873,N_1840,N_1848);
or U1874 (N_1874,N_1813,N_1810);
and U1875 (N_1875,N_1810,N_1809);
and U1876 (N_1876,N_1806,N_1834);
and U1877 (N_1877,N_1825,N_1805);
and U1878 (N_1878,N_1828,N_1812);
and U1879 (N_1879,N_1824,N_1846);
nor U1880 (N_1880,N_1806,N_1822);
and U1881 (N_1881,N_1841,N_1837);
and U1882 (N_1882,N_1826,N_1831);
or U1883 (N_1883,N_1845,N_1801);
and U1884 (N_1884,N_1829,N_1849);
or U1885 (N_1885,N_1820,N_1825);
nor U1886 (N_1886,N_1824,N_1832);
and U1887 (N_1887,N_1823,N_1816);
and U1888 (N_1888,N_1820,N_1817);
or U1889 (N_1889,N_1828,N_1839);
and U1890 (N_1890,N_1808,N_1815);
or U1891 (N_1891,N_1825,N_1828);
nor U1892 (N_1892,N_1828,N_1844);
nand U1893 (N_1893,N_1843,N_1831);
nor U1894 (N_1894,N_1817,N_1812);
or U1895 (N_1895,N_1819,N_1849);
nor U1896 (N_1896,N_1817,N_1805);
and U1897 (N_1897,N_1824,N_1849);
nor U1898 (N_1898,N_1813,N_1848);
and U1899 (N_1899,N_1802,N_1827);
or U1900 (N_1900,N_1879,N_1891);
nand U1901 (N_1901,N_1857,N_1860);
nor U1902 (N_1902,N_1858,N_1877);
and U1903 (N_1903,N_1853,N_1855);
or U1904 (N_1904,N_1887,N_1882);
nor U1905 (N_1905,N_1897,N_1890);
nand U1906 (N_1906,N_1868,N_1850);
nand U1907 (N_1907,N_1856,N_1863);
or U1908 (N_1908,N_1852,N_1867);
nor U1909 (N_1909,N_1885,N_1871);
nand U1910 (N_1910,N_1886,N_1872);
and U1911 (N_1911,N_1876,N_1892);
and U1912 (N_1912,N_1894,N_1875);
and U1913 (N_1913,N_1883,N_1866);
nand U1914 (N_1914,N_1864,N_1896);
or U1915 (N_1915,N_1873,N_1895);
nor U1916 (N_1916,N_1854,N_1869);
nor U1917 (N_1917,N_1884,N_1870);
nand U1918 (N_1918,N_1861,N_1880);
and U1919 (N_1919,N_1899,N_1881);
nand U1920 (N_1920,N_1851,N_1865);
nor U1921 (N_1921,N_1889,N_1898);
or U1922 (N_1922,N_1874,N_1888);
nand U1923 (N_1923,N_1859,N_1862);
nor U1924 (N_1924,N_1893,N_1878);
or U1925 (N_1925,N_1895,N_1852);
nand U1926 (N_1926,N_1851,N_1897);
or U1927 (N_1927,N_1876,N_1859);
or U1928 (N_1928,N_1894,N_1893);
nand U1929 (N_1929,N_1850,N_1875);
or U1930 (N_1930,N_1862,N_1867);
nor U1931 (N_1931,N_1898,N_1891);
and U1932 (N_1932,N_1881,N_1858);
and U1933 (N_1933,N_1855,N_1852);
or U1934 (N_1934,N_1891,N_1895);
and U1935 (N_1935,N_1867,N_1890);
nor U1936 (N_1936,N_1881,N_1895);
nor U1937 (N_1937,N_1881,N_1859);
and U1938 (N_1938,N_1852,N_1858);
nand U1939 (N_1939,N_1899,N_1892);
and U1940 (N_1940,N_1889,N_1896);
or U1941 (N_1941,N_1882,N_1872);
nor U1942 (N_1942,N_1862,N_1896);
and U1943 (N_1943,N_1897,N_1857);
and U1944 (N_1944,N_1874,N_1891);
or U1945 (N_1945,N_1884,N_1873);
nor U1946 (N_1946,N_1898,N_1874);
or U1947 (N_1947,N_1858,N_1882);
and U1948 (N_1948,N_1868,N_1857);
nand U1949 (N_1949,N_1856,N_1857);
and U1950 (N_1950,N_1914,N_1940);
or U1951 (N_1951,N_1900,N_1925);
nand U1952 (N_1952,N_1934,N_1935);
nand U1953 (N_1953,N_1917,N_1938);
nand U1954 (N_1954,N_1910,N_1939);
and U1955 (N_1955,N_1936,N_1928);
nor U1956 (N_1956,N_1937,N_1918);
nand U1957 (N_1957,N_1924,N_1926);
or U1958 (N_1958,N_1945,N_1944);
or U1959 (N_1959,N_1908,N_1904);
nor U1960 (N_1960,N_1946,N_1916);
or U1961 (N_1961,N_1920,N_1933);
nor U1962 (N_1962,N_1941,N_1948);
and U1963 (N_1963,N_1906,N_1922);
nand U1964 (N_1964,N_1947,N_1927);
nand U1965 (N_1965,N_1911,N_1905);
nand U1966 (N_1966,N_1931,N_1949);
nor U1967 (N_1967,N_1929,N_1915);
or U1968 (N_1968,N_1943,N_1932);
nand U1969 (N_1969,N_1907,N_1902);
nand U1970 (N_1970,N_1912,N_1909);
nand U1971 (N_1971,N_1921,N_1901);
nor U1972 (N_1972,N_1942,N_1919);
xor U1973 (N_1973,N_1913,N_1923);
and U1974 (N_1974,N_1930,N_1903);
nor U1975 (N_1975,N_1939,N_1913);
xnor U1976 (N_1976,N_1938,N_1904);
nor U1977 (N_1977,N_1906,N_1900);
or U1978 (N_1978,N_1925,N_1940);
nor U1979 (N_1979,N_1924,N_1905);
or U1980 (N_1980,N_1932,N_1917);
nor U1981 (N_1981,N_1901,N_1900);
nand U1982 (N_1982,N_1917,N_1923);
nor U1983 (N_1983,N_1930,N_1906);
nor U1984 (N_1984,N_1915,N_1949);
nor U1985 (N_1985,N_1921,N_1903);
xnor U1986 (N_1986,N_1904,N_1942);
nor U1987 (N_1987,N_1935,N_1944);
nand U1988 (N_1988,N_1935,N_1931);
or U1989 (N_1989,N_1934,N_1943);
or U1990 (N_1990,N_1917,N_1918);
nor U1991 (N_1991,N_1912,N_1906);
nand U1992 (N_1992,N_1929,N_1917);
and U1993 (N_1993,N_1945,N_1941);
or U1994 (N_1994,N_1948,N_1909);
nand U1995 (N_1995,N_1945,N_1949);
nor U1996 (N_1996,N_1930,N_1922);
nand U1997 (N_1997,N_1916,N_1904);
xnor U1998 (N_1998,N_1936,N_1919);
and U1999 (N_1999,N_1926,N_1904);
and U2000 (N_2000,N_1959,N_1972);
nand U2001 (N_2001,N_1988,N_1955);
nand U2002 (N_2002,N_1980,N_1984);
and U2003 (N_2003,N_1956,N_1957);
and U2004 (N_2004,N_1982,N_1964);
xor U2005 (N_2005,N_1998,N_1970);
nand U2006 (N_2006,N_1963,N_1960);
and U2007 (N_2007,N_1958,N_1950);
nand U2008 (N_2008,N_1994,N_1990);
nor U2009 (N_2009,N_1951,N_1997);
nand U2010 (N_2010,N_1953,N_1952);
nor U2011 (N_2011,N_1999,N_1996);
or U2012 (N_2012,N_1979,N_1976);
nand U2013 (N_2013,N_1962,N_1961);
and U2014 (N_2014,N_1966,N_1985);
nand U2015 (N_2015,N_1971,N_1967);
nand U2016 (N_2016,N_1983,N_1954);
or U2017 (N_2017,N_1974,N_1993);
or U2018 (N_2018,N_1986,N_1995);
or U2019 (N_2019,N_1969,N_1973);
and U2020 (N_2020,N_1975,N_1992);
nor U2021 (N_2021,N_1968,N_1977);
xnor U2022 (N_2022,N_1981,N_1965);
and U2023 (N_2023,N_1978,N_1991);
nor U2024 (N_2024,N_1987,N_1989);
and U2025 (N_2025,N_1964,N_1951);
and U2026 (N_2026,N_1988,N_1974);
or U2027 (N_2027,N_1992,N_1950);
nand U2028 (N_2028,N_1969,N_1966);
and U2029 (N_2029,N_1970,N_1980);
and U2030 (N_2030,N_1972,N_1953);
nor U2031 (N_2031,N_1973,N_1980);
nor U2032 (N_2032,N_1978,N_1975);
nand U2033 (N_2033,N_1971,N_1998);
and U2034 (N_2034,N_1982,N_1998);
or U2035 (N_2035,N_1969,N_1971);
nand U2036 (N_2036,N_1995,N_1952);
nand U2037 (N_2037,N_1993,N_1962);
or U2038 (N_2038,N_1966,N_1986);
and U2039 (N_2039,N_1953,N_1999);
or U2040 (N_2040,N_1986,N_1994);
nor U2041 (N_2041,N_1968,N_1965);
nand U2042 (N_2042,N_1967,N_1972);
nand U2043 (N_2043,N_1991,N_1962);
nor U2044 (N_2044,N_1989,N_1954);
and U2045 (N_2045,N_1960,N_1956);
xnor U2046 (N_2046,N_1955,N_1974);
nor U2047 (N_2047,N_1961,N_1993);
nor U2048 (N_2048,N_1973,N_1957);
or U2049 (N_2049,N_1970,N_1978);
and U2050 (N_2050,N_2013,N_2015);
nor U2051 (N_2051,N_2005,N_2012);
and U2052 (N_2052,N_2016,N_2039);
or U2053 (N_2053,N_2043,N_2019);
nor U2054 (N_2054,N_2007,N_2020);
or U2055 (N_2055,N_2008,N_2028);
and U2056 (N_2056,N_2034,N_2002);
nand U2057 (N_2057,N_2011,N_2029);
or U2058 (N_2058,N_2025,N_2040);
or U2059 (N_2059,N_2044,N_2010);
or U2060 (N_2060,N_2026,N_2018);
nand U2061 (N_2061,N_2009,N_2037);
or U2062 (N_2062,N_2006,N_2048);
or U2063 (N_2063,N_2047,N_2030);
nor U2064 (N_2064,N_2036,N_2035);
and U2065 (N_2065,N_2049,N_2038);
and U2066 (N_2066,N_2045,N_2004);
nor U2067 (N_2067,N_2032,N_2000);
or U2068 (N_2068,N_2042,N_2023);
and U2069 (N_2069,N_2031,N_2003);
and U2070 (N_2070,N_2021,N_2022);
or U2071 (N_2071,N_2033,N_2001);
and U2072 (N_2072,N_2027,N_2017);
nor U2073 (N_2073,N_2046,N_2041);
or U2074 (N_2074,N_2014,N_2024);
nor U2075 (N_2075,N_2042,N_2028);
and U2076 (N_2076,N_2020,N_2011);
and U2077 (N_2077,N_2027,N_2043);
nand U2078 (N_2078,N_2042,N_2037);
or U2079 (N_2079,N_2036,N_2009);
nand U2080 (N_2080,N_2016,N_2040);
nand U2081 (N_2081,N_2018,N_2016);
and U2082 (N_2082,N_2004,N_2002);
and U2083 (N_2083,N_2010,N_2012);
nor U2084 (N_2084,N_2009,N_2012);
or U2085 (N_2085,N_2023,N_2011);
nor U2086 (N_2086,N_2023,N_2035);
and U2087 (N_2087,N_2005,N_2038);
nor U2088 (N_2088,N_2024,N_2002);
nand U2089 (N_2089,N_2035,N_2022);
nand U2090 (N_2090,N_2044,N_2024);
xor U2091 (N_2091,N_2044,N_2037);
nand U2092 (N_2092,N_2013,N_2003);
and U2093 (N_2093,N_2015,N_2036);
and U2094 (N_2094,N_2015,N_2030);
nor U2095 (N_2095,N_2002,N_2046);
nand U2096 (N_2096,N_2042,N_2041);
nor U2097 (N_2097,N_2026,N_2008);
nand U2098 (N_2098,N_2010,N_2030);
and U2099 (N_2099,N_2028,N_2019);
nand U2100 (N_2100,N_2074,N_2085);
xnor U2101 (N_2101,N_2051,N_2082);
or U2102 (N_2102,N_2078,N_2055);
xnor U2103 (N_2103,N_2096,N_2073);
xnor U2104 (N_2104,N_2083,N_2068);
or U2105 (N_2105,N_2091,N_2097);
or U2106 (N_2106,N_2056,N_2067);
nand U2107 (N_2107,N_2066,N_2063);
or U2108 (N_2108,N_2098,N_2072);
and U2109 (N_2109,N_2095,N_2093);
nor U2110 (N_2110,N_2092,N_2065);
xnor U2111 (N_2111,N_2088,N_2086);
xnor U2112 (N_2112,N_2058,N_2079);
or U2113 (N_2113,N_2080,N_2069);
or U2114 (N_2114,N_2060,N_2081);
nor U2115 (N_2115,N_2094,N_2071);
or U2116 (N_2116,N_2084,N_2059);
nor U2117 (N_2117,N_2070,N_2076);
nor U2118 (N_2118,N_2057,N_2087);
and U2119 (N_2119,N_2090,N_2064);
nor U2120 (N_2120,N_2089,N_2062);
nor U2121 (N_2121,N_2054,N_2050);
and U2122 (N_2122,N_2075,N_2099);
and U2123 (N_2123,N_2053,N_2061);
xor U2124 (N_2124,N_2052,N_2077);
and U2125 (N_2125,N_2097,N_2059);
nand U2126 (N_2126,N_2063,N_2097);
or U2127 (N_2127,N_2082,N_2070);
nor U2128 (N_2128,N_2079,N_2070);
and U2129 (N_2129,N_2093,N_2077);
and U2130 (N_2130,N_2050,N_2061);
and U2131 (N_2131,N_2074,N_2075);
nand U2132 (N_2132,N_2076,N_2087);
or U2133 (N_2133,N_2086,N_2052);
or U2134 (N_2134,N_2066,N_2092);
nand U2135 (N_2135,N_2052,N_2099);
nand U2136 (N_2136,N_2072,N_2052);
and U2137 (N_2137,N_2053,N_2079);
nor U2138 (N_2138,N_2086,N_2096);
nand U2139 (N_2139,N_2066,N_2094);
and U2140 (N_2140,N_2095,N_2083);
and U2141 (N_2141,N_2051,N_2099);
nand U2142 (N_2142,N_2056,N_2077);
or U2143 (N_2143,N_2095,N_2055);
nand U2144 (N_2144,N_2071,N_2067);
and U2145 (N_2145,N_2091,N_2098);
xor U2146 (N_2146,N_2075,N_2078);
nand U2147 (N_2147,N_2069,N_2057);
nand U2148 (N_2148,N_2069,N_2094);
nand U2149 (N_2149,N_2060,N_2052);
nor U2150 (N_2150,N_2110,N_2114);
nand U2151 (N_2151,N_2109,N_2142);
nor U2152 (N_2152,N_2141,N_2148);
and U2153 (N_2153,N_2104,N_2107);
nand U2154 (N_2154,N_2130,N_2127);
nor U2155 (N_2155,N_2125,N_2146);
and U2156 (N_2156,N_2108,N_2118);
and U2157 (N_2157,N_2105,N_2120);
and U2158 (N_2158,N_2111,N_2133);
and U2159 (N_2159,N_2139,N_2138);
nor U2160 (N_2160,N_2135,N_2124);
nand U2161 (N_2161,N_2102,N_2117);
nand U2162 (N_2162,N_2128,N_2143);
and U2163 (N_2163,N_2129,N_2134);
nand U2164 (N_2164,N_2116,N_2149);
nor U2165 (N_2165,N_2106,N_2131);
nand U2166 (N_2166,N_2122,N_2147);
or U2167 (N_2167,N_2136,N_2101);
nand U2168 (N_2168,N_2140,N_2113);
and U2169 (N_2169,N_2119,N_2103);
and U2170 (N_2170,N_2145,N_2137);
or U2171 (N_2171,N_2126,N_2100);
or U2172 (N_2172,N_2132,N_2112);
or U2173 (N_2173,N_2144,N_2121);
nor U2174 (N_2174,N_2123,N_2115);
nand U2175 (N_2175,N_2110,N_2107);
and U2176 (N_2176,N_2126,N_2120);
nand U2177 (N_2177,N_2147,N_2130);
and U2178 (N_2178,N_2101,N_2123);
nand U2179 (N_2179,N_2120,N_2110);
and U2180 (N_2180,N_2137,N_2131);
and U2181 (N_2181,N_2120,N_2103);
nor U2182 (N_2182,N_2136,N_2114);
and U2183 (N_2183,N_2130,N_2135);
and U2184 (N_2184,N_2144,N_2135);
or U2185 (N_2185,N_2113,N_2117);
nor U2186 (N_2186,N_2102,N_2128);
nor U2187 (N_2187,N_2132,N_2127);
and U2188 (N_2188,N_2130,N_2107);
nand U2189 (N_2189,N_2134,N_2133);
or U2190 (N_2190,N_2109,N_2121);
nand U2191 (N_2191,N_2119,N_2142);
or U2192 (N_2192,N_2116,N_2123);
and U2193 (N_2193,N_2139,N_2105);
nand U2194 (N_2194,N_2127,N_2128);
or U2195 (N_2195,N_2130,N_2139);
and U2196 (N_2196,N_2111,N_2104);
xnor U2197 (N_2197,N_2105,N_2148);
or U2198 (N_2198,N_2141,N_2142);
and U2199 (N_2199,N_2144,N_2114);
nor U2200 (N_2200,N_2184,N_2153);
nor U2201 (N_2201,N_2154,N_2193);
and U2202 (N_2202,N_2158,N_2192);
nor U2203 (N_2203,N_2167,N_2197);
or U2204 (N_2204,N_2157,N_2182);
nand U2205 (N_2205,N_2170,N_2168);
nand U2206 (N_2206,N_2187,N_2162);
or U2207 (N_2207,N_2174,N_2172);
and U2208 (N_2208,N_2180,N_2173);
or U2209 (N_2209,N_2164,N_2181);
and U2210 (N_2210,N_2165,N_2183);
or U2211 (N_2211,N_2169,N_2185);
nand U2212 (N_2212,N_2155,N_2152);
nor U2213 (N_2213,N_2171,N_2156);
and U2214 (N_2214,N_2178,N_2198);
nor U2215 (N_2215,N_2175,N_2194);
or U2216 (N_2216,N_2190,N_2196);
nor U2217 (N_2217,N_2160,N_2191);
and U2218 (N_2218,N_2176,N_2151);
or U2219 (N_2219,N_2188,N_2150);
nand U2220 (N_2220,N_2159,N_2195);
or U2221 (N_2221,N_2189,N_2179);
and U2222 (N_2222,N_2166,N_2177);
or U2223 (N_2223,N_2199,N_2161);
and U2224 (N_2224,N_2163,N_2186);
nor U2225 (N_2225,N_2192,N_2170);
nor U2226 (N_2226,N_2157,N_2180);
nand U2227 (N_2227,N_2175,N_2153);
nand U2228 (N_2228,N_2194,N_2160);
or U2229 (N_2229,N_2182,N_2155);
nand U2230 (N_2230,N_2174,N_2154);
or U2231 (N_2231,N_2161,N_2166);
or U2232 (N_2232,N_2191,N_2154);
nand U2233 (N_2233,N_2152,N_2176);
nor U2234 (N_2234,N_2189,N_2178);
nor U2235 (N_2235,N_2187,N_2171);
and U2236 (N_2236,N_2167,N_2181);
or U2237 (N_2237,N_2181,N_2163);
nor U2238 (N_2238,N_2158,N_2191);
nor U2239 (N_2239,N_2189,N_2175);
and U2240 (N_2240,N_2191,N_2150);
or U2241 (N_2241,N_2188,N_2156);
nand U2242 (N_2242,N_2164,N_2198);
and U2243 (N_2243,N_2199,N_2197);
and U2244 (N_2244,N_2152,N_2153);
or U2245 (N_2245,N_2197,N_2156);
nand U2246 (N_2246,N_2153,N_2168);
nand U2247 (N_2247,N_2166,N_2151);
nand U2248 (N_2248,N_2164,N_2162);
and U2249 (N_2249,N_2185,N_2189);
or U2250 (N_2250,N_2240,N_2220);
and U2251 (N_2251,N_2211,N_2237);
nand U2252 (N_2252,N_2230,N_2216);
nor U2253 (N_2253,N_2248,N_2246);
nand U2254 (N_2254,N_2245,N_2242);
nor U2255 (N_2255,N_2236,N_2224);
nand U2256 (N_2256,N_2210,N_2204);
xnor U2257 (N_2257,N_2247,N_2207);
and U2258 (N_2258,N_2214,N_2202);
and U2259 (N_2259,N_2243,N_2209);
and U2260 (N_2260,N_2244,N_2231);
and U2261 (N_2261,N_2228,N_2200);
or U2262 (N_2262,N_2225,N_2229);
nand U2263 (N_2263,N_2232,N_2208);
and U2264 (N_2264,N_2235,N_2213);
nand U2265 (N_2265,N_2249,N_2218);
nor U2266 (N_2266,N_2239,N_2205);
and U2267 (N_2267,N_2215,N_2227);
and U2268 (N_2268,N_2219,N_2206);
or U2269 (N_2269,N_2201,N_2241);
xor U2270 (N_2270,N_2217,N_2212);
nor U2271 (N_2271,N_2238,N_2222);
or U2272 (N_2272,N_2226,N_2223);
nor U2273 (N_2273,N_2234,N_2221);
or U2274 (N_2274,N_2203,N_2233);
nand U2275 (N_2275,N_2243,N_2223);
nand U2276 (N_2276,N_2239,N_2219);
or U2277 (N_2277,N_2217,N_2246);
xnor U2278 (N_2278,N_2228,N_2203);
or U2279 (N_2279,N_2213,N_2217);
nor U2280 (N_2280,N_2234,N_2246);
and U2281 (N_2281,N_2235,N_2204);
or U2282 (N_2282,N_2203,N_2236);
nor U2283 (N_2283,N_2245,N_2205);
nand U2284 (N_2284,N_2201,N_2203);
and U2285 (N_2285,N_2239,N_2206);
nand U2286 (N_2286,N_2228,N_2227);
or U2287 (N_2287,N_2227,N_2246);
nand U2288 (N_2288,N_2240,N_2208);
nand U2289 (N_2289,N_2223,N_2211);
nor U2290 (N_2290,N_2233,N_2225);
or U2291 (N_2291,N_2239,N_2209);
nand U2292 (N_2292,N_2210,N_2202);
nor U2293 (N_2293,N_2221,N_2202);
and U2294 (N_2294,N_2209,N_2240);
nor U2295 (N_2295,N_2209,N_2201);
and U2296 (N_2296,N_2240,N_2237);
nand U2297 (N_2297,N_2204,N_2245);
nand U2298 (N_2298,N_2231,N_2243);
or U2299 (N_2299,N_2213,N_2208);
nor U2300 (N_2300,N_2258,N_2261);
nand U2301 (N_2301,N_2281,N_2289);
and U2302 (N_2302,N_2298,N_2286);
or U2303 (N_2303,N_2284,N_2293);
or U2304 (N_2304,N_2292,N_2271);
or U2305 (N_2305,N_2294,N_2297);
or U2306 (N_2306,N_2267,N_2296);
nand U2307 (N_2307,N_2268,N_2255);
nor U2308 (N_2308,N_2256,N_2250);
and U2309 (N_2309,N_2260,N_2278);
or U2310 (N_2310,N_2276,N_2299);
nand U2311 (N_2311,N_2264,N_2262);
or U2312 (N_2312,N_2266,N_2285);
or U2313 (N_2313,N_2291,N_2263);
and U2314 (N_2314,N_2269,N_2274);
nand U2315 (N_2315,N_2251,N_2280);
or U2316 (N_2316,N_2282,N_2277);
nand U2317 (N_2317,N_2273,N_2288);
and U2318 (N_2318,N_2287,N_2253);
nor U2319 (N_2319,N_2279,N_2283);
nor U2320 (N_2320,N_2290,N_2257);
or U2321 (N_2321,N_2275,N_2272);
nand U2322 (N_2322,N_2252,N_2295);
nand U2323 (N_2323,N_2259,N_2265);
or U2324 (N_2324,N_2270,N_2254);
or U2325 (N_2325,N_2274,N_2258);
nor U2326 (N_2326,N_2292,N_2259);
nor U2327 (N_2327,N_2252,N_2291);
nor U2328 (N_2328,N_2264,N_2275);
and U2329 (N_2329,N_2286,N_2274);
nor U2330 (N_2330,N_2269,N_2288);
or U2331 (N_2331,N_2299,N_2281);
and U2332 (N_2332,N_2256,N_2259);
or U2333 (N_2333,N_2288,N_2277);
nor U2334 (N_2334,N_2258,N_2254);
and U2335 (N_2335,N_2284,N_2276);
and U2336 (N_2336,N_2276,N_2265);
nand U2337 (N_2337,N_2299,N_2254);
or U2338 (N_2338,N_2268,N_2290);
or U2339 (N_2339,N_2252,N_2266);
nand U2340 (N_2340,N_2297,N_2275);
and U2341 (N_2341,N_2288,N_2261);
or U2342 (N_2342,N_2270,N_2284);
nand U2343 (N_2343,N_2288,N_2297);
nor U2344 (N_2344,N_2291,N_2280);
and U2345 (N_2345,N_2268,N_2289);
or U2346 (N_2346,N_2296,N_2270);
nand U2347 (N_2347,N_2268,N_2269);
nand U2348 (N_2348,N_2277,N_2286);
and U2349 (N_2349,N_2271,N_2296);
nand U2350 (N_2350,N_2328,N_2302);
nand U2351 (N_2351,N_2301,N_2323);
nand U2352 (N_2352,N_2349,N_2338);
nand U2353 (N_2353,N_2325,N_2315);
xor U2354 (N_2354,N_2342,N_2333);
nand U2355 (N_2355,N_2348,N_2334);
nor U2356 (N_2356,N_2322,N_2310);
and U2357 (N_2357,N_2320,N_2312);
or U2358 (N_2358,N_2300,N_2326);
or U2359 (N_2359,N_2308,N_2341);
nor U2360 (N_2360,N_2321,N_2305);
nand U2361 (N_2361,N_2309,N_2306);
nand U2362 (N_2362,N_2324,N_2329);
and U2363 (N_2363,N_2344,N_2318);
and U2364 (N_2364,N_2316,N_2313);
or U2365 (N_2365,N_2330,N_2340);
nand U2366 (N_2366,N_2343,N_2332);
nor U2367 (N_2367,N_2314,N_2303);
nand U2368 (N_2368,N_2327,N_2304);
nand U2369 (N_2369,N_2347,N_2307);
nand U2370 (N_2370,N_2336,N_2317);
and U2371 (N_2371,N_2345,N_2337);
nand U2372 (N_2372,N_2319,N_2335);
nor U2373 (N_2373,N_2346,N_2339);
and U2374 (N_2374,N_2311,N_2331);
nand U2375 (N_2375,N_2326,N_2331);
nand U2376 (N_2376,N_2313,N_2341);
nor U2377 (N_2377,N_2344,N_2315);
or U2378 (N_2378,N_2309,N_2340);
and U2379 (N_2379,N_2335,N_2314);
nor U2380 (N_2380,N_2337,N_2303);
or U2381 (N_2381,N_2302,N_2339);
or U2382 (N_2382,N_2320,N_2336);
nand U2383 (N_2383,N_2323,N_2329);
and U2384 (N_2384,N_2325,N_2317);
and U2385 (N_2385,N_2348,N_2331);
nor U2386 (N_2386,N_2314,N_2337);
and U2387 (N_2387,N_2303,N_2302);
nor U2388 (N_2388,N_2302,N_2342);
nor U2389 (N_2389,N_2318,N_2307);
and U2390 (N_2390,N_2321,N_2309);
or U2391 (N_2391,N_2310,N_2307);
and U2392 (N_2392,N_2317,N_2322);
or U2393 (N_2393,N_2348,N_2308);
and U2394 (N_2394,N_2300,N_2330);
nor U2395 (N_2395,N_2347,N_2317);
nand U2396 (N_2396,N_2316,N_2325);
or U2397 (N_2397,N_2314,N_2311);
and U2398 (N_2398,N_2309,N_2308);
and U2399 (N_2399,N_2301,N_2319);
xor U2400 (N_2400,N_2367,N_2360);
and U2401 (N_2401,N_2361,N_2358);
nand U2402 (N_2402,N_2389,N_2390);
and U2403 (N_2403,N_2366,N_2399);
and U2404 (N_2404,N_2392,N_2395);
nor U2405 (N_2405,N_2352,N_2377);
or U2406 (N_2406,N_2370,N_2378);
nand U2407 (N_2407,N_2380,N_2354);
nand U2408 (N_2408,N_2387,N_2359);
nand U2409 (N_2409,N_2397,N_2353);
and U2410 (N_2410,N_2371,N_2364);
nand U2411 (N_2411,N_2376,N_2355);
and U2412 (N_2412,N_2384,N_2396);
nor U2413 (N_2413,N_2374,N_2385);
and U2414 (N_2414,N_2350,N_2362);
or U2415 (N_2415,N_2381,N_2386);
nand U2416 (N_2416,N_2391,N_2394);
nor U2417 (N_2417,N_2365,N_2368);
nor U2418 (N_2418,N_2383,N_2356);
nor U2419 (N_2419,N_2398,N_2357);
nand U2420 (N_2420,N_2375,N_2351);
or U2421 (N_2421,N_2382,N_2373);
or U2422 (N_2422,N_2372,N_2393);
and U2423 (N_2423,N_2379,N_2388);
nor U2424 (N_2424,N_2363,N_2369);
nand U2425 (N_2425,N_2376,N_2383);
nor U2426 (N_2426,N_2359,N_2358);
or U2427 (N_2427,N_2377,N_2367);
or U2428 (N_2428,N_2384,N_2397);
or U2429 (N_2429,N_2398,N_2367);
nand U2430 (N_2430,N_2394,N_2386);
nor U2431 (N_2431,N_2358,N_2369);
nor U2432 (N_2432,N_2363,N_2367);
and U2433 (N_2433,N_2367,N_2376);
or U2434 (N_2434,N_2375,N_2376);
and U2435 (N_2435,N_2365,N_2390);
xnor U2436 (N_2436,N_2396,N_2370);
nor U2437 (N_2437,N_2370,N_2394);
nor U2438 (N_2438,N_2389,N_2364);
and U2439 (N_2439,N_2362,N_2354);
nand U2440 (N_2440,N_2353,N_2366);
or U2441 (N_2441,N_2375,N_2363);
nand U2442 (N_2442,N_2355,N_2357);
nor U2443 (N_2443,N_2399,N_2365);
nand U2444 (N_2444,N_2396,N_2392);
xnor U2445 (N_2445,N_2370,N_2387);
and U2446 (N_2446,N_2399,N_2384);
or U2447 (N_2447,N_2356,N_2351);
and U2448 (N_2448,N_2375,N_2362);
or U2449 (N_2449,N_2383,N_2386);
nor U2450 (N_2450,N_2417,N_2402);
nand U2451 (N_2451,N_2412,N_2434);
and U2452 (N_2452,N_2420,N_2437);
and U2453 (N_2453,N_2401,N_2411);
and U2454 (N_2454,N_2405,N_2445);
nand U2455 (N_2455,N_2442,N_2444);
or U2456 (N_2456,N_2426,N_2410);
and U2457 (N_2457,N_2421,N_2427);
and U2458 (N_2458,N_2416,N_2409);
and U2459 (N_2459,N_2422,N_2430);
or U2460 (N_2460,N_2406,N_2428);
nor U2461 (N_2461,N_2419,N_2413);
or U2462 (N_2462,N_2438,N_2439);
nand U2463 (N_2463,N_2418,N_2433);
nor U2464 (N_2464,N_2415,N_2414);
and U2465 (N_2465,N_2440,N_2425);
and U2466 (N_2466,N_2403,N_2407);
and U2467 (N_2467,N_2449,N_2446);
nand U2468 (N_2468,N_2443,N_2431);
nand U2469 (N_2469,N_2436,N_2423);
nor U2470 (N_2470,N_2424,N_2432);
nand U2471 (N_2471,N_2429,N_2448);
nor U2472 (N_2472,N_2408,N_2441);
nor U2473 (N_2473,N_2404,N_2435);
xor U2474 (N_2474,N_2447,N_2400);
nor U2475 (N_2475,N_2436,N_2407);
nor U2476 (N_2476,N_2407,N_2412);
or U2477 (N_2477,N_2400,N_2436);
or U2478 (N_2478,N_2403,N_2434);
and U2479 (N_2479,N_2423,N_2409);
nor U2480 (N_2480,N_2404,N_2436);
xnor U2481 (N_2481,N_2433,N_2425);
nand U2482 (N_2482,N_2406,N_2420);
and U2483 (N_2483,N_2429,N_2404);
or U2484 (N_2484,N_2400,N_2417);
nor U2485 (N_2485,N_2415,N_2446);
nand U2486 (N_2486,N_2413,N_2438);
or U2487 (N_2487,N_2443,N_2421);
and U2488 (N_2488,N_2419,N_2432);
nor U2489 (N_2489,N_2416,N_2446);
nand U2490 (N_2490,N_2432,N_2402);
or U2491 (N_2491,N_2433,N_2413);
and U2492 (N_2492,N_2411,N_2441);
and U2493 (N_2493,N_2409,N_2434);
nor U2494 (N_2494,N_2442,N_2429);
xnor U2495 (N_2495,N_2431,N_2435);
and U2496 (N_2496,N_2422,N_2435);
or U2497 (N_2497,N_2429,N_2414);
and U2498 (N_2498,N_2414,N_2441);
nor U2499 (N_2499,N_2411,N_2423);
nor U2500 (N_2500,N_2465,N_2461);
or U2501 (N_2501,N_2472,N_2475);
nor U2502 (N_2502,N_2454,N_2493);
and U2503 (N_2503,N_2457,N_2453);
nand U2504 (N_2504,N_2469,N_2485);
or U2505 (N_2505,N_2482,N_2451);
or U2506 (N_2506,N_2484,N_2478);
or U2507 (N_2507,N_2499,N_2455);
or U2508 (N_2508,N_2483,N_2464);
nand U2509 (N_2509,N_2456,N_2489);
or U2510 (N_2510,N_2452,N_2497);
or U2511 (N_2511,N_2486,N_2495);
and U2512 (N_2512,N_2463,N_2468);
nand U2513 (N_2513,N_2466,N_2458);
nor U2514 (N_2514,N_2498,N_2491);
or U2515 (N_2515,N_2467,N_2477);
or U2516 (N_2516,N_2470,N_2450);
nand U2517 (N_2517,N_2459,N_2476);
or U2518 (N_2518,N_2487,N_2473);
and U2519 (N_2519,N_2490,N_2460);
nand U2520 (N_2520,N_2480,N_2496);
nand U2521 (N_2521,N_2471,N_2494);
nand U2522 (N_2522,N_2462,N_2492);
nor U2523 (N_2523,N_2474,N_2488);
nor U2524 (N_2524,N_2479,N_2481);
nor U2525 (N_2525,N_2457,N_2464);
and U2526 (N_2526,N_2490,N_2464);
nand U2527 (N_2527,N_2495,N_2475);
nor U2528 (N_2528,N_2466,N_2453);
nor U2529 (N_2529,N_2472,N_2463);
nand U2530 (N_2530,N_2456,N_2453);
nand U2531 (N_2531,N_2475,N_2497);
nand U2532 (N_2532,N_2461,N_2451);
or U2533 (N_2533,N_2499,N_2463);
and U2534 (N_2534,N_2454,N_2460);
nor U2535 (N_2535,N_2499,N_2495);
nand U2536 (N_2536,N_2466,N_2465);
nand U2537 (N_2537,N_2498,N_2470);
or U2538 (N_2538,N_2468,N_2459);
nand U2539 (N_2539,N_2488,N_2491);
and U2540 (N_2540,N_2453,N_2492);
nor U2541 (N_2541,N_2463,N_2486);
and U2542 (N_2542,N_2456,N_2460);
and U2543 (N_2543,N_2488,N_2466);
nand U2544 (N_2544,N_2478,N_2450);
nor U2545 (N_2545,N_2485,N_2478);
nor U2546 (N_2546,N_2463,N_2476);
nor U2547 (N_2547,N_2452,N_2473);
nand U2548 (N_2548,N_2462,N_2468);
nor U2549 (N_2549,N_2460,N_2451);
or U2550 (N_2550,N_2544,N_2509);
or U2551 (N_2551,N_2535,N_2536);
or U2552 (N_2552,N_2541,N_2543);
nor U2553 (N_2553,N_2500,N_2545);
and U2554 (N_2554,N_2531,N_2527);
or U2555 (N_2555,N_2505,N_2518);
nor U2556 (N_2556,N_2539,N_2503);
nor U2557 (N_2557,N_2546,N_2526);
nand U2558 (N_2558,N_2525,N_2537);
nor U2559 (N_2559,N_2511,N_2532);
and U2560 (N_2560,N_2549,N_2510);
or U2561 (N_2561,N_2521,N_2506);
and U2562 (N_2562,N_2501,N_2522);
or U2563 (N_2563,N_2530,N_2529);
and U2564 (N_2564,N_2547,N_2542);
or U2565 (N_2565,N_2517,N_2524);
nand U2566 (N_2566,N_2538,N_2502);
nand U2567 (N_2567,N_2533,N_2512);
nand U2568 (N_2568,N_2520,N_2513);
nor U2569 (N_2569,N_2515,N_2548);
nor U2570 (N_2570,N_2504,N_2523);
nand U2571 (N_2571,N_2528,N_2519);
nor U2572 (N_2572,N_2534,N_2540);
or U2573 (N_2573,N_2507,N_2516);
and U2574 (N_2574,N_2514,N_2508);
nand U2575 (N_2575,N_2531,N_2543);
nor U2576 (N_2576,N_2514,N_2505);
nor U2577 (N_2577,N_2504,N_2529);
or U2578 (N_2578,N_2523,N_2532);
and U2579 (N_2579,N_2514,N_2518);
nand U2580 (N_2580,N_2540,N_2522);
or U2581 (N_2581,N_2548,N_2535);
nand U2582 (N_2582,N_2511,N_2533);
nor U2583 (N_2583,N_2517,N_2508);
and U2584 (N_2584,N_2536,N_2506);
or U2585 (N_2585,N_2527,N_2546);
or U2586 (N_2586,N_2522,N_2538);
nor U2587 (N_2587,N_2510,N_2536);
nand U2588 (N_2588,N_2528,N_2507);
and U2589 (N_2589,N_2547,N_2521);
nor U2590 (N_2590,N_2523,N_2516);
nor U2591 (N_2591,N_2521,N_2516);
nor U2592 (N_2592,N_2503,N_2521);
nor U2593 (N_2593,N_2514,N_2516);
nor U2594 (N_2594,N_2546,N_2537);
or U2595 (N_2595,N_2512,N_2540);
nor U2596 (N_2596,N_2508,N_2504);
nor U2597 (N_2597,N_2508,N_2532);
nand U2598 (N_2598,N_2500,N_2528);
or U2599 (N_2599,N_2535,N_2534);
or U2600 (N_2600,N_2587,N_2569);
nor U2601 (N_2601,N_2591,N_2595);
nor U2602 (N_2602,N_2565,N_2571);
and U2603 (N_2603,N_2588,N_2575);
nor U2604 (N_2604,N_2578,N_2554);
nand U2605 (N_2605,N_2564,N_2559);
nand U2606 (N_2606,N_2590,N_2584);
or U2607 (N_2607,N_2580,N_2560);
nand U2608 (N_2608,N_2550,N_2557);
nand U2609 (N_2609,N_2573,N_2563);
and U2610 (N_2610,N_2567,N_2576);
nand U2611 (N_2611,N_2551,N_2562);
nand U2612 (N_2612,N_2598,N_2586);
nor U2613 (N_2613,N_2558,N_2556);
and U2614 (N_2614,N_2577,N_2593);
nor U2615 (N_2615,N_2552,N_2599);
nor U2616 (N_2616,N_2561,N_2570);
nor U2617 (N_2617,N_2555,N_2566);
or U2618 (N_2618,N_2596,N_2594);
nand U2619 (N_2619,N_2583,N_2597);
nand U2620 (N_2620,N_2553,N_2568);
nor U2621 (N_2621,N_2592,N_2572);
or U2622 (N_2622,N_2589,N_2581);
nand U2623 (N_2623,N_2585,N_2582);
nand U2624 (N_2624,N_2579,N_2574);
nand U2625 (N_2625,N_2591,N_2580);
nor U2626 (N_2626,N_2596,N_2560);
and U2627 (N_2627,N_2568,N_2570);
nor U2628 (N_2628,N_2578,N_2562);
and U2629 (N_2629,N_2593,N_2574);
nor U2630 (N_2630,N_2553,N_2563);
or U2631 (N_2631,N_2563,N_2550);
nand U2632 (N_2632,N_2594,N_2591);
and U2633 (N_2633,N_2570,N_2589);
nor U2634 (N_2634,N_2561,N_2555);
and U2635 (N_2635,N_2551,N_2555);
and U2636 (N_2636,N_2561,N_2577);
nor U2637 (N_2637,N_2563,N_2551);
and U2638 (N_2638,N_2599,N_2585);
and U2639 (N_2639,N_2595,N_2576);
nand U2640 (N_2640,N_2579,N_2580);
nor U2641 (N_2641,N_2584,N_2576);
nand U2642 (N_2642,N_2564,N_2576);
and U2643 (N_2643,N_2577,N_2583);
and U2644 (N_2644,N_2594,N_2552);
or U2645 (N_2645,N_2551,N_2569);
nor U2646 (N_2646,N_2583,N_2563);
or U2647 (N_2647,N_2560,N_2594);
nor U2648 (N_2648,N_2575,N_2569);
nand U2649 (N_2649,N_2585,N_2552);
nand U2650 (N_2650,N_2648,N_2639);
nand U2651 (N_2651,N_2620,N_2629);
or U2652 (N_2652,N_2612,N_2605);
or U2653 (N_2653,N_2614,N_2628);
and U2654 (N_2654,N_2634,N_2638);
and U2655 (N_2655,N_2631,N_2608);
and U2656 (N_2656,N_2640,N_2645);
or U2657 (N_2657,N_2636,N_2601);
or U2658 (N_2658,N_2625,N_2610);
and U2659 (N_2659,N_2630,N_2621);
nand U2660 (N_2660,N_2626,N_2604);
nor U2661 (N_2661,N_2603,N_2618);
nor U2662 (N_2662,N_2643,N_2606);
and U2663 (N_2663,N_2649,N_2617);
nand U2664 (N_2664,N_2615,N_2635);
and U2665 (N_2665,N_2609,N_2637);
nand U2666 (N_2666,N_2642,N_2647);
or U2667 (N_2667,N_2627,N_2644);
or U2668 (N_2668,N_2641,N_2611);
or U2669 (N_2669,N_2623,N_2607);
nand U2670 (N_2670,N_2633,N_2632);
and U2671 (N_2671,N_2619,N_2616);
nand U2672 (N_2672,N_2613,N_2646);
or U2673 (N_2673,N_2600,N_2622);
or U2674 (N_2674,N_2624,N_2602);
or U2675 (N_2675,N_2635,N_2608);
or U2676 (N_2676,N_2633,N_2631);
or U2677 (N_2677,N_2648,N_2647);
or U2678 (N_2678,N_2615,N_2607);
and U2679 (N_2679,N_2600,N_2611);
nor U2680 (N_2680,N_2640,N_2626);
nand U2681 (N_2681,N_2623,N_2647);
or U2682 (N_2682,N_2603,N_2643);
nand U2683 (N_2683,N_2614,N_2637);
and U2684 (N_2684,N_2629,N_2618);
nor U2685 (N_2685,N_2626,N_2624);
nand U2686 (N_2686,N_2628,N_2625);
xnor U2687 (N_2687,N_2634,N_2635);
nand U2688 (N_2688,N_2638,N_2614);
nand U2689 (N_2689,N_2642,N_2601);
nand U2690 (N_2690,N_2624,N_2625);
xnor U2691 (N_2691,N_2639,N_2609);
nor U2692 (N_2692,N_2601,N_2621);
nand U2693 (N_2693,N_2624,N_2605);
nor U2694 (N_2694,N_2628,N_2621);
nand U2695 (N_2695,N_2602,N_2648);
nor U2696 (N_2696,N_2603,N_2606);
nor U2697 (N_2697,N_2637,N_2649);
or U2698 (N_2698,N_2643,N_2644);
nor U2699 (N_2699,N_2624,N_2620);
nor U2700 (N_2700,N_2674,N_2659);
nor U2701 (N_2701,N_2673,N_2665);
or U2702 (N_2702,N_2680,N_2672);
nand U2703 (N_2703,N_2668,N_2662);
or U2704 (N_2704,N_2692,N_2697);
or U2705 (N_2705,N_2690,N_2678);
and U2706 (N_2706,N_2663,N_2686);
and U2707 (N_2707,N_2683,N_2666);
xnor U2708 (N_2708,N_2691,N_2682);
or U2709 (N_2709,N_2676,N_2655);
or U2710 (N_2710,N_2685,N_2695);
nand U2711 (N_2711,N_2669,N_2699);
and U2712 (N_2712,N_2651,N_2670);
xor U2713 (N_2713,N_2652,N_2660);
nor U2714 (N_2714,N_2654,N_2664);
xor U2715 (N_2715,N_2658,N_2677);
nor U2716 (N_2716,N_2671,N_2681);
nand U2717 (N_2717,N_2650,N_2689);
and U2718 (N_2718,N_2693,N_2687);
and U2719 (N_2719,N_2698,N_2656);
nor U2720 (N_2720,N_2667,N_2657);
nand U2721 (N_2721,N_2675,N_2661);
or U2722 (N_2722,N_2653,N_2694);
or U2723 (N_2723,N_2684,N_2679);
nand U2724 (N_2724,N_2688,N_2696);
nand U2725 (N_2725,N_2673,N_2669);
nand U2726 (N_2726,N_2676,N_2656);
nor U2727 (N_2727,N_2665,N_2672);
nand U2728 (N_2728,N_2697,N_2662);
or U2729 (N_2729,N_2692,N_2661);
nor U2730 (N_2730,N_2695,N_2690);
and U2731 (N_2731,N_2688,N_2698);
and U2732 (N_2732,N_2680,N_2670);
or U2733 (N_2733,N_2699,N_2692);
nand U2734 (N_2734,N_2665,N_2656);
and U2735 (N_2735,N_2673,N_2686);
nor U2736 (N_2736,N_2669,N_2662);
and U2737 (N_2737,N_2661,N_2671);
nor U2738 (N_2738,N_2653,N_2690);
nand U2739 (N_2739,N_2678,N_2658);
or U2740 (N_2740,N_2676,N_2664);
nand U2741 (N_2741,N_2663,N_2665);
nor U2742 (N_2742,N_2699,N_2694);
and U2743 (N_2743,N_2671,N_2682);
nand U2744 (N_2744,N_2694,N_2654);
or U2745 (N_2745,N_2687,N_2663);
nor U2746 (N_2746,N_2685,N_2697);
nor U2747 (N_2747,N_2696,N_2687);
nor U2748 (N_2748,N_2680,N_2690);
or U2749 (N_2749,N_2693,N_2653);
nand U2750 (N_2750,N_2724,N_2722);
or U2751 (N_2751,N_2742,N_2705);
and U2752 (N_2752,N_2701,N_2710);
nor U2753 (N_2753,N_2737,N_2716);
nand U2754 (N_2754,N_2736,N_2709);
or U2755 (N_2755,N_2704,N_2727);
nor U2756 (N_2756,N_2717,N_2733);
and U2757 (N_2757,N_2711,N_2735);
nor U2758 (N_2758,N_2749,N_2743);
and U2759 (N_2759,N_2718,N_2726);
nand U2760 (N_2760,N_2703,N_2738);
nor U2761 (N_2761,N_2723,N_2708);
and U2762 (N_2762,N_2720,N_2702);
and U2763 (N_2763,N_2748,N_2721);
nor U2764 (N_2764,N_2715,N_2732);
or U2765 (N_2765,N_2706,N_2714);
nand U2766 (N_2766,N_2746,N_2725);
or U2767 (N_2767,N_2739,N_2707);
or U2768 (N_2768,N_2712,N_2730);
xnor U2769 (N_2769,N_2744,N_2734);
nor U2770 (N_2770,N_2729,N_2740);
or U2771 (N_2771,N_2731,N_2747);
or U2772 (N_2772,N_2700,N_2719);
nor U2773 (N_2773,N_2713,N_2728);
and U2774 (N_2774,N_2745,N_2741);
nor U2775 (N_2775,N_2718,N_2741);
nand U2776 (N_2776,N_2743,N_2741);
nor U2777 (N_2777,N_2729,N_2704);
or U2778 (N_2778,N_2727,N_2713);
nand U2779 (N_2779,N_2731,N_2736);
and U2780 (N_2780,N_2728,N_2740);
and U2781 (N_2781,N_2702,N_2709);
nor U2782 (N_2782,N_2710,N_2715);
and U2783 (N_2783,N_2706,N_2718);
and U2784 (N_2784,N_2728,N_2727);
or U2785 (N_2785,N_2732,N_2700);
nand U2786 (N_2786,N_2745,N_2722);
and U2787 (N_2787,N_2707,N_2725);
nor U2788 (N_2788,N_2734,N_2704);
nor U2789 (N_2789,N_2715,N_2748);
or U2790 (N_2790,N_2706,N_2740);
or U2791 (N_2791,N_2711,N_2746);
or U2792 (N_2792,N_2739,N_2712);
nand U2793 (N_2793,N_2710,N_2727);
nor U2794 (N_2794,N_2735,N_2736);
nand U2795 (N_2795,N_2727,N_2730);
or U2796 (N_2796,N_2713,N_2749);
nor U2797 (N_2797,N_2722,N_2731);
or U2798 (N_2798,N_2722,N_2714);
nor U2799 (N_2799,N_2713,N_2704);
nand U2800 (N_2800,N_2799,N_2798);
nor U2801 (N_2801,N_2762,N_2786);
nor U2802 (N_2802,N_2789,N_2780);
nor U2803 (N_2803,N_2795,N_2778);
and U2804 (N_2804,N_2754,N_2773);
and U2805 (N_2805,N_2761,N_2794);
xnor U2806 (N_2806,N_2775,N_2765);
nand U2807 (N_2807,N_2756,N_2758);
nand U2808 (N_2808,N_2782,N_2776);
and U2809 (N_2809,N_2768,N_2777);
nor U2810 (N_2810,N_2769,N_2788);
or U2811 (N_2811,N_2781,N_2760);
or U2812 (N_2812,N_2751,N_2791);
nand U2813 (N_2813,N_2787,N_2759);
or U2814 (N_2814,N_2750,N_2779);
nor U2815 (N_2815,N_2770,N_2767);
or U2816 (N_2816,N_2753,N_2796);
or U2817 (N_2817,N_2797,N_2784);
nand U2818 (N_2818,N_2752,N_2772);
nor U2819 (N_2819,N_2793,N_2790);
nand U2820 (N_2820,N_2755,N_2763);
and U2821 (N_2821,N_2757,N_2792);
xor U2822 (N_2822,N_2783,N_2774);
nor U2823 (N_2823,N_2764,N_2766);
nor U2824 (N_2824,N_2771,N_2785);
and U2825 (N_2825,N_2762,N_2797);
and U2826 (N_2826,N_2756,N_2786);
and U2827 (N_2827,N_2764,N_2778);
and U2828 (N_2828,N_2799,N_2752);
or U2829 (N_2829,N_2755,N_2781);
nor U2830 (N_2830,N_2790,N_2776);
and U2831 (N_2831,N_2792,N_2758);
or U2832 (N_2832,N_2772,N_2764);
nor U2833 (N_2833,N_2784,N_2758);
or U2834 (N_2834,N_2777,N_2775);
nor U2835 (N_2835,N_2791,N_2769);
and U2836 (N_2836,N_2783,N_2779);
nor U2837 (N_2837,N_2783,N_2772);
or U2838 (N_2838,N_2768,N_2755);
nor U2839 (N_2839,N_2772,N_2765);
nor U2840 (N_2840,N_2771,N_2766);
and U2841 (N_2841,N_2797,N_2789);
nor U2842 (N_2842,N_2774,N_2777);
nand U2843 (N_2843,N_2786,N_2765);
nor U2844 (N_2844,N_2781,N_2775);
nor U2845 (N_2845,N_2774,N_2763);
nor U2846 (N_2846,N_2774,N_2797);
nand U2847 (N_2847,N_2756,N_2778);
or U2848 (N_2848,N_2761,N_2799);
nand U2849 (N_2849,N_2756,N_2784);
or U2850 (N_2850,N_2844,N_2808);
and U2851 (N_2851,N_2835,N_2803);
and U2852 (N_2852,N_2827,N_2846);
or U2853 (N_2853,N_2848,N_2801);
nor U2854 (N_2854,N_2838,N_2837);
nor U2855 (N_2855,N_2819,N_2834);
and U2856 (N_2856,N_2829,N_2816);
or U2857 (N_2857,N_2840,N_2800);
nor U2858 (N_2858,N_2815,N_2812);
and U2859 (N_2859,N_2820,N_2807);
and U2860 (N_2860,N_2824,N_2806);
nand U2861 (N_2861,N_2813,N_2818);
nor U2862 (N_2862,N_2810,N_2843);
and U2863 (N_2863,N_2802,N_2831);
nor U2864 (N_2864,N_2845,N_2833);
nor U2865 (N_2865,N_2811,N_2825);
nor U2866 (N_2866,N_2822,N_2842);
nand U2867 (N_2867,N_2823,N_2832);
and U2868 (N_2868,N_2839,N_2821);
or U2869 (N_2869,N_2814,N_2804);
and U2870 (N_2870,N_2817,N_2841);
nor U2871 (N_2871,N_2836,N_2830);
or U2872 (N_2872,N_2805,N_2847);
nor U2873 (N_2873,N_2826,N_2809);
nand U2874 (N_2874,N_2828,N_2849);
nand U2875 (N_2875,N_2844,N_2806);
nor U2876 (N_2876,N_2815,N_2846);
and U2877 (N_2877,N_2816,N_2825);
and U2878 (N_2878,N_2829,N_2815);
nor U2879 (N_2879,N_2815,N_2811);
or U2880 (N_2880,N_2800,N_2837);
or U2881 (N_2881,N_2805,N_2822);
and U2882 (N_2882,N_2823,N_2849);
or U2883 (N_2883,N_2815,N_2837);
and U2884 (N_2884,N_2820,N_2837);
nand U2885 (N_2885,N_2804,N_2843);
and U2886 (N_2886,N_2829,N_2822);
nor U2887 (N_2887,N_2818,N_2809);
and U2888 (N_2888,N_2838,N_2820);
and U2889 (N_2889,N_2840,N_2833);
nor U2890 (N_2890,N_2843,N_2823);
or U2891 (N_2891,N_2847,N_2829);
nand U2892 (N_2892,N_2803,N_2805);
xnor U2893 (N_2893,N_2817,N_2824);
nand U2894 (N_2894,N_2829,N_2800);
or U2895 (N_2895,N_2839,N_2813);
or U2896 (N_2896,N_2841,N_2815);
nor U2897 (N_2897,N_2844,N_2828);
and U2898 (N_2898,N_2828,N_2835);
nand U2899 (N_2899,N_2828,N_2804);
nor U2900 (N_2900,N_2884,N_2851);
or U2901 (N_2901,N_2878,N_2885);
nor U2902 (N_2902,N_2858,N_2877);
nand U2903 (N_2903,N_2859,N_2891);
nand U2904 (N_2904,N_2850,N_2867);
and U2905 (N_2905,N_2861,N_2887);
nand U2906 (N_2906,N_2886,N_2873);
nor U2907 (N_2907,N_2868,N_2894);
nor U2908 (N_2908,N_2897,N_2865);
and U2909 (N_2909,N_2899,N_2875);
nor U2910 (N_2910,N_2896,N_2888);
nor U2911 (N_2911,N_2876,N_2898);
nor U2912 (N_2912,N_2857,N_2871);
or U2913 (N_2913,N_2874,N_2863);
nand U2914 (N_2914,N_2890,N_2853);
or U2915 (N_2915,N_2889,N_2895);
and U2916 (N_2916,N_2870,N_2862);
nand U2917 (N_2917,N_2883,N_2880);
nor U2918 (N_2918,N_2872,N_2893);
or U2919 (N_2919,N_2881,N_2860);
and U2920 (N_2920,N_2879,N_2892);
and U2921 (N_2921,N_2852,N_2854);
nor U2922 (N_2922,N_2864,N_2856);
xor U2923 (N_2923,N_2855,N_2882);
nor U2924 (N_2924,N_2866,N_2869);
nor U2925 (N_2925,N_2868,N_2867);
nand U2926 (N_2926,N_2875,N_2871);
nor U2927 (N_2927,N_2892,N_2871);
nor U2928 (N_2928,N_2871,N_2879);
or U2929 (N_2929,N_2888,N_2876);
and U2930 (N_2930,N_2885,N_2886);
and U2931 (N_2931,N_2867,N_2877);
nor U2932 (N_2932,N_2862,N_2867);
or U2933 (N_2933,N_2869,N_2892);
or U2934 (N_2934,N_2871,N_2895);
and U2935 (N_2935,N_2876,N_2894);
nor U2936 (N_2936,N_2857,N_2860);
nand U2937 (N_2937,N_2884,N_2856);
or U2938 (N_2938,N_2898,N_2886);
xnor U2939 (N_2939,N_2854,N_2871);
nand U2940 (N_2940,N_2857,N_2854);
nand U2941 (N_2941,N_2865,N_2881);
nand U2942 (N_2942,N_2899,N_2860);
or U2943 (N_2943,N_2866,N_2868);
nor U2944 (N_2944,N_2886,N_2893);
or U2945 (N_2945,N_2855,N_2894);
or U2946 (N_2946,N_2891,N_2852);
and U2947 (N_2947,N_2868,N_2856);
nand U2948 (N_2948,N_2874,N_2881);
nor U2949 (N_2949,N_2878,N_2884);
and U2950 (N_2950,N_2929,N_2923);
or U2951 (N_2951,N_2927,N_2915);
nand U2952 (N_2952,N_2932,N_2931);
nor U2953 (N_2953,N_2913,N_2934);
nand U2954 (N_2954,N_2947,N_2902);
nor U2955 (N_2955,N_2921,N_2906);
and U2956 (N_2956,N_2948,N_2909);
nor U2957 (N_2957,N_2928,N_2903);
or U2958 (N_2958,N_2924,N_2937);
nor U2959 (N_2959,N_2940,N_2916);
nand U2960 (N_2960,N_2925,N_2933);
or U2961 (N_2961,N_2941,N_2900);
nand U2962 (N_2962,N_2938,N_2935);
xnor U2963 (N_2963,N_2911,N_2901);
nand U2964 (N_2964,N_2926,N_2908);
nand U2965 (N_2965,N_2946,N_2942);
nor U2966 (N_2966,N_2919,N_2914);
or U2967 (N_2967,N_2944,N_2907);
nor U2968 (N_2968,N_2930,N_2910);
or U2969 (N_2969,N_2939,N_2920);
nand U2970 (N_2970,N_2943,N_2949);
nor U2971 (N_2971,N_2912,N_2917);
nand U2972 (N_2972,N_2945,N_2922);
or U2973 (N_2973,N_2936,N_2905);
or U2974 (N_2974,N_2904,N_2918);
nor U2975 (N_2975,N_2946,N_2931);
xor U2976 (N_2976,N_2928,N_2938);
and U2977 (N_2977,N_2924,N_2900);
and U2978 (N_2978,N_2926,N_2932);
and U2979 (N_2979,N_2923,N_2911);
and U2980 (N_2980,N_2928,N_2919);
nand U2981 (N_2981,N_2902,N_2929);
nor U2982 (N_2982,N_2901,N_2943);
or U2983 (N_2983,N_2930,N_2936);
nand U2984 (N_2984,N_2928,N_2941);
or U2985 (N_2985,N_2940,N_2943);
and U2986 (N_2986,N_2934,N_2939);
or U2987 (N_2987,N_2912,N_2913);
nand U2988 (N_2988,N_2934,N_2902);
nand U2989 (N_2989,N_2900,N_2938);
nand U2990 (N_2990,N_2922,N_2926);
nand U2991 (N_2991,N_2940,N_2935);
nand U2992 (N_2992,N_2949,N_2910);
or U2993 (N_2993,N_2919,N_2947);
or U2994 (N_2994,N_2915,N_2914);
or U2995 (N_2995,N_2922,N_2930);
or U2996 (N_2996,N_2943,N_2927);
or U2997 (N_2997,N_2916,N_2923);
nand U2998 (N_2998,N_2908,N_2914);
nand U2999 (N_2999,N_2910,N_2936);
nand UO_0 (O_0,N_2980,N_2979);
nand UO_1 (O_1,N_2995,N_2951);
nand UO_2 (O_2,N_2999,N_2993);
and UO_3 (O_3,N_2956,N_2977);
and UO_4 (O_4,N_2970,N_2971);
nor UO_5 (O_5,N_2955,N_2958);
nand UO_6 (O_6,N_2962,N_2989);
nand UO_7 (O_7,N_2965,N_2997);
or UO_8 (O_8,N_2981,N_2954);
or UO_9 (O_9,N_2998,N_2990);
nand UO_10 (O_10,N_2992,N_2957);
and UO_11 (O_11,N_2969,N_2987);
nor UO_12 (O_12,N_2983,N_2985);
or UO_13 (O_13,N_2972,N_2982);
nor UO_14 (O_14,N_2963,N_2953);
nand UO_15 (O_15,N_2996,N_2984);
and UO_16 (O_16,N_2994,N_2960);
or UO_17 (O_17,N_2986,N_2968);
and UO_18 (O_18,N_2974,N_2959);
nor UO_19 (O_19,N_2975,N_2973);
and UO_20 (O_20,N_2991,N_2967);
and UO_21 (O_21,N_2950,N_2952);
nor UO_22 (O_22,N_2964,N_2988);
and UO_23 (O_23,N_2961,N_2976);
and UO_24 (O_24,N_2978,N_2966);
or UO_25 (O_25,N_2996,N_2954);
nand UO_26 (O_26,N_2998,N_2966);
and UO_27 (O_27,N_2987,N_2988);
nor UO_28 (O_28,N_2968,N_2992);
and UO_29 (O_29,N_2981,N_2952);
nor UO_30 (O_30,N_2957,N_2993);
and UO_31 (O_31,N_2966,N_2975);
or UO_32 (O_32,N_2956,N_2983);
nand UO_33 (O_33,N_2973,N_2980);
nand UO_34 (O_34,N_2951,N_2954);
nand UO_35 (O_35,N_2984,N_2989);
and UO_36 (O_36,N_2963,N_2979);
or UO_37 (O_37,N_2952,N_2996);
nand UO_38 (O_38,N_2973,N_2957);
or UO_39 (O_39,N_2991,N_2956);
and UO_40 (O_40,N_2983,N_2959);
and UO_41 (O_41,N_2979,N_2960);
and UO_42 (O_42,N_2976,N_2971);
nor UO_43 (O_43,N_2970,N_2960);
nand UO_44 (O_44,N_2971,N_2989);
or UO_45 (O_45,N_2967,N_2986);
or UO_46 (O_46,N_2976,N_2962);
nor UO_47 (O_47,N_2967,N_2995);
nor UO_48 (O_48,N_2996,N_2997);
and UO_49 (O_49,N_2991,N_2989);
or UO_50 (O_50,N_2955,N_2976);
or UO_51 (O_51,N_2993,N_2981);
nor UO_52 (O_52,N_2957,N_2979);
nor UO_53 (O_53,N_2978,N_2999);
nor UO_54 (O_54,N_2951,N_2989);
or UO_55 (O_55,N_2980,N_2974);
or UO_56 (O_56,N_2958,N_2964);
nand UO_57 (O_57,N_2987,N_2982);
nor UO_58 (O_58,N_2989,N_2979);
nor UO_59 (O_59,N_2975,N_2954);
or UO_60 (O_60,N_2985,N_2999);
or UO_61 (O_61,N_2964,N_2986);
xnor UO_62 (O_62,N_2972,N_2988);
and UO_63 (O_63,N_2980,N_2986);
or UO_64 (O_64,N_2962,N_2978);
nand UO_65 (O_65,N_2998,N_2986);
or UO_66 (O_66,N_2977,N_2973);
nand UO_67 (O_67,N_2955,N_2970);
and UO_68 (O_68,N_2968,N_2957);
nand UO_69 (O_69,N_2967,N_2966);
nand UO_70 (O_70,N_2985,N_2980);
nand UO_71 (O_71,N_2966,N_2982);
and UO_72 (O_72,N_2980,N_2991);
xor UO_73 (O_73,N_2966,N_2996);
and UO_74 (O_74,N_2958,N_2995);
nor UO_75 (O_75,N_2984,N_2967);
nand UO_76 (O_76,N_2958,N_2963);
nor UO_77 (O_77,N_2950,N_2958);
and UO_78 (O_78,N_2986,N_2992);
and UO_79 (O_79,N_2964,N_2974);
or UO_80 (O_80,N_2992,N_2987);
or UO_81 (O_81,N_2965,N_2951);
and UO_82 (O_82,N_2999,N_2961);
nor UO_83 (O_83,N_2995,N_2984);
and UO_84 (O_84,N_2996,N_2951);
or UO_85 (O_85,N_2950,N_2994);
nand UO_86 (O_86,N_2977,N_2953);
and UO_87 (O_87,N_2979,N_2994);
nor UO_88 (O_88,N_2982,N_2954);
nor UO_89 (O_89,N_2966,N_2976);
or UO_90 (O_90,N_2990,N_2951);
nor UO_91 (O_91,N_2973,N_2960);
nor UO_92 (O_92,N_2974,N_2985);
nand UO_93 (O_93,N_2992,N_2999);
xnor UO_94 (O_94,N_2954,N_2976);
nand UO_95 (O_95,N_2971,N_2993);
and UO_96 (O_96,N_2967,N_2961);
nor UO_97 (O_97,N_2978,N_2984);
and UO_98 (O_98,N_2956,N_2994);
nand UO_99 (O_99,N_2975,N_2968);
nor UO_100 (O_100,N_2955,N_2968);
nor UO_101 (O_101,N_2975,N_2976);
or UO_102 (O_102,N_2963,N_2961);
and UO_103 (O_103,N_2953,N_2990);
and UO_104 (O_104,N_2950,N_2995);
nand UO_105 (O_105,N_2976,N_2979);
or UO_106 (O_106,N_2951,N_2956);
and UO_107 (O_107,N_2961,N_2986);
and UO_108 (O_108,N_2952,N_2999);
nor UO_109 (O_109,N_2989,N_2963);
nor UO_110 (O_110,N_2960,N_2986);
nand UO_111 (O_111,N_2990,N_2973);
or UO_112 (O_112,N_2982,N_2995);
or UO_113 (O_113,N_2997,N_2999);
nand UO_114 (O_114,N_2968,N_2969);
or UO_115 (O_115,N_2965,N_2988);
nor UO_116 (O_116,N_2979,N_2967);
and UO_117 (O_117,N_2972,N_2968);
nor UO_118 (O_118,N_2977,N_2992);
nand UO_119 (O_119,N_2984,N_2957);
nand UO_120 (O_120,N_2985,N_2965);
nand UO_121 (O_121,N_2964,N_2989);
nand UO_122 (O_122,N_2991,N_2957);
nand UO_123 (O_123,N_2961,N_2975);
or UO_124 (O_124,N_2978,N_2973);
nor UO_125 (O_125,N_2971,N_2956);
and UO_126 (O_126,N_2973,N_2984);
nand UO_127 (O_127,N_2971,N_2978);
nand UO_128 (O_128,N_2956,N_2984);
nor UO_129 (O_129,N_2998,N_2959);
or UO_130 (O_130,N_2989,N_2972);
nor UO_131 (O_131,N_2964,N_2994);
nor UO_132 (O_132,N_2997,N_2956);
nand UO_133 (O_133,N_2977,N_2961);
nor UO_134 (O_134,N_2977,N_2964);
and UO_135 (O_135,N_2971,N_2968);
or UO_136 (O_136,N_2958,N_2975);
and UO_137 (O_137,N_2954,N_2978);
nor UO_138 (O_138,N_2958,N_2996);
nand UO_139 (O_139,N_2986,N_2974);
and UO_140 (O_140,N_2972,N_2951);
or UO_141 (O_141,N_2973,N_2997);
nor UO_142 (O_142,N_2964,N_2961);
or UO_143 (O_143,N_2951,N_2953);
nand UO_144 (O_144,N_2978,N_2995);
or UO_145 (O_145,N_2961,N_2995);
or UO_146 (O_146,N_2957,N_2969);
and UO_147 (O_147,N_2967,N_2950);
nand UO_148 (O_148,N_2983,N_2984);
or UO_149 (O_149,N_2979,N_2998);
nor UO_150 (O_150,N_2975,N_2997);
nand UO_151 (O_151,N_2974,N_2996);
nor UO_152 (O_152,N_2966,N_2962);
or UO_153 (O_153,N_2960,N_2991);
and UO_154 (O_154,N_2970,N_2969);
or UO_155 (O_155,N_2961,N_2971);
or UO_156 (O_156,N_2956,N_2972);
nand UO_157 (O_157,N_2993,N_2973);
or UO_158 (O_158,N_2972,N_2979);
nand UO_159 (O_159,N_2974,N_2988);
nor UO_160 (O_160,N_2994,N_2965);
nor UO_161 (O_161,N_2964,N_2998);
nor UO_162 (O_162,N_2960,N_2995);
nor UO_163 (O_163,N_2952,N_2980);
or UO_164 (O_164,N_2954,N_2966);
nand UO_165 (O_165,N_2964,N_2981);
or UO_166 (O_166,N_2994,N_2971);
nand UO_167 (O_167,N_2965,N_2982);
nand UO_168 (O_168,N_2990,N_2982);
and UO_169 (O_169,N_2988,N_2992);
or UO_170 (O_170,N_2989,N_2974);
nor UO_171 (O_171,N_2958,N_2983);
nor UO_172 (O_172,N_2959,N_2960);
or UO_173 (O_173,N_2998,N_2989);
or UO_174 (O_174,N_2951,N_2973);
nand UO_175 (O_175,N_2959,N_2951);
and UO_176 (O_176,N_2970,N_2988);
and UO_177 (O_177,N_2997,N_2961);
nor UO_178 (O_178,N_2960,N_2950);
and UO_179 (O_179,N_2993,N_2975);
nor UO_180 (O_180,N_2954,N_2987);
nor UO_181 (O_181,N_2957,N_2950);
and UO_182 (O_182,N_2993,N_2986);
or UO_183 (O_183,N_2958,N_2986);
nor UO_184 (O_184,N_2951,N_2999);
and UO_185 (O_185,N_2952,N_2958);
and UO_186 (O_186,N_2995,N_2998);
and UO_187 (O_187,N_2998,N_2970);
and UO_188 (O_188,N_2965,N_2959);
nand UO_189 (O_189,N_2959,N_2989);
nand UO_190 (O_190,N_2991,N_2953);
nor UO_191 (O_191,N_2965,N_2981);
nor UO_192 (O_192,N_2980,N_2990);
or UO_193 (O_193,N_2958,N_2968);
xor UO_194 (O_194,N_2951,N_2981);
nand UO_195 (O_195,N_2964,N_2982);
or UO_196 (O_196,N_2950,N_2955);
and UO_197 (O_197,N_2984,N_2964);
or UO_198 (O_198,N_2957,N_2999);
nor UO_199 (O_199,N_2987,N_2964);
nor UO_200 (O_200,N_2978,N_2957);
nor UO_201 (O_201,N_2986,N_2977);
xnor UO_202 (O_202,N_2972,N_2958);
nand UO_203 (O_203,N_2986,N_2950);
nor UO_204 (O_204,N_2960,N_2974);
and UO_205 (O_205,N_2955,N_2978);
nor UO_206 (O_206,N_2976,N_2951);
xnor UO_207 (O_207,N_2952,N_2973);
nor UO_208 (O_208,N_2970,N_2993);
and UO_209 (O_209,N_2997,N_2969);
nand UO_210 (O_210,N_2998,N_2991);
or UO_211 (O_211,N_2977,N_2978);
nor UO_212 (O_212,N_2976,N_2988);
nand UO_213 (O_213,N_2962,N_2973);
and UO_214 (O_214,N_2966,N_2999);
nor UO_215 (O_215,N_2951,N_2991);
or UO_216 (O_216,N_2983,N_2962);
or UO_217 (O_217,N_2992,N_2994);
nor UO_218 (O_218,N_2953,N_2995);
or UO_219 (O_219,N_2960,N_2972);
or UO_220 (O_220,N_2978,N_2963);
nor UO_221 (O_221,N_2998,N_2975);
nor UO_222 (O_222,N_2995,N_2988);
xnor UO_223 (O_223,N_2950,N_2981);
nand UO_224 (O_224,N_2988,N_2989);
or UO_225 (O_225,N_2998,N_2951);
nand UO_226 (O_226,N_2965,N_2998);
or UO_227 (O_227,N_2955,N_2989);
nand UO_228 (O_228,N_2980,N_2996);
nand UO_229 (O_229,N_2990,N_2974);
nor UO_230 (O_230,N_2967,N_2985);
or UO_231 (O_231,N_2991,N_2979);
and UO_232 (O_232,N_2950,N_2991);
nor UO_233 (O_233,N_2977,N_2982);
nor UO_234 (O_234,N_2959,N_2953);
nor UO_235 (O_235,N_2984,N_2975);
and UO_236 (O_236,N_2983,N_2978);
nand UO_237 (O_237,N_2983,N_2954);
and UO_238 (O_238,N_2960,N_2990);
or UO_239 (O_239,N_2963,N_2954);
and UO_240 (O_240,N_2977,N_2985);
nand UO_241 (O_241,N_2996,N_2991);
and UO_242 (O_242,N_2952,N_2956);
and UO_243 (O_243,N_2951,N_2975);
and UO_244 (O_244,N_2994,N_2983);
or UO_245 (O_245,N_2997,N_2990);
nor UO_246 (O_246,N_2961,N_2958);
or UO_247 (O_247,N_2986,N_2984);
nand UO_248 (O_248,N_2965,N_2954);
nor UO_249 (O_249,N_2982,N_2963);
nand UO_250 (O_250,N_2996,N_2964);
nor UO_251 (O_251,N_2982,N_2961);
nand UO_252 (O_252,N_2971,N_2959);
or UO_253 (O_253,N_2969,N_2972);
and UO_254 (O_254,N_2986,N_2955);
nand UO_255 (O_255,N_2954,N_2993);
or UO_256 (O_256,N_2997,N_2970);
xor UO_257 (O_257,N_2951,N_2997);
nand UO_258 (O_258,N_2976,N_2963);
or UO_259 (O_259,N_2975,N_2990);
nor UO_260 (O_260,N_2976,N_2989);
and UO_261 (O_261,N_2963,N_2999);
and UO_262 (O_262,N_2968,N_2959);
nor UO_263 (O_263,N_2986,N_2953);
nor UO_264 (O_264,N_2985,N_2951);
or UO_265 (O_265,N_2963,N_2966);
nand UO_266 (O_266,N_2950,N_2965);
or UO_267 (O_267,N_2969,N_2966);
or UO_268 (O_268,N_2994,N_2990);
or UO_269 (O_269,N_2954,N_2986);
nor UO_270 (O_270,N_2975,N_2955);
or UO_271 (O_271,N_2987,N_2999);
or UO_272 (O_272,N_2987,N_2995);
nor UO_273 (O_273,N_2972,N_2993);
or UO_274 (O_274,N_2954,N_2990);
and UO_275 (O_275,N_2950,N_2962);
and UO_276 (O_276,N_2960,N_2955);
nor UO_277 (O_277,N_2990,N_2965);
nor UO_278 (O_278,N_2980,N_2989);
nand UO_279 (O_279,N_2973,N_2996);
nor UO_280 (O_280,N_2952,N_2966);
or UO_281 (O_281,N_2993,N_2980);
or UO_282 (O_282,N_2999,N_2959);
or UO_283 (O_283,N_2960,N_2961);
nand UO_284 (O_284,N_2979,N_2986);
nor UO_285 (O_285,N_2968,N_2989);
nand UO_286 (O_286,N_2977,N_2954);
nor UO_287 (O_287,N_2967,N_2996);
and UO_288 (O_288,N_2959,N_2978);
nand UO_289 (O_289,N_2979,N_2981);
and UO_290 (O_290,N_2996,N_2950);
or UO_291 (O_291,N_2952,N_2970);
or UO_292 (O_292,N_2995,N_2975);
nand UO_293 (O_293,N_2952,N_2964);
or UO_294 (O_294,N_2951,N_2983);
nor UO_295 (O_295,N_2971,N_2983);
nand UO_296 (O_296,N_2978,N_2950);
or UO_297 (O_297,N_2988,N_2990);
nand UO_298 (O_298,N_2972,N_2999);
or UO_299 (O_299,N_2963,N_2985);
or UO_300 (O_300,N_2984,N_2987);
and UO_301 (O_301,N_2993,N_2962);
nor UO_302 (O_302,N_2976,N_2993);
nor UO_303 (O_303,N_2989,N_2952);
or UO_304 (O_304,N_2968,N_2976);
and UO_305 (O_305,N_2976,N_2965);
or UO_306 (O_306,N_2968,N_2990);
nand UO_307 (O_307,N_2972,N_2952);
or UO_308 (O_308,N_2969,N_2996);
nor UO_309 (O_309,N_2977,N_2951);
nand UO_310 (O_310,N_2985,N_2988);
and UO_311 (O_311,N_2964,N_2978);
nor UO_312 (O_312,N_2977,N_2970);
nor UO_313 (O_313,N_2989,N_2985);
or UO_314 (O_314,N_2991,N_2984);
nor UO_315 (O_315,N_2991,N_2992);
nor UO_316 (O_316,N_2977,N_2995);
or UO_317 (O_317,N_2953,N_2975);
and UO_318 (O_318,N_2979,N_2961);
nor UO_319 (O_319,N_2998,N_2953);
and UO_320 (O_320,N_2993,N_2992);
or UO_321 (O_321,N_2995,N_2952);
and UO_322 (O_322,N_2983,N_2982);
or UO_323 (O_323,N_2992,N_2973);
or UO_324 (O_324,N_2983,N_2981);
nor UO_325 (O_325,N_2961,N_2959);
nand UO_326 (O_326,N_2991,N_2988);
or UO_327 (O_327,N_2996,N_2960);
nand UO_328 (O_328,N_2973,N_2989);
nand UO_329 (O_329,N_2956,N_2987);
and UO_330 (O_330,N_2959,N_2963);
or UO_331 (O_331,N_2960,N_2956);
or UO_332 (O_332,N_2990,N_2984);
nand UO_333 (O_333,N_2987,N_2989);
and UO_334 (O_334,N_2972,N_2954);
nor UO_335 (O_335,N_2953,N_2956);
nor UO_336 (O_336,N_2970,N_2964);
xor UO_337 (O_337,N_2979,N_2983);
and UO_338 (O_338,N_2972,N_2975);
nand UO_339 (O_339,N_2957,N_2960);
nor UO_340 (O_340,N_2961,N_2956);
nand UO_341 (O_341,N_2996,N_2956);
nand UO_342 (O_342,N_2984,N_2998);
and UO_343 (O_343,N_2971,N_2999);
xor UO_344 (O_344,N_2971,N_2964);
xnor UO_345 (O_345,N_2967,N_2987);
nand UO_346 (O_346,N_2957,N_2956);
and UO_347 (O_347,N_2969,N_2974);
nor UO_348 (O_348,N_2997,N_2994);
and UO_349 (O_349,N_2964,N_2993);
nor UO_350 (O_350,N_2962,N_2964);
and UO_351 (O_351,N_2991,N_2961);
and UO_352 (O_352,N_2953,N_2952);
nor UO_353 (O_353,N_2956,N_2963);
or UO_354 (O_354,N_2985,N_2975);
xor UO_355 (O_355,N_2991,N_2990);
and UO_356 (O_356,N_2978,N_2982);
or UO_357 (O_357,N_2951,N_2971);
nor UO_358 (O_358,N_2975,N_2996);
nor UO_359 (O_359,N_2994,N_2955);
and UO_360 (O_360,N_2952,N_2992);
nor UO_361 (O_361,N_2950,N_2964);
nor UO_362 (O_362,N_2960,N_2963);
or UO_363 (O_363,N_2956,N_2979);
nand UO_364 (O_364,N_2988,N_2959);
nand UO_365 (O_365,N_2956,N_2992);
xnor UO_366 (O_366,N_2975,N_2977);
nand UO_367 (O_367,N_2972,N_2985);
nor UO_368 (O_368,N_2994,N_2986);
and UO_369 (O_369,N_2987,N_2985);
or UO_370 (O_370,N_2957,N_2967);
or UO_371 (O_371,N_2981,N_2996);
nor UO_372 (O_372,N_2997,N_2982);
and UO_373 (O_373,N_2994,N_2989);
nand UO_374 (O_374,N_2958,N_2998);
nor UO_375 (O_375,N_2967,N_2974);
nor UO_376 (O_376,N_2968,N_2977);
or UO_377 (O_377,N_2961,N_2980);
and UO_378 (O_378,N_2952,N_2975);
and UO_379 (O_379,N_2984,N_2988);
nor UO_380 (O_380,N_2980,N_2958);
nand UO_381 (O_381,N_2964,N_2966);
xor UO_382 (O_382,N_2969,N_2985);
nand UO_383 (O_383,N_2988,N_2952);
nor UO_384 (O_384,N_2978,N_2996);
or UO_385 (O_385,N_2999,N_2964);
nand UO_386 (O_386,N_2977,N_2952);
or UO_387 (O_387,N_2981,N_2962);
nand UO_388 (O_388,N_2981,N_2982);
or UO_389 (O_389,N_2970,N_2967);
and UO_390 (O_390,N_2983,N_2992);
and UO_391 (O_391,N_2975,N_2999);
or UO_392 (O_392,N_2958,N_2953);
and UO_393 (O_393,N_2976,N_2981);
and UO_394 (O_394,N_2989,N_2969);
nor UO_395 (O_395,N_2997,N_2957);
and UO_396 (O_396,N_2970,N_2950);
and UO_397 (O_397,N_2963,N_2988);
or UO_398 (O_398,N_2966,N_2995);
nand UO_399 (O_399,N_2983,N_2986);
nand UO_400 (O_400,N_2951,N_2950);
and UO_401 (O_401,N_2976,N_2983);
nand UO_402 (O_402,N_2960,N_2966);
nor UO_403 (O_403,N_2970,N_2978);
and UO_404 (O_404,N_2952,N_2959);
xor UO_405 (O_405,N_2950,N_2966);
and UO_406 (O_406,N_2954,N_2964);
nand UO_407 (O_407,N_2971,N_2986);
nand UO_408 (O_408,N_2968,N_2965);
nor UO_409 (O_409,N_2985,N_2952);
or UO_410 (O_410,N_2957,N_2955);
or UO_411 (O_411,N_2984,N_2992);
or UO_412 (O_412,N_2963,N_2996);
nor UO_413 (O_413,N_2955,N_2990);
nor UO_414 (O_414,N_2978,N_2968);
and UO_415 (O_415,N_2977,N_2996);
and UO_416 (O_416,N_2957,N_2961);
nor UO_417 (O_417,N_2955,N_2998);
or UO_418 (O_418,N_2989,N_2993);
or UO_419 (O_419,N_2963,N_2998);
nor UO_420 (O_420,N_2964,N_2972);
nor UO_421 (O_421,N_2964,N_2951);
and UO_422 (O_422,N_2981,N_2958);
nand UO_423 (O_423,N_2963,N_2975);
nor UO_424 (O_424,N_2984,N_2952);
or UO_425 (O_425,N_2963,N_2983);
or UO_426 (O_426,N_2963,N_2992);
and UO_427 (O_427,N_2996,N_2988);
nand UO_428 (O_428,N_2997,N_2954);
nand UO_429 (O_429,N_2963,N_2952);
nand UO_430 (O_430,N_2992,N_2971);
nor UO_431 (O_431,N_2983,N_2997);
nor UO_432 (O_432,N_2966,N_2997);
and UO_433 (O_433,N_2987,N_2974);
nor UO_434 (O_434,N_2979,N_2968);
or UO_435 (O_435,N_2952,N_2987);
nor UO_436 (O_436,N_2969,N_2962);
or UO_437 (O_437,N_2968,N_2994);
nor UO_438 (O_438,N_2976,N_2987);
and UO_439 (O_439,N_2973,N_2987);
nand UO_440 (O_440,N_2966,N_2957);
or UO_441 (O_441,N_2997,N_2962);
or UO_442 (O_442,N_2989,N_2992);
nor UO_443 (O_443,N_2997,N_2979);
nor UO_444 (O_444,N_2961,N_2994);
or UO_445 (O_445,N_2990,N_2970);
nor UO_446 (O_446,N_2961,N_2968);
nand UO_447 (O_447,N_2967,N_2998);
or UO_448 (O_448,N_2975,N_2978);
nor UO_449 (O_449,N_2951,N_2987);
xor UO_450 (O_450,N_2993,N_2977);
and UO_451 (O_451,N_2983,N_2953);
or UO_452 (O_452,N_2959,N_2956);
nand UO_453 (O_453,N_2997,N_2971);
and UO_454 (O_454,N_2959,N_2979);
and UO_455 (O_455,N_2967,N_2975);
xor UO_456 (O_456,N_2955,N_2992);
or UO_457 (O_457,N_2981,N_2955);
nand UO_458 (O_458,N_2986,N_2959);
nor UO_459 (O_459,N_2963,N_2973);
nor UO_460 (O_460,N_2965,N_2964);
nor UO_461 (O_461,N_2967,N_2997);
nor UO_462 (O_462,N_2999,N_2958);
nor UO_463 (O_463,N_2953,N_2973);
nand UO_464 (O_464,N_2999,N_2968);
nor UO_465 (O_465,N_2968,N_2997);
and UO_466 (O_466,N_2987,N_2996);
nand UO_467 (O_467,N_2989,N_2975);
and UO_468 (O_468,N_2999,N_2979);
nand UO_469 (O_469,N_2979,N_2985);
or UO_470 (O_470,N_2953,N_2962);
nor UO_471 (O_471,N_2960,N_2976);
and UO_472 (O_472,N_2969,N_2954);
nor UO_473 (O_473,N_2992,N_2954);
nand UO_474 (O_474,N_2960,N_2967);
nand UO_475 (O_475,N_2983,N_2960);
nand UO_476 (O_476,N_2984,N_2982);
or UO_477 (O_477,N_2986,N_2970);
nand UO_478 (O_478,N_2991,N_2983);
or UO_479 (O_479,N_2965,N_2966);
nand UO_480 (O_480,N_2980,N_2957);
or UO_481 (O_481,N_2978,N_2976);
or UO_482 (O_482,N_2970,N_2958);
or UO_483 (O_483,N_2963,N_2986);
nor UO_484 (O_484,N_2980,N_2978);
and UO_485 (O_485,N_2970,N_2959);
nor UO_486 (O_486,N_2967,N_2978);
and UO_487 (O_487,N_2999,N_2995);
nand UO_488 (O_488,N_2952,N_2994);
nand UO_489 (O_489,N_2997,N_2980);
or UO_490 (O_490,N_2981,N_2990);
nor UO_491 (O_491,N_2966,N_2985);
nand UO_492 (O_492,N_2970,N_2991);
nor UO_493 (O_493,N_2980,N_2968);
and UO_494 (O_494,N_2980,N_2984);
or UO_495 (O_495,N_2998,N_2968);
or UO_496 (O_496,N_2997,N_2953);
or UO_497 (O_497,N_2986,N_2995);
nand UO_498 (O_498,N_2950,N_2954);
nor UO_499 (O_499,N_2956,N_2958);
endmodule