module basic_750_5000_1000_10_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_356,In_172);
nor U1 (N_1,In_724,In_312);
or U2 (N_2,In_640,In_41);
nor U3 (N_3,In_630,In_10);
nand U4 (N_4,In_326,In_639);
nor U5 (N_5,In_106,In_484);
and U6 (N_6,In_60,In_345);
nor U7 (N_7,In_252,In_352);
and U8 (N_8,In_350,In_121);
and U9 (N_9,In_66,In_288);
and U10 (N_10,In_522,In_478);
nor U11 (N_11,In_569,In_310);
nand U12 (N_12,In_470,In_155);
or U13 (N_13,In_464,In_582);
nor U14 (N_14,In_289,In_163);
and U15 (N_15,In_670,In_315);
or U16 (N_16,In_131,In_87);
nand U17 (N_17,In_114,In_229);
and U18 (N_18,In_319,In_605);
or U19 (N_19,In_634,In_578);
nor U20 (N_20,In_604,In_526);
nand U21 (N_21,In_94,In_328);
and U22 (N_22,In_437,In_553);
or U23 (N_23,In_392,In_727);
or U24 (N_24,In_378,In_462);
or U25 (N_25,In_151,In_199);
or U26 (N_26,In_46,In_287);
and U27 (N_27,In_258,In_255);
nand U28 (N_28,In_446,In_689);
nor U29 (N_29,In_124,In_203);
or U30 (N_30,In_701,In_644);
and U31 (N_31,In_54,In_20);
and U32 (N_32,In_428,In_188);
nor U33 (N_33,In_308,In_683);
and U34 (N_34,In_561,In_589);
nor U35 (N_35,In_463,In_50);
or U36 (N_36,In_195,In_190);
nand U37 (N_37,In_460,In_362);
xor U38 (N_38,In_682,In_196);
nand U39 (N_39,In_520,In_548);
or U40 (N_40,In_506,In_280);
nand U41 (N_41,In_129,In_442);
nand U42 (N_42,In_127,In_562);
and U43 (N_43,In_135,In_403);
and U44 (N_44,In_435,In_343);
nand U45 (N_45,In_646,In_304);
or U46 (N_46,In_427,In_735);
nand U47 (N_47,In_498,In_744);
nor U48 (N_48,In_448,In_104);
and U49 (N_49,In_268,In_438);
nand U50 (N_50,In_489,In_603);
nor U51 (N_51,In_278,In_545);
nand U52 (N_52,In_309,In_47);
nand U53 (N_53,In_598,In_500);
and U54 (N_54,In_574,In_714);
nand U55 (N_55,In_523,In_33);
or U56 (N_56,In_338,In_390);
or U57 (N_57,In_633,In_732);
nor U58 (N_58,In_361,In_314);
and U59 (N_59,In_414,In_141);
or U60 (N_60,In_445,In_547);
nor U61 (N_61,In_111,In_524);
or U62 (N_62,In_185,In_697);
nor U63 (N_63,In_595,In_167);
nand U64 (N_64,In_486,In_510);
and U65 (N_65,In_576,In_730);
and U66 (N_66,In_406,In_453);
or U67 (N_67,In_371,In_681);
nand U68 (N_68,In_231,In_596);
and U69 (N_69,In_243,In_126);
and U70 (N_70,In_704,In_497);
nor U71 (N_71,In_409,In_80);
nand U72 (N_72,In_159,In_7);
or U73 (N_73,In_81,In_337);
nor U74 (N_74,In_713,In_236);
nand U75 (N_75,In_148,In_24);
and U76 (N_76,In_330,In_291);
nor U77 (N_77,In_105,In_218);
nor U78 (N_78,In_217,In_327);
nor U79 (N_79,In_721,In_147);
and U80 (N_80,In_373,In_139);
nor U81 (N_81,In_23,In_62);
and U82 (N_82,In_279,In_737);
nand U83 (N_83,In_723,In_251);
nand U84 (N_84,In_495,In_230);
nand U85 (N_85,In_662,In_469);
or U86 (N_86,In_181,In_137);
nor U87 (N_87,In_96,In_663);
and U88 (N_88,In_55,In_257);
or U89 (N_89,In_26,In_125);
and U90 (N_90,In_581,In_281);
or U91 (N_91,In_655,In_742);
and U92 (N_92,In_164,In_197);
nand U93 (N_93,In_38,In_465);
or U94 (N_94,In_136,In_563);
nand U95 (N_95,In_717,In_3);
and U96 (N_96,In_690,In_146);
nor U97 (N_97,In_4,In_535);
and U98 (N_98,In_696,In_456);
xor U99 (N_99,In_206,In_511);
nand U100 (N_100,In_570,In_408);
and U101 (N_101,In_75,In_193);
nor U102 (N_102,In_567,In_397);
or U103 (N_103,In_573,In_450);
and U104 (N_104,In_283,In_31);
nor U105 (N_105,In_64,In_360);
nor U106 (N_106,In_659,In_566);
and U107 (N_107,In_99,In_457);
nor U108 (N_108,In_198,In_443);
xnor U109 (N_109,In_529,In_669);
or U110 (N_110,In_439,In_29);
and U111 (N_111,In_241,In_6);
nor U112 (N_112,In_128,In_739);
nor U113 (N_113,In_564,In_297);
and U114 (N_114,In_142,In_364);
and U115 (N_115,In_179,In_487);
nor U116 (N_116,In_607,In_57);
or U117 (N_117,In_592,In_447);
nand U118 (N_118,In_347,In_368);
nand U119 (N_119,In_219,In_533);
and U120 (N_120,In_194,In_247);
or U121 (N_121,In_377,In_132);
nor U122 (N_122,In_317,In_693);
or U123 (N_123,In_554,In_176);
nand U124 (N_124,In_558,In_461);
or U125 (N_125,In_245,In_534);
or U126 (N_126,In_264,In_538);
or U127 (N_127,In_149,In_215);
or U128 (N_128,In_45,In_119);
nand U129 (N_129,In_358,In_402);
nor U130 (N_130,In_40,In_5);
xor U131 (N_131,In_216,In_299);
or U132 (N_132,In_665,In_286);
nand U133 (N_133,In_606,In_521);
or U134 (N_134,In_676,In_134);
and U135 (N_135,In_441,In_674);
and U136 (N_136,In_587,In_260);
nor U137 (N_137,In_494,In_560);
or U138 (N_138,In_452,In_16);
and U139 (N_139,In_375,In_440);
and U140 (N_140,In_168,In_161);
or U141 (N_141,In_583,In_635);
xor U142 (N_142,In_749,In_282);
or U143 (N_143,In_232,In_374);
nand U144 (N_144,In_747,In_515);
or U145 (N_145,In_539,In_579);
nand U146 (N_146,In_459,In_333);
nor U147 (N_147,In_242,In_746);
nor U148 (N_148,In_708,In_37);
nand U149 (N_149,In_525,In_228);
and U150 (N_150,In_22,In_209);
nand U151 (N_151,In_654,In_399);
nand U152 (N_152,In_89,In_725);
or U153 (N_153,In_156,In_340);
or U154 (N_154,In_543,In_184);
and U155 (N_155,In_458,In_613);
or U156 (N_156,In_711,In_101);
or U157 (N_157,In_656,In_542);
and U158 (N_158,In_324,In_472);
or U159 (N_159,In_366,In_12);
nand U160 (N_160,In_468,In_76);
nand U161 (N_161,In_369,In_187);
or U162 (N_162,In_715,In_741);
or U163 (N_163,In_51,In_290);
nor U164 (N_164,In_731,In_158);
and U165 (N_165,In_413,In_651);
and U166 (N_166,In_244,In_175);
nor U167 (N_167,In_471,In_429);
and U168 (N_168,In_536,In_444);
nor U169 (N_169,In_387,In_295);
and U170 (N_170,In_449,In_201);
and U171 (N_171,In_417,In_718);
or U172 (N_172,In_313,In_454);
and U173 (N_173,In_380,In_19);
nor U174 (N_174,In_227,In_35);
nand U175 (N_175,In_680,In_671);
and U176 (N_176,In_572,In_138);
and U177 (N_177,In_467,In_678);
nand U178 (N_178,In_590,In_699);
nand U179 (N_179,In_367,In_30);
and U180 (N_180,In_733,In_17);
and U181 (N_181,In_505,In_389);
nor U182 (N_182,In_70,In_27);
nor U183 (N_183,In_637,In_621);
nand U184 (N_184,In_615,In_165);
nand U185 (N_185,In_152,In_745);
nor U186 (N_186,In_234,In_379);
nor U187 (N_187,In_157,In_239);
nand U188 (N_188,In_113,In_476);
or U189 (N_189,In_95,In_349);
nor U190 (N_190,In_226,In_684);
nand U191 (N_191,In_48,In_11);
and U192 (N_192,In_36,In_477);
or U193 (N_193,In_643,In_618);
or U194 (N_194,In_544,In_346);
or U195 (N_195,In_632,In_394);
and U196 (N_196,In_357,In_180);
and U197 (N_197,In_620,In_102);
or U198 (N_198,In_235,In_556);
and U199 (N_199,In_39,In_650);
or U200 (N_200,In_586,In_68);
and U201 (N_201,In_479,In_200);
or U202 (N_202,In_423,In_424);
nor U203 (N_203,In_381,In_58);
or U204 (N_204,In_174,In_551);
and U205 (N_205,In_117,In_336);
xor U206 (N_206,In_648,In_116);
nand U207 (N_207,In_677,In_455);
or U208 (N_208,In_254,In_153);
or U209 (N_209,In_483,In_485);
nor U210 (N_210,In_514,In_303);
and U211 (N_211,In_609,In_416);
xor U212 (N_212,In_720,In_473);
nand U213 (N_213,In_599,In_593);
or U214 (N_214,In_436,In_395);
nor U215 (N_215,In_425,In_559);
nor U216 (N_216,In_496,In_658);
or U217 (N_217,In_594,In_318);
and U218 (N_218,In_667,In_186);
and U219 (N_219,In_32,In_143);
and U220 (N_220,In_173,In_610);
nor U221 (N_221,In_237,In_355);
xnor U222 (N_222,In_382,In_531);
nor U223 (N_223,In_202,In_528);
and U224 (N_224,In_332,In_178);
and U225 (N_225,In_97,In_600);
and U226 (N_226,In_365,In_335);
nand U227 (N_227,In_384,In_133);
and U228 (N_228,In_518,In_666);
nand U229 (N_229,In_614,In_123);
and U230 (N_230,In_616,In_706);
and U231 (N_231,In_657,In_246);
and U232 (N_232,In_171,In_433);
and U233 (N_233,In_169,In_224);
nor U234 (N_234,In_293,In_591);
xor U235 (N_235,In_418,In_284);
and U236 (N_236,In_623,In_44);
nor U237 (N_237,In_405,In_679);
and U238 (N_238,In_700,In_385);
nand U239 (N_239,In_555,In_67);
and U240 (N_240,In_398,In_625);
nand U241 (N_241,In_546,In_59);
or U242 (N_242,In_311,In_517);
nand U243 (N_243,In_348,In_624);
and U244 (N_244,In_557,In_503);
or U245 (N_245,In_65,In_519);
nand U246 (N_246,In_601,In_72);
nor U247 (N_247,In_210,In_419);
nand U248 (N_248,In_636,In_370);
nor U249 (N_249,In_617,In_69);
xnor U250 (N_250,In_276,In_56);
and U251 (N_251,In_103,In_363);
nand U252 (N_252,In_166,In_144);
nand U253 (N_253,In_645,In_302);
nor U254 (N_254,In_233,In_28);
nor U255 (N_255,In_507,In_73);
nand U256 (N_256,In_339,In_1);
nand U257 (N_257,In_647,In_292);
nand U258 (N_258,In_716,In_63);
or U259 (N_259,In_743,In_710);
nand U260 (N_260,In_513,In_294);
nor U261 (N_261,In_552,In_422);
nor U262 (N_262,In_100,In_25);
and U263 (N_263,In_488,In_92);
nand U264 (N_264,In_703,In_359);
and U265 (N_265,In_316,In_480);
nand U266 (N_266,In_493,In_376);
and U267 (N_267,In_83,In_688);
or U268 (N_268,In_736,In_150);
or U269 (N_269,In_602,In_627);
nand U270 (N_270,In_532,In_432);
nand U271 (N_271,In_722,In_274);
nand U272 (N_272,In_430,In_296);
nor U273 (N_273,In_325,In_298);
nand U274 (N_274,In_410,In_481);
nor U275 (N_275,In_222,In_388);
nand U276 (N_276,In_431,In_391);
nand U277 (N_277,In_492,In_262);
nand U278 (N_278,In_619,In_734);
nand U279 (N_279,In_502,In_334);
nand U280 (N_280,In_110,In_565);
nand U281 (N_281,In_691,In_191);
and U282 (N_282,In_628,In_482);
nand U283 (N_283,In_275,In_162);
nand U284 (N_284,In_189,In_154);
and U285 (N_285,In_629,In_49);
nor U286 (N_286,In_698,In_223);
nor U287 (N_287,In_214,In_675);
or U288 (N_288,In_273,In_568);
or U289 (N_289,In_145,In_9);
nand U290 (N_290,In_71,In_306);
or U291 (N_291,In_537,In_709);
and U292 (N_292,In_15,In_277);
nand U293 (N_293,In_98,In_571);
nor U294 (N_294,In_401,In_74);
xor U295 (N_295,In_322,In_263);
and U296 (N_296,In_673,In_272);
or U297 (N_297,In_331,In_52);
or U298 (N_298,In_88,In_78);
nand U299 (N_299,In_420,In_211);
nand U300 (N_300,In_323,In_386);
nor U301 (N_301,In_740,In_383);
nand U302 (N_302,In_354,In_466);
nand U303 (N_303,In_549,In_649);
nand U304 (N_304,In_412,In_240);
nor U305 (N_305,In_626,In_160);
and U306 (N_306,In_695,In_42);
and U307 (N_307,In_259,In_719);
and U308 (N_308,In_192,In_305);
nand U309 (N_309,In_491,In_585);
or U310 (N_310,In_170,In_90);
nor U311 (N_311,In_307,In_0);
nand U312 (N_312,In_652,In_238);
xnor U313 (N_313,In_748,In_269);
nor U314 (N_314,In_641,In_653);
xnor U315 (N_315,In_256,In_415);
and U316 (N_316,In_501,In_597);
nor U317 (N_317,In_738,In_271);
or U318 (N_318,In_253,In_120);
nor U319 (N_319,In_13,In_660);
nand U320 (N_320,In_270,In_301);
and U321 (N_321,In_182,In_85);
and U322 (N_322,In_109,In_248);
nor U323 (N_323,In_686,In_407);
nand U324 (N_324,In_611,In_115);
and U325 (N_325,In_588,In_329);
nor U326 (N_326,In_122,In_729);
or U327 (N_327,In_250,In_207);
nor U328 (N_328,In_266,In_685);
nand U329 (N_329,In_661,In_212);
nor U330 (N_330,In_475,In_14);
nor U331 (N_331,In_622,In_396);
nor U332 (N_332,In_61,In_404);
nor U333 (N_333,In_177,In_261);
nor U334 (N_334,In_93,In_208);
or U335 (N_335,In_687,In_107);
or U336 (N_336,In_130,In_638);
nand U337 (N_337,In_541,In_584);
or U338 (N_338,In_265,In_577);
nor U339 (N_339,In_118,In_712);
and U340 (N_340,In_580,In_504);
nor U341 (N_341,In_575,In_411);
and U342 (N_342,In_426,In_393);
nor U343 (N_343,In_77,In_672);
or U344 (N_344,In_267,In_474);
nand U345 (N_345,In_344,In_21);
and U346 (N_346,In_82,In_53);
and U347 (N_347,In_2,In_509);
nor U348 (N_348,In_8,In_527);
and U349 (N_349,In_285,In_702);
and U350 (N_350,In_530,In_512);
or U351 (N_351,In_726,In_351);
xnor U352 (N_352,In_668,In_300);
nand U353 (N_353,In_540,In_372);
nand U354 (N_354,In_707,In_490);
or U355 (N_355,In_108,In_642);
nor U356 (N_356,In_320,In_353);
or U357 (N_357,In_728,In_608);
nor U358 (N_358,In_112,In_213);
and U359 (N_359,In_84,In_221);
nand U360 (N_360,In_220,In_204);
or U361 (N_361,In_341,In_664);
and U362 (N_362,In_225,In_140);
or U363 (N_363,In_550,In_421);
or U364 (N_364,In_86,In_451);
nor U365 (N_365,In_692,In_91);
nor U366 (N_366,In_342,In_18);
or U367 (N_367,In_705,In_43);
or U368 (N_368,In_249,In_321);
or U369 (N_369,In_499,In_205);
xnor U370 (N_370,In_400,In_694);
nand U371 (N_371,In_612,In_508);
and U372 (N_372,In_34,In_434);
nand U373 (N_373,In_183,In_631);
and U374 (N_374,In_516,In_79);
and U375 (N_375,In_150,In_586);
nand U376 (N_376,In_399,In_423);
and U377 (N_377,In_56,In_559);
xnor U378 (N_378,In_322,In_312);
nor U379 (N_379,In_690,In_551);
and U380 (N_380,In_549,In_64);
nor U381 (N_381,In_45,In_360);
nand U382 (N_382,In_144,In_338);
nor U383 (N_383,In_482,In_169);
nand U384 (N_384,In_596,In_64);
nand U385 (N_385,In_543,In_464);
or U386 (N_386,In_247,In_650);
nand U387 (N_387,In_615,In_127);
and U388 (N_388,In_268,In_263);
or U389 (N_389,In_403,In_324);
nor U390 (N_390,In_639,In_244);
nand U391 (N_391,In_568,In_330);
and U392 (N_392,In_330,In_591);
or U393 (N_393,In_470,In_425);
nor U394 (N_394,In_724,In_323);
or U395 (N_395,In_469,In_715);
nor U396 (N_396,In_541,In_397);
and U397 (N_397,In_440,In_234);
and U398 (N_398,In_221,In_635);
nor U399 (N_399,In_20,In_428);
nand U400 (N_400,In_337,In_382);
and U401 (N_401,In_12,In_308);
and U402 (N_402,In_340,In_746);
or U403 (N_403,In_200,In_63);
nand U404 (N_404,In_241,In_402);
nand U405 (N_405,In_440,In_729);
nand U406 (N_406,In_19,In_165);
nor U407 (N_407,In_674,In_166);
nand U408 (N_408,In_258,In_204);
and U409 (N_409,In_55,In_439);
and U410 (N_410,In_505,In_7);
and U411 (N_411,In_658,In_570);
nor U412 (N_412,In_21,In_628);
xor U413 (N_413,In_427,In_650);
xor U414 (N_414,In_514,In_283);
nand U415 (N_415,In_2,In_642);
nand U416 (N_416,In_150,In_261);
or U417 (N_417,In_414,In_221);
nand U418 (N_418,In_269,In_141);
or U419 (N_419,In_136,In_724);
or U420 (N_420,In_572,In_217);
or U421 (N_421,In_671,In_298);
and U422 (N_422,In_7,In_498);
and U423 (N_423,In_337,In_637);
or U424 (N_424,In_2,In_282);
or U425 (N_425,In_652,In_672);
and U426 (N_426,In_518,In_124);
nor U427 (N_427,In_190,In_136);
nor U428 (N_428,In_633,In_691);
nor U429 (N_429,In_186,In_153);
nand U430 (N_430,In_222,In_88);
nor U431 (N_431,In_436,In_401);
nor U432 (N_432,In_47,In_577);
and U433 (N_433,In_541,In_420);
nand U434 (N_434,In_215,In_503);
and U435 (N_435,In_446,In_383);
nand U436 (N_436,In_174,In_645);
and U437 (N_437,In_239,In_337);
or U438 (N_438,In_650,In_372);
nand U439 (N_439,In_608,In_430);
nand U440 (N_440,In_261,In_512);
nor U441 (N_441,In_708,In_305);
and U442 (N_442,In_315,In_351);
nor U443 (N_443,In_380,In_529);
nor U444 (N_444,In_707,In_293);
nand U445 (N_445,In_20,In_162);
nand U446 (N_446,In_327,In_622);
and U447 (N_447,In_407,In_742);
nand U448 (N_448,In_254,In_571);
and U449 (N_449,In_473,In_56);
or U450 (N_450,In_370,In_126);
and U451 (N_451,In_562,In_551);
or U452 (N_452,In_214,In_555);
nor U453 (N_453,In_270,In_108);
nor U454 (N_454,In_206,In_311);
and U455 (N_455,In_615,In_136);
nor U456 (N_456,In_3,In_5);
nor U457 (N_457,In_401,In_502);
and U458 (N_458,In_198,In_291);
or U459 (N_459,In_564,In_63);
nand U460 (N_460,In_134,In_407);
nand U461 (N_461,In_478,In_588);
or U462 (N_462,In_588,In_637);
nor U463 (N_463,In_444,In_51);
and U464 (N_464,In_66,In_145);
nand U465 (N_465,In_458,In_595);
and U466 (N_466,In_224,In_138);
or U467 (N_467,In_341,In_268);
nand U468 (N_468,In_180,In_171);
or U469 (N_469,In_664,In_492);
and U470 (N_470,In_742,In_49);
or U471 (N_471,In_655,In_392);
or U472 (N_472,In_501,In_48);
nor U473 (N_473,In_354,In_595);
and U474 (N_474,In_213,In_143);
or U475 (N_475,In_108,In_180);
or U476 (N_476,In_321,In_62);
nor U477 (N_477,In_558,In_349);
xnor U478 (N_478,In_113,In_378);
or U479 (N_479,In_142,In_379);
nor U480 (N_480,In_200,In_127);
nor U481 (N_481,In_51,In_607);
or U482 (N_482,In_96,In_656);
or U483 (N_483,In_212,In_283);
or U484 (N_484,In_242,In_218);
or U485 (N_485,In_176,In_680);
and U486 (N_486,In_395,In_644);
nor U487 (N_487,In_290,In_271);
nor U488 (N_488,In_310,In_10);
and U489 (N_489,In_680,In_242);
nor U490 (N_490,In_215,In_659);
or U491 (N_491,In_544,In_550);
nor U492 (N_492,In_429,In_641);
nand U493 (N_493,In_259,In_735);
and U494 (N_494,In_700,In_278);
nor U495 (N_495,In_163,In_292);
nor U496 (N_496,In_183,In_215);
or U497 (N_497,In_591,In_4);
nand U498 (N_498,In_214,In_553);
and U499 (N_499,In_690,In_652);
nor U500 (N_500,N_59,N_343);
nand U501 (N_501,N_131,N_492);
nor U502 (N_502,N_295,N_222);
or U503 (N_503,N_266,N_341);
and U504 (N_504,N_57,N_221);
nor U505 (N_505,N_172,N_108);
nor U506 (N_506,N_361,N_237);
nor U507 (N_507,N_356,N_477);
nand U508 (N_508,N_335,N_283);
or U509 (N_509,N_475,N_324);
or U510 (N_510,N_365,N_58);
and U511 (N_511,N_248,N_163);
or U512 (N_512,N_480,N_269);
or U513 (N_513,N_357,N_85);
nand U514 (N_514,N_88,N_438);
or U515 (N_515,N_265,N_91);
nand U516 (N_516,N_26,N_408);
xnor U517 (N_517,N_359,N_35);
and U518 (N_518,N_473,N_472);
and U519 (N_519,N_351,N_194);
and U520 (N_520,N_141,N_417);
nand U521 (N_521,N_465,N_282);
nand U522 (N_522,N_39,N_214);
nand U523 (N_523,N_232,N_441);
nor U524 (N_524,N_268,N_235);
nand U525 (N_525,N_130,N_3);
nor U526 (N_526,N_411,N_211);
nor U527 (N_527,N_174,N_491);
or U528 (N_528,N_354,N_116);
or U529 (N_529,N_117,N_393);
nand U530 (N_530,N_318,N_281);
or U531 (N_531,N_405,N_421);
or U532 (N_532,N_476,N_319);
or U533 (N_533,N_423,N_159);
nor U534 (N_534,N_449,N_120);
nor U535 (N_535,N_305,N_121);
and U536 (N_536,N_327,N_245);
nor U537 (N_537,N_100,N_155);
nand U538 (N_538,N_320,N_350);
and U539 (N_539,N_311,N_5);
or U540 (N_540,N_161,N_24);
nor U541 (N_541,N_382,N_242);
nand U542 (N_542,N_30,N_276);
nand U543 (N_543,N_12,N_287);
xnor U544 (N_544,N_367,N_176);
and U545 (N_545,N_96,N_387);
nand U546 (N_546,N_13,N_239);
nand U547 (N_547,N_455,N_160);
or U548 (N_548,N_450,N_360);
nor U549 (N_549,N_252,N_389);
nor U550 (N_550,N_209,N_499);
or U551 (N_551,N_256,N_427);
and U552 (N_552,N_437,N_136);
nand U553 (N_553,N_412,N_383);
and U554 (N_554,N_369,N_33);
and U555 (N_555,N_145,N_115);
or U556 (N_556,N_386,N_302);
and U557 (N_557,N_123,N_177);
nor U558 (N_558,N_90,N_200);
and U559 (N_559,N_1,N_229);
or U560 (N_560,N_373,N_485);
nor U561 (N_561,N_346,N_309);
or U562 (N_562,N_67,N_328);
nand U563 (N_563,N_173,N_468);
or U564 (N_564,N_192,N_493);
nand U565 (N_565,N_169,N_395);
xor U566 (N_566,N_271,N_363);
nand U567 (N_567,N_81,N_352);
or U568 (N_568,N_144,N_203);
nor U569 (N_569,N_128,N_340);
nand U570 (N_570,N_488,N_315);
and U571 (N_571,N_394,N_40);
and U572 (N_572,N_261,N_213);
xnor U573 (N_573,N_9,N_253);
nand U574 (N_574,N_288,N_375);
xnor U575 (N_575,N_385,N_380);
and U576 (N_576,N_304,N_11);
or U577 (N_577,N_7,N_279);
or U578 (N_578,N_443,N_110);
nor U579 (N_579,N_138,N_204);
and U580 (N_580,N_22,N_48);
nor U581 (N_581,N_378,N_422);
and U582 (N_582,N_399,N_482);
xnor U583 (N_583,N_93,N_95);
nand U584 (N_584,N_436,N_366);
or U585 (N_585,N_274,N_300);
or U586 (N_586,N_409,N_339);
nand U587 (N_587,N_381,N_296);
or U588 (N_588,N_151,N_153);
and U589 (N_589,N_36,N_379);
nand U590 (N_590,N_0,N_218);
nand U591 (N_591,N_18,N_495);
nand U592 (N_592,N_255,N_27);
nand U593 (N_593,N_165,N_162);
nand U594 (N_594,N_466,N_303);
and U595 (N_595,N_196,N_202);
and U596 (N_596,N_215,N_267);
nor U597 (N_597,N_69,N_77);
nand U598 (N_598,N_34,N_38);
nand U599 (N_599,N_306,N_164);
and U600 (N_600,N_212,N_29);
nor U601 (N_601,N_259,N_16);
and U602 (N_602,N_28,N_78);
and U603 (N_603,N_56,N_19);
xnor U604 (N_604,N_23,N_25);
nand U605 (N_605,N_246,N_126);
or U606 (N_606,N_206,N_316);
and U607 (N_607,N_406,N_481);
and U608 (N_608,N_483,N_486);
or U609 (N_609,N_157,N_80);
or U610 (N_610,N_452,N_122);
and U611 (N_611,N_413,N_461);
nand U612 (N_612,N_178,N_73);
and U613 (N_613,N_10,N_228);
or U614 (N_614,N_97,N_111);
or U615 (N_615,N_314,N_462);
nand U616 (N_616,N_396,N_390);
or U617 (N_617,N_453,N_220);
xnor U618 (N_618,N_479,N_407);
or U619 (N_619,N_113,N_496);
or U620 (N_620,N_275,N_330);
or U621 (N_621,N_82,N_249);
and U622 (N_622,N_277,N_197);
nor U623 (N_623,N_227,N_105);
nand U624 (N_624,N_109,N_101);
or U625 (N_625,N_250,N_43);
nand U626 (N_626,N_258,N_41);
or U627 (N_627,N_338,N_273);
nand U628 (N_628,N_332,N_290);
nor U629 (N_629,N_297,N_47);
or U630 (N_630,N_460,N_182);
or U631 (N_631,N_429,N_284);
nor U632 (N_632,N_185,N_294);
and U633 (N_633,N_31,N_166);
and U634 (N_634,N_447,N_345);
or U635 (N_635,N_124,N_428);
nand U636 (N_636,N_60,N_133);
and U637 (N_637,N_474,N_127);
nand U638 (N_638,N_326,N_310);
nand U639 (N_639,N_293,N_175);
xnor U640 (N_640,N_167,N_53);
or U641 (N_641,N_299,N_333);
and U642 (N_642,N_112,N_189);
nand U643 (N_643,N_317,N_168);
or U644 (N_644,N_156,N_377);
or U645 (N_645,N_334,N_397);
and U646 (N_646,N_125,N_454);
or U647 (N_647,N_42,N_420);
or U648 (N_648,N_52,N_8);
or U649 (N_649,N_187,N_102);
or U650 (N_650,N_191,N_439);
nor U651 (N_651,N_17,N_464);
nor U652 (N_652,N_87,N_402);
and U653 (N_653,N_83,N_329);
nor U654 (N_654,N_65,N_372);
nand U655 (N_655,N_376,N_118);
nand U656 (N_656,N_446,N_463);
nand U657 (N_657,N_348,N_150);
and U658 (N_658,N_219,N_431);
or U659 (N_659,N_226,N_490);
and U660 (N_660,N_289,N_414);
or U661 (N_661,N_171,N_233);
nor U662 (N_662,N_236,N_254);
or U663 (N_663,N_45,N_15);
xor U664 (N_664,N_199,N_139);
and U665 (N_665,N_240,N_32);
nor U666 (N_666,N_364,N_494);
nand U667 (N_667,N_181,N_99);
xor U668 (N_668,N_404,N_50);
or U669 (N_669,N_238,N_331);
or U670 (N_670,N_49,N_119);
nor U671 (N_671,N_426,N_400);
or U672 (N_672,N_68,N_79);
or U673 (N_673,N_358,N_312);
and U674 (N_674,N_484,N_2);
nand U675 (N_675,N_291,N_134);
and U676 (N_676,N_370,N_86);
nand U677 (N_677,N_457,N_37);
and U678 (N_678,N_264,N_241);
nand U679 (N_679,N_70,N_243);
or U680 (N_680,N_280,N_132);
or U681 (N_681,N_51,N_64);
nand U682 (N_682,N_244,N_21);
nor U683 (N_683,N_489,N_442);
nor U684 (N_684,N_63,N_391);
nand U685 (N_685,N_349,N_445);
nor U686 (N_686,N_292,N_46);
nand U687 (N_687,N_301,N_190);
nor U688 (N_688,N_403,N_75);
nand U689 (N_689,N_129,N_216);
xor U690 (N_690,N_247,N_223);
nor U691 (N_691,N_322,N_440);
nor U692 (N_692,N_234,N_179);
nand U693 (N_693,N_362,N_323);
nand U694 (N_694,N_217,N_398);
or U695 (N_695,N_61,N_207);
nor U696 (N_696,N_307,N_106);
nand U697 (N_697,N_195,N_342);
or U698 (N_698,N_84,N_135);
nor U699 (N_699,N_210,N_321);
and U700 (N_700,N_231,N_154);
nand U701 (N_701,N_251,N_107);
or U702 (N_702,N_66,N_262);
and U703 (N_703,N_478,N_142);
nor U704 (N_704,N_392,N_419);
and U705 (N_705,N_434,N_469);
or U706 (N_706,N_208,N_140);
or U707 (N_707,N_487,N_415);
or U708 (N_708,N_143,N_225);
or U709 (N_709,N_470,N_98);
nand U710 (N_710,N_344,N_149);
and U711 (N_711,N_355,N_180);
nor U712 (N_712,N_201,N_471);
or U713 (N_713,N_336,N_92);
or U714 (N_714,N_146,N_325);
nor U715 (N_715,N_298,N_71);
or U716 (N_716,N_497,N_76);
nor U717 (N_717,N_152,N_263);
and U718 (N_718,N_451,N_44);
or U719 (N_719,N_384,N_347);
and U720 (N_720,N_147,N_4);
or U721 (N_721,N_104,N_416);
or U722 (N_722,N_94,N_270);
and U723 (N_723,N_278,N_114);
nand U724 (N_724,N_170,N_257);
or U725 (N_725,N_425,N_186);
or U726 (N_726,N_435,N_433);
nor U727 (N_727,N_418,N_424);
and U728 (N_728,N_148,N_14);
or U729 (N_729,N_158,N_410);
nand U730 (N_730,N_272,N_458);
nand U731 (N_731,N_137,N_459);
nor U732 (N_732,N_353,N_401);
nand U733 (N_733,N_188,N_193);
xnor U734 (N_734,N_371,N_103);
or U735 (N_735,N_374,N_183);
or U736 (N_736,N_498,N_205);
or U737 (N_737,N_260,N_368);
nor U738 (N_738,N_456,N_285);
and U739 (N_739,N_20,N_430);
and U740 (N_740,N_313,N_55);
nand U741 (N_741,N_444,N_184);
nor U742 (N_742,N_337,N_388);
nand U743 (N_743,N_448,N_62);
nand U744 (N_744,N_432,N_224);
nand U745 (N_745,N_89,N_6);
and U746 (N_746,N_308,N_230);
or U747 (N_747,N_467,N_198);
nor U748 (N_748,N_54,N_286);
nor U749 (N_749,N_74,N_72);
or U750 (N_750,N_284,N_223);
nor U751 (N_751,N_319,N_62);
or U752 (N_752,N_33,N_159);
nor U753 (N_753,N_150,N_108);
nor U754 (N_754,N_203,N_214);
and U755 (N_755,N_435,N_383);
and U756 (N_756,N_472,N_336);
nand U757 (N_757,N_418,N_327);
or U758 (N_758,N_92,N_182);
nor U759 (N_759,N_55,N_173);
nor U760 (N_760,N_266,N_126);
and U761 (N_761,N_191,N_435);
nand U762 (N_762,N_238,N_386);
and U763 (N_763,N_9,N_483);
and U764 (N_764,N_337,N_497);
and U765 (N_765,N_111,N_357);
nand U766 (N_766,N_436,N_456);
nand U767 (N_767,N_104,N_167);
nand U768 (N_768,N_200,N_117);
nand U769 (N_769,N_85,N_259);
and U770 (N_770,N_325,N_436);
nand U771 (N_771,N_230,N_167);
nand U772 (N_772,N_67,N_433);
nand U773 (N_773,N_212,N_237);
or U774 (N_774,N_181,N_37);
and U775 (N_775,N_186,N_114);
and U776 (N_776,N_8,N_225);
nand U777 (N_777,N_420,N_253);
and U778 (N_778,N_473,N_109);
nand U779 (N_779,N_143,N_239);
nor U780 (N_780,N_388,N_36);
or U781 (N_781,N_291,N_409);
nand U782 (N_782,N_163,N_266);
nor U783 (N_783,N_61,N_3);
or U784 (N_784,N_69,N_237);
nor U785 (N_785,N_490,N_375);
xor U786 (N_786,N_388,N_173);
or U787 (N_787,N_387,N_252);
and U788 (N_788,N_339,N_493);
or U789 (N_789,N_175,N_300);
nor U790 (N_790,N_409,N_121);
nand U791 (N_791,N_257,N_87);
nand U792 (N_792,N_101,N_208);
nand U793 (N_793,N_335,N_422);
nor U794 (N_794,N_187,N_120);
and U795 (N_795,N_470,N_362);
nand U796 (N_796,N_157,N_319);
or U797 (N_797,N_219,N_493);
nand U798 (N_798,N_19,N_138);
or U799 (N_799,N_180,N_129);
nor U800 (N_800,N_1,N_158);
or U801 (N_801,N_50,N_458);
or U802 (N_802,N_143,N_244);
or U803 (N_803,N_48,N_305);
nand U804 (N_804,N_69,N_15);
nand U805 (N_805,N_196,N_367);
nor U806 (N_806,N_200,N_301);
or U807 (N_807,N_392,N_386);
and U808 (N_808,N_470,N_359);
or U809 (N_809,N_131,N_329);
nand U810 (N_810,N_187,N_301);
xnor U811 (N_811,N_434,N_30);
nand U812 (N_812,N_480,N_202);
nor U813 (N_813,N_492,N_368);
nor U814 (N_814,N_378,N_199);
nor U815 (N_815,N_403,N_2);
or U816 (N_816,N_88,N_259);
nand U817 (N_817,N_317,N_104);
nand U818 (N_818,N_246,N_163);
nor U819 (N_819,N_252,N_458);
or U820 (N_820,N_19,N_275);
nand U821 (N_821,N_305,N_412);
and U822 (N_822,N_3,N_132);
nor U823 (N_823,N_222,N_160);
and U824 (N_824,N_11,N_140);
and U825 (N_825,N_232,N_56);
or U826 (N_826,N_187,N_198);
and U827 (N_827,N_12,N_473);
nand U828 (N_828,N_103,N_136);
nor U829 (N_829,N_288,N_17);
or U830 (N_830,N_472,N_428);
and U831 (N_831,N_130,N_255);
and U832 (N_832,N_91,N_5);
nor U833 (N_833,N_332,N_435);
nand U834 (N_834,N_161,N_431);
and U835 (N_835,N_172,N_208);
nand U836 (N_836,N_137,N_388);
nand U837 (N_837,N_395,N_316);
or U838 (N_838,N_106,N_95);
or U839 (N_839,N_127,N_252);
or U840 (N_840,N_250,N_48);
or U841 (N_841,N_71,N_482);
or U842 (N_842,N_13,N_89);
and U843 (N_843,N_121,N_455);
and U844 (N_844,N_20,N_442);
nor U845 (N_845,N_167,N_428);
or U846 (N_846,N_182,N_371);
and U847 (N_847,N_481,N_111);
or U848 (N_848,N_287,N_66);
and U849 (N_849,N_265,N_270);
nand U850 (N_850,N_136,N_402);
nand U851 (N_851,N_121,N_144);
or U852 (N_852,N_340,N_131);
or U853 (N_853,N_213,N_405);
or U854 (N_854,N_86,N_332);
or U855 (N_855,N_177,N_86);
nor U856 (N_856,N_282,N_347);
or U857 (N_857,N_104,N_31);
and U858 (N_858,N_267,N_429);
nor U859 (N_859,N_402,N_443);
nor U860 (N_860,N_398,N_32);
nand U861 (N_861,N_59,N_358);
and U862 (N_862,N_424,N_336);
nor U863 (N_863,N_172,N_61);
and U864 (N_864,N_382,N_109);
or U865 (N_865,N_396,N_98);
and U866 (N_866,N_102,N_337);
or U867 (N_867,N_477,N_229);
nand U868 (N_868,N_70,N_259);
nor U869 (N_869,N_407,N_51);
nor U870 (N_870,N_290,N_250);
and U871 (N_871,N_339,N_438);
nand U872 (N_872,N_110,N_63);
and U873 (N_873,N_116,N_40);
nor U874 (N_874,N_344,N_421);
nor U875 (N_875,N_449,N_244);
and U876 (N_876,N_90,N_405);
nor U877 (N_877,N_426,N_133);
and U878 (N_878,N_444,N_317);
nor U879 (N_879,N_185,N_163);
xor U880 (N_880,N_336,N_485);
and U881 (N_881,N_55,N_101);
and U882 (N_882,N_265,N_108);
and U883 (N_883,N_139,N_430);
nor U884 (N_884,N_393,N_150);
and U885 (N_885,N_115,N_423);
nor U886 (N_886,N_27,N_130);
nor U887 (N_887,N_361,N_161);
and U888 (N_888,N_102,N_136);
and U889 (N_889,N_218,N_388);
nand U890 (N_890,N_276,N_455);
and U891 (N_891,N_256,N_343);
nor U892 (N_892,N_171,N_52);
xnor U893 (N_893,N_457,N_47);
or U894 (N_894,N_416,N_389);
and U895 (N_895,N_462,N_358);
or U896 (N_896,N_394,N_331);
or U897 (N_897,N_424,N_154);
or U898 (N_898,N_480,N_445);
nand U899 (N_899,N_403,N_66);
nand U900 (N_900,N_468,N_90);
nand U901 (N_901,N_242,N_385);
and U902 (N_902,N_182,N_467);
and U903 (N_903,N_250,N_17);
and U904 (N_904,N_497,N_444);
and U905 (N_905,N_411,N_228);
or U906 (N_906,N_127,N_417);
nor U907 (N_907,N_85,N_312);
nand U908 (N_908,N_292,N_162);
nand U909 (N_909,N_473,N_497);
nor U910 (N_910,N_251,N_15);
nand U911 (N_911,N_399,N_233);
nand U912 (N_912,N_132,N_395);
nor U913 (N_913,N_354,N_60);
or U914 (N_914,N_353,N_390);
and U915 (N_915,N_349,N_397);
nor U916 (N_916,N_321,N_272);
xnor U917 (N_917,N_82,N_28);
and U918 (N_918,N_48,N_164);
or U919 (N_919,N_161,N_299);
nor U920 (N_920,N_379,N_101);
nor U921 (N_921,N_34,N_430);
nor U922 (N_922,N_166,N_463);
or U923 (N_923,N_128,N_322);
nand U924 (N_924,N_114,N_296);
nor U925 (N_925,N_186,N_159);
or U926 (N_926,N_337,N_434);
and U927 (N_927,N_351,N_106);
nand U928 (N_928,N_179,N_388);
xnor U929 (N_929,N_451,N_436);
or U930 (N_930,N_117,N_261);
nor U931 (N_931,N_480,N_171);
nand U932 (N_932,N_56,N_499);
nor U933 (N_933,N_32,N_298);
nand U934 (N_934,N_438,N_490);
and U935 (N_935,N_372,N_62);
nor U936 (N_936,N_251,N_456);
nand U937 (N_937,N_193,N_178);
and U938 (N_938,N_430,N_394);
or U939 (N_939,N_142,N_355);
and U940 (N_940,N_117,N_432);
and U941 (N_941,N_259,N_83);
nor U942 (N_942,N_285,N_291);
nor U943 (N_943,N_5,N_319);
or U944 (N_944,N_155,N_47);
nor U945 (N_945,N_333,N_173);
and U946 (N_946,N_242,N_341);
or U947 (N_947,N_407,N_98);
and U948 (N_948,N_329,N_305);
or U949 (N_949,N_352,N_58);
or U950 (N_950,N_440,N_336);
nand U951 (N_951,N_212,N_135);
nor U952 (N_952,N_483,N_406);
nand U953 (N_953,N_94,N_464);
nor U954 (N_954,N_119,N_439);
and U955 (N_955,N_347,N_133);
and U956 (N_956,N_469,N_238);
nand U957 (N_957,N_400,N_153);
nand U958 (N_958,N_116,N_124);
nor U959 (N_959,N_152,N_366);
nand U960 (N_960,N_447,N_33);
and U961 (N_961,N_79,N_360);
nand U962 (N_962,N_151,N_229);
nor U963 (N_963,N_213,N_197);
nand U964 (N_964,N_329,N_169);
nand U965 (N_965,N_23,N_67);
nor U966 (N_966,N_41,N_223);
and U967 (N_967,N_332,N_402);
or U968 (N_968,N_24,N_439);
and U969 (N_969,N_301,N_105);
nor U970 (N_970,N_412,N_421);
and U971 (N_971,N_352,N_431);
nand U972 (N_972,N_159,N_277);
nand U973 (N_973,N_422,N_372);
nand U974 (N_974,N_124,N_101);
nand U975 (N_975,N_490,N_294);
or U976 (N_976,N_498,N_420);
or U977 (N_977,N_453,N_374);
nor U978 (N_978,N_406,N_382);
and U979 (N_979,N_235,N_34);
or U980 (N_980,N_118,N_347);
or U981 (N_981,N_420,N_277);
and U982 (N_982,N_232,N_165);
nor U983 (N_983,N_405,N_219);
nor U984 (N_984,N_85,N_329);
nor U985 (N_985,N_486,N_63);
xor U986 (N_986,N_115,N_21);
nor U987 (N_987,N_239,N_145);
nand U988 (N_988,N_151,N_70);
nor U989 (N_989,N_45,N_460);
or U990 (N_990,N_197,N_431);
nand U991 (N_991,N_379,N_369);
or U992 (N_992,N_145,N_25);
and U993 (N_993,N_202,N_331);
or U994 (N_994,N_201,N_489);
nand U995 (N_995,N_375,N_333);
nor U996 (N_996,N_302,N_454);
nor U997 (N_997,N_103,N_184);
nand U998 (N_998,N_13,N_143);
or U999 (N_999,N_111,N_409);
or U1000 (N_1000,N_597,N_971);
and U1001 (N_1001,N_998,N_838);
or U1002 (N_1002,N_809,N_978);
nor U1003 (N_1003,N_933,N_717);
nor U1004 (N_1004,N_648,N_864);
xnor U1005 (N_1005,N_728,N_736);
nand U1006 (N_1006,N_907,N_512);
or U1007 (N_1007,N_955,N_990);
or U1008 (N_1008,N_820,N_901);
nand U1009 (N_1009,N_531,N_965);
or U1010 (N_1010,N_787,N_614);
and U1011 (N_1011,N_945,N_560);
nand U1012 (N_1012,N_631,N_724);
xor U1013 (N_1013,N_924,N_942);
and U1014 (N_1014,N_869,N_959);
nor U1015 (N_1015,N_984,N_659);
nand U1016 (N_1016,N_992,N_503);
nor U1017 (N_1017,N_879,N_610);
or U1018 (N_1018,N_985,N_528);
nor U1019 (N_1019,N_582,N_700);
nor U1020 (N_1020,N_989,N_943);
or U1021 (N_1021,N_516,N_583);
nand U1022 (N_1022,N_609,N_630);
nand U1023 (N_1023,N_876,N_977);
nor U1024 (N_1024,N_602,N_702);
or U1025 (N_1025,N_675,N_592);
nand U1026 (N_1026,N_829,N_756);
nand U1027 (N_1027,N_634,N_904);
and U1028 (N_1028,N_510,N_673);
nor U1029 (N_1029,N_680,N_605);
nor U1030 (N_1030,N_727,N_735);
nand U1031 (N_1031,N_967,N_962);
nor U1032 (N_1032,N_543,N_914);
and U1033 (N_1033,N_637,N_890);
nor U1034 (N_1034,N_733,N_851);
or U1035 (N_1035,N_612,N_797);
and U1036 (N_1036,N_526,N_807);
nand U1037 (N_1037,N_784,N_645);
xnor U1038 (N_1038,N_628,N_931);
and U1039 (N_1039,N_906,N_939);
or U1040 (N_1040,N_867,N_881);
or U1041 (N_1041,N_566,N_611);
or U1042 (N_1042,N_655,N_948);
nand U1043 (N_1043,N_969,N_885);
nor U1044 (N_1044,N_828,N_830);
nand U1045 (N_1045,N_649,N_753);
nand U1046 (N_1046,N_685,N_875);
and U1047 (N_1047,N_552,N_619);
nor U1048 (N_1048,N_672,N_987);
nand U1049 (N_1049,N_690,N_658);
or U1050 (N_1050,N_932,N_520);
nand U1051 (N_1051,N_922,N_589);
or U1052 (N_1052,N_849,N_621);
xor U1053 (N_1053,N_535,N_586);
or U1054 (N_1054,N_646,N_693);
nor U1055 (N_1055,N_796,N_755);
nand U1056 (N_1056,N_670,N_816);
nor U1057 (N_1057,N_776,N_683);
and U1058 (N_1058,N_994,N_719);
or U1059 (N_1059,N_622,N_633);
or U1060 (N_1060,N_979,N_928);
and U1061 (N_1061,N_749,N_635);
and U1062 (N_1062,N_781,N_926);
nand U1063 (N_1063,N_530,N_811);
and U1064 (N_1064,N_911,N_506);
nor U1065 (N_1065,N_529,N_833);
nor U1066 (N_1066,N_620,N_825);
nor U1067 (N_1067,N_587,N_910);
nand U1068 (N_1068,N_862,N_661);
or U1069 (N_1069,N_815,N_803);
nand U1070 (N_1070,N_522,N_832);
nand U1071 (N_1071,N_903,N_762);
and U1072 (N_1072,N_854,N_738);
nand U1073 (N_1073,N_714,N_773);
and U1074 (N_1074,N_871,N_938);
and U1075 (N_1075,N_786,N_653);
and U1076 (N_1076,N_523,N_580);
and U1077 (N_1077,N_766,N_791);
nand U1078 (N_1078,N_537,N_663);
or U1079 (N_1079,N_853,N_555);
and U1080 (N_1080,N_944,N_843);
nor U1081 (N_1081,N_794,N_823);
or U1082 (N_1082,N_940,N_930);
or U1083 (N_1083,N_720,N_841);
and U1084 (N_1084,N_742,N_684);
and U1085 (N_1085,N_826,N_750);
or U1086 (N_1086,N_629,N_565);
nand U1087 (N_1087,N_761,N_613);
and U1088 (N_1088,N_793,N_568);
nor U1089 (N_1089,N_827,N_704);
nand U1090 (N_1090,N_790,N_958);
and U1091 (N_1091,N_961,N_687);
nor U1092 (N_1092,N_688,N_866);
or U1093 (N_1093,N_639,N_997);
or U1094 (N_1094,N_554,N_647);
or U1095 (N_1095,N_991,N_974);
and U1096 (N_1096,N_918,N_559);
and U1097 (N_1097,N_842,N_596);
and U1098 (N_1098,N_970,N_578);
nand U1099 (N_1099,N_547,N_763);
nand U1100 (N_1100,N_892,N_627);
and U1101 (N_1101,N_908,N_674);
nand U1102 (N_1102,N_860,N_544);
or U1103 (N_1103,N_575,N_590);
nor U1104 (N_1104,N_817,N_725);
nor U1105 (N_1105,N_946,N_777);
xor U1106 (N_1106,N_935,N_534);
nand U1107 (N_1107,N_744,N_874);
nor U1108 (N_1108,N_912,N_599);
nor U1109 (N_1109,N_723,N_746);
and U1110 (N_1110,N_643,N_950);
nor U1111 (N_1111,N_505,N_561);
nand U1112 (N_1112,N_972,N_863);
or U1113 (N_1113,N_713,N_595);
or U1114 (N_1114,N_898,N_508);
or U1115 (N_1115,N_995,N_837);
xor U1116 (N_1116,N_600,N_999);
nor U1117 (N_1117,N_515,N_665);
nor U1118 (N_1118,N_546,N_752);
nor U1119 (N_1119,N_701,N_868);
or U1120 (N_1120,N_834,N_802);
nand U1121 (N_1121,N_934,N_657);
and U1122 (N_1122,N_651,N_801);
nor U1123 (N_1123,N_988,N_986);
nor U1124 (N_1124,N_740,N_859);
and U1125 (N_1125,N_699,N_968);
or U1126 (N_1126,N_536,N_981);
and U1127 (N_1127,N_588,N_694);
nor U1128 (N_1128,N_897,N_716);
nor U1129 (N_1129,N_800,N_812);
nor U1130 (N_1130,N_920,N_877);
or U1131 (N_1131,N_973,N_564);
nand U1132 (N_1132,N_601,N_598);
and U1133 (N_1133,N_677,N_654);
or U1134 (N_1134,N_818,N_804);
and U1135 (N_1135,N_513,N_913);
and U1136 (N_1136,N_521,N_636);
or U1137 (N_1137,N_840,N_887);
or U1138 (N_1138,N_993,N_916);
nor U1139 (N_1139,N_921,N_792);
nand U1140 (N_1140,N_509,N_632);
nor U1141 (N_1141,N_896,N_872);
nor U1142 (N_1142,N_626,N_567);
nor U1143 (N_1143,N_710,N_532);
nand U1144 (N_1144,N_511,N_855);
or U1145 (N_1145,N_571,N_795);
nor U1146 (N_1146,N_782,N_617);
nor U1147 (N_1147,N_712,N_810);
xnor U1148 (N_1148,N_765,N_551);
nor U1149 (N_1149,N_669,N_715);
nor U1150 (N_1150,N_572,N_960);
nor U1151 (N_1151,N_861,N_718);
and U1152 (N_1152,N_603,N_808);
nor U1153 (N_1153,N_917,N_604);
and U1154 (N_1154,N_865,N_905);
nor U1155 (N_1155,N_697,N_780);
nand U1156 (N_1156,N_731,N_642);
or U1157 (N_1157,N_774,N_982);
xor U1158 (N_1158,N_562,N_668);
nand U1159 (N_1159,N_707,N_739);
nor U1160 (N_1160,N_574,N_754);
and U1161 (N_1161,N_557,N_660);
nand U1162 (N_1162,N_788,N_770);
nand U1163 (N_1163,N_726,N_734);
nand U1164 (N_1164,N_732,N_949);
nor U1165 (N_1165,N_751,N_846);
and U1166 (N_1166,N_764,N_813);
or U1167 (N_1167,N_757,N_937);
nand U1168 (N_1168,N_593,N_856);
and U1169 (N_1169,N_689,N_504);
nor U1170 (N_1170,N_667,N_692);
nand U1171 (N_1171,N_894,N_640);
nor U1172 (N_1172,N_524,N_963);
nand U1173 (N_1173,N_679,N_570);
or U1174 (N_1174,N_553,N_721);
nor U1175 (N_1175,N_591,N_616);
and U1176 (N_1176,N_666,N_691);
or U1177 (N_1177,N_549,N_775);
nor U1178 (N_1178,N_835,N_641);
nor U1179 (N_1179,N_839,N_759);
or U1180 (N_1180,N_698,N_569);
nor U1181 (N_1181,N_623,N_947);
or U1182 (N_1182,N_706,N_915);
or U1183 (N_1183,N_548,N_929);
nand U1184 (N_1184,N_686,N_664);
or U1185 (N_1185,N_883,N_880);
and U1186 (N_1186,N_767,N_644);
or U1187 (N_1187,N_507,N_606);
or U1188 (N_1188,N_848,N_518);
and U1189 (N_1189,N_953,N_743);
or U1190 (N_1190,N_671,N_824);
and U1191 (N_1191,N_585,N_836);
and U1192 (N_1192,N_577,N_747);
or U1193 (N_1193,N_941,N_996);
nand U1194 (N_1194,N_656,N_500);
and U1195 (N_1195,N_760,N_709);
or U1196 (N_1196,N_847,N_579);
or U1197 (N_1197,N_975,N_772);
or U1198 (N_1198,N_638,N_729);
and U1199 (N_1199,N_805,N_983);
nand U1200 (N_1200,N_966,N_514);
nor U1201 (N_1201,N_618,N_819);
and U1202 (N_1202,N_711,N_799);
and U1203 (N_1203,N_519,N_576);
nand U1204 (N_1204,N_541,N_878);
nand U1205 (N_1205,N_769,N_745);
nand U1206 (N_1206,N_852,N_703);
nor U1207 (N_1207,N_539,N_785);
and U1208 (N_1208,N_925,N_730);
and U1209 (N_1209,N_558,N_678);
nand U1210 (N_1210,N_936,N_771);
or U1211 (N_1211,N_798,N_889);
nand U1212 (N_1212,N_741,N_822);
and U1213 (N_1213,N_676,N_682);
nand U1214 (N_1214,N_951,N_884);
or U1215 (N_1215,N_844,N_895);
or U1216 (N_1216,N_882,N_550);
nor U1217 (N_1217,N_758,N_527);
and U1218 (N_1218,N_594,N_737);
nor U1219 (N_1219,N_909,N_814);
and U1220 (N_1220,N_545,N_584);
or U1221 (N_1221,N_538,N_722);
or U1222 (N_1222,N_783,N_650);
and U1223 (N_1223,N_517,N_705);
nor U1224 (N_1224,N_573,N_857);
nor U1225 (N_1225,N_886,N_831);
nor U1226 (N_1226,N_540,N_789);
or U1227 (N_1227,N_533,N_581);
and U1228 (N_1228,N_608,N_964);
or U1229 (N_1229,N_888,N_607);
nor U1230 (N_1230,N_768,N_624);
xor U1231 (N_1231,N_806,N_927);
nor U1232 (N_1232,N_748,N_957);
or U1233 (N_1233,N_899,N_525);
nor U1234 (N_1234,N_542,N_980);
nor U1235 (N_1235,N_858,N_696);
and U1236 (N_1236,N_956,N_708);
nor U1237 (N_1237,N_952,N_919);
nor U1238 (N_1238,N_976,N_891);
nand U1239 (N_1239,N_954,N_662);
nor U1240 (N_1240,N_845,N_873);
or U1241 (N_1241,N_900,N_779);
or U1242 (N_1242,N_563,N_695);
or U1243 (N_1243,N_850,N_652);
nand U1244 (N_1244,N_625,N_778);
nor U1245 (N_1245,N_821,N_923);
nor U1246 (N_1246,N_502,N_681);
or U1247 (N_1247,N_893,N_615);
nor U1248 (N_1248,N_501,N_902);
nand U1249 (N_1249,N_556,N_870);
nand U1250 (N_1250,N_591,N_500);
and U1251 (N_1251,N_899,N_866);
or U1252 (N_1252,N_805,N_737);
and U1253 (N_1253,N_862,N_659);
and U1254 (N_1254,N_643,N_730);
or U1255 (N_1255,N_973,N_865);
and U1256 (N_1256,N_505,N_629);
nand U1257 (N_1257,N_729,N_840);
nand U1258 (N_1258,N_972,N_925);
nor U1259 (N_1259,N_904,N_716);
nand U1260 (N_1260,N_761,N_660);
or U1261 (N_1261,N_955,N_925);
or U1262 (N_1262,N_513,N_505);
nand U1263 (N_1263,N_597,N_867);
and U1264 (N_1264,N_873,N_604);
nand U1265 (N_1265,N_605,N_649);
nand U1266 (N_1266,N_698,N_805);
nor U1267 (N_1267,N_744,N_960);
nand U1268 (N_1268,N_693,N_744);
and U1269 (N_1269,N_887,N_701);
or U1270 (N_1270,N_809,N_544);
and U1271 (N_1271,N_959,N_835);
or U1272 (N_1272,N_954,N_578);
nor U1273 (N_1273,N_699,N_682);
and U1274 (N_1274,N_782,N_507);
nand U1275 (N_1275,N_751,N_739);
nand U1276 (N_1276,N_787,N_961);
and U1277 (N_1277,N_566,N_797);
or U1278 (N_1278,N_513,N_880);
and U1279 (N_1279,N_963,N_842);
and U1280 (N_1280,N_536,N_942);
nor U1281 (N_1281,N_721,N_921);
nand U1282 (N_1282,N_694,N_507);
nand U1283 (N_1283,N_952,N_912);
nor U1284 (N_1284,N_631,N_643);
nor U1285 (N_1285,N_722,N_708);
or U1286 (N_1286,N_794,N_919);
or U1287 (N_1287,N_501,N_944);
nor U1288 (N_1288,N_503,N_786);
and U1289 (N_1289,N_793,N_504);
or U1290 (N_1290,N_866,N_521);
nor U1291 (N_1291,N_581,N_793);
or U1292 (N_1292,N_519,N_990);
and U1293 (N_1293,N_948,N_641);
nand U1294 (N_1294,N_935,N_514);
or U1295 (N_1295,N_958,N_994);
and U1296 (N_1296,N_862,N_619);
nor U1297 (N_1297,N_625,N_556);
and U1298 (N_1298,N_667,N_737);
or U1299 (N_1299,N_823,N_667);
or U1300 (N_1300,N_502,N_521);
or U1301 (N_1301,N_772,N_603);
nor U1302 (N_1302,N_600,N_886);
or U1303 (N_1303,N_913,N_936);
and U1304 (N_1304,N_815,N_821);
or U1305 (N_1305,N_860,N_924);
and U1306 (N_1306,N_549,N_846);
nor U1307 (N_1307,N_637,N_593);
xor U1308 (N_1308,N_974,N_736);
or U1309 (N_1309,N_710,N_625);
or U1310 (N_1310,N_632,N_961);
or U1311 (N_1311,N_561,N_697);
and U1312 (N_1312,N_778,N_910);
nor U1313 (N_1313,N_682,N_745);
nand U1314 (N_1314,N_996,N_790);
and U1315 (N_1315,N_934,N_959);
nand U1316 (N_1316,N_999,N_604);
or U1317 (N_1317,N_940,N_827);
nor U1318 (N_1318,N_701,N_856);
nor U1319 (N_1319,N_944,N_851);
or U1320 (N_1320,N_814,N_740);
nand U1321 (N_1321,N_950,N_613);
and U1322 (N_1322,N_531,N_566);
nor U1323 (N_1323,N_500,N_676);
or U1324 (N_1324,N_637,N_847);
and U1325 (N_1325,N_720,N_699);
nor U1326 (N_1326,N_998,N_565);
and U1327 (N_1327,N_718,N_509);
nor U1328 (N_1328,N_659,N_578);
xnor U1329 (N_1329,N_516,N_953);
and U1330 (N_1330,N_924,N_943);
nand U1331 (N_1331,N_970,N_881);
xnor U1332 (N_1332,N_857,N_815);
nand U1333 (N_1333,N_831,N_616);
and U1334 (N_1334,N_922,N_787);
xor U1335 (N_1335,N_762,N_815);
and U1336 (N_1336,N_593,N_872);
or U1337 (N_1337,N_860,N_833);
and U1338 (N_1338,N_701,N_816);
xor U1339 (N_1339,N_663,N_949);
or U1340 (N_1340,N_812,N_653);
or U1341 (N_1341,N_934,N_609);
nand U1342 (N_1342,N_587,N_986);
nand U1343 (N_1343,N_903,N_613);
nor U1344 (N_1344,N_697,N_989);
and U1345 (N_1345,N_892,N_914);
and U1346 (N_1346,N_946,N_762);
nor U1347 (N_1347,N_906,N_509);
nand U1348 (N_1348,N_749,N_859);
or U1349 (N_1349,N_933,N_729);
nand U1350 (N_1350,N_537,N_810);
nor U1351 (N_1351,N_682,N_661);
or U1352 (N_1352,N_750,N_821);
nor U1353 (N_1353,N_940,N_751);
xor U1354 (N_1354,N_729,N_985);
and U1355 (N_1355,N_929,N_660);
xnor U1356 (N_1356,N_528,N_732);
nand U1357 (N_1357,N_663,N_635);
nand U1358 (N_1358,N_747,N_513);
or U1359 (N_1359,N_878,N_993);
or U1360 (N_1360,N_746,N_675);
nand U1361 (N_1361,N_612,N_768);
nand U1362 (N_1362,N_603,N_618);
or U1363 (N_1363,N_514,N_875);
or U1364 (N_1364,N_547,N_709);
and U1365 (N_1365,N_570,N_877);
and U1366 (N_1366,N_626,N_949);
nor U1367 (N_1367,N_666,N_977);
and U1368 (N_1368,N_626,N_579);
nand U1369 (N_1369,N_646,N_907);
and U1370 (N_1370,N_690,N_853);
or U1371 (N_1371,N_968,N_638);
or U1372 (N_1372,N_885,N_850);
nor U1373 (N_1373,N_932,N_919);
nor U1374 (N_1374,N_536,N_914);
or U1375 (N_1375,N_871,N_944);
nand U1376 (N_1376,N_631,N_827);
nand U1377 (N_1377,N_789,N_794);
xor U1378 (N_1378,N_573,N_812);
nand U1379 (N_1379,N_828,N_811);
nand U1380 (N_1380,N_906,N_609);
nor U1381 (N_1381,N_686,N_919);
and U1382 (N_1382,N_500,N_797);
nand U1383 (N_1383,N_950,N_511);
nand U1384 (N_1384,N_755,N_937);
nand U1385 (N_1385,N_879,N_713);
nand U1386 (N_1386,N_910,N_560);
or U1387 (N_1387,N_629,N_817);
and U1388 (N_1388,N_710,N_547);
nand U1389 (N_1389,N_623,N_775);
nand U1390 (N_1390,N_839,N_738);
and U1391 (N_1391,N_511,N_859);
and U1392 (N_1392,N_603,N_501);
nor U1393 (N_1393,N_829,N_539);
and U1394 (N_1394,N_510,N_689);
or U1395 (N_1395,N_570,N_958);
nand U1396 (N_1396,N_685,N_848);
nand U1397 (N_1397,N_602,N_745);
or U1398 (N_1398,N_912,N_720);
nand U1399 (N_1399,N_570,N_573);
and U1400 (N_1400,N_601,N_554);
nand U1401 (N_1401,N_779,N_976);
nand U1402 (N_1402,N_963,N_867);
xor U1403 (N_1403,N_842,N_892);
nor U1404 (N_1404,N_553,N_788);
and U1405 (N_1405,N_914,N_722);
nand U1406 (N_1406,N_929,N_839);
xor U1407 (N_1407,N_556,N_803);
nor U1408 (N_1408,N_670,N_578);
nand U1409 (N_1409,N_936,N_615);
and U1410 (N_1410,N_595,N_596);
nand U1411 (N_1411,N_704,N_830);
nand U1412 (N_1412,N_627,N_534);
and U1413 (N_1413,N_509,N_524);
nand U1414 (N_1414,N_794,N_712);
nor U1415 (N_1415,N_779,N_892);
nor U1416 (N_1416,N_706,N_579);
and U1417 (N_1417,N_860,N_647);
or U1418 (N_1418,N_649,N_506);
and U1419 (N_1419,N_726,N_982);
nor U1420 (N_1420,N_604,N_732);
nor U1421 (N_1421,N_851,N_576);
nor U1422 (N_1422,N_939,N_797);
or U1423 (N_1423,N_782,N_542);
nand U1424 (N_1424,N_687,N_823);
and U1425 (N_1425,N_892,N_669);
or U1426 (N_1426,N_790,N_601);
and U1427 (N_1427,N_952,N_959);
and U1428 (N_1428,N_755,N_716);
nor U1429 (N_1429,N_793,N_869);
nand U1430 (N_1430,N_771,N_931);
or U1431 (N_1431,N_974,N_972);
and U1432 (N_1432,N_862,N_925);
and U1433 (N_1433,N_975,N_777);
and U1434 (N_1434,N_771,N_630);
nor U1435 (N_1435,N_713,N_677);
nand U1436 (N_1436,N_929,N_703);
and U1437 (N_1437,N_739,N_554);
nand U1438 (N_1438,N_557,N_684);
or U1439 (N_1439,N_958,N_582);
and U1440 (N_1440,N_701,N_707);
and U1441 (N_1441,N_584,N_991);
nand U1442 (N_1442,N_636,N_659);
or U1443 (N_1443,N_682,N_513);
nand U1444 (N_1444,N_743,N_776);
nor U1445 (N_1445,N_662,N_858);
or U1446 (N_1446,N_687,N_688);
or U1447 (N_1447,N_865,N_683);
or U1448 (N_1448,N_699,N_898);
nor U1449 (N_1449,N_648,N_829);
nor U1450 (N_1450,N_561,N_892);
or U1451 (N_1451,N_776,N_614);
or U1452 (N_1452,N_985,N_767);
or U1453 (N_1453,N_531,N_623);
and U1454 (N_1454,N_900,N_860);
nor U1455 (N_1455,N_862,N_769);
xnor U1456 (N_1456,N_702,N_535);
nand U1457 (N_1457,N_914,N_792);
and U1458 (N_1458,N_652,N_710);
nor U1459 (N_1459,N_804,N_860);
xnor U1460 (N_1460,N_634,N_942);
or U1461 (N_1461,N_900,N_708);
nand U1462 (N_1462,N_685,N_510);
nor U1463 (N_1463,N_990,N_775);
or U1464 (N_1464,N_908,N_842);
and U1465 (N_1465,N_518,N_879);
and U1466 (N_1466,N_735,N_917);
nand U1467 (N_1467,N_666,N_624);
nor U1468 (N_1468,N_828,N_820);
nor U1469 (N_1469,N_647,N_977);
nor U1470 (N_1470,N_997,N_539);
and U1471 (N_1471,N_939,N_650);
or U1472 (N_1472,N_764,N_715);
and U1473 (N_1473,N_550,N_938);
and U1474 (N_1474,N_535,N_936);
or U1475 (N_1475,N_610,N_758);
and U1476 (N_1476,N_571,N_576);
nand U1477 (N_1477,N_701,N_998);
or U1478 (N_1478,N_725,N_804);
and U1479 (N_1479,N_719,N_733);
or U1480 (N_1480,N_776,N_515);
or U1481 (N_1481,N_600,N_576);
nor U1482 (N_1482,N_857,N_692);
nor U1483 (N_1483,N_785,N_782);
and U1484 (N_1484,N_862,N_746);
or U1485 (N_1485,N_658,N_607);
nor U1486 (N_1486,N_668,N_744);
and U1487 (N_1487,N_997,N_738);
and U1488 (N_1488,N_635,N_975);
nand U1489 (N_1489,N_666,N_725);
nor U1490 (N_1490,N_862,N_513);
and U1491 (N_1491,N_771,N_930);
nand U1492 (N_1492,N_612,N_564);
nand U1493 (N_1493,N_611,N_923);
nor U1494 (N_1494,N_881,N_985);
nor U1495 (N_1495,N_829,N_522);
nand U1496 (N_1496,N_803,N_514);
nand U1497 (N_1497,N_801,N_561);
or U1498 (N_1498,N_791,N_654);
or U1499 (N_1499,N_651,N_959);
nand U1500 (N_1500,N_1172,N_1440);
nor U1501 (N_1501,N_1334,N_1108);
nor U1502 (N_1502,N_1078,N_1408);
and U1503 (N_1503,N_1236,N_1422);
nor U1504 (N_1504,N_1030,N_1074);
or U1505 (N_1505,N_1162,N_1188);
xnor U1506 (N_1506,N_1059,N_1204);
nor U1507 (N_1507,N_1446,N_1023);
and U1508 (N_1508,N_1160,N_1038);
nor U1509 (N_1509,N_1146,N_1185);
or U1510 (N_1510,N_1098,N_1212);
xnor U1511 (N_1511,N_1274,N_1497);
or U1512 (N_1512,N_1429,N_1327);
or U1513 (N_1513,N_1383,N_1371);
nor U1514 (N_1514,N_1073,N_1045);
nor U1515 (N_1515,N_1254,N_1243);
and U1516 (N_1516,N_1256,N_1178);
nand U1517 (N_1517,N_1436,N_1443);
or U1518 (N_1518,N_1181,N_1275);
nand U1519 (N_1519,N_1495,N_1482);
nor U1520 (N_1520,N_1329,N_1092);
nand U1521 (N_1521,N_1381,N_1084);
or U1522 (N_1522,N_1117,N_1069);
or U1523 (N_1523,N_1259,N_1199);
nand U1524 (N_1524,N_1270,N_1324);
or U1525 (N_1525,N_1039,N_1197);
and U1526 (N_1526,N_1114,N_1096);
nand U1527 (N_1527,N_1437,N_1289);
nand U1528 (N_1528,N_1113,N_1018);
and U1529 (N_1529,N_1124,N_1339);
nor U1530 (N_1530,N_1128,N_1261);
nor U1531 (N_1531,N_1413,N_1017);
nor U1532 (N_1532,N_1224,N_1161);
and U1533 (N_1533,N_1307,N_1347);
nor U1534 (N_1534,N_1077,N_1125);
and U1535 (N_1535,N_1239,N_1228);
nand U1536 (N_1536,N_1299,N_1068);
nand U1537 (N_1537,N_1200,N_1325);
nor U1538 (N_1538,N_1163,N_1321);
nand U1539 (N_1539,N_1390,N_1460);
or U1540 (N_1540,N_1029,N_1216);
or U1541 (N_1541,N_1341,N_1235);
nand U1542 (N_1542,N_1374,N_1145);
or U1543 (N_1543,N_1222,N_1474);
or U1544 (N_1544,N_1166,N_1496);
and U1545 (N_1545,N_1143,N_1001);
and U1546 (N_1546,N_1294,N_1221);
or U1547 (N_1547,N_1486,N_1396);
or U1548 (N_1548,N_1019,N_1317);
nor U1549 (N_1549,N_1282,N_1064);
or U1550 (N_1550,N_1070,N_1388);
and U1551 (N_1551,N_1491,N_1298);
nor U1552 (N_1552,N_1404,N_1449);
and U1553 (N_1553,N_1398,N_1310);
or U1554 (N_1554,N_1182,N_1387);
and U1555 (N_1555,N_1263,N_1135);
nand U1556 (N_1556,N_1157,N_1260);
or U1557 (N_1557,N_1229,N_1418);
and U1558 (N_1558,N_1444,N_1223);
nand U1559 (N_1559,N_1384,N_1269);
or U1560 (N_1560,N_1133,N_1332);
nand U1561 (N_1561,N_1129,N_1392);
nand U1562 (N_1562,N_1461,N_1245);
nor U1563 (N_1563,N_1369,N_1462);
nor U1564 (N_1564,N_1085,N_1126);
or U1565 (N_1565,N_1463,N_1237);
and U1566 (N_1566,N_1025,N_1430);
nand U1567 (N_1567,N_1112,N_1206);
and U1568 (N_1568,N_1366,N_1424);
nor U1569 (N_1569,N_1058,N_1044);
or U1570 (N_1570,N_1407,N_1082);
nand U1571 (N_1571,N_1072,N_1258);
nor U1572 (N_1572,N_1301,N_1149);
or U1573 (N_1573,N_1006,N_1217);
nand U1574 (N_1574,N_1159,N_1426);
nor U1575 (N_1575,N_1265,N_1210);
nor U1576 (N_1576,N_1350,N_1008);
and U1577 (N_1577,N_1148,N_1304);
xor U1578 (N_1578,N_1293,N_1296);
nand U1579 (N_1579,N_1292,N_1309);
nor U1580 (N_1580,N_1016,N_1391);
or U1581 (N_1581,N_1477,N_1499);
nor U1582 (N_1582,N_1055,N_1331);
or U1583 (N_1583,N_1196,N_1470);
nand U1584 (N_1584,N_1138,N_1397);
nand U1585 (N_1585,N_1238,N_1028);
or U1586 (N_1586,N_1484,N_1107);
or U1587 (N_1587,N_1140,N_1454);
or U1588 (N_1588,N_1090,N_1032);
or U1589 (N_1589,N_1376,N_1343);
nand U1590 (N_1590,N_1231,N_1319);
nor U1591 (N_1591,N_1132,N_1177);
xnor U1592 (N_1592,N_1315,N_1403);
nor U1593 (N_1593,N_1004,N_1455);
or U1594 (N_1594,N_1356,N_1050);
nor U1595 (N_1595,N_1414,N_1399);
and U1596 (N_1596,N_1232,N_1338);
and U1597 (N_1597,N_1021,N_1280);
or U1598 (N_1598,N_1419,N_1036);
nor U1599 (N_1599,N_1027,N_1433);
nor U1600 (N_1600,N_1358,N_1240);
nand U1601 (N_1601,N_1284,N_1186);
and U1602 (N_1602,N_1322,N_1170);
nand U1603 (N_1603,N_1067,N_1119);
nor U1604 (N_1604,N_1115,N_1087);
nor U1605 (N_1605,N_1441,N_1066);
nand U1606 (N_1606,N_1137,N_1445);
nor U1607 (N_1607,N_1155,N_1362);
and U1608 (N_1608,N_1105,N_1102);
or U1609 (N_1609,N_1233,N_1279);
nand U1610 (N_1610,N_1187,N_1048);
nand U1611 (N_1611,N_1230,N_1213);
and U1612 (N_1612,N_1219,N_1352);
or U1613 (N_1613,N_1054,N_1031);
nand U1614 (N_1614,N_1011,N_1337);
nand U1615 (N_1615,N_1435,N_1041);
or U1616 (N_1616,N_1302,N_1227);
xnor U1617 (N_1617,N_1173,N_1361);
nor U1618 (N_1618,N_1106,N_1425);
and U1619 (N_1619,N_1053,N_1349);
nand U1620 (N_1620,N_1333,N_1421);
nand U1621 (N_1621,N_1167,N_1409);
nand U1622 (N_1622,N_1395,N_1348);
and U1623 (N_1623,N_1377,N_1257);
nor U1624 (N_1624,N_1262,N_1379);
nor U1625 (N_1625,N_1415,N_1453);
and U1626 (N_1626,N_1264,N_1225);
nor U1627 (N_1627,N_1340,N_1427);
or U1628 (N_1628,N_1290,N_1479);
or U1629 (N_1629,N_1323,N_1357);
nand U1630 (N_1630,N_1131,N_1364);
or U1631 (N_1631,N_1447,N_1189);
nand U1632 (N_1632,N_1373,N_1056);
or U1633 (N_1633,N_1060,N_1104);
nor U1634 (N_1634,N_1368,N_1130);
nand U1635 (N_1635,N_1351,N_1450);
nand U1636 (N_1636,N_1116,N_1095);
nor U1637 (N_1637,N_1014,N_1168);
or U1638 (N_1638,N_1022,N_1483);
and U1639 (N_1639,N_1393,N_1336);
and U1640 (N_1640,N_1005,N_1089);
and U1641 (N_1641,N_1111,N_1075);
or U1642 (N_1642,N_1291,N_1305);
or U1643 (N_1643,N_1083,N_1490);
or U1644 (N_1644,N_1375,N_1246);
or U1645 (N_1645,N_1494,N_1448);
and U1646 (N_1646,N_1015,N_1320);
xor U1647 (N_1647,N_1266,N_1151);
nand U1648 (N_1648,N_1241,N_1152);
nand U1649 (N_1649,N_1099,N_1451);
nor U1650 (N_1650,N_1311,N_1110);
nand U1651 (N_1651,N_1209,N_1047);
or U1652 (N_1652,N_1285,N_1389);
and U1653 (N_1653,N_1201,N_1150);
and U1654 (N_1654,N_1382,N_1147);
nand U1655 (N_1655,N_1498,N_1295);
nand U1656 (N_1656,N_1158,N_1314);
or U1657 (N_1657,N_1080,N_1434);
nor U1658 (N_1658,N_1024,N_1417);
or U1659 (N_1659,N_1198,N_1492);
nand U1660 (N_1660,N_1308,N_1416);
nor U1661 (N_1661,N_1288,N_1208);
and U1662 (N_1662,N_1442,N_1037);
nor U1663 (N_1663,N_1169,N_1464);
nand U1664 (N_1664,N_1267,N_1247);
or U1665 (N_1665,N_1194,N_1205);
nand U1666 (N_1666,N_1218,N_1471);
nand U1667 (N_1667,N_1481,N_1438);
and U1668 (N_1668,N_1252,N_1202);
or U1669 (N_1669,N_1278,N_1303);
nor U1670 (N_1670,N_1176,N_1093);
or U1671 (N_1671,N_1086,N_1043);
nand U1672 (N_1672,N_1370,N_1156);
and U1673 (N_1673,N_1042,N_1485);
and U1674 (N_1674,N_1428,N_1277);
nand U1675 (N_1675,N_1120,N_1255);
or U1676 (N_1676,N_1183,N_1326);
nor U1677 (N_1677,N_1051,N_1052);
or U1678 (N_1678,N_1091,N_1242);
nor U1679 (N_1679,N_1100,N_1071);
or U1680 (N_1680,N_1012,N_1286);
nand U1681 (N_1681,N_1431,N_1121);
nor U1682 (N_1682,N_1330,N_1355);
nor U1683 (N_1683,N_1345,N_1405);
nand U1684 (N_1684,N_1401,N_1088);
nor U1685 (N_1685,N_1297,N_1476);
nor U1686 (N_1686,N_1040,N_1175);
nor U1687 (N_1687,N_1380,N_1020);
and U1688 (N_1688,N_1094,N_1211);
nor U1689 (N_1689,N_1473,N_1195);
nor U1690 (N_1690,N_1457,N_1142);
nor U1691 (N_1691,N_1010,N_1316);
nand U1692 (N_1692,N_1033,N_1122);
nor U1693 (N_1693,N_1271,N_1180);
xnor U1694 (N_1694,N_1478,N_1003);
nor U1695 (N_1695,N_1400,N_1363);
or U1696 (N_1696,N_1081,N_1207);
and U1697 (N_1697,N_1184,N_1372);
nand U1698 (N_1698,N_1378,N_1359);
nor U1699 (N_1699,N_1057,N_1079);
and U1700 (N_1700,N_1097,N_1179);
nand U1701 (N_1701,N_1469,N_1234);
nor U1702 (N_1702,N_1153,N_1063);
nand U1703 (N_1703,N_1250,N_1062);
and U1704 (N_1704,N_1488,N_1214);
nor U1705 (N_1705,N_1360,N_1367);
nand U1706 (N_1706,N_1439,N_1313);
or U1707 (N_1707,N_1385,N_1215);
nand U1708 (N_1708,N_1287,N_1141);
and U1709 (N_1709,N_1127,N_1467);
nor U1710 (N_1710,N_1076,N_1251);
nand U1711 (N_1711,N_1065,N_1456);
and U1712 (N_1712,N_1101,N_1342);
or U1713 (N_1713,N_1344,N_1139);
and U1714 (N_1714,N_1244,N_1335);
nand U1715 (N_1715,N_1423,N_1034);
or U1716 (N_1716,N_1253,N_1489);
or U1717 (N_1717,N_1480,N_1049);
nand U1718 (N_1718,N_1458,N_1283);
nor U1719 (N_1719,N_1203,N_1365);
nand U1720 (N_1720,N_1061,N_1026);
nor U1721 (N_1721,N_1171,N_1420);
nand U1722 (N_1722,N_1190,N_1154);
nand U1723 (N_1723,N_1248,N_1406);
or U1724 (N_1724,N_1386,N_1472);
nand U1725 (N_1725,N_1273,N_1459);
and U1726 (N_1726,N_1268,N_1000);
and U1727 (N_1727,N_1009,N_1402);
nand U1728 (N_1728,N_1007,N_1475);
and U1729 (N_1729,N_1354,N_1346);
nor U1730 (N_1730,N_1410,N_1312);
and U1731 (N_1731,N_1164,N_1165);
nand U1732 (N_1732,N_1272,N_1328);
or U1733 (N_1733,N_1412,N_1046);
nor U1734 (N_1734,N_1468,N_1276);
nor U1735 (N_1735,N_1432,N_1394);
or U1736 (N_1736,N_1002,N_1466);
or U1737 (N_1737,N_1411,N_1109);
or U1738 (N_1738,N_1353,N_1193);
and U1739 (N_1739,N_1134,N_1013);
and U1740 (N_1740,N_1035,N_1318);
nor U1741 (N_1741,N_1191,N_1192);
or U1742 (N_1742,N_1465,N_1300);
or U1743 (N_1743,N_1249,N_1123);
nor U1744 (N_1744,N_1226,N_1118);
nor U1745 (N_1745,N_1144,N_1136);
and U1746 (N_1746,N_1103,N_1487);
nor U1747 (N_1747,N_1174,N_1306);
nor U1748 (N_1748,N_1493,N_1452);
or U1749 (N_1749,N_1220,N_1281);
or U1750 (N_1750,N_1432,N_1039);
xnor U1751 (N_1751,N_1291,N_1259);
nand U1752 (N_1752,N_1273,N_1145);
xor U1753 (N_1753,N_1451,N_1207);
and U1754 (N_1754,N_1381,N_1012);
nand U1755 (N_1755,N_1462,N_1481);
or U1756 (N_1756,N_1019,N_1465);
nor U1757 (N_1757,N_1387,N_1145);
xor U1758 (N_1758,N_1293,N_1032);
or U1759 (N_1759,N_1173,N_1038);
nor U1760 (N_1760,N_1032,N_1201);
and U1761 (N_1761,N_1021,N_1184);
or U1762 (N_1762,N_1335,N_1379);
nand U1763 (N_1763,N_1400,N_1351);
nor U1764 (N_1764,N_1285,N_1077);
or U1765 (N_1765,N_1019,N_1353);
or U1766 (N_1766,N_1000,N_1077);
nand U1767 (N_1767,N_1377,N_1394);
and U1768 (N_1768,N_1310,N_1253);
or U1769 (N_1769,N_1023,N_1355);
nand U1770 (N_1770,N_1365,N_1172);
or U1771 (N_1771,N_1362,N_1314);
or U1772 (N_1772,N_1068,N_1256);
nor U1773 (N_1773,N_1453,N_1187);
nand U1774 (N_1774,N_1150,N_1392);
xnor U1775 (N_1775,N_1094,N_1001);
or U1776 (N_1776,N_1460,N_1196);
nand U1777 (N_1777,N_1030,N_1457);
or U1778 (N_1778,N_1242,N_1313);
and U1779 (N_1779,N_1204,N_1438);
and U1780 (N_1780,N_1474,N_1089);
nand U1781 (N_1781,N_1442,N_1189);
nor U1782 (N_1782,N_1196,N_1321);
nand U1783 (N_1783,N_1306,N_1037);
nand U1784 (N_1784,N_1085,N_1058);
nor U1785 (N_1785,N_1180,N_1441);
nand U1786 (N_1786,N_1309,N_1419);
nor U1787 (N_1787,N_1447,N_1409);
and U1788 (N_1788,N_1186,N_1149);
xor U1789 (N_1789,N_1452,N_1201);
or U1790 (N_1790,N_1415,N_1367);
and U1791 (N_1791,N_1387,N_1457);
nor U1792 (N_1792,N_1115,N_1130);
nor U1793 (N_1793,N_1217,N_1219);
nand U1794 (N_1794,N_1153,N_1205);
nor U1795 (N_1795,N_1216,N_1090);
nor U1796 (N_1796,N_1145,N_1415);
nor U1797 (N_1797,N_1212,N_1231);
and U1798 (N_1798,N_1448,N_1453);
nor U1799 (N_1799,N_1480,N_1401);
xnor U1800 (N_1800,N_1062,N_1093);
nand U1801 (N_1801,N_1155,N_1429);
nor U1802 (N_1802,N_1205,N_1075);
and U1803 (N_1803,N_1260,N_1007);
or U1804 (N_1804,N_1029,N_1217);
nor U1805 (N_1805,N_1171,N_1388);
nand U1806 (N_1806,N_1104,N_1162);
nor U1807 (N_1807,N_1452,N_1272);
or U1808 (N_1808,N_1387,N_1006);
or U1809 (N_1809,N_1223,N_1042);
or U1810 (N_1810,N_1296,N_1244);
nor U1811 (N_1811,N_1214,N_1337);
nor U1812 (N_1812,N_1068,N_1361);
or U1813 (N_1813,N_1379,N_1084);
nor U1814 (N_1814,N_1245,N_1070);
or U1815 (N_1815,N_1003,N_1355);
nor U1816 (N_1816,N_1067,N_1159);
nand U1817 (N_1817,N_1103,N_1454);
nand U1818 (N_1818,N_1049,N_1246);
nor U1819 (N_1819,N_1018,N_1414);
nor U1820 (N_1820,N_1436,N_1439);
or U1821 (N_1821,N_1002,N_1402);
and U1822 (N_1822,N_1311,N_1277);
nand U1823 (N_1823,N_1163,N_1373);
or U1824 (N_1824,N_1448,N_1284);
nand U1825 (N_1825,N_1288,N_1021);
xor U1826 (N_1826,N_1399,N_1205);
nand U1827 (N_1827,N_1459,N_1105);
nand U1828 (N_1828,N_1240,N_1006);
xnor U1829 (N_1829,N_1441,N_1354);
nand U1830 (N_1830,N_1059,N_1330);
nand U1831 (N_1831,N_1349,N_1228);
xor U1832 (N_1832,N_1001,N_1403);
nand U1833 (N_1833,N_1078,N_1116);
or U1834 (N_1834,N_1189,N_1198);
xor U1835 (N_1835,N_1127,N_1063);
nand U1836 (N_1836,N_1135,N_1038);
nor U1837 (N_1837,N_1293,N_1347);
nand U1838 (N_1838,N_1009,N_1086);
and U1839 (N_1839,N_1331,N_1376);
or U1840 (N_1840,N_1411,N_1138);
nand U1841 (N_1841,N_1472,N_1011);
nand U1842 (N_1842,N_1448,N_1368);
and U1843 (N_1843,N_1369,N_1124);
and U1844 (N_1844,N_1065,N_1314);
nand U1845 (N_1845,N_1053,N_1109);
nand U1846 (N_1846,N_1184,N_1425);
or U1847 (N_1847,N_1312,N_1164);
or U1848 (N_1848,N_1453,N_1300);
or U1849 (N_1849,N_1238,N_1249);
nor U1850 (N_1850,N_1199,N_1079);
nor U1851 (N_1851,N_1072,N_1354);
nand U1852 (N_1852,N_1420,N_1377);
or U1853 (N_1853,N_1190,N_1257);
nor U1854 (N_1854,N_1066,N_1463);
or U1855 (N_1855,N_1345,N_1277);
nor U1856 (N_1856,N_1141,N_1447);
and U1857 (N_1857,N_1185,N_1092);
and U1858 (N_1858,N_1463,N_1376);
nor U1859 (N_1859,N_1493,N_1008);
or U1860 (N_1860,N_1326,N_1115);
nand U1861 (N_1861,N_1457,N_1361);
and U1862 (N_1862,N_1197,N_1142);
or U1863 (N_1863,N_1002,N_1029);
xnor U1864 (N_1864,N_1214,N_1087);
or U1865 (N_1865,N_1393,N_1060);
nand U1866 (N_1866,N_1131,N_1407);
nand U1867 (N_1867,N_1217,N_1026);
nor U1868 (N_1868,N_1192,N_1090);
or U1869 (N_1869,N_1401,N_1259);
and U1870 (N_1870,N_1111,N_1257);
or U1871 (N_1871,N_1467,N_1104);
nor U1872 (N_1872,N_1340,N_1248);
nor U1873 (N_1873,N_1379,N_1134);
or U1874 (N_1874,N_1028,N_1239);
and U1875 (N_1875,N_1404,N_1244);
and U1876 (N_1876,N_1022,N_1492);
xor U1877 (N_1877,N_1497,N_1474);
nor U1878 (N_1878,N_1489,N_1185);
nand U1879 (N_1879,N_1147,N_1209);
or U1880 (N_1880,N_1373,N_1496);
or U1881 (N_1881,N_1477,N_1014);
or U1882 (N_1882,N_1193,N_1343);
nand U1883 (N_1883,N_1280,N_1055);
nand U1884 (N_1884,N_1087,N_1464);
and U1885 (N_1885,N_1020,N_1112);
and U1886 (N_1886,N_1205,N_1106);
or U1887 (N_1887,N_1291,N_1470);
nor U1888 (N_1888,N_1116,N_1233);
or U1889 (N_1889,N_1214,N_1123);
nor U1890 (N_1890,N_1099,N_1212);
nand U1891 (N_1891,N_1020,N_1138);
and U1892 (N_1892,N_1251,N_1167);
or U1893 (N_1893,N_1421,N_1155);
or U1894 (N_1894,N_1253,N_1440);
nand U1895 (N_1895,N_1346,N_1095);
or U1896 (N_1896,N_1045,N_1157);
nand U1897 (N_1897,N_1146,N_1014);
nand U1898 (N_1898,N_1292,N_1388);
or U1899 (N_1899,N_1275,N_1431);
nor U1900 (N_1900,N_1067,N_1178);
nand U1901 (N_1901,N_1226,N_1402);
or U1902 (N_1902,N_1353,N_1159);
nor U1903 (N_1903,N_1219,N_1415);
nor U1904 (N_1904,N_1345,N_1162);
and U1905 (N_1905,N_1163,N_1498);
xor U1906 (N_1906,N_1318,N_1256);
nand U1907 (N_1907,N_1348,N_1444);
xnor U1908 (N_1908,N_1370,N_1137);
nor U1909 (N_1909,N_1312,N_1095);
nand U1910 (N_1910,N_1045,N_1173);
nand U1911 (N_1911,N_1233,N_1404);
and U1912 (N_1912,N_1095,N_1124);
and U1913 (N_1913,N_1442,N_1052);
nand U1914 (N_1914,N_1169,N_1165);
xnor U1915 (N_1915,N_1338,N_1270);
or U1916 (N_1916,N_1120,N_1480);
nor U1917 (N_1917,N_1021,N_1435);
nor U1918 (N_1918,N_1226,N_1104);
nand U1919 (N_1919,N_1297,N_1423);
and U1920 (N_1920,N_1368,N_1254);
or U1921 (N_1921,N_1331,N_1044);
nor U1922 (N_1922,N_1355,N_1147);
and U1923 (N_1923,N_1222,N_1266);
or U1924 (N_1924,N_1039,N_1128);
nor U1925 (N_1925,N_1436,N_1067);
nor U1926 (N_1926,N_1311,N_1057);
nand U1927 (N_1927,N_1072,N_1391);
or U1928 (N_1928,N_1297,N_1047);
or U1929 (N_1929,N_1313,N_1104);
or U1930 (N_1930,N_1017,N_1085);
nor U1931 (N_1931,N_1407,N_1305);
nand U1932 (N_1932,N_1183,N_1235);
and U1933 (N_1933,N_1392,N_1078);
and U1934 (N_1934,N_1233,N_1316);
and U1935 (N_1935,N_1150,N_1214);
or U1936 (N_1936,N_1475,N_1013);
nor U1937 (N_1937,N_1323,N_1079);
nor U1938 (N_1938,N_1428,N_1053);
nand U1939 (N_1939,N_1165,N_1321);
or U1940 (N_1940,N_1101,N_1090);
and U1941 (N_1941,N_1214,N_1460);
or U1942 (N_1942,N_1142,N_1261);
nand U1943 (N_1943,N_1442,N_1357);
or U1944 (N_1944,N_1447,N_1351);
nor U1945 (N_1945,N_1013,N_1116);
nand U1946 (N_1946,N_1326,N_1161);
or U1947 (N_1947,N_1156,N_1094);
nor U1948 (N_1948,N_1157,N_1461);
nor U1949 (N_1949,N_1484,N_1370);
nand U1950 (N_1950,N_1448,N_1066);
nand U1951 (N_1951,N_1429,N_1034);
or U1952 (N_1952,N_1368,N_1445);
xnor U1953 (N_1953,N_1188,N_1033);
or U1954 (N_1954,N_1353,N_1006);
and U1955 (N_1955,N_1052,N_1183);
nor U1956 (N_1956,N_1476,N_1189);
and U1957 (N_1957,N_1470,N_1209);
or U1958 (N_1958,N_1498,N_1124);
or U1959 (N_1959,N_1220,N_1350);
nand U1960 (N_1960,N_1498,N_1159);
nor U1961 (N_1961,N_1468,N_1425);
nor U1962 (N_1962,N_1255,N_1273);
xor U1963 (N_1963,N_1287,N_1128);
nor U1964 (N_1964,N_1433,N_1394);
nor U1965 (N_1965,N_1303,N_1367);
and U1966 (N_1966,N_1320,N_1086);
nor U1967 (N_1967,N_1404,N_1020);
nor U1968 (N_1968,N_1207,N_1073);
and U1969 (N_1969,N_1342,N_1477);
or U1970 (N_1970,N_1183,N_1344);
nor U1971 (N_1971,N_1444,N_1093);
xor U1972 (N_1972,N_1472,N_1465);
or U1973 (N_1973,N_1178,N_1140);
nand U1974 (N_1974,N_1061,N_1257);
or U1975 (N_1975,N_1179,N_1356);
or U1976 (N_1976,N_1265,N_1144);
and U1977 (N_1977,N_1469,N_1116);
and U1978 (N_1978,N_1364,N_1000);
or U1979 (N_1979,N_1301,N_1093);
or U1980 (N_1980,N_1181,N_1286);
nand U1981 (N_1981,N_1377,N_1250);
nor U1982 (N_1982,N_1151,N_1369);
nand U1983 (N_1983,N_1352,N_1093);
nor U1984 (N_1984,N_1009,N_1212);
and U1985 (N_1985,N_1254,N_1044);
nor U1986 (N_1986,N_1063,N_1008);
and U1987 (N_1987,N_1295,N_1255);
xnor U1988 (N_1988,N_1083,N_1207);
or U1989 (N_1989,N_1190,N_1059);
and U1990 (N_1990,N_1491,N_1046);
nor U1991 (N_1991,N_1017,N_1143);
xnor U1992 (N_1992,N_1201,N_1311);
and U1993 (N_1993,N_1238,N_1165);
and U1994 (N_1994,N_1011,N_1288);
or U1995 (N_1995,N_1356,N_1308);
and U1996 (N_1996,N_1217,N_1279);
and U1997 (N_1997,N_1098,N_1206);
nand U1998 (N_1998,N_1224,N_1205);
or U1999 (N_1999,N_1306,N_1409);
nor U2000 (N_2000,N_1971,N_1747);
nor U2001 (N_2001,N_1639,N_1546);
nand U2002 (N_2002,N_1663,N_1679);
nand U2003 (N_2003,N_1753,N_1505);
nand U2004 (N_2004,N_1963,N_1518);
or U2005 (N_2005,N_1784,N_1981);
nor U2006 (N_2006,N_1863,N_1590);
nand U2007 (N_2007,N_1579,N_1956);
or U2008 (N_2008,N_1597,N_1754);
nand U2009 (N_2009,N_1924,N_1884);
or U2010 (N_2010,N_1990,N_1900);
and U2011 (N_2011,N_1858,N_1929);
or U2012 (N_2012,N_1841,N_1680);
or U2013 (N_2013,N_1816,N_1714);
nand U2014 (N_2014,N_1643,N_1550);
nand U2015 (N_2015,N_1813,N_1585);
and U2016 (N_2016,N_1659,N_1996);
or U2017 (N_2017,N_1959,N_1684);
and U2018 (N_2018,N_1622,N_1601);
nor U2019 (N_2019,N_1961,N_1834);
nand U2020 (N_2020,N_1548,N_1756);
nand U2021 (N_2021,N_1811,N_1503);
and U2022 (N_2022,N_1611,N_1665);
nor U2023 (N_2023,N_1551,N_1874);
or U2024 (N_2024,N_1802,N_1575);
nor U2025 (N_2025,N_1570,N_1772);
nor U2026 (N_2026,N_1750,N_1689);
and U2027 (N_2027,N_1629,N_1693);
nor U2028 (N_2028,N_1952,N_1891);
or U2029 (N_2029,N_1835,N_1796);
or U2030 (N_2030,N_1846,N_1702);
nand U2031 (N_2031,N_1562,N_1602);
nand U2032 (N_2032,N_1778,N_1736);
or U2033 (N_2033,N_1882,N_1529);
nor U2034 (N_2034,N_1661,N_1587);
and U2035 (N_2035,N_1890,N_1708);
nand U2036 (N_2036,N_1692,N_1568);
nand U2037 (N_2037,N_1888,N_1901);
nand U2038 (N_2038,N_1892,N_1598);
or U2039 (N_2039,N_1742,N_1628);
nor U2040 (N_2040,N_1905,N_1848);
nand U2041 (N_2041,N_1873,N_1508);
nor U2042 (N_2042,N_1928,N_1715);
nand U2043 (N_2043,N_1589,N_1524);
nor U2044 (N_2044,N_1856,N_1818);
xnor U2045 (N_2045,N_1703,N_1648);
nand U2046 (N_2046,N_1849,N_1682);
nand U2047 (N_2047,N_1509,N_1902);
nor U2048 (N_2048,N_1539,N_1870);
nor U2049 (N_2049,N_1506,N_1886);
nand U2050 (N_2050,N_1515,N_1545);
nand U2051 (N_2051,N_1604,N_1623);
and U2052 (N_2052,N_1710,N_1526);
nor U2053 (N_2053,N_1867,N_1554);
nor U2054 (N_2054,N_1790,N_1542);
nor U2055 (N_2055,N_1957,N_1766);
nor U2056 (N_2056,N_1519,N_1711);
or U2057 (N_2057,N_1855,N_1584);
nor U2058 (N_2058,N_1748,N_1922);
or U2059 (N_2059,N_1713,N_1945);
or U2060 (N_2060,N_1982,N_1883);
or U2061 (N_2061,N_1919,N_1899);
nand U2062 (N_2062,N_1989,N_1953);
nor U2063 (N_2063,N_1740,N_1885);
nor U2064 (N_2064,N_1707,N_1752);
and U2065 (N_2065,N_1785,N_1534);
and U2066 (N_2066,N_1719,N_1552);
nor U2067 (N_2067,N_1718,N_1591);
nor U2068 (N_2068,N_1763,N_1838);
nand U2069 (N_2069,N_1522,N_1943);
nor U2070 (N_2070,N_1691,N_1560);
nor U2071 (N_2071,N_1572,N_1857);
nor U2072 (N_2072,N_1675,N_1864);
nor U2073 (N_2073,N_1843,N_1949);
and U2074 (N_2074,N_1781,N_1859);
and U2075 (N_2075,N_1898,N_1828);
and U2076 (N_2076,N_1523,N_1653);
or U2077 (N_2077,N_1946,N_1993);
or U2078 (N_2078,N_1700,N_1842);
and U2079 (N_2079,N_1836,N_1638);
and U2080 (N_2080,N_1851,N_1532);
or U2081 (N_2081,N_1581,N_1617);
nor U2082 (N_2082,N_1549,N_1869);
nor U2083 (N_2083,N_1516,N_1951);
or U2084 (N_2084,N_1765,N_1705);
or U2085 (N_2085,N_1862,N_1938);
or U2086 (N_2086,N_1616,N_1970);
and U2087 (N_2087,N_1757,N_1582);
nand U2088 (N_2088,N_1930,N_1944);
nor U2089 (N_2089,N_1773,N_1668);
nand U2090 (N_2090,N_1521,N_1916);
nor U2091 (N_2091,N_1879,N_1729);
nor U2092 (N_2092,N_1776,N_1725);
or U2093 (N_2093,N_1988,N_1803);
and U2094 (N_2094,N_1738,N_1676);
nand U2095 (N_2095,N_1914,N_1845);
or U2096 (N_2096,N_1935,N_1671);
or U2097 (N_2097,N_1656,N_1887);
and U2098 (N_2098,N_1793,N_1644);
and U2099 (N_2099,N_1866,N_1975);
and U2100 (N_2100,N_1543,N_1701);
nand U2101 (N_2101,N_1502,N_1730);
nand U2102 (N_2102,N_1674,N_1972);
or U2103 (N_2103,N_1646,N_1614);
and U2104 (N_2104,N_1619,N_1699);
or U2105 (N_2105,N_1755,N_1673);
nor U2106 (N_2106,N_1651,N_1758);
nand U2107 (N_2107,N_1973,N_1969);
and U2108 (N_2108,N_1564,N_1947);
or U2109 (N_2109,N_1939,N_1712);
or U2110 (N_2110,N_1829,N_1652);
nor U2111 (N_2111,N_1985,N_1995);
or U2112 (N_2112,N_1706,N_1530);
nand U2113 (N_2113,N_1909,N_1799);
and U2114 (N_2114,N_1775,N_1955);
nand U2115 (N_2115,N_1615,N_1868);
nor U2116 (N_2116,N_1797,N_1788);
or U2117 (N_2117,N_1717,N_1561);
and U2118 (N_2118,N_1832,N_1686);
nor U2119 (N_2119,N_1726,N_1932);
or U2120 (N_2120,N_1721,N_1809);
nand U2121 (N_2121,N_1595,N_1594);
nor U2122 (N_2122,N_1852,N_1931);
and U2123 (N_2123,N_1606,N_1583);
and U2124 (N_2124,N_1837,N_1517);
nand U2125 (N_2125,N_1540,N_1812);
nand U2126 (N_2126,N_1626,N_1620);
nand U2127 (N_2127,N_1724,N_1830);
nand U2128 (N_2128,N_1817,N_1940);
nor U2129 (N_2129,N_1920,N_1994);
nor U2130 (N_2130,N_1897,N_1926);
or U2131 (N_2131,N_1798,N_1685);
nor U2132 (N_2132,N_1915,N_1823);
nor U2133 (N_2133,N_1513,N_1681);
nand U2134 (N_2134,N_1672,N_1536);
nand U2135 (N_2135,N_1670,N_1563);
and U2136 (N_2136,N_1520,N_1768);
nor U2137 (N_2137,N_1556,N_1878);
nand U2138 (N_2138,N_1677,N_1553);
nand U2139 (N_2139,N_1635,N_1918);
nor U2140 (N_2140,N_1801,N_1815);
nor U2141 (N_2141,N_1744,N_1669);
and U2142 (N_2142,N_1732,N_1633);
or U2143 (N_2143,N_1625,N_1840);
and U2144 (N_2144,N_1877,N_1997);
nor U2145 (N_2145,N_1737,N_1965);
nor U2146 (N_2146,N_1998,N_1774);
xor U2147 (N_2147,N_1658,N_1824);
nor U2148 (N_2148,N_1647,N_1983);
and U2149 (N_2149,N_1903,N_1722);
nor U2150 (N_2150,N_1610,N_1704);
nand U2151 (N_2151,N_1966,N_1777);
and U2152 (N_2152,N_1865,N_1573);
nand U2153 (N_2153,N_1746,N_1807);
nand U2154 (N_2154,N_1787,N_1979);
nor U2155 (N_2155,N_1872,N_1537);
nand U2156 (N_2156,N_1531,N_1547);
nand U2157 (N_2157,N_1637,N_1667);
nand U2158 (N_2158,N_1745,N_1767);
and U2159 (N_2159,N_1504,N_1805);
and U2160 (N_2160,N_1645,N_1861);
nand U2161 (N_2161,N_1860,N_1723);
or U2162 (N_2162,N_1779,N_1806);
and U2163 (N_2163,N_1751,N_1688);
nand U2164 (N_2164,N_1850,N_1881);
nand U2165 (N_2165,N_1566,N_1749);
nand U2166 (N_2166,N_1716,N_1795);
and U2167 (N_2167,N_1720,N_1769);
and U2168 (N_2168,N_1618,N_1627);
or U2169 (N_2169,N_1895,N_1599);
and U2170 (N_2170,N_1839,N_1603);
or U2171 (N_2171,N_1569,N_1950);
and U2172 (N_2172,N_1600,N_1664);
and U2173 (N_2173,N_1780,N_1655);
nor U2174 (N_2174,N_1762,N_1967);
nand U2175 (N_2175,N_1789,N_1733);
or U2176 (N_2176,N_1612,N_1921);
and U2177 (N_2177,N_1650,N_1974);
nand U2178 (N_2178,N_1962,N_1854);
or U2179 (N_2179,N_1596,N_1609);
nand U2180 (N_2180,N_1694,N_1889);
nor U2181 (N_2181,N_1907,N_1820);
and U2182 (N_2182,N_1927,N_1605);
nor U2183 (N_2183,N_1913,N_1634);
and U2184 (N_2184,N_1786,N_1734);
nor U2185 (N_2185,N_1976,N_1586);
and U2186 (N_2186,N_1814,N_1608);
and U2187 (N_2187,N_1654,N_1535);
nand U2188 (N_2188,N_1968,N_1514);
or U2189 (N_2189,N_1528,N_1739);
and U2190 (N_2190,N_1741,N_1690);
or U2191 (N_2191,N_1678,N_1687);
nor U2192 (N_2192,N_1986,N_1574);
nor U2193 (N_2193,N_1941,N_1808);
nor U2194 (N_2194,N_1771,N_1984);
xnor U2195 (N_2195,N_1925,N_1743);
and U2196 (N_2196,N_1880,N_1875);
nand U2197 (N_2197,N_1933,N_1695);
and U2198 (N_2198,N_1791,N_1657);
nand U2199 (N_2199,N_1571,N_1770);
nand U2200 (N_2200,N_1511,N_1510);
nor U2201 (N_2201,N_1696,N_1666);
xor U2202 (N_2202,N_1592,N_1764);
nand U2203 (N_2203,N_1844,N_1735);
or U2204 (N_2204,N_1960,N_1992);
nand U2205 (N_2205,N_1821,N_1507);
or U2206 (N_2206,N_1588,N_1567);
and U2207 (N_2207,N_1565,N_1819);
and U2208 (N_2208,N_1825,N_1501);
or U2209 (N_2209,N_1662,N_1783);
nand U2210 (N_2210,N_1906,N_1593);
xor U2211 (N_2211,N_1810,N_1761);
nand U2212 (N_2212,N_1964,N_1728);
and U2213 (N_2213,N_1512,N_1912);
and U2214 (N_2214,N_1853,N_1613);
nor U2215 (N_2215,N_1937,N_1917);
nor U2216 (N_2216,N_1580,N_1630);
and U2217 (N_2217,N_1760,N_1893);
nor U2218 (N_2218,N_1904,N_1987);
nand U2219 (N_2219,N_1683,N_1936);
and U2220 (N_2220,N_1709,N_1800);
and U2221 (N_2221,N_1578,N_1557);
xor U2222 (N_2222,N_1804,N_1831);
or U2223 (N_2223,N_1636,N_1500);
nor U2224 (N_2224,N_1794,N_1576);
nor U2225 (N_2225,N_1991,N_1876);
or U2226 (N_2226,N_1980,N_1942);
and U2227 (N_2227,N_1731,N_1977);
or U2228 (N_2228,N_1541,N_1911);
and U2229 (N_2229,N_1822,N_1538);
and U2230 (N_2230,N_1631,N_1954);
nand U2231 (N_2231,N_1558,N_1827);
xnor U2232 (N_2232,N_1759,N_1559);
nand U2233 (N_2233,N_1833,N_1525);
and U2234 (N_2234,N_1782,N_1649);
nor U2235 (N_2235,N_1792,N_1894);
or U2236 (N_2236,N_1544,N_1641);
nor U2237 (N_2237,N_1621,N_1978);
or U2238 (N_2238,N_1642,N_1948);
and U2239 (N_2239,N_1934,N_1826);
nand U2240 (N_2240,N_1697,N_1896);
and U2241 (N_2241,N_1624,N_1958);
nand U2242 (N_2242,N_1527,N_1847);
nor U2243 (N_2243,N_1632,N_1698);
nand U2244 (N_2244,N_1640,N_1910);
and U2245 (N_2245,N_1871,N_1607);
nor U2246 (N_2246,N_1533,N_1923);
or U2247 (N_2247,N_1727,N_1555);
nor U2248 (N_2248,N_1908,N_1660);
nand U2249 (N_2249,N_1577,N_1999);
and U2250 (N_2250,N_1503,N_1922);
nor U2251 (N_2251,N_1893,N_1870);
and U2252 (N_2252,N_1660,N_1621);
or U2253 (N_2253,N_1816,N_1576);
nor U2254 (N_2254,N_1823,N_1989);
nor U2255 (N_2255,N_1800,N_1966);
nor U2256 (N_2256,N_1776,N_1893);
or U2257 (N_2257,N_1863,N_1827);
nor U2258 (N_2258,N_1713,N_1821);
and U2259 (N_2259,N_1697,N_1929);
xnor U2260 (N_2260,N_1559,N_1948);
or U2261 (N_2261,N_1892,N_1889);
or U2262 (N_2262,N_1858,N_1572);
and U2263 (N_2263,N_1508,N_1552);
or U2264 (N_2264,N_1552,N_1539);
nand U2265 (N_2265,N_1667,N_1547);
nand U2266 (N_2266,N_1631,N_1630);
and U2267 (N_2267,N_1602,N_1754);
nand U2268 (N_2268,N_1691,N_1694);
nand U2269 (N_2269,N_1774,N_1672);
xor U2270 (N_2270,N_1633,N_1684);
nand U2271 (N_2271,N_1588,N_1963);
nand U2272 (N_2272,N_1977,N_1743);
or U2273 (N_2273,N_1699,N_1782);
and U2274 (N_2274,N_1874,N_1678);
nand U2275 (N_2275,N_1508,N_1526);
nand U2276 (N_2276,N_1712,N_1723);
nand U2277 (N_2277,N_1874,N_1675);
and U2278 (N_2278,N_1761,N_1719);
and U2279 (N_2279,N_1657,N_1504);
and U2280 (N_2280,N_1530,N_1718);
or U2281 (N_2281,N_1923,N_1725);
nor U2282 (N_2282,N_1642,N_1576);
and U2283 (N_2283,N_1680,N_1729);
xnor U2284 (N_2284,N_1711,N_1951);
and U2285 (N_2285,N_1903,N_1509);
and U2286 (N_2286,N_1725,N_1893);
or U2287 (N_2287,N_1684,N_1950);
and U2288 (N_2288,N_1630,N_1649);
nand U2289 (N_2289,N_1571,N_1598);
nor U2290 (N_2290,N_1907,N_1802);
and U2291 (N_2291,N_1791,N_1827);
nand U2292 (N_2292,N_1868,N_1739);
and U2293 (N_2293,N_1576,N_1709);
nor U2294 (N_2294,N_1985,N_1931);
nand U2295 (N_2295,N_1567,N_1865);
and U2296 (N_2296,N_1816,N_1821);
or U2297 (N_2297,N_1905,N_1964);
or U2298 (N_2298,N_1682,N_1769);
nor U2299 (N_2299,N_1620,N_1716);
nand U2300 (N_2300,N_1763,N_1900);
or U2301 (N_2301,N_1890,N_1736);
nand U2302 (N_2302,N_1948,N_1850);
nand U2303 (N_2303,N_1622,N_1914);
or U2304 (N_2304,N_1525,N_1764);
xnor U2305 (N_2305,N_1766,N_1646);
nor U2306 (N_2306,N_1832,N_1544);
or U2307 (N_2307,N_1666,N_1678);
or U2308 (N_2308,N_1612,N_1667);
nand U2309 (N_2309,N_1956,N_1703);
nor U2310 (N_2310,N_1684,N_1906);
and U2311 (N_2311,N_1652,N_1625);
nand U2312 (N_2312,N_1582,N_1697);
and U2313 (N_2313,N_1760,N_1566);
and U2314 (N_2314,N_1777,N_1710);
nor U2315 (N_2315,N_1700,N_1854);
nand U2316 (N_2316,N_1862,N_1984);
and U2317 (N_2317,N_1584,N_1688);
and U2318 (N_2318,N_1939,N_1761);
nand U2319 (N_2319,N_1908,N_1658);
and U2320 (N_2320,N_1695,N_1634);
nor U2321 (N_2321,N_1566,N_1690);
and U2322 (N_2322,N_1631,N_1995);
nor U2323 (N_2323,N_1535,N_1536);
or U2324 (N_2324,N_1722,N_1671);
or U2325 (N_2325,N_1730,N_1970);
nand U2326 (N_2326,N_1532,N_1507);
nor U2327 (N_2327,N_1562,N_1913);
and U2328 (N_2328,N_1768,N_1815);
nand U2329 (N_2329,N_1919,N_1819);
nand U2330 (N_2330,N_1806,N_1932);
nor U2331 (N_2331,N_1638,N_1905);
and U2332 (N_2332,N_1607,N_1720);
nand U2333 (N_2333,N_1734,N_1620);
nand U2334 (N_2334,N_1643,N_1953);
and U2335 (N_2335,N_1567,N_1521);
xor U2336 (N_2336,N_1728,N_1616);
nand U2337 (N_2337,N_1797,N_1537);
and U2338 (N_2338,N_1721,N_1857);
and U2339 (N_2339,N_1870,N_1739);
nand U2340 (N_2340,N_1685,N_1721);
or U2341 (N_2341,N_1920,N_1782);
nor U2342 (N_2342,N_1803,N_1584);
nor U2343 (N_2343,N_1746,N_1769);
nor U2344 (N_2344,N_1952,N_1976);
nor U2345 (N_2345,N_1699,N_1503);
or U2346 (N_2346,N_1532,N_1538);
nor U2347 (N_2347,N_1514,N_1820);
and U2348 (N_2348,N_1707,N_1713);
nor U2349 (N_2349,N_1925,N_1868);
or U2350 (N_2350,N_1650,N_1748);
nor U2351 (N_2351,N_1808,N_1549);
nand U2352 (N_2352,N_1761,N_1911);
nand U2353 (N_2353,N_1534,N_1803);
or U2354 (N_2354,N_1578,N_1776);
nor U2355 (N_2355,N_1587,N_1761);
nor U2356 (N_2356,N_1848,N_1658);
or U2357 (N_2357,N_1864,N_1643);
nor U2358 (N_2358,N_1728,N_1540);
nor U2359 (N_2359,N_1647,N_1673);
nand U2360 (N_2360,N_1704,N_1908);
nand U2361 (N_2361,N_1620,N_1940);
xor U2362 (N_2362,N_1768,N_1983);
and U2363 (N_2363,N_1709,N_1637);
or U2364 (N_2364,N_1538,N_1613);
or U2365 (N_2365,N_1503,N_1510);
and U2366 (N_2366,N_1912,N_1706);
nand U2367 (N_2367,N_1929,N_1984);
and U2368 (N_2368,N_1895,N_1875);
and U2369 (N_2369,N_1601,N_1875);
nand U2370 (N_2370,N_1990,N_1875);
nand U2371 (N_2371,N_1678,N_1784);
nand U2372 (N_2372,N_1818,N_1993);
nor U2373 (N_2373,N_1868,N_1614);
nor U2374 (N_2374,N_1595,N_1883);
and U2375 (N_2375,N_1747,N_1636);
and U2376 (N_2376,N_1968,N_1954);
nand U2377 (N_2377,N_1815,N_1598);
xnor U2378 (N_2378,N_1990,N_1572);
xnor U2379 (N_2379,N_1616,N_1571);
and U2380 (N_2380,N_1820,N_1870);
and U2381 (N_2381,N_1956,N_1558);
nand U2382 (N_2382,N_1685,N_1728);
or U2383 (N_2383,N_1509,N_1975);
xor U2384 (N_2384,N_1845,N_1515);
nor U2385 (N_2385,N_1827,N_1689);
nand U2386 (N_2386,N_1523,N_1654);
xor U2387 (N_2387,N_1841,N_1646);
or U2388 (N_2388,N_1800,N_1870);
or U2389 (N_2389,N_1555,N_1783);
nor U2390 (N_2390,N_1650,N_1877);
and U2391 (N_2391,N_1948,N_1553);
or U2392 (N_2392,N_1725,N_1855);
nand U2393 (N_2393,N_1696,N_1745);
and U2394 (N_2394,N_1602,N_1879);
and U2395 (N_2395,N_1595,N_1778);
and U2396 (N_2396,N_1786,N_1627);
nand U2397 (N_2397,N_1609,N_1923);
xnor U2398 (N_2398,N_1625,N_1644);
nand U2399 (N_2399,N_1603,N_1661);
and U2400 (N_2400,N_1681,N_1769);
nor U2401 (N_2401,N_1904,N_1510);
or U2402 (N_2402,N_1573,N_1994);
nor U2403 (N_2403,N_1597,N_1811);
or U2404 (N_2404,N_1709,N_1729);
and U2405 (N_2405,N_1879,N_1712);
or U2406 (N_2406,N_1875,N_1897);
nand U2407 (N_2407,N_1656,N_1626);
and U2408 (N_2408,N_1506,N_1943);
nand U2409 (N_2409,N_1823,N_1640);
and U2410 (N_2410,N_1824,N_1728);
nand U2411 (N_2411,N_1622,N_1924);
and U2412 (N_2412,N_1984,N_1743);
nand U2413 (N_2413,N_1704,N_1514);
nor U2414 (N_2414,N_1608,N_1664);
nor U2415 (N_2415,N_1513,N_1774);
or U2416 (N_2416,N_1570,N_1751);
and U2417 (N_2417,N_1923,N_1634);
xor U2418 (N_2418,N_1933,N_1834);
and U2419 (N_2419,N_1856,N_1798);
and U2420 (N_2420,N_1889,N_1816);
nand U2421 (N_2421,N_1537,N_1870);
nor U2422 (N_2422,N_1615,N_1534);
nor U2423 (N_2423,N_1675,N_1892);
or U2424 (N_2424,N_1760,N_1661);
nand U2425 (N_2425,N_1750,N_1635);
and U2426 (N_2426,N_1676,N_1557);
or U2427 (N_2427,N_1591,N_1914);
or U2428 (N_2428,N_1962,N_1766);
nor U2429 (N_2429,N_1548,N_1696);
nand U2430 (N_2430,N_1916,N_1880);
nand U2431 (N_2431,N_1903,N_1993);
nand U2432 (N_2432,N_1693,N_1595);
xnor U2433 (N_2433,N_1909,N_1544);
and U2434 (N_2434,N_1582,N_1564);
or U2435 (N_2435,N_1605,N_1730);
or U2436 (N_2436,N_1672,N_1575);
nand U2437 (N_2437,N_1848,N_1602);
nand U2438 (N_2438,N_1950,N_1644);
nor U2439 (N_2439,N_1808,N_1924);
nand U2440 (N_2440,N_1711,N_1870);
nor U2441 (N_2441,N_1694,N_1586);
nor U2442 (N_2442,N_1676,N_1805);
or U2443 (N_2443,N_1815,N_1800);
and U2444 (N_2444,N_1917,N_1506);
nor U2445 (N_2445,N_1627,N_1522);
nor U2446 (N_2446,N_1652,N_1948);
nor U2447 (N_2447,N_1611,N_1802);
nand U2448 (N_2448,N_1526,N_1886);
nand U2449 (N_2449,N_1938,N_1808);
nor U2450 (N_2450,N_1553,N_1905);
or U2451 (N_2451,N_1766,N_1864);
and U2452 (N_2452,N_1656,N_1640);
nor U2453 (N_2453,N_1508,N_1688);
or U2454 (N_2454,N_1792,N_1596);
xor U2455 (N_2455,N_1643,N_1748);
nor U2456 (N_2456,N_1792,N_1640);
nor U2457 (N_2457,N_1646,N_1849);
nand U2458 (N_2458,N_1549,N_1502);
nor U2459 (N_2459,N_1554,N_1952);
or U2460 (N_2460,N_1831,N_1776);
and U2461 (N_2461,N_1502,N_1665);
and U2462 (N_2462,N_1777,N_1729);
nor U2463 (N_2463,N_1623,N_1705);
and U2464 (N_2464,N_1539,N_1697);
nand U2465 (N_2465,N_1870,N_1622);
and U2466 (N_2466,N_1692,N_1506);
nand U2467 (N_2467,N_1805,N_1932);
and U2468 (N_2468,N_1660,N_1750);
nor U2469 (N_2469,N_1582,N_1848);
nand U2470 (N_2470,N_1538,N_1634);
and U2471 (N_2471,N_1994,N_1786);
or U2472 (N_2472,N_1890,N_1960);
nor U2473 (N_2473,N_1502,N_1525);
and U2474 (N_2474,N_1886,N_1598);
nor U2475 (N_2475,N_1788,N_1611);
nand U2476 (N_2476,N_1535,N_1880);
and U2477 (N_2477,N_1596,N_1788);
nand U2478 (N_2478,N_1521,N_1655);
nor U2479 (N_2479,N_1894,N_1717);
nand U2480 (N_2480,N_1664,N_1516);
nor U2481 (N_2481,N_1522,N_1717);
nand U2482 (N_2482,N_1594,N_1523);
and U2483 (N_2483,N_1895,N_1801);
nor U2484 (N_2484,N_1862,N_1909);
nor U2485 (N_2485,N_1919,N_1854);
and U2486 (N_2486,N_1881,N_1956);
or U2487 (N_2487,N_1688,N_1998);
and U2488 (N_2488,N_1754,N_1616);
nor U2489 (N_2489,N_1734,N_1821);
nand U2490 (N_2490,N_1876,N_1986);
and U2491 (N_2491,N_1677,N_1842);
nor U2492 (N_2492,N_1514,N_1538);
and U2493 (N_2493,N_1948,N_1873);
nor U2494 (N_2494,N_1581,N_1953);
nor U2495 (N_2495,N_1776,N_1557);
and U2496 (N_2496,N_1917,N_1899);
xnor U2497 (N_2497,N_1700,N_1881);
nand U2498 (N_2498,N_1972,N_1976);
and U2499 (N_2499,N_1577,N_1854);
nor U2500 (N_2500,N_2103,N_2083);
xnor U2501 (N_2501,N_2479,N_2478);
or U2502 (N_2502,N_2014,N_2249);
xnor U2503 (N_2503,N_2127,N_2205);
or U2504 (N_2504,N_2402,N_2257);
nor U2505 (N_2505,N_2338,N_2178);
nor U2506 (N_2506,N_2405,N_2432);
nor U2507 (N_2507,N_2238,N_2355);
and U2508 (N_2508,N_2477,N_2277);
nand U2509 (N_2509,N_2363,N_2487);
or U2510 (N_2510,N_2379,N_2275);
or U2511 (N_2511,N_2396,N_2198);
or U2512 (N_2512,N_2326,N_2380);
and U2513 (N_2513,N_2137,N_2063);
or U2514 (N_2514,N_2320,N_2086);
and U2515 (N_2515,N_2241,N_2407);
and U2516 (N_2516,N_2029,N_2260);
nand U2517 (N_2517,N_2498,N_2066);
nand U2518 (N_2518,N_2124,N_2138);
or U2519 (N_2519,N_2291,N_2025);
or U2520 (N_2520,N_2077,N_2049);
or U2521 (N_2521,N_2195,N_2167);
nand U2522 (N_2522,N_2236,N_2343);
and U2523 (N_2523,N_2356,N_2162);
xor U2524 (N_2524,N_2362,N_2327);
or U2525 (N_2525,N_2449,N_2147);
xnor U2526 (N_2526,N_2372,N_2213);
and U2527 (N_2527,N_2068,N_2459);
and U2528 (N_2528,N_2388,N_2136);
nand U2529 (N_2529,N_2353,N_2149);
nor U2530 (N_2530,N_2280,N_2473);
and U2531 (N_2531,N_2112,N_2331);
and U2532 (N_2532,N_2001,N_2187);
nor U2533 (N_2533,N_2446,N_2134);
or U2534 (N_2534,N_2116,N_2090);
nor U2535 (N_2535,N_2299,N_2039);
nand U2536 (N_2536,N_2429,N_2357);
or U2537 (N_2537,N_2129,N_2024);
nor U2538 (N_2538,N_2110,N_2161);
or U2539 (N_2539,N_2219,N_2007);
nor U2540 (N_2540,N_2344,N_2413);
or U2541 (N_2541,N_2102,N_2227);
and U2542 (N_2542,N_2211,N_2093);
nand U2543 (N_2543,N_2259,N_2101);
and U2544 (N_2544,N_2398,N_2109);
or U2545 (N_2545,N_2113,N_2144);
nand U2546 (N_2546,N_2471,N_2223);
or U2547 (N_2547,N_2329,N_2239);
nor U2548 (N_2548,N_2425,N_2181);
nand U2549 (N_2549,N_2108,N_2071);
nand U2550 (N_2550,N_2294,N_2119);
or U2551 (N_2551,N_2180,N_2079);
nand U2552 (N_2552,N_2266,N_2319);
nor U2553 (N_2553,N_2295,N_2250);
nor U2554 (N_2554,N_2455,N_2315);
xnor U2555 (N_2555,N_2058,N_2106);
and U2556 (N_2556,N_2349,N_2378);
nor U2557 (N_2557,N_2439,N_2158);
nand U2558 (N_2558,N_2153,N_2284);
nor U2559 (N_2559,N_2465,N_2381);
and U2560 (N_2560,N_2050,N_2210);
nand U2561 (N_2561,N_2186,N_2423);
or U2562 (N_2562,N_2217,N_2006);
nor U2563 (N_2563,N_2251,N_2428);
nor U2564 (N_2564,N_2300,N_2476);
xor U2565 (N_2565,N_2323,N_2482);
and U2566 (N_2566,N_2496,N_2494);
or U2567 (N_2567,N_2033,N_2164);
nand U2568 (N_2568,N_2325,N_2027);
nand U2569 (N_2569,N_2472,N_2155);
nor U2570 (N_2570,N_2069,N_2202);
and U2571 (N_2571,N_2031,N_2092);
nand U2572 (N_2572,N_2267,N_2287);
and U2573 (N_2573,N_2206,N_2375);
nand U2574 (N_2574,N_2240,N_2096);
nor U2575 (N_2575,N_2281,N_2453);
nor U2576 (N_2576,N_2056,N_2261);
and U2577 (N_2577,N_2456,N_2305);
nor U2578 (N_2578,N_2021,N_2059);
and U2579 (N_2579,N_2133,N_2188);
nand U2580 (N_2580,N_2207,N_2171);
nor U2581 (N_2581,N_2190,N_2156);
nand U2582 (N_2582,N_2182,N_2491);
nor U2583 (N_2583,N_2070,N_2234);
and U2584 (N_2584,N_2414,N_2409);
or U2585 (N_2585,N_2034,N_2037);
nand U2586 (N_2586,N_2032,N_2154);
or U2587 (N_2587,N_2040,N_2159);
nand U2588 (N_2588,N_2192,N_2364);
and U2589 (N_2589,N_2023,N_2334);
nand U2590 (N_2590,N_2463,N_2309);
xnor U2591 (N_2591,N_2324,N_2216);
or U2592 (N_2592,N_2225,N_2082);
or U2593 (N_2593,N_2229,N_2076);
or U2594 (N_2594,N_2061,N_2497);
nand U2595 (N_2595,N_2157,N_2486);
nand U2596 (N_2596,N_2395,N_2072);
nand U2597 (N_2597,N_2427,N_2448);
and U2598 (N_2598,N_2107,N_2218);
nor U2599 (N_2599,N_2354,N_2399);
or U2600 (N_2600,N_2098,N_2437);
and U2601 (N_2601,N_2314,N_2183);
nand U2602 (N_2602,N_2495,N_2330);
nor U2603 (N_2603,N_2417,N_2328);
nor U2604 (N_2604,N_2146,N_2335);
or U2605 (N_2605,N_2013,N_2262);
nor U2606 (N_2606,N_2081,N_2151);
nor U2607 (N_2607,N_2390,N_2252);
nand U2608 (N_2608,N_2336,N_2018);
or U2609 (N_2609,N_2470,N_2150);
nand U2610 (N_2610,N_2253,N_2304);
nand U2611 (N_2611,N_2469,N_2360);
nand U2612 (N_2612,N_2318,N_2274);
and U2613 (N_2613,N_2481,N_2060);
or U2614 (N_2614,N_2002,N_2493);
nor U2615 (N_2615,N_2163,N_2369);
nor U2616 (N_2616,N_2004,N_2135);
or U2617 (N_2617,N_2194,N_2283);
nand U2618 (N_2618,N_2115,N_2139);
and U2619 (N_2619,N_2176,N_2172);
xnor U2620 (N_2620,N_2140,N_2293);
nor U2621 (N_2621,N_2298,N_2411);
xnor U2622 (N_2622,N_2288,N_2272);
or U2623 (N_2623,N_2036,N_2204);
nor U2624 (N_2624,N_2475,N_2265);
nor U2625 (N_2625,N_2244,N_2200);
and U2626 (N_2626,N_2333,N_2447);
and U2627 (N_2627,N_2384,N_2087);
or U2628 (N_2628,N_2278,N_2243);
or U2629 (N_2629,N_2292,N_2185);
nand U2630 (N_2630,N_2394,N_2410);
or U2631 (N_2631,N_2008,N_2175);
nor U2632 (N_2632,N_2285,N_2412);
or U2633 (N_2633,N_2038,N_2080);
nor U2634 (N_2634,N_2422,N_2317);
or U2635 (N_2635,N_2121,N_2351);
nor U2636 (N_2636,N_2128,N_2208);
nor U2637 (N_2637,N_2230,N_2464);
or U2638 (N_2638,N_2342,N_2114);
nor U2639 (N_2639,N_2053,N_2169);
nand U2640 (N_2640,N_2166,N_2254);
nor U2641 (N_2641,N_2094,N_2370);
nor U2642 (N_2642,N_2256,N_2452);
nand U2643 (N_2643,N_2196,N_2145);
nand U2644 (N_2644,N_2377,N_2421);
and U2645 (N_2645,N_2088,N_2026);
nand U2646 (N_2646,N_2431,N_2074);
or U2647 (N_2647,N_2242,N_2052);
nand U2648 (N_2648,N_2221,N_2485);
and U2649 (N_2649,N_2480,N_2345);
nor U2650 (N_2650,N_2468,N_2433);
and U2651 (N_2651,N_2445,N_2359);
and U2652 (N_2652,N_2451,N_2048);
and U2653 (N_2653,N_2035,N_2458);
nor U2654 (N_2654,N_2130,N_2201);
or U2655 (N_2655,N_2095,N_2228);
or U2656 (N_2656,N_2235,N_2313);
and U2657 (N_2657,N_2415,N_2308);
and U2658 (N_2658,N_2075,N_2264);
nor U2659 (N_2659,N_2184,N_2368);
and U2660 (N_2660,N_2019,N_2332);
or U2661 (N_2661,N_2111,N_2212);
and U2662 (N_2662,N_2030,N_2022);
and U2663 (N_2663,N_2215,N_2043);
nor U2664 (N_2664,N_2419,N_2142);
nor U2665 (N_2665,N_2011,N_2105);
and U2666 (N_2666,N_2177,N_2269);
or U2667 (N_2667,N_2416,N_2276);
or U2668 (N_2668,N_2322,N_2404);
nor U2669 (N_2669,N_2191,N_2165);
nand U2670 (N_2670,N_2499,N_2400);
and U2671 (N_2671,N_2347,N_2091);
nand U2672 (N_2672,N_2462,N_2016);
or U2673 (N_2673,N_2255,N_2125);
or U2674 (N_2674,N_2461,N_2492);
or U2675 (N_2675,N_2012,N_2382);
nand U2676 (N_2676,N_2055,N_2339);
or U2677 (N_2677,N_2420,N_2141);
nor U2678 (N_2678,N_2220,N_2312);
nand U2679 (N_2679,N_2391,N_2279);
and U2680 (N_2680,N_2385,N_2454);
or U2681 (N_2681,N_2442,N_2245);
nand U2682 (N_2682,N_2376,N_2065);
nand U2683 (N_2683,N_2387,N_2393);
nand U2684 (N_2684,N_2231,N_2436);
or U2685 (N_2685,N_2078,N_2403);
or U2686 (N_2686,N_2440,N_2297);
or U2687 (N_2687,N_2148,N_2406);
and U2688 (N_2688,N_2131,N_2289);
and U2689 (N_2689,N_2099,N_2044);
or U2690 (N_2690,N_2341,N_2020);
nor U2691 (N_2691,N_2232,N_2003);
nor U2692 (N_2692,N_2466,N_2017);
and U2693 (N_2693,N_2046,N_2100);
or U2694 (N_2694,N_2435,N_2045);
or U2695 (N_2695,N_2348,N_2000);
nand U2696 (N_2696,N_2270,N_2047);
and U2697 (N_2697,N_2246,N_2430);
nor U2698 (N_2698,N_2042,N_2361);
and U2699 (N_2699,N_2089,N_2358);
or U2700 (N_2700,N_2397,N_2434);
nand U2701 (N_2701,N_2340,N_2054);
nor U2702 (N_2702,N_2474,N_2160);
nand U2703 (N_2703,N_2005,N_2271);
nand U2704 (N_2704,N_2209,N_2365);
nor U2705 (N_2705,N_2441,N_2389);
or U2706 (N_2706,N_2189,N_2123);
or U2707 (N_2707,N_2484,N_2041);
and U2708 (N_2708,N_2010,N_2450);
nor U2709 (N_2709,N_2302,N_2179);
or U2710 (N_2710,N_2371,N_2489);
and U2711 (N_2711,N_2321,N_2418);
xnor U2712 (N_2712,N_2122,N_2226);
and U2713 (N_2713,N_2401,N_2303);
nor U2714 (N_2714,N_2120,N_2483);
and U2715 (N_2715,N_2132,N_2366);
xor U2716 (N_2716,N_2214,N_2367);
nand U2717 (N_2717,N_2237,N_2170);
xnor U2718 (N_2718,N_2490,N_2273);
xnor U2719 (N_2719,N_2064,N_2443);
nand U2720 (N_2720,N_2290,N_2222);
nand U2721 (N_2721,N_2203,N_2350);
xor U2722 (N_2722,N_2386,N_2311);
nand U2723 (N_2723,N_2152,N_2424);
and U2724 (N_2724,N_2197,N_2009);
and U2725 (N_2725,N_2248,N_2457);
nor U2726 (N_2726,N_2373,N_2352);
and U2727 (N_2727,N_2168,N_2392);
nor U2728 (N_2728,N_2438,N_2301);
or U2729 (N_2729,N_2199,N_2028);
nand U2730 (N_2730,N_2118,N_2282);
and U2731 (N_2731,N_2460,N_2085);
nand U2732 (N_2732,N_2258,N_2346);
or U2733 (N_2733,N_2488,N_2307);
nand U2734 (N_2734,N_2104,N_2073);
or U2735 (N_2735,N_2233,N_2084);
nor U2736 (N_2736,N_2143,N_2173);
or U2737 (N_2737,N_2374,N_2296);
or U2738 (N_2738,N_2015,N_2057);
and U2739 (N_2739,N_2426,N_2263);
nor U2740 (N_2740,N_2408,N_2051);
or U2741 (N_2741,N_2383,N_2117);
nand U2742 (N_2742,N_2286,N_2310);
nor U2743 (N_2743,N_2067,N_2247);
or U2744 (N_2744,N_2268,N_2306);
nor U2745 (N_2745,N_2467,N_2193);
and U2746 (N_2746,N_2097,N_2224);
nor U2747 (N_2747,N_2126,N_2316);
nand U2748 (N_2748,N_2337,N_2174);
nor U2749 (N_2749,N_2062,N_2444);
nor U2750 (N_2750,N_2008,N_2308);
nor U2751 (N_2751,N_2284,N_2358);
or U2752 (N_2752,N_2399,N_2302);
or U2753 (N_2753,N_2229,N_2149);
and U2754 (N_2754,N_2283,N_2430);
and U2755 (N_2755,N_2166,N_2414);
nand U2756 (N_2756,N_2013,N_2061);
nand U2757 (N_2757,N_2025,N_2218);
and U2758 (N_2758,N_2292,N_2316);
or U2759 (N_2759,N_2483,N_2496);
and U2760 (N_2760,N_2225,N_2274);
xnor U2761 (N_2761,N_2359,N_2181);
nand U2762 (N_2762,N_2207,N_2394);
nand U2763 (N_2763,N_2085,N_2070);
nand U2764 (N_2764,N_2445,N_2471);
and U2765 (N_2765,N_2257,N_2114);
or U2766 (N_2766,N_2116,N_2305);
and U2767 (N_2767,N_2376,N_2039);
and U2768 (N_2768,N_2453,N_2228);
nand U2769 (N_2769,N_2414,N_2235);
and U2770 (N_2770,N_2221,N_2045);
and U2771 (N_2771,N_2129,N_2089);
nand U2772 (N_2772,N_2343,N_2316);
or U2773 (N_2773,N_2250,N_2336);
nand U2774 (N_2774,N_2292,N_2194);
nor U2775 (N_2775,N_2400,N_2066);
or U2776 (N_2776,N_2122,N_2159);
or U2777 (N_2777,N_2011,N_2213);
and U2778 (N_2778,N_2252,N_2345);
nand U2779 (N_2779,N_2025,N_2040);
and U2780 (N_2780,N_2162,N_2131);
and U2781 (N_2781,N_2308,N_2217);
and U2782 (N_2782,N_2373,N_2071);
nor U2783 (N_2783,N_2179,N_2136);
nand U2784 (N_2784,N_2471,N_2437);
and U2785 (N_2785,N_2222,N_2100);
and U2786 (N_2786,N_2404,N_2214);
and U2787 (N_2787,N_2267,N_2459);
nand U2788 (N_2788,N_2078,N_2307);
nor U2789 (N_2789,N_2175,N_2480);
nand U2790 (N_2790,N_2233,N_2135);
and U2791 (N_2791,N_2068,N_2339);
nand U2792 (N_2792,N_2110,N_2277);
nand U2793 (N_2793,N_2378,N_2148);
nor U2794 (N_2794,N_2272,N_2179);
and U2795 (N_2795,N_2217,N_2068);
xnor U2796 (N_2796,N_2020,N_2188);
nand U2797 (N_2797,N_2017,N_2069);
or U2798 (N_2798,N_2203,N_2345);
nand U2799 (N_2799,N_2271,N_2291);
and U2800 (N_2800,N_2399,N_2069);
nand U2801 (N_2801,N_2054,N_2399);
nand U2802 (N_2802,N_2080,N_2458);
and U2803 (N_2803,N_2263,N_2306);
nor U2804 (N_2804,N_2455,N_2323);
nand U2805 (N_2805,N_2025,N_2176);
or U2806 (N_2806,N_2167,N_2423);
or U2807 (N_2807,N_2119,N_2029);
nand U2808 (N_2808,N_2321,N_2103);
xor U2809 (N_2809,N_2067,N_2488);
nand U2810 (N_2810,N_2047,N_2115);
nor U2811 (N_2811,N_2417,N_2307);
nand U2812 (N_2812,N_2344,N_2244);
nor U2813 (N_2813,N_2143,N_2099);
and U2814 (N_2814,N_2153,N_2003);
or U2815 (N_2815,N_2178,N_2295);
nor U2816 (N_2816,N_2243,N_2454);
or U2817 (N_2817,N_2458,N_2189);
nand U2818 (N_2818,N_2180,N_2011);
or U2819 (N_2819,N_2287,N_2194);
or U2820 (N_2820,N_2344,N_2411);
nand U2821 (N_2821,N_2359,N_2104);
and U2822 (N_2822,N_2476,N_2101);
and U2823 (N_2823,N_2437,N_2449);
and U2824 (N_2824,N_2148,N_2264);
nand U2825 (N_2825,N_2312,N_2392);
nor U2826 (N_2826,N_2462,N_2231);
nor U2827 (N_2827,N_2390,N_2177);
or U2828 (N_2828,N_2065,N_2338);
and U2829 (N_2829,N_2439,N_2354);
and U2830 (N_2830,N_2405,N_2167);
and U2831 (N_2831,N_2391,N_2406);
and U2832 (N_2832,N_2155,N_2082);
nand U2833 (N_2833,N_2084,N_2268);
and U2834 (N_2834,N_2200,N_2463);
and U2835 (N_2835,N_2486,N_2452);
and U2836 (N_2836,N_2299,N_2191);
xnor U2837 (N_2837,N_2481,N_2032);
xnor U2838 (N_2838,N_2004,N_2182);
nor U2839 (N_2839,N_2200,N_2214);
and U2840 (N_2840,N_2392,N_2095);
and U2841 (N_2841,N_2319,N_2392);
xor U2842 (N_2842,N_2485,N_2309);
nor U2843 (N_2843,N_2433,N_2342);
and U2844 (N_2844,N_2164,N_2438);
or U2845 (N_2845,N_2327,N_2037);
nand U2846 (N_2846,N_2017,N_2001);
and U2847 (N_2847,N_2192,N_2379);
and U2848 (N_2848,N_2219,N_2402);
xnor U2849 (N_2849,N_2219,N_2063);
xnor U2850 (N_2850,N_2336,N_2069);
and U2851 (N_2851,N_2332,N_2147);
and U2852 (N_2852,N_2375,N_2396);
nor U2853 (N_2853,N_2195,N_2299);
and U2854 (N_2854,N_2493,N_2157);
and U2855 (N_2855,N_2072,N_2083);
nor U2856 (N_2856,N_2008,N_2218);
or U2857 (N_2857,N_2367,N_2449);
nand U2858 (N_2858,N_2180,N_2056);
nor U2859 (N_2859,N_2436,N_2285);
nor U2860 (N_2860,N_2090,N_2301);
nand U2861 (N_2861,N_2285,N_2201);
nand U2862 (N_2862,N_2400,N_2413);
nand U2863 (N_2863,N_2145,N_2340);
nor U2864 (N_2864,N_2347,N_2399);
nand U2865 (N_2865,N_2284,N_2470);
or U2866 (N_2866,N_2033,N_2126);
and U2867 (N_2867,N_2399,N_2165);
or U2868 (N_2868,N_2403,N_2000);
nand U2869 (N_2869,N_2032,N_2422);
or U2870 (N_2870,N_2322,N_2141);
and U2871 (N_2871,N_2276,N_2351);
nor U2872 (N_2872,N_2318,N_2401);
nand U2873 (N_2873,N_2103,N_2098);
xor U2874 (N_2874,N_2408,N_2483);
and U2875 (N_2875,N_2128,N_2407);
nor U2876 (N_2876,N_2284,N_2150);
or U2877 (N_2877,N_2206,N_2359);
or U2878 (N_2878,N_2362,N_2401);
or U2879 (N_2879,N_2176,N_2274);
or U2880 (N_2880,N_2315,N_2256);
nor U2881 (N_2881,N_2462,N_2050);
nor U2882 (N_2882,N_2030,N_2297);
and U2883 (N_2883,N_2420,N_2431);
and U2884 (N_2884,N_2451,N_2340);
and U2885 (N_2885,N_2472,N_2381);
nand U2886 (N_2886,N_2150,N_2133);
nor U2887 (N_2887,N_2458,N_2115);
nor U2888 (N_2888,N_2081,N_2428);
xnor U2889 (N_2889,N_2152,N_2167);
or U2890 (N_2890,N_2337,N_2021);
nor U2891 (N_2891,N_2050,N_2426);
nand U2892 (N_2892,N_2361,N_2144);
nor U2893 (N_2893,N_2332,N_2178);
and U2894 (N_2894,N_2150,N_2229);
and U2895 (N_2895,N_2405,N_2336);
nor U2896 (N_2896,N_2413,N_2236);
and U2897 (N_2897,N_2351,N_2268);
nor U2898 (N_2898,N_2215,N_2462);
nor U2899 (N_2899,N_2258,N_2155);
nand U2900 (N_2900,N_2257,N_2318);
nor U2901 (N_2901,N_2163,N_2469);
and U2902 (N_2902,N_2459,N_2318);
nor U2903 (N_2903,N_2295,N_2362);
or U2904 (N_2904,N_2257,N_2352);
nor U2905 (N_2905,N_2386,N_2490);
or U2906 (N_2906,N_2310,N_2213);
and U2907 (N_2907,N_2204,N_2075);
nor U2908 (N_2908,N_2250,N_2107);
nand U2909 (N_2909,N_2114,N_2458);
nand U2910 (N_2910,N_2206,N_2384);
nand U2911 (N_2911,N_2168,N_2367);
nor U2912 (N_2912,N_2225,N_2318);
nand U2913 (N_2913,N_2000,N_2484);
and U2914 (N_2914,N_2444,N_2498);
or U2915 (N_2915,N_2348,N_2365);
nor U2916 (N_2916,N_2236,N_2209);
and U2917 (N_2917,N_2348,N_2292);
nand U2918 (N_2918,N_2441,N_2211);
and U2919 (N_2919,N_2042,N_2117);
or U2920 (N_2920,N_2434,N_2419);
nand U2921 (N_2921,N_2435,N_2159);
or U2922 (N_2922,N_2457,N_2012);
nor U2923 (N_2923,N_2415,N_2108);
nand U2924 (N_2924,N_2151,N_2003);
nand U2925 (N_2925,N_2362,N_2420);
or U2926 (N_2926,N_2212,N_2206);
nor U2927 (N_2927,N_2025,N_2399);
or U2928 (N_2928,N_2303,N_2293);
and U2929 (N_2929,N_2433,N_2398);
nor U2930 (N_2930,N_2164,N_2409);
and U2931 (N_2931,N_2496,N_2333);
nand U2932 (N_2932,N_2103,N_2024);
or U2933 (N_2933,N_2295,N_2284);
or U2934 (N_2934,N_2127,N_2152);
and U2935 (N_2935,N_2125,N_2353);
or U2936 (N_2936,N_2314,N_2001);
and U2937 (N_2937,N_2059,N_2101);
or U2938 (N_2938,N_2497,N_2314);
and U2939 (N_2939,N_2254,N_2426);
nand U2940 (N_2940,N_2472,N_2150);
nor U2941 (N_2941,N_2272,N_2400);
nand U2942 (N_2942,N_2107,N_2359);
nor U2943 (N_2943,N_2292,N_2289);
nor U2944 (N_2944,N_2449,N_2331);
nor U2945 (N_2945,N_2026,N_2460);
and U2946 (N_2946,N_2197,N_2497);
nand U2947 (N_2947,N_2482,N_2446);
or U2948 (N_2948,N_2281,N_2164);
nor U2949 (N_2949,N_2037,N_2105);
and U2950 (N_2950,N_2439,N_2212);
nand U2951 (N_2951,N_2443,N_2320);
or U2952 (N_2952,N_2061,N_2005);
and U2953 (N_2953,N_2264,N_2073);
or U2954 (N_2954,N_2206,N_2302);
and U2955 (N_2955,N_2285,N_2075);
or U2956 (N_2956,N_2364,N_2009);
or U2957 (N_2957,N_2312,N_2230);
and U2958 (N_2958,N_2458,N_2338);
nand U2959 (N_2959,N_2451,N_2240);
nor U2960 (N_2960,N_2311,N_2227);
nand U2961 (N_2961,N_2410,N_2311);
and U2962 (N_2962,N_2480,N_2126);
nor U2963 (N_2963,N_2008,N_2345);
and U2964 (N_2964,N_2424,N_2321);
xnor U2965 (N_2965,N_2471,N_2059);
nor U2966 (N_2966,N_2373,N_2476);
nand U2967 (N_2967,N_2293,N_2168);
nor U2968 (N_2968,N_2257,N_2411);
or U2969 (N_2969,N_2110,N_2321);
or U2970 (N_2970,N_2088,N_2322);
or U2971 (N_2971,N_2451,N_2165);
or U2972 (N_2972,N_2057,N_2005);
or U2973 (N_2973,N_2286,N_2002);
nor U2974 (N_2974,N_2054,N_2212);
nand U2975 (N_2975,N_2206,N_2298);
nand U2976 (N_2976,N_2097,N_2418);
nor U2977 (N_2977,N_2033,N_2399);
nor U2978 (N_2978,N_2092,N_2104);
and U2979 (N_2979,N_2263,N_2354);
or U2980 (N_2980,N_2109,N_2040);
nor U2981 (N_2981,N_2401,N_2041);
nand U2982 (N_2982,N_2483,N_2435);
nor U2983 (N_2983,N_2431,N_2253);
or U2984 (N_2984,N_2144,N_2183);
nand U2985 (N_2985,N_2353,N_2252);
nor U2986 (N_2986,N_2190,N_2493);
xnor U2987 (N_2987,N_2209,N_2206);
and U2988 (N_2988,N_2189,N_2025);
or U2989 (N_2989,N_2038,N_2329);
nand U2990 (N_2990,N_2323,N_2261);
nor U2991 (N_2991,N_2330,N_2430);
and U2992 (N_2992,N_2202,N_2429);
or U2993 (N_2993,N_2487,N_2284);
or U2994 (N_2994,N_2357,N_2077);
nand U2995 (N_2995,N_2371,N_2223);
nand U2996 (N_2996,N_2389,N_2329);
and U2997 (N_2997,N_2240,N_2275);
and U2998 (N_2998,N_2106,N_2097);
nand U2999 (N_2999,N_2152,N_2081);
nand U3000 (N_3000,N_2790,N_2656);
nand U3001 (N_3001,N_2984,N_2542);
nor U3002 (N_3002,N_2761,N_2543);
and U3003 (N_3003,N_2769,N_2808);
or U3004 (N_3004,N_2986,N_2563);
nand U3005 (N_3005,N_2521,N_2886);
or U3006 (N_3006,N_2929,N_2576);
nand U3007 (N_3007,N_2503,N_2983);
and U3008 (N_3008,N_2988,N_2575);
nand U3009 (N_3009,N_2847,N_2533);
and U3010 (N_3010,N_2978,N_2574);
or U3011 (N_3011,N_2914,N_2906);
nand U3012 (N_3012,N_2952,N_2505);
nand U3013 (N_3013,N_2958,N_2806);
nand U3014 (N_3014,N_2719,N_2512);
and U3015 (N_3015,N_2705,N_2820);
or U3016 (N_3016,N_2697,N_2941);
and U3017 (N_3017,N_2608,N_2579);
or U3018 (N_3018,N_2541,N_2682);
nor U3019 (N_3019,N_2582,N_2909);
nand U3020 (N_3020,N_2686,N_2736);
and U3021 (N_3021,N_2974,N_2931);
and U3022 (N_3022,N_2973,N_2710);
and U3023 (N_3023,N_2902,N_2774);
nand U3024 (N_3024,N_2823,N_2896);
nand U3025 (N_3025,N_2751,N_2725);
and U3026 (N_3026,N_2753,N_2711);
or U3027 (N_3027,N_2803,N_2894);
and U3028 (N_3028,N_2900,N_2739);
and U3029 (N_3029,N_2773,N_2922);
or U3030 (N_3030,N_2530,N_2712);
nand U3031 (N_3031,N_2923,N_2917);
nand U3032 (N_3032,N_2972,N_2737);
nand U3033 (N_3033,N_2675,N_2891);
and U3034 (N_3034,N_2805,N_2507);
or U3035 (N_3035,N_2870,N_2634);
and U3036 (N_3036,N_2968,N_2564);
or U3037 (N_3037,N_2932,N_2584);
and U3038 (N_3038,N_2910,N_2752);
nor U3039 (N_3039,N_2933,N_2573);
and U3040 (N_3040,N_2846,N_2556);
or U3041 (N_3041,N_2545,N_2966);
nand U3042 (N_3042,N_2963,N_2943);
and U3043 (N_3043,N_2755,N_2690);
and U3044 (N_3044,N_2625,N_2523);
and U3045 (N_3045,N_2946,N_2904);
or U3046 (N_3046,N_2525,N_2801);
nand U3047 (N_3047,N_2536,N_2691);
nand U3048 (N_3048,N_2758,N_2514);
and U3049 (N_3049,N_2621,N_2982);
nor U3050 (N_3050,N_2819,N_2813);
nor U3051 (N_3051,N_2568,N_2701);
nand U3052 (N_3052,N_2727,N_2729);
and U3053 (N_3053,N_2700,N_2674);
xnor U3054 (N_3054,N_2793,N_2889);
or U3055 (N_3055,N_2558,N_2760);
or U3056 (N_3056,N_2692,N_2854);
nand U3057 (N_3057,N_2708,N_2681);
and U3058 (N_3058,N_2626,N_2669);
or U3059 (N_3059,N_2785,N_2672);
and U3060 (N_3060,N_2955,N_2893);
or U3061 (N_3061,N_2744,N_2586);
and U3062 (N_3062,N_2880,N_2853);
nor U3063 (N_3063,N_2513,N_2577);
and U3064 (N_3064,N_2726,N_2651);
xor U3065 (N_3065,N_2509,N_2835);
xnor U3066 (N_3066,N_2949,N_2531);
nor U3067 (N_3067,N_2925,N_2845);
nor U3068 (N_3068,N_2501,N_2567);
nor U3069 (N_3069,N_2856,N_2927);
nand U3070 (N_3070,N_2954,N_2799);
nor U3071 (N_3071,N_2762,N_2520);
nand U3072 (N_3072,N_2680,N_2809);
or U3073 (N_3073,N_2770,N_2524);
and U3074 (N_3074,N_2864,N_2571);
and U3075 (N_3075,N_2779,N_2868);
xnor U3076 (N_3076,N_2640,N_2679);
or U3077 (N_3077,N_2637,N_2662);
and U3078 (N_3078,N_2605,N_2839);
and U3079 (N_3079,N_2783,N_2713);
nor U3080 (N_3080,N_2738,N_2863);
and U3081 (N_3081,N_2628,N_2555);
nor U3082 (N_3082,N_2825,N_2549);
or U3083 (N_3083,N_2882,N_2976);
and U3084 (N_3084,N_2585,N_2551);
nor U3085 (N_3085,N_2554,N_2862);
nor U3086 (N_3086,N_2926,N_2791);
nor U3087 (N_3087,N_2877,N_2604);
nor U3088 (N_3088,N_2598,N_2782);
nand U3089 (N_3089,N_2648,N_2993);
nor U3090 (N_3090,N_2590,N_2668);
and U3091 (N_3091,N_2630,N_2559);
or U3092 (N_3092,N_2694,N_2595);
nor U3093 (N_3093,N_2935,N_2616);
nand U3094 (N_3094,N_2750,N_2560);
nand U3095 (N_3095,N_2996,N_2588);
nand U3096 (N_3096,N_2607,N_2735);
nand U3097 (N_3097,N_2995,N_2898);
nand U3098 (N_3098,N_2504,N_2873);
nor U3099 (N_3099,N_2600,N_2592);
and U3100 (N_3100,N_2642,N_2627);
or U3101 (N_3101,N_2544,N_2714);
or U3102 (N_3102,N_2540,N_2765);
or U3103 (N_3103,N_2756,N_2947);
nor U3104 (N_3104,N_2665,N_2824);
or U3105 (N_3105,N_2731,N_2658);
xnor U3106 (N_3106,N_2561,N_2798);
nand U3107 (N_3107,N_2807,N_2644);
nand U3108 (N_3108,N_2659,N_2733);
nor U3109 (N_3109,N_2992,N_2657);
nand U3110 (N_3110,N_2606,N_2580);
nand U3111 (N_3111,N_2620,N_2962);
nand U3112 (N_3112,N_2800,N_2757);
nand U3113 (N_3113,N_2775,N_2818);
and U3114 (N_3114,N_2876,N_2817);
and U3115 (N_3115,N_2602,N_2609);
and U3116 (N_3116,N_2812,N_2622);
nand U3117 (N_3117,N_2895,N_2546);
nor U3118 (N_3118,N_2810,N_2772);
nor U3119 (N_3119,N_2934,N_2875);
and U3120 (N_3120,N_2615,N_2532);
and U3121 (N_3121,N_2646,N_2589);
nand U3122 (N_3122,N_2899,N_2897);
nand U3123 (N_3123,N_2715,N_2961);
nand U3124 (N_3124,N_2937,N_2901);
or U3125 (N_3125,N_2594,N_2912);
and U3126 (N_3126,N_2861,N_2908);
and U3127 (N_3127,N_2892,N_2841);
nor U3128 (N_3128,N_2612,N_2591);
xor U3129 (N_3129,N_2850,N_2948);
or U3130 (N_3130,N_2506,N_2730);
and U3131 (N_3131,N_2650,N_2953);
or U3132 (N_3132,N_2538,N_2519);
and U3133 (N_3133,N_2684,N_2911);
and U3134 (N_3134,N_2887,N_2639);
nor U3135 (N_3135,N_2718,N_2918);
nand U3136 (N_3136,N_2618,N_2928);
and U3137 (N_3137,N_2670,N_2689);
nor U3138 (N_3138,N_2534,N_2814);
or U3139 (N_3139,N_2977,N_2759);
xor U3140 (N_3140,N_2641,N_2678);
nand U3141 (N_3141,N_2732,N_2572);
or U3142 (N_3142,N_2619,N_2516);
or U3143 (N_3143,N_2771,N_2967);
or U3144 (N_3144,N_2858,N_2510);
and U3145 (N_3145,N_2921,N_2740);
nor U3146 (N_3146,N_2587,N_2916);
nor U3147 (N_3147,N_2844,N_2865);
or U3148 (N_3148,N_2788,N_2971);
nor U3149 (N_3149,N_2964,N_2528);
nor U3150 (N_3150,N_2522,N_2826);
and U3151 (N_3151,N_2890,N_2614);
or U3152 (N_3152,N_2849,N_2830);
and U3153 (N_3153,N_2989,N_2944);
nor U3154 (N_3154,N_2950,N_2647);
nor U3155 (N_3155,N_2633,N_2557);
nor U3156 (N_3156,N_2994,N_2831);
nand U3157 (N_3157,N_2763,N_2802);
and U3158 (N_3158,N_2913,N_2789);
and U3159 (N_3159,N_2696,N_2578);
nor U3160 (N_3160,N_2720,N_2749);
and U3161 (N_3161,N_2747,N_2645);
or U3162 (N_3162,N_2951,N_2673);
nand U3163 (N_3163,N_2610,N_2529);
nor U3164 (N_3164,N_2613,N_2666);
and U3165 (N_3165,N_2722,N_2624);
nand U3166 (N_3166,N_2938,N_2838);
or U3167 (N_3167,N_2742,N_2537);
and U3168 (N_3168,N_2716,N_2667);
nor U3169 (N_3169,N_2717,N_2631);
and U3170 (N_3170,N_2878,N_2723);
and U3171 (N_3171,N_2920,N_2939);
or U3172 (N_3172,N_2872,N_2811);
and U3173 (N_3173,N_2695,N_2981);
and U3174 (N_3174,N_2991,N_2767);
xnor U3175 (N_3175,N_2784,N_2698);
nor U3176 (N_3176,N_2985,N_2687);
or U3177 (N_3177,N_2570,N_2748);
nor U3178 (N_3178,N_2743,N_2797);
and U3179 (N_3179,N_2764,N_2874);
nand U3180 (N_3180,N_2857,N_2833);
nor U3181 (N_3181,N_2550,N_2704);
nor U3182 (N_3182,N_2676,N_2535);
and U3183 (N_3183,N_2885,N_2821);
nand U3184 (N_3184,N_2688,N_2871);
and U3185 (N_3185,N_2884,N_2975);
or U3186 (N_3186,N_2778,N_2671);
and U3187 (N_3187,N_2508,N_2795);
xnor U3188 (N_3188,N_2754,N_2888);
and U3189 (N_3189,N_2832,N_2611);
or U3190 (N_3190,N_2566,N_2728);
nor U3191 (N_3191,N_2822,N_2517);
or U3192 (N_3192,N_2636,N_2734);
nor U3193 (N_3193,N_2721,N_2652);
or U3194 (N_3194,N_2649,N_2623);
nand U3195 (N_3195,N_2816,N_2706);
and U3196 (N_3196,N_2829,N_2539);
nand U3197 (N_3197,N_2548,N_2804);
nand U3198 (N_3198,N_2518,N_2781);
nand U3199 (N_3199,N_2746,N_2699);
and U3200 (N_3200,N_2959,N_2834);
nor U3201 (N_3201,N_2960,N_2547);
and U3202 (N_3202,N_2970,N_2999);
nand U3203 (N_3203,N_2990,N_2987);
nor U3204 (N_3204,N_2741,N_2945);
and U3205 (N_3205,N_2500,N_2794);
nand U3206 (N_3206,N_2664,N_2940);
and U3207 (N_3207,N_2654,N_2552);
or U3208 (N_3208,N_2969,N_2869);
nand U3209 (N_3209,N_2724,N_2957);
xor U3210 (N_3210,N_2511,N_2827);
nor U3211 (N_3211,N_2815,N_2924);
nor U3212 (N_3212,N_2629,N_2836);
or U3213 (N_3213,N_2792,N_2956);
nand U3214 (N_3214,N_2881,N_2603);
nor U3215 (N_3215,N_2930,N_2780);
xor U3216 (N_3216,N_2709,N_2677);
or U3217 (N_3217,N_2843,N_2766);
nand U3218 (N_3218,N_2569,N_2786);
nand U3219 (N_3219,N_2965,N_2693);
nor U3220 (N_3220,N_2683,N_2562);
nand U3221 (N_3221,N_2919,N_2903);
nor U3222 (N_3222,N_2685,N_2581);
nor U3223 (N_3223,N_2915,N_2768);
and U3224 (N_3224,N_2828,N_2998);
or U3225 (N_3225,N_2565,N_2593);
nor U3226 (N_3226,N_2866,N_2855);
nand U3227 (N_3227,N_2907,N_2980);
or U3228 (N_3228,N_2527,N_2655);
or U3229 (N_3229,N_2776,N_2777);
nand U3230 (N_3230,N_2852,N_2660);
xnor U3231 (N_3231,N_2883,N_2848);
or U3232 (N_3232,N_2617,N_2643);
and U3233 (N_3233,N_2707,N_2638);
nor U3234 (N_3234,N_2859,N_2942);
or U3235 (N_3235,N_2860,N_2635);
nand U3236 (N_3236,N_2702,N_2905);
nor U3237 (N_3237,N_2936,N_2703);
xor U3238 (N_3238,N_2553,N_2583);
or U3239 (N_3239,N_2502,N_2840);
nand U3240 (N_3240,N_2879,N_2632);
nor U3241 (N_3241,N_2796,N_2599);
nor U3242 (N_3242,N_2851,N_2837);
nor U3243 (N_3243,N_2745,N_2663);
nor U3244 (N_3244,N_2787,N_2653);
or U3245 (N_3245,N_2601,N_2979);
nor U3246 (N_3246,N_2597,N_2867);
nand U3247 (N_3247,N_2661,N_2596);
nor U3248 (N_3248,N_2515,N_2997);
nand U3249 (N_3249,N_2526,N_2842);
and U3250 (N_3250,N_2584,N_2684);
nand U3251 (N_3251,N_2932,N_2929);
or U3252 (N_3252,N_2518,N_2598);
and U3253 (N_3253,N_2933,N_2836);
and U3254 (N_3254,N_2528,N_2614);
and U3255 (N_3255,N_2567,N_2857);
or U3256 (N_3256,N_2719,N_2969);
nor U3257 (N_3257,N_2699,N_2606);
nand U3258 (N_3258,N_2512,N_2751);
xnor U3259 (N_3259,N_2623,N_2773);
nor U3260 (N_3260,N_2780,N_2777);
nand U3261 (N_3261,N_2638,N_2595);
nand U3262 (N_3262,N_2979,N_2701);
or U3263 (N_3263,N_2597,N_2894);
and U3264 (N_3264,N_2869,N_2948);
nand U3265 (N_3265,N_2640,N_2527);
or U3266 (N_3266,N_2907,N_2670);
nor U3267 (N_3267,N_2765,N_2944);
nor U3268 (N_3268,N_2731,N_2587);
and U3269 (N_3269,N_2537,N_2927);
or U3270 (N_3270,N_2772,N_2501);
and U3271 (N_3271,N_2765,N_2595);
nor U3272 (N_3272,N_2751,N_2787);
xnor U3273 (N_3273,N_2852,N_2785);
or U3274 (N_3274,N_2719,N_2771);
nor U3275 (N_3275,N_2573,N_2594);
or U3276 (N_3276,N_2946,N_2621);
nor U3277 (N_3277,N_2546,N_2798);
and U3278 (N_3278,N_2514,N_2899);
nand U3279 (N_3279,N_2834,N_2536);
and U3280 (N_3280,N_2520,N_2582);
nand U3281 (N_3281,N_2663,N_2637);
nor U3282 (N_3282,N_2660,N_2974);
nor U3283 (N_3283,N_2684,N_2700);
or U3284 (N_3284,N_2976,N_2936);
or U3285 (N_3285,N_2973,N_2756);
nand U3286 (N_3286,N_2949,N_2893);
or U3287 (N_3287,N_2658,N_2552);
nor U3288 (N_3288,N_2927,N_2530);
nand U3289 (N_3289,N_2680,N_2954);
nor U3290 (N_3290,N_2857,N_2837);
and U3291 (N_3291,N_2817,N_2501);
and U3292 (N_3292,N_2750,N_2892);
nand U3293 (N_3293,N_2874,N_2684);
and U3294 (N_3294,N_2698,N_2756);
and U3295 (N_3295,N_2765,N_2601);
or U3296 (N_3296,N_2749,N_2801);
nand U3297 (N_3297,N_2618,N_2656);
nor U3298 (N_3298,N_2537,N_2662);
or U3299 (N_3299,N_2600,N_2617);
and U3300 (N_3300,N_2977,N_2979);
or U3301 (N_3301,N_2825,N_2537);
or U3302 (N_3302,N_2823,N_2616);
and U3303 (N_3303,N_2651,N_2614);
or U3304 (N_3304,N_2936,N_2628);
and U3305 (N_3305,N_2761,N_2995);
nor U3306 (N_3306,N_2706,N_2733);
nand U3307 (N_3307,N_2782,N_2893);
and U3308 (N_3308,N_2778,N_2819);
and U3309 (N_3309,N_2961,N_2907);
or U3310 (N_3310,N_2861,N_2668);
nor U3311 (N_3311,N_2984,N_2867);
and U3312 (N_3312,N_2541,N_2986);
and U3313 (N_3313,N_2633,N_2809);
and U3314 (N_3314,N_2996,N_2707);
nor U3315 (N_3315,N_2701,N_2502);
nor U3316 (N_3316,N_2539,N_2857);
nand U3317 (N_3317,N_2510,N_2690);
or U3318 (N_3318,N_2695,N_2839);
nand U3319 (N_3319,N_2551,N_2523);
xnor U3320 (N_3320,N_2823,N_2838);
or U3321 (N_3321,N_2766,N_2517);
nor U3322 (N_3322,N_2576,N_2740);
or U3323 (N_3323,N_2668,N_2578);
and U3324 (N_3324,N_2954,N_2831);
nand U3325 (N_3325,N_2682,N_2969);
nor U3326 (N_3326,N_2991,N_2828);
nand U3327 (N_3327,N_2509,N_2840);
nor U3328 (N_3328,N_2880,N_2754);
nand U3329 (N_3329,N_2563,N_2714);
nor U3330 (N_3330,N_2707,N_2637);
or U3331 (N_3331,N_2805,N_2799);
nand U3332 (N_3332,N_2663,N_2703);
or U3333 (N_3333,N_2972,N_2513);
or U3334 (N_3334,N_2539,N_2641);
nor U3335 (N_3335,N_2751,N_2881);
nor U3336 (N_3336,N_2681,N_2702);
and U3337 (N_3337,N_2587,N_2635);
nor U3338 (N_3338,N_2878,N_2942);
nor U3339 (N_3339,N_2514,N_2917);
nor U3340 (N_3340,N_2652,N_2503);
and U3341 (N_3341,N_2527,N_2565);
nand U3342 (N_3342,N_2632,N_2506);
nand U3343 (N_3343,N_2745,N_2657);
or U3344 (N_3344,N_2981,N_2601);
nor U3345 (N_3345,N_2950,N_2804);
or U3346 (N_3346,N_2532,N_2985);
nand U3347 (N_3347,N_2576,N_2537);
nor U3348 (N_3348,N_2907,N_2741);
and U3349 (N_3349,N_2851,N_2573);
or U3350 (N_3350,N_2977,N_2620);
nor U3351 (N_3351,N_2986,N_2790);
nand U3352 (N_3352,N_2855,N_2774);
nor U3353 (N_3353,N_2648,N_2596);
or U3354 (N_3354,N_2563,N_2885);
nor U3355 (N_3355,N_2625,N_2541);
nor U3356 (N_3356,N_2831,N_2899);
nor U3357 (N_3357,N_2518,N_2594);
or U3358 (N_3358,N_2851,N_2849);
or U3359 (N_3359,N_2536,N_2788);
nor U3360 (N_3360,N_2583,N_2925);
and U3361 (N_3361,N_2987,N_2780);
or U3362 (N_3362,N_2603,N_2726);
nor U3363 (N_3363,N_2944,N_2564);
nand U3364 (N_3364,N_2887,N_2795);
and U3365 (N_3365,N_2857,N_2945);
or U3366 (N_3366,N_2987,N_2877);
nand U3367 (N_3367,N_2711,N_2651);
or U3368 (N_3368,N_2855,N_2945);
and U3369 (N_3369,N_2555,N_2632);
and U3370 (N_3370,N_2921,N_2749);
or U3371 (N_3371,N_2553,N_2881);
nor U3372 (N_3372,N_2930,N_2629);
nand U3373 (N_3373,N_2530,N_2858);
nor U3374 (N_3374,N_2805,N_2858);
nor U3375 (N_3375,N_2860,N_2756);
nand U3376 (N_3376,N_2842,N_2772);
nor U3377 (N_3377,N_2743,N_2594);
nand U3378 (N_3378,N_2891,N_2687);
or U3379 (N_3379,N_2575,N_2889);
nor U3380 (N_3380,N_2717,N_2583);
nand U3381 (N_3381,N_2561,N_2961);
nor U3382 (N_3382,N_2871,N_2824);
or U3383 (N_3383,N_2736,N_2911);
nor U3384 (N_3384,N_2986,N_2979);
nor U3385 (N_3385,N_2633,N_2650);
and U3386 (N_3386,N_2918,N_2877);
or U3387 (N_3387,N_2917,N_2984);
and U3388 (N_3388,N_2682,N_2909);
nor U3389 (N_3389,N_2667,N_2630);
and U3390 (N_3390,N_2850,N_2666);
nand U3391 (N_3391,N_2863,N_2891);
nor U3392 (N_3392,N_2983,N_2778);
nand U3393 (N_3393,N_2855,N_2934);
or U3394 (N_3394,N_2790,N_2551);
and U3395 (N_3395,N_2846,N_2571);
or U3396 (N_3396,N_2594,N_2860);
or U3397 (N_3397,N_2977,N_2501);
nor U3398 (N_3398,N_2559,N_2840);
and U3399 (N_3399,N_2744,N_2589);
nand U3400 (N_3400,N_2788,N_2705);
nand U3401 (N_3401,N_2850,N_2667);
nor U3402 (N_3402,N_2523,N_2905);
nand U3403 (N_3403,N_2569,N_2893);
nand U3404 (N_3404,N_2927,N_2626);
or U3405 (N_3405,N_2931,N_2655);
and U3406 (N_3406,N_2901,N_2653);
nand U3407 (N_3407,N_2708,N_2895);
nor U3408 (N_3408,N_2897,N_2638);
and U3409 (N_3409,N_2824,N_2654);
or U3410 (N_3410,N_2711,N_2879);
nand U3411 (N_3411,N_2963,N_2951);
nand U3412 (N_3412,N_2765,N_2972);
and U3413 (N_3413,N_2826,N_2590);
nor U3414 (N_3414,N_2721,N_2879);
nand U3415 (N_3415,N_2518,N_2718);
or U3416 (N_3416,N_2899,N_2695);
nor U3417 (N_3417,N_2835,N_2515);
nand U3418 (N_3418,N_2907,N_2942);
nand U3419 (N_3419,N_2762,N_2893);
xnor U3420 (N_3420,N_2544,N_2857);
or U3421 (N_3421,N_2889,N_2632);
or U3422 (N_3422,N_2973,N_2923);
and U3423 (N_3423,N_2872,N_2826);
or U3424 (N_3424,N_2678,N_2785);
or U3425 (N_3425,N_2917,N_2819);
or U3426 (N_3426,N_2750,N_2801);
and U3427 (N_3427,N_2617,N_2894);
or U3428 (N_3428,N_2803,N_2544);
or U3429 (N_3429,N_2970,N_2891);
and U3430 (N_3430,N_2954,N_2736);
nand U3431 (N_3431,N_2600,N_2578);
and U3432 (N_3432,N_2904,N_2775);
nor U3433 (N_3433,N_2765,N_2905);
and U3434 (N_3434,N_2855,N_2635);
nor U3435 (N_3435,N_2978,N_2560);
and U3436 (N_3436,N_2809,N_2891);
or U3437 (N_3437,N_2976,N_2937);
nand U3438 (N_3438,N_2796,N_2983);
or U3439 (N_3439,N_2878,N_2791);
or U3440 (N_3440,N_2552,N_2868);
or U3441 (N_3441,N_2737,N_2664);
and U3442 (N_3442,N_2935,N_2977);
nor U3443 (N_3443,N_2615,N_2948);
nand U3444 (N_3444,N_2671,N_2913);
xor U3445 (N_3445,N_2934,N_2968);
or U3446 (N_3446,N_2599,N_2669);
or U3447 (N_3447,N_2826,N_2842);
and U3448 (N_3448,N_2555,N_2640);
nor U3449 (N_3449,N_2645,N_2870);
nand U3450 (N_3450,N_2970,N_2786);
or U3451 (N_3451,N_2616,N_2517);
nand U3452 (N_3452,N_2619,N_2918);
and U3453 (N_3453,N_2717,N_2633);
nor U3454 (N_3454,N_2594,N_2515);
nand U3455 (N_3455,N_2920,N_2572);
and U3456 (N_3456,N_2725,N_2546);
and U3457 (N_3457,N_2756,N_2789);
and U3458 (N_3458,N_2552,N_2641);
nor U3459 (N_3459,N_2851,N_2545);
xor U3460 (N_3460,N_2992,N_2915);
and U3461 (N_3461,N_2720,N_2890);
nand U3462 (N_3462,N_2700,N_2562);
nand U3463 (N_3463,N_2561,N_2630);
xor U3464 (N_3464,N_2841,N_2859);
nand U3465 (N_3465,N_2588,N_2664);
and U3466 (N_3466,N_2955,N_2891);
nor U3467 (N_3467,N_2752,N_2888);
nand U3468 (N_3468,N_2734,N_2567);
nand U3469 (N_3469,N_2540,N_2684);
nor U3470 (N_3470,N_2937,N_2648);
nand U3471 (N_3471,N_2927,N_2921);
nand U3472 (N_3472,N_2741,N_2736);
nand U3473 (N_3473,N_2865,N_2615);
nor U3474 (N_3474,N_2778,N_2708);
nand U3475 (N_3475,N_2822,N_2948);
nand U3476 (N_3476,N_2748,N_2898);
nand U3477 (N_3477,N_2610,N_2724);
and U3478 (N_3478,N_2728,N_2956);
and U3479 (N_3479,N_2631,N_2875);
or U3480 (N_3480,N_2506,N_2743);
nor U3481 (N_3481,N_2922,N_2701);
or U3482 (N_3482,N_2864,N_2851);
or U3483 (N_3483,N_2944,N_2930);
and U3484 (N_3484,N_2926,N_2794);
and U3485 (N_3485,N_2900,N_2710);
or U3486 (N_3486,N_2971,N_2955);
xor U3487 (N_3487,N_2552,N_2811);
and U3488 (N_3488,N_2508,N_2992);
nand U3489 (N_3489,N_2511,N_2858);
or U3490 (N_3490,N_2857,N_2713);
nor U3491 (N_3491,N_2629,N_2797);
nand U3492 (N_3492,N_2501,N_2633);
and U3493 (N_3493,N_2541,N_2810);
or U3494 (N_3494,N_2857,N_2903);
nor U3495 (N_3495,N_2620,N_2859);
nor U3496 (N_3496,N_2931,N_2537);
and U3497 (N_3497,N_2732,N_2795);
nor U3498 (N_3498,N_2871,N_2940);
nand U3499 (N_3499,N_2511,N_2535);
nor U3500 (N_3500,N_3091,N_3328);
nand U3501 (N_3501,N_3352,N_3251);
nor U3502 (N_3502,N_3240,N_3196);
and U3503 (N_3503,N_3306,N_3057);
and U3504 (N_3504,N_3066,N_3464);
and U3505 (N_3505,N_3233,N_3408);
and U3506 (N_3506,N_3148,N_3474);
or U3507 (N_3507,N_3270,N_3247);
or U3508 (N_3508,N_3465,N_3107);
nor U3509 (N_3509,N_3297,N_3495);
or U3510 (N_3510,N_3095,N_3365);
nor U3511 (N_3511,N_3001,N_3074);
nor U3512 (N_3512,N_3183,N_3228);
or U3513 (N_3513,N_3372,N_3103);
nor U3514 (N_3514,N_3382,N_3337);
nand U3515 (N_3515,N_3113,N_3271);
nor U3516 (N_3516,N_3283,N_3087);
nor U3517 (N_3517,N_3301,N_3244);
or U3518 (N_3518,N_3289,N_3304);
nand U3519 (N_3519,N_3193,N_3295);
xor U3520 (N_3520,N_3092,N_3303);
or U3521 (N_3521,N_3286,N_3361);
or U3522 (N_3522,N_3349,N_3419);
and U3523 (N_3523,N_3315,N_3359);
nand U3524 (N_3524,N_3348,N_3025);
or U3525 (N_3525,N_3053,N_3498);
or U3526 (N_3526,N_3438,N_3085);
and U3527 (N_3527,N_3044,N_3344);
or U3528 (N_3528,N_3215,N_3032);
nand U3529 (N_3529,N_3071,N_3437);
nand U3530 (N_3530,N_3406,N_3015);
nand U3531 (N_3531,N_3209,N_3332);
and U3532 (N_3532,N_3230,N_3040);
or U3533 (N_3533,N_3075,N_3358);
or U3534 (N_3534,N_3170,N_3083);
nor U3535 (N_3535,N_3314,N_3214);
or U3536 (N_3536,N_3211,N_3429);
nand U3537 (N_3537,N_3168,N_3064);
or U3538 (N_3538,N_3355,N_3364);
or U3539 (N_3539,N_3011,N_3018);
and U3540 (N_3540,N_3448,N_3341);
or U3541 (N_3541,N_3246,N_3147);
nand U3542 (N_3542,N_3176,N_3141);
and U3543 (N_3543,N_3418,N_3264);
xnor U3544 (N_3544,N_3117,N_3178);
nand U3545 (N_3545,N_3009,N_3310);
nand U3546 (N_3546,N_3299,N_3456);
and U3547 (N_3547,N_3427,N_3200);
nor U3548 (N_3548,N_3035,N_3252);
or U3549 (N_3549,N_3030,N_3114);
or U3550 (N_3550,N_3256,N_3182);
nand U3551 (N_3551,N_3201,N_3106);
xnor U3552 (N_3552,N_3157,N_3098);
nand U3553 (N_3553,N_3399,N_3278);
nand U3554 (N_3554,N_3353,N_3043);
nand U3555 (N_3555,N_3369,N_3296);
nor U3556 (N_3556,N_3088,N_3130);
and U3557 (N_3557,N_3363,N_3167);
nor U3558 (N_3558,N_3312,N_3234);
or U3559 (N_3559,N_3006,N_3056);
nand U3560 (N_3560,N_3439,N_3414);
and U3561 (N_3561,N_3477,N_3145);
nand U3562 (N_3562,N_3253,N_3041);
and U3563 (N_3563,N_3089,N_3330);
nand U3564 (N_3564,N_3135,N_3104);
nand U3565 (N_3565,N_3346,N_3119);
nor U3566 (N_3566,N_3449,N_3409);
nand U3567 (N_3567,N_3150,N_3245);
nor U3568 (N_3568,N_3415,N_3423);
nand U3569 (N_3569,N_3189,N_3061);
nand U3570 (N_3570,N_3275,N_3054);
nand U3571 (N_3571,N_3156,N_3421);
and U3572 (N_3572,N_3229,N_3360);
and U3573 (N_3573,N_3146,N_3093);
and U3574 (N_3574,N_3453,N_3099);
nand U3575 (N_3575,N_3466,N_3460);
and U3576 (N_3576,N_3037,N_3070);
nand U3577 (N_3577,N_3120,N_3134);
nand U3578 (N_3578,N_3475,N_3327);
nor U3579 (N_3579,N_3462,N_3187);
xor U3580 (N_3580,N_3012,N_3254);
nand U3581 (N_3581,N_3160,N_3339);
nor U3582 (N_3582,N_3013,N_3375);
and U3583 (N_3583,N_3084,N_3351);
nor U3584 (N_3584,N_3067,N_3463);
nor U3585 (N_3585,N_3292,N_3342);
nor U3586 (N_3586,N_3016,N_3046);
nand U3587 (N_3587,N_3380,N_3336);
and U3588 (N_3588,N_3482,N_3123);
nand U3589 (N_3589,N_3118,N_3020);
and U3590 (N_3590,N_3058,N_3322);
and U3591 (N_3591,N_3468,N_3432);
xor U3592 (N_3592,N_3003,N_3115);
and U3593 (N_3593,N_3285,N_3082);
or U3594 (N_3594,N_3396,N_3192);
nand U3595 (N_3595,N_3371,N_3316);
nor U3596 (N_3596,N_3321,N_3329);
and U3597 (N_3597,N_3195,N_3100);
nor U3598 (N_3598,N_3131,N_3052);
nand U3599 (N_3599,N_3220,N_3065);
nand U3600 (N_3600,N_3048,N_3407);
nor U3601 (N_3601,N_3425,N_3305);
and U3602 (N_3602,N_3362,N_3478);
nand U3603 (N_3603,N_3174,N_3413);
nor U3604 (N_3604,N_3036,N_3129);
or U3605 (N_3605,N_3207,N_3300);
or U3606 (N_3606,N_3203,N_3441);
and U3607 (N_3607,N_3333,N_3491);
and U3608 (N_3608,N_3481,N_3444);
and U3609 (N_3609,N_3451,N_3005);
and U3610 (N_3610,N_3487,N_3402);
nand U3611 (N_3611,N_3259,N_3469);
nor U3612 (N_3612,N_3267,N_3266);
nand U3613 (N_3613,N_3105,N_3279);
or U3614 (N_3614,N_3242,N_3412);
or U3615 (N_3615,N_3436,N_3197);
xor U3616 (N_3616,N_3260,N_3488);
and U3617 (N_3617,N_3384,N_3308);
and U3618 (N_3618,N_3169,N_3010);
nor U3619 (N_3619,N_3383,N_3216);
and U3620 (N_3620,N_3389,N_3378);
and U3621 (N_3621,N_3411,N_3094);
or U3622 (N_3622,N_3161,N_3325);
and U3623 (N_3623,N_3345,N_3077);
nand U3624 (N_3624,N_3096,N_3366);
xnor U3625 (N_3625,N_3493,N_3347);
or U3626 (N_3626,N_3318,N_3155);
and U3627 (N_3627,N_3097,N_3068);
and U3628 (N_3628,N_3014,N_3374);
and U3629 (N_3629,N_3248,N_3250);
nand U3630 (N_3630,N_3177,N_3467);
nand U3631 (N_3631,N_3079,N_3442);
or U3632 (N_3632,N_3231,N_3224);
nor U3633 (N_3633,N_3000,N_3401);
and U3634 (N_3634,N_3357,N_3241);
nor U3635 (N_3635,N_3479,N_3494);
and U3636 (N_3636,N_3072,N_3208);
nor U3637 (N_3637,N_3368,N_3073);
and U3638 (N_3638,N_3027,N_3403);
nand U3639 (N_3639,N_3039,N_3446);
and U3640 (N_3640,N_3078,N_3454);
or U3641 (N_3641,N_3002,N_3116);
and U3642 (N_3642,N_3317,N_3268);
nor U3643 (N_3643,N_3017,N_3294);
and U3644 (N_3644,N_3434,N_3435);
nor U3645 (N_3645,N_3338,N_3038);
and U3646 (N_3646,N_3159,N_3138);
or U3647 (N_3647,N_3142,N_3485);
nor U3648 (N_3648,N_3239,N_3184);
or U3649 (N_3649,N_3210,N_3045);
or U3650 (N_3650,N_3205,N_3221);
and U3651 (N_3651,N_3219,N_3356);
or U3652 (N_3652,N_3171,N_3126);
xnor U3653 (N_3653,N_3143,N_3023);
nor U3654 (N_3654,N_3154,N_3455);
nor U3655 (N_3655,N_3019,N_3175);
nor U3656 (N_3656,N_3133,N_3059);
and U3657 (N_3657,N_3062,N_3188);
nor U3658 (N_3658,N_3029,N_3452);
and U3659 (N_3659,N_3461,N_3125);
or U3660 (N_3660,N_3472,N_3280);
and U3661 (N_3661,N_3202,N_3108);
or U3662 (N_3662,N_3471,N_3139);
or U3663 (N_3663,N_3185,N_3031);
nand U3664 (N_3664,N_3324,N_3144);
nand U3665 (N_3665,N_3024,N_3284);
nand U3666 (N_3666,N_3354,N_3319);
and U3667 (N_3667,N_3377,N_3213);
and U3668 (N_3668,N_3033,N_3217);
nor U3669 (N_3669,N_3163,N_3034);
and U3670 (N_3670,N_3291,N_3249);
or U3671 (N_3671,N_3181,N_3225);
and U3672 (N_3672,N_3186,N_3483);
and U3673 (N_3673,N_3237,N_3026);
nand U3674 (N_3674,N_3496,N_3109);
and U3675 (N_3675,N_3398,N_3343);
or U3676 (N_3676,N_3261,N_3090);
and U3677 (N_3677,N_3121,N_3497);
or U3678 (N_3678,N_3334,N_3004);
nor U3679 (N_3679,N_3257,N_3424);
or U3680 (N_3680,N_3445,N_3152);
and U3681 (N_3681,N_3350,N_3122);
nand U3682 (N_3682,N_3222,N_3243);
nand U3683 (N_3683,N_3111,N_3028);
nor U3684 (N_3684,N_3290,N_3484);
and U3685 (N_3685,N_3367,N_3262);
nor U3686 (N_3686,N_3320,N_3391);
and U3687 (N_3687,N_3051,N_3081);
and U3688 (N_3688,N_3486,N_3166);
and U3689 (N_3689,N_3307,N_3311);
or U3690 (N_3690,N_3255,N_3489);
xnor U3691 (N_3691,N_3263,N_3470);
nand U3692 (N_3692,N_3063,N_3236);
nor U3693 (N_3693,N_3218,N_3450);
nand U3694 (N_3694,N_3400,N_3323);
or U3695 (N_3695,N_3370,N_3232);
nand U3696 (N_3696,N_3490,N_3430);
nor U3697 (N_3697,N_3373,N_3393);
nor U3698 (N_3698,N_3136,N_3404);
nand U3699 (N_3699,N_3459,N_3313);
nor U3700 (N_3700,N_3179,N_3492);
or U3701 (N_3701,N_3394,N_3128);
or U3702 (N_3702,N_3416,N_3173);
nor U3703 (N_3703,N_3458,N_3457);
and U3704 (N_3704,N_3055,N_3381);
and U3705 (N_3705,N_3151,N_3238);
or U3706 (N_3706,N_3410,N_3417);
or U3707 (N_3707,N_3326,N_3110);
or U3708 (N_3708,N_3235,N_3190);
nor U3709 (N_3709,N_3433,N_3282);
nand U3710 (N_3710,N_3276,N_3049);
or U3711 (N_3711,N_3340,N_3265);
nand U3712 (N_3712,N_3101,N_3165);
and U3713 (N_3713,N_3387,N_3153);
and U3714 (N_3714,N_3199,N_3331);
or U3715 (N_3715,N_3180,N_3080);
or U3716 (N_3716,N_3277,N_3140);
nor U3717 (N_3717,N_3223,N_3440);
nand U3718 (N_3718,N_3162,N_3047);
nand U3719 (N_3719,N_3388,N_3395);
or U3720 (N_3720,N_3422,N_3132);
nand U3721 (N_3721,N_3204,N_3273);
or U3722 (N_3722,N_3287,N_3212);
or U3723 (N_3723,N_3386,N_3428);
nor U3724 (N_3724,N_3022,N_3473);
nand U3725 (N_3725,N_3443,N_3480);
and U3726 (N_3726,N_3302,N_3127);
or U3727 (N_3727,N_3258,N_3112);
nand U3728 (N_3728,N_3269,N_3102);
and U3729 (N_3729,N_3379,N_3164);
nand U3730 (N_3730,N_3206,N_3191);
and U3731 (N_3731,N_3499,N_3272);
and U3732 (N_3732,N_3060,N_3069);
and U3733 (N_3733,N_3021,N_3042);
or U3734 (N_3734,N_3281,N_3124);
and U3735 (N_3735,N_3149,N_3392);
nand U3736 (N_3736,N_3431,N_3376);
nor U3737 (N_3737,N_3390,N_3194);
or U3738 (N_3738,N_3007,N_3172);
or U3739 (N_3739,N_3420,N_3226);
nor U3740 (N_3740,N_3050,N_3076);
or U3741 (N_3741,N_3288,N_3405);
and U3742 (N_3742,N_3198,N_3309);
and U3743 (N_3743,N_3086,N_3426);
and U3744 (N_3744,N_3335,N_3476);
nand U3745 (N_3745,N_3298,N_3274);
and U3746 (N_3746,N_3008,N_3447);
or U3747 (N_3747,N_3397,N_3158);
nand U3748 (N_3748,N_3293,N_3137);
nand U3749 (N_3749,N_3227,N_3385);
and U3750 (N_3750,N_3217,N_3281);
nand U3751 (N_3751,N_3359,N_3433);
nand U3752 (N_3752,N_3370,N_3192);
nor U3753 (N_3753,N_3425,N_3231);
and U3754 (N_3754,N_3286,N_3195);
or U3755 (N_3755,N_3467,N_3213);
and U3756 (N_3756,N_3459,N_3369);
nor U3757 (N_3757,N_3265,N_3427);
nand U3758 (N_3758,N_3249,N_3293);
nor U3759 (N_3759,N_3158,N_3454);
nand U3760 (N_3760,N_3207,N_3377);
or U3761 (N_3761,N_3148,N_3496);
nand U3762 (N_3762,N_3246,N_3310);
and U3763 (N_3763,N_3137,N_3246);
nor U3764 (N_3764,N_3401,N_3376);
or U3765 (N_3765,N_3030,N_3249);
or U3766 (N_3766,N_3268,N_3092);
and U3767 (N_3767,N_3353,N_3074);
and U3768 (N_3768,N_3071,N_3249);
xnor U3769 (N_3769,N_3170,N_3321);
or U3770 (N_3770,N_3144,N_3243);
nand U3771 (N_3771,N_3239,N_3195);
and U3772 (N_3772,N_3066,N_3237);
nand U3773 (N_3773,N_3087,N_3112);
or U3774 (N_3774,N_3353,N_3141);
nand U3775 (N_3775,N_3457,N_3119);
nor U3776 (N_3776,N_3172,N_3069);
or U3777 (N_3777,N_3297,N_3367);
nand U3778 (N_3778,N_3133,N_3231);
and U3779 (N_3779,N_3037,N_3019);
nand U3780 (N_3780,N_3376,N_3330);
and U3781 (N_3781,N_3179,N_3054);
or U3782 (N_3782,N_3164,N_3426);
nand U3783 (N_3783,N_3360,N_3211);
and U3784 (N_3784,N_3062,N_3318);
nand U3785 (N_3785,N_3439,N_3464);
nand U3786 (N_3786,N_3290,N_3380);
nor U3787 (N_3787,N_3070,N_3247);
nor U3788 (N_3788,N_3131,N_3227);
nand U3789 (N_3789,N_3236,N_3160);
and U3790 (N_3790,N_3323,N_3113);
and U3791 (N_3791,N_3140,N_3156);
nor U3792 (N_3792,N_3290,N_3038);
nand U3793 (N_3793,N_3143,N_3438);
nand U3794 (N_3794,N_3181,N_3082);
or U3795 (N_3795,N_3375,N_3251);
and U3796 (N_3796,N_3391,N_3203);
nand U3797 (N_3797,N_3329,N_3080);
and U3798 (N_3798,N_3395,N_3327);
or U3799 (N_3799,N_3315,N_3021);
or U3800 (N_3800,N_3304,N_3468);
nor U3801 (N_3801,N_3125,N_3091);
and U3802 (N_3802,N_3402,N_3056);
nor U3803 (N_3803,N_3359,N_3065);
or U3804 (N_3804,N_3473,N_3493);
or U3805 (N_3805,N_3154,N_3035);
or U3806 (N_3806,N_3050,N_3352);
or U3807 (N_3807,N_3131,N_3356);
or U3808 (N_3808,N_3224,N_3170);
or U3809 (N_3809,N_3154,N_3118);
or U3810 (N_3810,N_3072,N_3295);
nand U3811 (N_3811,N_3333,N_3021);
nor U3812 (N_3812,N_3311,N_3459);
and U3813 (N_3813,N_3430,N_3004);
and U3814 (N_3814,N_3495,N_3393);
and U3815 (N_3815,N_3228,N_3193);
nor U3816 (N_3816,N_3288,N_3446);
nand U3817 (N_3817,N_3258,N_3297);
or U3818 (N_3818,N_3170,N_3446);
nand U3819 (N_3819,N_3454,N_3388);
and U3820 (N_3820,N_3280,N_3267);
and U3821 (N_3821,N_3371,N_3329);
nand U3822 (N_3822,N_3294,N_3360);
nand U3823 (N_3823,N_3023,N_3223);
nor U3824 (N_3824,N_3376,N_3329);
nand U3825 (N_3825,N_3168,N_3035);
nor U3826 (N_3826,N_3294,N_3194);
nand U3827 (N_3827,N_3404,N_3162);
nor U3828 (N_3828,N_3338,N_3260);
and U3829 (N_3829,N_3461,N_3246);
nand U3830 (N_3830,N_3315,N_3026);
nor U3831 (N_3831,N_3249,N_3416);
nor U3832 (N_3832,N_3330,N_3477);
or U3833 (N_3833,N_3480,N_3413);
nor U3834 (N_3834,N_3033,N_3392);
nand U3835 (N_3835,N_3198,N_3168);
nor U3836 (N_3836,N_3250,N_3330);
nand U3837 (N_3837,N_3203,N_3414);
nand U3838 (N_3838,N_3202,N_3245);
nand U3839 (N_3839,N_3232,N_3251);
nand U3840 (N_3840,N_3193,N_3108);
or U3841 (N_3841,N_3174,N_3203);
nand U3842 (N_3842,N_3252,N_3277);
nand U3843 (N_3843,N_3134,N_3428);
nor U3844 (N_3844,N_3383,N_3147);
nor U3845 (N_3845,N_3065,N_3082);
nor U3846 (N_3846,N_3465,N_3334);
nor U3847 (N_3847,N_3105,N_3290);
and U3848 (N_3848,N_3408,N_3154);
nor U3849 (N_3849,N_3366,N_3233);
nand U3850 (N_3850,N_3389,N_3391);
or U3851 (N_3851,N_3161,N_3443);
nand U3852 (N_3852,N_3028,N_3334);
nand U3853 (N_3853,N_3239,N_3155);
and U3854 (N_3854,N_3270,N_3067);
nand U3855 (N_3855,N_3312,N_3215);
and U3856 (N_3856,N_3129,N_3427);
nor U3857 (N_3857,N_3079,N_3301);
nor U3858 (N_3858,N_3383,N_3344);
nor U3859 (N_3859,N_3225,N_3325);
nand U3860 (N_3860,N_3291,N_3426);
nand U3861 (N_3861,N_3365,N_3249);
nand U3862 (N_3862,N_3235,N_3421);
and U3863 (N_3863,N_3385,N_3357);
or U3864 (N_3864,N_3355,N_3058);
nand U3865 (N_3865,N_3201,N_3171);
nor U3866 (N_3866,N_3463,N_3035);
nor U3867 (N_3867,N_3207,N_3450);
nand U3868 (N_3868,N_3482,N_3345);
nand U3869 (N_3869,N_3056,N_3455);
or U3870 (N_3870,N_3249,N_3358);
nor U3871 (N_3871,N_3488,N_3113);
nor U3872 (N_3872,N_3384,N_3149);
nand U3873 (N_3873,N_3267,N_3008);
nor U3874 (N_3874,N_3392,N_3459);
nand U3875 (N_3875,N_3346,N_3479);
and U3876 (N_3876,N_3435,N_3302);
nand U3877 (N_3877,N_3370,N_3150);
and U3878 (N_3878,N_3282,N_3399);
xor U3879 (N_3879,N_3193,N_3236);
or U3880 (N_3880,N_3039,N_3178);
or U3881 (N_3881,N_3338,N_3257);
nor U3882 (N_3882,N_3342,N_3241);
or U3883 (N_3883,N_3081,N_3381);
and U3884 (N_3884,N_3178,N_3342);
and U3885 (N_3885,N_3460,N_3217);
nor U3886 (N_3886,N_3251,N_3409);
and U3887 (N_3887,N_3001,N_3139);
or U3888 (N_3888,N_3161,N_3227);
or U3889 (N_3889,N_3128,N_3402);
nor U3890 (N_3890,N_3433,N_3048);
nor U3891 (N_3891,N_3007,N_3262);
or U3892 (N_3892,N_3242,N_3241);
nand U3893 (N_3893,N_3146,N_3366);
or U3894 (N_3894,N_3036,N_3172);
and U3895 (N_3895,N_3430,N_3107);
xor U3896 (N_3896,N_3126,N_3436);
and U3897 (N_3897,N_3346,N_3484);
nand U3898 (N_3898,N_3230,N_3488);
nand U3899 (N_3899,N_3104,N_3180);
nand U3900 (N_3900,N_3057,N_3115);
or U3901 (N_3901,N_3483,N_3007);
and U3902 (N_3902,N_3346,N_3252);
nand U3903 (N_3903,N_3433,N_3361);
and U3904 (N_3904,N_3430,N_3495);
or U3905 (N_3905,N_3469,N_3051);
nor U3906 (N_3906,N_3021,N_3249);
nand U3907 (N_3907,N_3058,N_3137);
nand U3908 (N_3908,N_3404,N_3031);
and U3909 (N_3909,N_3176,N_3257);
nand U3910 (N_3910,N_3445,N_3139);
nor U3911 (N_3911,N_3444,N_3073);
and U3912 (N_3912,N_3463,N_3454);
nor U3913 (N_3913,N_3182,N_3450);
nand U3914 (N_3914,N_3245,N_3111);
and U3915 (N_3915,N_3050,N_3054);
or U3916 (N_3916,N_3342,N_3334);
nor U3917 (N_3917,N_3232,N_3006);
nor U3918 (N_3918,N_3139,N_3415);
or U3919 (N_3919,N_3022,N_3402);
and U3920 (N_3920,N_3078,N_3307);
or U3921 (N_3921,N_3108,N_3245);
and U3922 (N_3922,N_3026,N_3313);
or U3923 (N_3923,N_3016,N_3469);
nor U3924 (N_3924,N_3047,N_3469);
nor U3925 (N_3925,N_3265,N_3238);
or U3926 (N_3926,N_3071,N_3345);
nand U3927 (N_3927,N_3497,N_3109);
and U3928 (N_3928,N_3417,N_3428);
nor U3929 (N_3929,N_3354,N_3045);
nor U3930 (N_3930,N_3232,N_3135);
nor U3931 (N_3931,N_3120,N_3041);
nor U3932 (N_3932,N_3076,N_3040);
nand U3933 (N_3933,N_3011,N_3297);
and U3934 (N_3934,N_3182,N_3318);
nor U3935 (N_3935,N_3334,N_3249);
xor U3936 (N_3936,N_3061,N_3100);
or U3937 (N_3937,N_3393,N_3205);
nand U3938 (N_3938,N_3314,N_3277);
or U3939 (N_3939,N_3022,N_3263);
and U3940 (N_3940,N_3069,N_3010);
nor U3941 (N_3941,N_3352,N_3073);
or U3942 (N_3942,N_3383,N_3197);
nand U3943 (N_3943,N_3119,N_3098);
and U3944 (N_3944,N_3285,N_3201);
nor U3945 (N_3945,N_3234,N_3090);
nand U3946 (N_3946,N_3333,N_3470);
or U3947 (N_3947,N_3411,N_3327);
nor U3948 (N_3948,N_3390,N_3151);
nand U3949 (N_3949,N_3336,N_3265);
nor U3950 (N_3950,N_3135,N_3097);
nand U3951 (N_3951,N_3351,N_3417);
or U3952 (N_3952,N_3373,N_3449);
nor U3953 (N_3953,N_3489,N_3387);
xnor U3954 (N_3954,N_3106,N_3326);
nand U3955 (N_3955,N_3027,N_3209);
nand U3956 (N_3956,N_3383,N_3475);
and U3957 (N_3957,N_3423,N_3384);
nor U3958 (N_3958,N_3212,N_3216);
or U3959 (N_3959,N_3108,N_3475);
and U3960 (N_3960,N_3208,N_3235);
nand U3961 (N_3961,N_3141,N_3097);
nand U3962 (N_3962,N_3119,N_3419);
nand U3963 (N_3963,N_3285,N_3127);
nor U3964 (N_3964,N_3011,N_3439);
xnor U3965 (N_3965,N_3350,N_3184);
nor U3966 (N_3966,N_3394,N_3026);
nor U3967 (N_3967,N_3352,N_3121);
nand U3968 (N_3968,N_3486,N_3373);
nor U3969 (N_3969,N_3290,N_3143);
or U3970 (N_3970,N_3415,N_3323);
nand U3971 (N_3971,N_3317,N_3149);
or U3972 (N_3972,N_3349,N_3372);
or U3973 (N_3973,N_3117,N_3048);
or U3974 (N_3974,N_3274,N_3403);
nor U3975 (N_3975,N_3118,N_3420);
nor U3976 (N_3976,N_3024,N_3123);
and U3977 (N_3977,N_3441,N_3192);
and U3978 (N_3978,N_3064,N_3343);
or U3979 (N_3979,N_3051,N_3281);
nor U3980 (N_3980,N_3436,N_3443);
or U3981 (N_3981,N_3001,N_3217);
nor U3982 (N_3982,N_3057,N_3089);
nor U3983 (N_3983,N_3130,N_3264);
nor U3984 (N_3984,N_3208,N_3187);
or U3985 (N_3985,N_3411,N_3160);
or U3986 (N_3986,N_3460,N_3470);
or U3987 (N_3987,N_3229,N_3201);
or U3988 (N_3988,N_3415,N_3086);
or U3989 (N_3989,N_3000,N_3121);
nor U3990 (N_3990,N_3198,N_3479);
and U3991 (N_3991,N_3460,N_3368);
nand U3992 (N_3992,N_3398,N_3383);
and U3993 (N_3993,N_3402,N_3179);
nand U3994 (N_3994,N_3031,N_3447);
nor U3995 (N_3995,N_3314,N_3293);
and U3996 (N_3996,N_3179,N_3065);
and U3997 (N_3997,N_3068,N_3006);
nand U3998 (N_3998,N_3023,N_3040);
xor U3999 (N_3999,N_3374,N_3315);
nor U4000 (N_4000,N_3908,N_3674);
or U4001 (N_4001,N_3869,N_3958);
nand U4002 (N_4002,N_3868,N_3986);
nand U4003 (N_4003,N_3858,N_3837);
nand U4004 (N_4004,N_3712,N_3609);
or U4005 (N_4005,N_3607,N_3900);
or U4006 (N_4006,N_3553,N_3894);
nand U4007 (N_4007,N_3801,N_3875);
nand U4008 (N_4008,N_3642,N_3898);
and U4009 (N_4009,N_3663,N_3807);
nand U4010 (N_4010,N_3647,N_3742);
nor U4011 (N_4011,N_3655,N_3882);
and U4012 (N_4012,N_3561,N_3501);
and U4013 (N_4013,N_3667,N_3690);
nand U4014 (N_4014,N_3987,N_3773);
nand U4015 (N_4015,N_3595,N_3623);
nor U4016 (N_4016,N_3866,N_3877);
nor U4017 (N_4017,N_3852,N_3989);
nor U4018 (N_4018,N_3550,N_3648);
and U4019 (N_4019,N_3565,N_3618);
and U4020 (N_4020,N_3803,N_3927);
and U4021 (N_4021,N_3760,N_3765);
and U4022 (N_4022,N_3814,N_3694);
and U4023 (N_4023,N_3670,N_3810);
or U4024 (N_4024,N_3676,N_3686);
nor U4025 (N_4025,N_3794,N_3833);
nor U4026 (N_4026,N_3622,N_3872);
and U4027 (N_4027,N_3813,N_3800);
nand U4028 (N_4028,N_3685,N_3588);
nand U4029 (N_4029,N_3909,N_3562);
nand U4030 (N_4030,N_3612,N_3913);
and U4031 (N_4031,N_3996,N_3579);
or U4032 (N_4032,N_3717,N_3665);
and U4033 (N_4033,N_3834,N_3584);
and U4034 (N_4034,N_3608,N_3515);
and U4035 (N_4035,N_3727,N_3829);
or U4036 (N_4036,N_3785,N_3977);
and U4037 (N_4037,N_3514,N_3723);
nor U4038 (N_4038,N_3518,N_3692);
nand U4039 (N_4039,N_3981,N_3512);
and U4040 (N_4040,N_3527,N_3681);
or U4041 (N_4041,N_3855,N_3994);
nor U4042 (N_4042,N_3632,N_3629);
or U4043 (N_4043,N_3583,N_3611);
and U4044 (N_4044,N_3574,N_3902);
nor U4045 (N_4045,N_3990,N_3641);
xor U4046 (N_4046,N_3534,N_3741);
or U4047 (N_4047,N_3532,N_3923);
or U4048 (N_4048,N_3839,N_3624);
nor U4049 (N_4049,N_3957,N_3998);
nor U4050 (N_4050,N_3896,N_3802);
and U4051 (N_4051,N_3503,N_3854);
nor U4052 (N_4052,N_3976,N_3770);
nor U4053 (N_4053,N_3747,N_3911);
and U4054 (N_4054,N_3951,N_3587);
nand U4055 (N_4055,N_3576,N_3700);
xor U4056 (N_4056,N_3889,N_3711);
and U4057 (N_4057,N_3787,N_3573);
and U4058 (N_4058,N_3556,N_3649);
and U4059 (N_4059,N_3631,N_3728);
nor U4060 (N_4060,N_3606,N_3945);
nor U4061 (N_4061,N_3849,N_3703);
or U4062 (N_4062,N_3755,N_3654);
or U4063 (N_4063,N_3821,N_3640);
nand U4064 (N_4064,N_3566,N_3823);
or U4065 (N_4065,N_3984,N_3962);
or U4066 (N_4066,N_3835,N_3726);
nand U4067 (N_4067,N_3838,N_3548);
and U4068 (N_4068,N_3751,N_3825);
and U4069 (N_4069,N_3888,N_3819);
nor U4070 (N_4070,N_3521,N_3954);
and U4071 (N_4071,N_3666,N_3675);
or U4072 (N_4072,N_3560,N_3806);
nor U4073 (N_4073,N_3828,N_3682);
nand U4074 (N_4074,N_3955,N_3589);
xor U4075 (N_4075,N_3792,N_3740);
and U4076 (N_4076,N_3997,N_3644);
nor U4077 (N_4077,N_3856,N_3526);
and U4078 (N_4078,N_3972,N_3547);
nor U4079 (N_4079,N_3847,N_3953);
nand U4080 (N_4080,N_3914,N_3893);
and U4081 (N_4081,N_3926,N_3643);
nand U4082 (N_4082,N_3591,N_3536);
or U4083 (N_4083,N_3774,N_3830);
nand U4084 (N_4084,N_3567,N_3704);
nor U4085 (N_4085,N_3967,N_3795);
nand U4086 (N_4086,N_3702,N_3918);
nor U4087 (N_4087,N_3621,N_3636);
nor U4088 (N_4088,N_3693,N_3883);
nand U4089 (N_4089,N_3523,N_3516);
nand U4090 (N_4090,N_3988,N_3777);
and U4091 (N_4091,N_3948,N_3797);
or U4092 (N_4092,N_3615,N_3610);
or U4093 (N_4093,N_3840,N_3881);
or U4094 (N_4094,N_3944,N_3769);
nand U4095 (N_4095,N_3921,N_3544);
or U4096 (N_4096,N_3818,N_3710);
and U4097 (N_4097,N_3890,N_3511);
and U4098 (N_4098,N_3718,N_3980);
or U4099 (N_4099,N_3793,N_3558);
and U4100 (N_4100,N_3942,N_3708);
or U4101 (N_4101,N_3683,N_3705);
or U4102 (N_4102,N_3815,N_3738);
and U4103 (N_4103,N_3920,N_3651);
nor U4104 (N_4104,N_3906,N_3910);
and U4105 (N_4105,N_3721,N_3941);
nor U4106 (N_4106,N_3940,N_3687);
or U4107 (N_4107,N_3634,N_3846);
xnor U4108 (N_4108,N_3713,N_3983);
and U4109 (N_4109,N_3791,N_3932);
xnor U4110 (N_4110,N_3824,N_3851);
or U4111 (N_4111,N_3778,N_3677);
nor U4112 (N_4112,N_3645,N_3873);
or U4113 (N_4113,N_3720,N_3772);
nand U4114 (N_4114,N_3684,N_3762);
nand U4115 (N_4115,N_3656,N_3575);
nand U4116 (N_4116,N_3991,N_3968);
and U4117 (N_4117,N_3580,N_3780);
nor U4118 (N_4118,N_3943,N_3689);
nand U4119 (N_4119,N_3601,N_3659);
or U4120 (N_4120,N_3695,N_3733);
nor U4121 (N_4121,N_3520,N_3500);
or U4122 (N_4122,N_3904,N_3593);
nand U4123 (N_4123,N_3749,N_3603);
and U4124 (N_4124,N_3820,N_3935);
nand U4125 (N_4125,N_3731,N_3581);
nor U4126 (N_4126,N_3864,N_3964);
nor U4127 (N_4127,N_3844,N_3826);
nor U4128 (N_4128,N_3892,N_3979);
and U4129 (N_4129,N_3812,N_3771);
nor U4130 (N_4130,N_3756,N_3734);
and U4131 (N_4131,N_3714,N_3633);
nand U4132 (N_4132,N_3706,N_3563);
nor U4133 (N_4133,N_3775,N_3750);
or U4134 (N_4134,N_3568,N_3571);
nand U4135 (N_4135,N_3860,N_3763);
nor U4136 (N_4136,N_3845,N_3551);
nand U4137 (N_4137,N_3745,N_3817);
or U4138 (N_4138,N_3669,N_3937);
nor U4139 (N_4139,N_3691,N_3969);
and U4140 (N_4140,N_3585,N_3946);
nand U4141 (N_4141,N_3552,N_3688);
or U4142 (N_4142,N_3639,N_3907);
and U4143 (N_4143,N_3759,N_3668);
nor U4144 (N_4144,N_3799,N_3886);
nand U4145 (N_4145,N_3798,N_3730);
and U4146 (N_4146,N_3614,N_3549);
and U4147 (N_4147,N_3832,N_3657);
or U4148 (N_4148,N_3925,N_3535);
nand U4149 (N_4149,N_3808,N_3528);
or U4150 (N_4150,N_3600,N_3978);
nand U4151 (N_4151,N_3783,N_3929);
nor U4152 (N_4152,N_3732,N_3861);
nand U4153 (N_4153,N_3960,N_3754);
xor U4154 (N_4154,N_3782,N_3796);
and U4155 (N_4155,N_3930,N_3905);
or U4156 (N_4156,N_3533,N_3934);
and U4157 (N_4157,N_3933,N_3507);
or U4158 (N_4158,N_3959,N_3707);
nor U4159 (N_4159,N_3891,N_3963);
or U4160 (N_4160,N_3776,N_3637);
xnor U4161 (N_4161,N_3874,N_3850);
nand U4162 (N_4162,N_3961,N_3592);
nand U4163 (N_4163,N_3788,N_3862);
or U4164 (N_4164,N_3790,N_3901);
nor U4165 (N_4165,N_3748,N_3950);
nand U4166 (N_4166,N_3922,N_3506);
nand U4167 (N_4167,N_3537,N_3816);
and U4168 (N_4168,N_3540,N_3671);
or U4169 (N_4169,N_3966,N_3938);
and U4170 (N_4170,N_3903,N_3982);
and U4171 (N_4171,N_3519,N_3764);
and U4172 (N_4172,N_3616,N_3586);
or U4173 (N_4173,N_3928,N_3917);
nand U4174 (N_4174,N_3661,N_3857);
nand U4175 (N_4175,N_3993,N_3784);
nor U4176 (N_4176,N_3572,N_3952);
or U4177 (N_4177,N_3646,N_3582);
nor U4178 (N_4178,N_3545,N_3753);
nand U4179 (N_4179,N_3912,N_3919);
xnor U4180 (N_4180,N_3590,N_3696);
and U4181 (N_4181,N_3627,N_3766);
or U4182 (N_4182,N_3811,N_3542);
or U4183 (N_4183,N_3719,N_3779);
nand U4184 (N_4184,N_3508,N_3768);
nor U4185 (N_4185,N_3736,N_3831);
or U4186 (N_4186,N_3554,N_3635);
xor U4187 (N_4187,N_3716,N_3975);
and U4188 (N_4188,N_3505,N_3625);
or U4189 (N_4189,N_3569,N_3504);
nand U4190 (N_4190,N_3529,N_3722);
and U4191 (N_4191,N_3758,N_3539);
nor U4192 (N_4192,N_3638,N_3739);
nand U4193 (N_4193,N_3956,N_3744);
or U4194 (N_4194,N_3680,N_3767);
nand U4195 (N_4195,N_3658,N_3510);
and U4196 (N_4196,N_3939,N_3971);
or U4197 (N_4197,N_3789,N_3842);
or U4198 (N_4198,N_3604,N_3848);
nor U4199 (N_4199,N_3502,N_3822);
or U4200 (N_4200,N_3619,N_3827);
or U4201 (N_4201,N_3679,N_3781);
or U4202 (N_4202,N_3884,N_3598);
nor U4203 (N_4203,N_3859,N_3757);
nor U4204 (N_4204,N_3660,N_3867);
and U4205 (N_4205,N_3973,N_3599);
nor U4206 (N_4206,N_3628,N_3517);
nor U4207 (N_4207,N_3613,N_3701);
nor U4208 (N_4208,N_3559,N_3678);
xnor U4209 (N_4209,N_3602,N_3897);
and U4210 (N_4210,N_3786,N_3931);
nor U4211 (N_4211,N_3617,N_3715);
nand U4212 (N_4212,N_3672,N_3879);
or U4213 (N_4213,N_3924,N_3531);
nand U4214 (N_4214,N_3853,N_3887);
nor U4215 (N_4215,N_3876,N_3836);
or U4216 (N_4216,N_3570,N_3916);
nand U4217 (N_4217,N_3809,N_3538);
nand U4218 (N_4218,N_3863,N_3985);
nand U4219 (N_4219,N_3737,N_3509);
nand U4220 (N_4220,N_3578,N_3743);
nor U4221 (N_4221,N_3564,N_3804);
or U4222 (N_4222,N_3999,N_3974);
and U4223 (N_4223,N_3513,N_3662);
nand U4224 (N_4224,N_3597,N_3577);
and U4225 (N_4225,N_3949,N_3843);
or U4226 (N_4226,N_3841,N_3995);
nor U4227 (N_4227,N_3880,N_3992);
xnor U4228 (N_4228,N_3546,N_3805);
and U4229 (N_4229,N_3871,N_3895);
or U4230 (N_4230,N_3725,N_3620);
nor U4231 (N_4231,N_3965,N_3936);
and U4232 (N_4232,N_3522,N_3605);
and U4233 (N_4233,N_3530,N_3524);
or U4234 (N_4234,N_3709,N_3915);
nand U4235 (N_4235,N_3870,N_3865);
nor U4236 (N_4236,N_3596,N_3735);
and U4237 (N_4237,N_3761,N_3752);
nand U4238 (N_4238,N_3947,N_3555);
and U4239 (N_4239,N_3541,N_3698);
xnor U4240 (N_4240,N_3557,N_3673);
and U4241 (N_4241,N_3697,N_3878);
or U4242 (N_4242,N_3729,N_3899);
or U4243 (N_4243,N_3653,N_3746);
xor U4244 (N_4244,N_3543,N_3724);
or U4245 (N_4245,N_3626,N_3652);
and U4246 (N_4246,N_3885,N_3630);
nand U4247 (N_4247,N_3525,N_3594);
nand U4248 (N_4248,N_3664,N_3650);
nand U4249 (N_4249,N_3699,N_3970);
or U4250 (N_4250,N_3879,N_3827);
nor U4251 (N_4251,N_3530,N_3807);
and U4252 (N_4252,N_3937,N_3646);
and U4253 (N_4253,N_3961,N_3896);
nor U4254 (N_4254,N_3836,N_3922);
nand U4255 (N_4255,N_3803,N_3636);
and U4256 (N_4256,N_3861,N_3739);
and U4257 (N_4257,N_3827,N_3672);
and U4258 (N_4258,N_3616,N_3802);
nor U4259 (N_4259,N_3582,N_3595);
nand U4260 (N_4260,N_3529,N_3769);
and U4261 (N_4261,N_3824,N_3785);
and U4262 (N_4262,N_3885,N_3838);
or U4263 (N_4263,N_3526,N_3701);
xor U4264 (N_4264,N_3560,N_3703);
and U4265 (N_4265,N_3936,N_3840);
and U4266 (N_4266,N_3812,N_3585);
or U4267 (N_4267,N_3922,N_3714);
nor U4268 (N_4268,N_3846,N_3865);
or U4269 (N_4269,N_3642,N_3682);
or U4270 (N_4270,N_3559,N_3896);
and U4271 (N_4271,N_3814,N_3620);
or U4272 (N_4272,N_3515,N_3665);
or U4273 (N_4273,N_3653,N_3940);
nor U4274 (N_4274,N_3516,N_3517);
and U4275 (N_4275,N_3526,N_3830);
or U4276 (N_4276,N_3862,N_3787);
nor U4277 (N_4277,N_3760,N_3985);
nand U4278 (N_4278,N_3836,N_3863);
nand U4279 (N_4279,N_3918,N_3508);
nor U4280 (N_4280,N_3718,N_3734);
nand U4281 (N_4281,N_3811,N_3924);
and U4282 (N_4282,N_3988,N_3687);
or U4283 (N_4283,N_3851,N_3817);
or U4284 (N_4284,N_3690,N_3698);
or U4285 (N_4285,N_3813,N_3530);
nand U4286 (N_4286,N_3869,N_3663);
nand U4287 (N_4287,N_3562,N_3923);
nand U4288 (N_4288,N_3516,N_3624);
and U4289 (N_4289,N_3711,N_3717);
nor U4290 (N_4290,N_3508,N_3775);
or U4291 (N_4291,N_3933,N_3777);
xor U4292 (N_4292,N_3894,N_3691);
and U4293 (N_4293,N_3552,N_3871);
nand U4294 (N_4294,N_3745,N_3513);
nand U4295 (N_4295,N_3769,N_3797);
nor U4296 (N_4296,N_3708,N_3915);
or U4297 (N_4297,N_3773,N_3577);
nand U4298 (N_4298,N_3681,N_3819);
and U4299 (N_4299,N_3917,N_3978);
and U4300 (N_4300,N_3779,N_3821);
nand U4301 (N_4301,N_3702,N_3563);
nand U4302 (N_4302,N_3950,N_3764);
and U4303 (N_4303,N_3930,N_3818);
nand U4304 (N_4304,N_3535,N_3618);
and U4305 (N_4305,N_3835,N_3624);
and U4306 (N_4306,N_3510,N_3885);
nor U4307 (N_4307,N_3644,N_3958);
or U4308 (N_4308,N_3778,N_3986);
and U4309 (N_4309,N_3881,N_3538);
nand U4310 (N_4310,N_3749,N_3693);
nand U4311 (N_4311,N_3719,N_3583);
and U4312 (N_4312,N_3980,N_3821);
nor U4313 (N_4313,N_3955,N_3985);
nand U4314 (N_4314,N_3727,N_3931);
nand U4315 (N_4315,N_3624,N_3790);
nor U4316 (N_4316,N_3978,N_3878);
and U4317 (N_4317,N_3756,N_3677);
or U4318 (N_4318,N_3890,N_3694);
and U4319 (N_4319,N_3614,N_3917);
and U4320 (N_4320,N_3935,N_3662);
nand U4321 (N_4321,N_3547,N_3672);
nor U4322 (N_4322,N_3838,N_3940);
nor U4323 (N_4323,N_3812,N_3779);
nor U4324 (N_4324,N_3562,N_3718);
nand U4325 (N_4325,N_3568,N_3976);
nor U4326 (N_4326,N_3552,N_3668);
nor U4327 (N_4327,N_3500,N_3539);
or U4328 (N_4328,N_3999,N_3764);
and U4329 (N_4329,N_3685,N_3912);
nand U4330 (N_4330,N_3561,N_3615);
or U4331 (N_4331,N_3907,N_3633);
and U4332 (N_4332,N_3835,N_3500);
and U4333 (N_4333,N_3900,N_3779);
and U4334 (N_4334,N_3672,N_3711);
or U4335 (N_4335,N_3543,N_3522);
nor U4336 (N_4336,N_3771,N_3864);
or U4337 (N_4337,N_3980,N_3904);
nand U4338 (N_4338,N_3741,N_3779);
and U4339 (N_4339,N_3982,N_3773);
nand U4340 (N_4340,N_3625,N_3657);
and U4341 (N_4341,N_3846,N_3963);
nand U4342 (N_4342,N_3986,N_3759);
and U4343 (N_4343,N_3693,N_3981);
and U4344 (N_4344,N_3859,N_3777);
nand U4345 (N_4345,N_3764,N_3921);
or U4346 (N_4346,N_3596,N_3788);
nor U4347 (N_4347,N_3669,N_3680);
and U4348 (N_4348,N_3641,N_3584);
nand U4349 (N_4349,N_3841,N_3819);
and U4350 (N_4350,N_3639,N_3521);
xnor U4351 (N_4351,N_3500,N_3567);
or U4352 (N_4352,N_3642,N_3620);
nor U4353 (N_4353,N_3933,N_3894);
nand U4354 (N_4354,N_3779,N_3695);
nor U4355 (N_4355,N_3724,N_3805);
nand U4356 (N_4356,N_3756,N_3732);
and U4357 (N_4357,N_3998,N_3835);
nor U4358 (N_4358,N_3549,N_3674);
or U4359 (N_4359,N_3810,N_3678);
nor U4360 (N_4360,N_3974,N_3917);
and U4361 (N_4361,N_3693,N_3516);
or U4362 (N_4362,N_3658,N_3662);
nor U4363 (N_4363,N_3605,N_3847);
xor U4364 (N_4364,N_3904,N_3819);
or U4365 (N_4365,N_3530,N_3598);
nor U4366 (N_4366,N_3811,N_3981);
nand U4367 (N_4367,N_3688,N_3889);
nand U4368 (N_4368,N_3595,N_3788);
or U4369 (N_4369,N_3563,N_3782);
and U4370 (N_4370,N_3961,N_3630);
or U4371 (N_4371,N_3656,N_3982);
and U4372 (N_4372,N_3602,N_3728);
and U4373 (N_4373,N_3783,N_3955);
nor U4374 (N_4374,N_3689,N_3988);
nor U4375 (N_4375,N_3529,N_3852);
and U4376 (N_4376,N_3950,N_3741);
nor U4377 (N_4377,N_3918,N_3853);
nor U4378 (N_4378,N_3751,N_3974);
xnor U4379 (N_4379,N_3817,N_3720);
and U4380 (N_4380,N_3799,N_3731);
nor U4381 (N_4381,N_3727,N_3772);
nand U4382 (N_4382,N_3581,N_3827);
nor U4383 (N_4383,N_3710,N_3770);
and U4384 (N_4384,N_3747,N_3792);
and U4385 (N_4385,N_3926,N_3786);
or U4386 (N_4386,N_3876,N_3522);
and U4387 (N_4387,N_3636,N_3579);
nand U4388 (N_4388,N_3878,N_3722);
nor U4389 (N_4389,N_3797,N_3981);
nand U4390 (N_4390,N_3565,N_3980);
nor U4391 (N_4391,N_3548,N_3861);
nor U4392 (N_4392,N_3778,N_3739);
xnor U4393 (N_4393,N_3921,N_3768);
or U4394 (N_4394,N_3963,N_3822);
nor U4395 (N_4395,N_3504,N_3677);
nand U4396 (N_4396,N_3607,N_3537);
nand U4397 (N_4397,N_3577,N_3706);
nand U4398 (N_4398,N_3621,N_3789);
or U4399 (N_4399,N_3613,N_3966);
nand U4400 (N_4400,N_3589,N_3817);
nand U4401 (N_4401,N_3568,N_3531);
nor U4402 (N_4402,N_3863,N_3517);
and U4403 (N_4403,N_3588,N_3629);
or U4404 (N_4404,N_3556,N_3912);
nor U4405 (N_4405,N_3924,N_3745);
xor U4406 (N_4406,N_3787,N_3501);
or U4407 (N_4407,N_3593,N_3896);
or U4408 (N_4408,N_3751,N_3645);
and U4409 (N_4409,N_3797,N_3873);
and U4410 (N_4410,N_3522,N_3966);
or U4411 (N_4411,N_3649,N_3867);
and U4412 (N_4412,N_3722,N_3874);
nor U4413 (N_4413,N_3822,N_3562);
and U4414 (N_4414,N_3678,N_3992);
nor U4415 (N_4415,N_3772,N_3877);
and U4416 (N_4416,N_3774,N_3881);
nand U4417 (N_4417,N_3583,N_3849);
nand U4418 (N_4418,N_3629,N_3724);
nand U4419 (N_4419,N_3753,N_3627);
and U4420 (N_4420,N_3956,N_3793);
and U4421 (N_4421,N_3884,N_3680);
nor U4422 (N_4422,N_3594,N_3704);
nand U4423 (N_4423,N_3870,N_3819);
or U4424 (N_4424,N_3703,N_3570);
and U4425 (N_4425,N_3625,N_3900);
nor U4426 (N_4426,N_3507,N_3800);
nor U4427 (N_4427,N_3884,N_3636);
nand U4428 (N_4428,N_3892,N_3688);
nor U4429 (N_4429,N_3615,N_3638);
nor U4430 (N_4430,N_3669,N_3735);
and U4431 (N_4431,N_3919,N_3665);
or U4432 (N_4432,N_3951,N_3942);
nand U4433 (N_4433,N_3603,N_3804);
nor U4434 (N_4434,N_3944,N_3641);
nand U4435 (N_4435,N_3917,N_3718);
nand U4436 (N_4436,N_3811,N_3653);
nand U4437 (N_4437,N_3837,N_3682);
nand U4438 (N_4438,N_3781,N_3866);
or U4439 (N_4439,N_3859,N_3529);
or U4440 (N_4440,N_3922,N_3983);
nor U4441 (N_4441,N_3757,N_3505);
and U4442 (N_4442,N_3818,N_3987);
nand U4443 (N_4443,N_3991,N_3618);
and U4444 (N_4444,N_3935,N_3595);
and U4445 (N_4445,N_3932,N_3608);
nand U4446 (N_4446,N_3697,N_3859);
or U4447 (N_4447,N_3568,N_3748);
nand U4448 (N_4448,N_3849,N_3762);
or U4449 (N_4449,N_3908,N_3553);
and U4450 (N_4450,N_3777,N_3639);
nand U4451 (N_4451,N_3573,N_3910);
nor U4452 (N_4452,N_3848,N_3912);
or U4453 (N_4453,N_3808,N_3702);
nand U4454 (N_4454,N_3929,N_3728);
nor U4455 (N_4455,N_3601,N_3524);
and U4456 (N_4456,N_3581,N_3777);
or U4457 (N_4457,N_3830,N_3815);
nand U4458 (N_4458,N_3676,N_3917);
or U4459 (N_4459,N_3775,N_3685);
nor U4460 (N_4460,N_3623,N_3985);
or U4461 (N_4461,N_3576,N_3627);
nand U4462 (N_4462,N_3529,N_3825);
nor U4463 (N_4463,N_3933,N_3587);
and U4464 (N_4464,N_3859,N_3880);
nand U4465 (N_4465,N_3537,N_3534);
nor U4466 (N_4466,N_3672,N_3645);
nand U4467 (N_4467,N_3565,N_3853);
nand U4468 (N_4468,N_3844,N_3681);
and U4469 (N_4469,N_3534,N_3766);
and U4470 (N_4470,N_3609,N_3708);
nand U4471 (N_4471,N_3751,N_3964);
and U4472 (N_4472,N_3518,N_3981);
nor U4473 (N_4473,N_3876,N_3649);
and U4474 (N_4474,N_3974,N_3685);
or U4475 (N_4475,N_3563,N_3653);
nand U4476 (N_4476,N_3816,N_3645);
xor U4477 (N_4477,N_3779,N_3865);
and U4478 (N_4478,N_3514,N_3810);
and U4479 (N_4479,N_3832,N_3855);
nor U4480 (N_4480,N_3758,N_3611);
or U4481 (N_4481,N_3630,N_3575);
or U4482 (N_4482,N_3959,N_3503);
nand U4483 (N_4483,N_3667,N_3896);
or U4484 (N_4484,N_3967,N_3740);
and U4485 (N_4485,N_3925,N_3545);
or U4486 (N_4486,N_3637,N_3709);
and U4487 (N_4487,N_3683,N_3667);
nand U4488 (N_4488,N_3558,N_3765);
nor U4489 (N_4489,N_3516,N_3839);
nand U4490 (N_4490,N_3894,N_3500);
nor U4491 (N_4491,N_3802,N_3729);
or U4492 (N_4492,N_3909,N_3845);
and U4493 (N_4493,N_3651,N_3682);
nor U4494 (N_4494,N_3603,N_3974);
or U4495 (N_4495,N_3815,N_3655);
and U4496 (N_4496,N_3964,N_3730);
or U4497 (N_4497,N_3757,N_3693);
or U4498 (N_4498,N_3847,N_3981);
and U4499 (N_4499,N_3573,N_3952);
nor U4500 (N_4500,N_4228,N_4165);
nor U4501 (N_4501,N_4101,N_4168);
or U4502 (N_4502,N_4176,N_4156);
or U4503 (N_4503,N_4230,N_4059);
nand U4504 (N_4504,N_4316,N_4409);
nor U4505 (N_4505,N_4272,N_4240);
or U4506 (N_4506,N_4390,N_4401);
nor U4507 (N_4507,N_4427,N_4103);
or U4508 (N_4508,N_4119,N_4046);
and U4509 (N_4509,N_4030,N_4471);
xor U4510 (N_4510,N_4411,N_4436);
nand U4511 (N_4511,N_4431,N_4134);
nand U4512 (N_4512,N_4155,N_4258);
nor U4513 (N_4513,N_4381,N_4294);
or U4514 (N_4514,N_4472,N_4335);
nand U4515 (N_4515,N_4445,N_4434);
nand U4516 (N_4516,N_4148,N_4279);
and U4517 (N_4517,N_4011,N_4125);
and U4518 (N_4518,N_4372,N_4102);
xnor U4519 (N_4519,N_4391,N_4211);
and U4520 (N_4520,N_4475,N_4243);
nand U4521 (N_4521,N_4301,N_4205);
and U4522 (N_4522,N_4019,N_4058);
nand U4523 (N_4523,N_4321,N_4362);
or U4524 (N_4524,N_4378,N_4139);
or U4525 (N_4525,N_4489,N_4353);
nand U4526 (N_4526,N_4450,N_4288);
nor U4527 (N_4527,N_4478,N_4226);
nand U4528 (N_4528,N_4220,N_4078);
or U4529 (N_4529,N_4157,N_4067);
or U4530 (N_4530,N_4105,N_4389);
and U4531 (N_4531,N_4474,N_4425);
and U4532 (N_4532,N_4460,N_4284);
nand U4533 (N_4533,N_4273,N_4479);
nor U4534 (N_4534,N_4376,N_4447);
or U4535 (N_4535,N_4229,N_4166);
or U4536 (N_4536,N_4051,N_4458);
nor U4537 (N_4537,N_4128,N_4412);
nor U4538 (N_4538,N_4375,N_4034);
or U4539 (N_4539,N_4063,N_4145);
nor U4540 (N_4540,N_4441,N_4295);
nand U4541 (N_4541,N_4498,N_4440);
nand U4542 (N_4542,N_4260,N_4071);
and U4543 (N_4543,N_4215,N_4363);
or U4544 (N_4544,N_4332,N_4266);
nor U4545 (N_4545,N_4488,N_4159);
or U4546 (N_4546,N_4268,N_4365);
nand U4547 (N_4547,N_4042,N_4347);
and U4548 (N_4548,N_4015,N_4449);
nand U4549 (N_4549,N_4120,N_4309);
nor U4550 (N_4550,N_4457,N_4461);
or U4551 (N_4551,N_4388,N_4278);
and U4552 (N_4552,N_4462,N_4081);
and U4553 (N_4553,N_4213,N_4257);
nor U4554 (N_4554,N_4334,N_4238);
and U4555 (N_4555,N_4031,N_4432);
and U4556 (N_4556,N_4181,N_4012);
nand U4557 (N_4557,N_4223,N_4323);
nor U4558 (N_4558,N_4056,N_4146);
nor U4559 (N_4559,N_4280,N_4190);
nor U4560 (N_4560,N_4452,N_4312);
nor U4561 (N_4561,N_4454,N_4173);
nor U4562 (N_4562,N_4355,N_4481);
and U4563 (N_4563,N_4195,N_4069);
nor U4564 (N_4564,N_4016,N_4466);
and U4565 (N_4565,N_4338,N_4027);
nor U4566 (N_4566,N_4249,N_4193);
or U4567 (N_4567,N_4467,N_4379);
and U4568 (N_4568,N_4403,N_4351);
nand U4569 (N_4569,N_4126,N_4402);
nor U4570 (N_4570,N_4065,N_4043);
and U4571 (N_4571,N_4404,N_4072);
nor U4572 (N_4572,N_4446,N_4453);
nand U4573 (N_4573,N_4331,N_4070);
nor U4574 (N_4574,N_4061,N_4209);
or U4575 (N_4575,N_4036,N_4191);
nand U4576 (N_4576,N_4340,N_4393);
nor U4577 (N_4577,N_4097,N_4261);
nor U4578 (N_4578,N_4000,N_4026);
nand U4579 (N_4579,N_4068,N_4304);
nand U4580 (N_4580,N_4368,N_4004);
nor U4581 (N_4581,N_4132,N_4217);
and U4582 (N_4582,N_4091,N_4151);
and U4583 (N_4583,N_4005,N_4109);
or U4584 (N_4584,N_4039,N_4192);
nor U4585 (N_4585,N_4199,N_4080);
and U4586 (N_4586,N_4374,N_4222);
nand U4587 (N_4587,N_4066,N_4345);
nor U4588 (N_4588,N_4326,N_4395);
or U4589 (N_4589,N_4428,N_4121);
nor U4590 (N_4590,N_4342,N_4171);
nand U4591 (N_4591,N_4003,N_4169);
nand U4592 (N_4592,N_4032,N_4164);
and U4593 (N_4593,N_4025,N_4140);
or U4594 (N_4594,N_4484,N_4253);
nor U4595 (N_4595,N_4439,N_4297);
nor U4596 (N_4596,N_4277,N_4414);
and U4597 (N_4597,N_4100,N_4406);
or U4598 (N_4598,N_4141,N_4413);
nand U4599 (N_4599,N_4341,N_4194);
or U4600 (N_4600,N_4186,N_4291);
nand U4601 (N_4601,N_4170,N_4179);
or U4602 (N_4602,N_4382,N_4408);
or U4603 (N_4603,N_4133,N_4089);
and U4604 (N_4604,N_4380,N_4189);
xnor U4605 (N_4605,N_4396,N_4269);
nor U4606 (N_4606,N_4443,N_4028);
nor U4607 (N_4607,N_4465,N_4485);
or U4608 (N_4608,N_4184,N_4469);
or U4609 (N_4609,N_4142,N_4200);
nand U4610 (N_4610,N_4442,N_4054);
and U4611 (N_4611,N_4163,N_4255);
nand U4612 (N_4612,N_4033,N_4483);
nand U4613 (N_4613,N_4429,N_4111);
or U4614 (N_4614,N_4104,N_4143);
and U4615 (N_4615,N_4468,N_4287);
nor U4616 (N_4616,N_4009,N_4496);
and U4617 (N_4617,N_4373,N_4343);
or U4618 (N_4618,N_4313,N_4399);
and U4619 (N_4619,N_4098,N_4197);
and U4620 (N_4620,N_4196,N_4346);
or U4621 (N_4621,N_4040,N_4377);
or U4622 (N_4622,N_4281,N_4292);
nand U4623 (N_4623,N_4085,N_4310);
nor U4624 (N_4624,N_4092,N_4049);
nand U4625 (N_4625,N_4497,N_4048);
and U4626 (N_4626,N_4177,N_4052);
and U4627 (N_4627,N_4094,N_4149);
and U4628 (N_4628,N_4088,N_4493);
nand U4629 (N_4629,N_4473,N_4327);
nor U4630 (N_4630,N_4053,N_4264);
xor U4631 (N_4631,N_4152,N_4250);
nor U4632 (N_4632,N_4150,N_4203);
nor U4633 (N_4633,N_4160,N_4320);
nand U4634 (N_4634,N_4010,N_4055);
xor U4635 (N_4635,N_4041,N_4114);
nand U4636 (N_4636,N_4463,N_4293);
and U4637 (N_4637,N_4419,N_4214);
or U4638 (N_4638,N_4456,N_4001);
and U4639 (N_4639,N_4083,N_4239);
and U4640 (N_4640,N_4175,N_4022);
xor U4641 (N_4641,N_4286,N_4477);
xnor U4642 (N_4642,N_4242,N_4137);
or U4643 (N_4643,N_4108,N_4337);
and U4644 (N_4644,N_4487,N_4305);
xor U4645 (N_4645,N_4259,N_4082);
or U4646 (N_4646,N_4167,N_4383);
nand U4647 (N_4647,N_4218,N_4147);
nor U4648 (N_4648,N_4117,N_4110);
nor U4649 (N_4649,N_4113,N_4495);
or U4650 (N_4650,N_4386,N_4492);
nor U4651 (N_4651,N_4020,N_4037);
and U4652 (N_4652,N_4210,N_4418);
and U4653 (N_4653,N_4002,N_4247);
nand U4654 (N_4654,N_4013,N_4023);
or U4655 (N_4655,N_4480,N_4336);
or U4656 (N_4656,N_4262,N_4017);
xor U4657 (N_4657,N_4106,N_4099);
nand U4658 (N_4658,N_4251,N_4035);
nand U4659 (N_4659,N_4322,N_4285);
nand U4660 (N_4660,N_4415,N_4241);
and U4661 (N_4661,N_4187,N_4451);
and U4662 (N_4662,N_4073,N_4127);
nor U4663 (N_4663,N_4296,N_4116);
or U4664 (N_4664,N_4158,N_4306);
nor U4665 (N_4665,N_4135,N_4317);
and U4666 (N_4666,N_4400,N_4090);
nor U4667 (N_4667,N_4499,N_4276);
or U4668 (N_4668,N_4038,N_4062);
nor U4669 (N_4669,N_4424,N_4369);
and U4670 (N_4670,N_4315,N_4221);
and U4671 (N_4671,N_4248,N_4093);
nand U4672 (N_4672,N_4314,N_4330);
nor U4673 (N_4673,N_4118,N_4459);
nor U4674 (N_4674,N_4208,N_4174);
or U4675 (N_4675,N_4282,N_4267);
or U4676 (N_4676,N_4256,N_4394);
and U4677 (N_4677,N_4339,N_4207);
or U4678 (N_4678,N_4131,N_4254);
and U4679 (N_4679,N_4201,N_4265);
or U4680 (N_4680,N_4178,N_4435);
and U4681 (N_4681,N_4245,N_4233);
nor U4682 (N_4682,N_4237,N_4044);
nand U4683 (N_4683,N_4448,N_4438);
nand U4684 (N_4684,N_4319,N_4354);
and U4685 (N_4685,N_4349,N_4324);
nor U4686 (N_4686,N_4227,N_4350);
and U4687 (N_4687,N_4057,N_4416);
and U4688 (N_4688,N_4270,N_4074);
nand U4689 (N_4689,N_4423,N_4107);
and U4690 (N_4690,N_4154,N_4482);
nor U4691 (N_4691,N_4014,N_4289);
and U4692 (N_4692,N_4444,N_4018);
or U4693 (N_4693,N_4206,N_4356);
or U4694 (N_4694,N_4318,N_4357);
nand U4695 (N_4695,N_4437,N_4311);
and U4696 (N_4696,N_4129,N_4328);
and U4697 (N_4697,N_4138,N_4172);
nand U4698 (N_4698,N_4352,N_4333);
nand U4699 (N_4699,N_4006,N_4360);
or U4700 (N_4700,N_4162,N_4244);
nand U4701 (N_4701,N_4077,N_4182);
and U4702 (N_4702,N_4366,N_4124);
nand U4703 (N_4703,N_4430,N_4290);
or U4704 (N_4704,N_4112,N_4246);
nor U4705 (N_4705,N_4422,N_4348);
nor U4706 (N_4706,N_4252,N_4325);
nand U4707 (N_4707,N_4204,N_4302);
or U4708 (N_4708,N_4476,N_4385);
and U4709 (N_4709,N_4405,N_4232);
and U4710 (N_4710,N_4299,N_4047);
or U4711 (N_4711,N_4307,N_4486);
nor U4712 (N_4712,N_4060,N_4421);
nand U4713 (N_4713,N_4216,N_4064);
or U4714 (N_4714,N_4225,N_4410);
nor U4715 (N_4715,N_4397,N_4130);
nand U4716 (N_4716,N_4426,N_4455);
or U4717 (N_4717,N_4096,N_4300);
nand U4718 (N_4718,N_4076,N_4029);
or U4719 (N_4719,N_4361,N_4231);
and U4720 (N_4720,N_4161,N_4271);
nor U4721 (N_4721,N_4274,N_4417);
or U4722 (N_4722,N_4358,N_4234);
and U4723 (N_4723,N_4235,N_4387);
and U4724 (N_4724,N_4359,N_4470);
nor U4725 (N_4725,N_4370,N_4144);
or U4726 (N_4726,N_4398,N_4153);
and U4727 (N_4727,N_4263,N_4050);
nor U4728 (N_4728,N_4123,N_4185);
nor U4729 (N_4729,N_4087,N_4007);
nor U4730 (N_4730,N_4188,N_4183);
nor U4731 (N_4731,N_4298,N_4420);
nor U4732 (N_4732,N_4008,N_4079);
or U4733 (N_4733,N_4371,N_4086);
xnor U4734 (N_4734,N_4024,N_4115);
or U4735 (N_4735,N_4224,N_4198);
and U4736 (N_4736,N_4308,N_4491);
nor U4737 (N_4737,N_4384,N_4202);
nor U4738 (N_4738,N_4344,N_4494);
and U4739 (N_4739,N_4021,N_4219);
and U4740 (N_4740,N_4490,N_4180);
or U4741 (N_4741,N_4433,N_4236);
nor U4742 (N_4742,N_4095,N_4407);
nand U4743 (N_4743,N_4329,N_4075);
nand U4744 (N_4744,N_4367,N_4084);
xnor U4745 (N_4745,N_4303,N_4275);
or U4746 (N_4746,N_4045,N_4392);
nand U4747 (N_4747,N_4464,N_4122);
and U4748 (N_4748,N_4283,N_4364);
nor U4749 (N_4749,N_4212,N_4136);
nand U4750 (N_4750,N_4092,N_4034);
nand U4751 (N_4751,N_4174,N_4013);
or U4752 (N_4752,N_4325,N_4277);
nor U4753 (N_4753,N_4170,N_4069);
and U4754 (N_4754,N_4325,N_4033);
nand U4755 (N_4755,N_4010,N_4232);
nand U4756 (N_4756,N_4333,N_4305);
xor U4757 (N_4757,N_4290,N_4439);
nor U4758 (N_4758,N_4498,N_4116);
nor U4759 (N_4759,N_4336,N_4264);
and U4760 (N_4760,N_4310,N_4472);
or U4761 (N_4761,N_4425,N_4121);
and U4762 (N_4762,N_4178,N_4174);
nand U4763 (N_4763,N_4424,N_4408);
or U4764 (N_4764,N_4213,N_4333);
and U4765 (N_4765,N_4263,N_4290);
or U4766 (N_4766,N_4045,N_4110);
and U4767 (N_4767,N_4471,N_4209);
or U4768 (N_4768,N_4488,N_4155);
xnor U4769 (N_4769,N_4271,N_4440);
nor U4770 (N_4770,N_4226,N_4157);
nand U4771 (N_4771,N_4380,N_4462);
or U4772 (N_4772,N_4240,N_4477);
and U4773 (N_4773,N_4001,N_4269);
nor U4774 (N_4774,N_4097,N_4073);
or U4775 (N_4775,N_4323,N_4232);
or U4776 (N_4776,N_4459,N_4031);
nand U4777 (N_4777,N_4305,N_4456);
and U4778 (N_4778,N_4047,N_4102);
nand U4779 (N_4779,N_4028,N_4099);
nor U4780 (N_4780,N_4266,N_4363);
nor U4781 (N_4781,N_4314,N_4184);
nand U4782 (N_4782,N_4073,N_4322);
or U4783 (N_4783,N_4210,N_4144);
or U4784 (N_4784,N_4336,N_4153);
xnor U4785 (N_4785,N_4253,N_4025);
and U4786 (N_4786,N_4037,N_4321);
nor U4787 (N_4787,N_4001,N_4049);
nor U4788 (N_4788,N_4259,N_4005);
or U4789 (N_4789,N_4268,N_4494);
nor U4790 (N_4790,N_4441,N_4152);
or U4791 (N_4791,N_4215,N_4188);
nand U4792 (N_4792,N_4155,N_4256);
nor U4793 (N_4793,N_4106,N_4223);
nor U4794 (N_4794,N_4245,N_4374);
nor U4795 (N_4795,N_4257,N_4300);
xnor U4796 (N_4796,N_4111,N_4401);
or U4797 (N_4797,N_4360,N_4213);
nand U4798 (N_4798,N_4386,N_4280);
nand U4799 (N_4799,N_4220,N_4311);
and U4800 (N_4800,N_4125,N_4266);
nor U4801 (N_4801,N_4261,N_4293);
and U4802 (N_4802,N_4035,N_4287);
and U4803 (N_4803,N_4446,N_4162);
or U4804 (N_4804,N_4369,N_4444);
or U4805 (N_4805,N_4056,N_4175);
or U4806 (N_4806,N_4281,N_4410);
nand U4807 (N_4807,N_4306,N_4090);
and U4808 (N_4808,N_4431,N_4214);
and U4809 (N_4809,N_4099,N_4049);
and U4810 (N_4810,N_4124,N_4203);
and U4811 (N_4811,N_4214,N_4420);
nand U4812 (N_4812,N_4081,N_4291);
nand U4813 (N_4813,N_4323,N_4246);
or U4814 (N_4814,N_4007,N_4116);
nand U4815 (N_4815,N_4301,N_4036);
nor U4816 (N_4816,N_4274,N_4375);
and U4817 (N_4817,N_4367,N_4096);
nor U4818 (N_4818,N_4296,N_4436);
or U4819 (N_4819,N_4448,N_4087);
nand U4820 (N_4820,N_4441,N_4196);
nor U4821 (N_4821,N_4264,N_4207);
and U4822 (N_4822,N_4352,N_4047);
nand U4823 (N_4823,N_4340,N_4209);
xor U4824 (N_4824,N_4350,N_4495);
nand U4825 (N_4825,N_4196,N_4078);
and U4826 (N_4826,N_4262,N_4498);
nor U4827 (N_4827,N_4274,N_4142);
xor U4828 (N_4828,N_4257,N_4194);
and U4829 (N_4829,N_4313,N_4015);
nand U4830 (N_4830,N_4212,N_4132);
and U4831 (N_4831,N_4092,N_4014);
and U4832 (N_4832,N_4258,N_4221);
nand U4833 (N_4833,N_4185,N_4446);
nor U4834 (N_4834,N_4260,N_4023);
nand U4835 (N_4835,N_4283,N_4326);
or U4836 (N_4836,N_4279,N_4327);
nor U4837 (N_4837,N_4422,N_4423);
or U4838 (N_4838,N_4401,N_4291);
or U4839 (N_4839,N_4454,N_4232);
nand U4840 (N_4840,N_4438,N_4246);
nand U4841 (N_4841,N_4469,N_4392);
or U4842 (N_4842,N_4001,N_4462);
nand U4843 (N_4843,N_4451,N_4335);
nand U4844 (N_4844,N_4489,N_4068);
nor U4845 (N_4845,N_4262,N_4479);
or U4846 (N_4846,N_4032,N_4491);
nand U4847 (N_4847,N_4266,N_4426);
nand U4848 (N_4848,N_4059,N_4017);
or U4849 (N_4849,N_4040,N_4296);
nand U4850 (N_4850,N_4348,N_4372);
xor U4851 (N_4851,N_4005,N_4225);
nand U4852 (N_4852,N_4195,N_4319);
nand U4853 (N_4853,N_4326,N_4253);
nor U4854 (N_4854,N_4287,N_4233);
or U4855 (N_4855,N_4336,N_4248);
xor U4856 (N_4856,N_4491,N_4315);
and U4857 (N_4857,N_4321,N_4158);
xnor U4858 (N_4858,N_4254,N_4186);
nor U4859 (N_4859,N_4264,N_4243);
and U4860 (N_4860,N_4206,N_4258);
nand U4861 (N_4861,N_4223,N_4280);
or U4862 (N_4862,N_4183,N_4320);
nand U4863 (N_4863,N_4371,N_4199);
or U4864 (N_4864,N_4187,N_4264);
or U4865 (N_4865,N_4231,N_4472);
nor U4866 (N_4866,N_4412,N_4337);
and U4867 (N_4867,N_4164,N_4095);
or U4868 (N_4868,N_4272,N_4139);
or U4869 (N_4869,N_4144,N_4199);
nor U4870 (N_4870,N_4118,N_4148);
nand U4871 (N_4871,N_4407,N_4011);
or U4872 (N_4872,N_4470,N_4177);
or U4873 (N_4873,N_4363,N_4271);
nand U4874 (N_4874,N_4414,N_4056);
nor U4875 (N_4875,N_4118,N_4067);
nor U4876 (N_4876,N_4473,N_4446);
nor U4877 (N_4877,N_4037,N_4153);
nor U4878 (N_4878,N_4230,N_4042);
nor U4879 (N_4879,N_4307,N_4208);
nand U4880 (N_4880,N_4242,N_4483);
nor U4881 (N_4881,N_4139,N_4478);
and U4882 (N_4882,N_4364,N_4339);
nand U4883 (N_4883,N_4172,N_4204);
nor U4884 (N_4884,N_4309,N_4237);
and U4885 (N_4885,N_4001,N_4149);
and U4886 (N_4886,N_4019,N_4317);
nor U4887 (N_4887,N_4320,N_4292);
and U4888 (N_4888,N_4155,N_4192);
nand U4889 (N_4889,N_4176,N_4422);
xor U4890 (N_4890,N_4059,N_4181);
or U4891 (N_4891,N_4069,N_4051);
nor U4892 (N_4892,N_4284,N_4133);
and U4893 (N_4893,N_4030,N_4003);
nand U4894 (N_4894,N_4049,N_4267);
and U4895 (N_4895,N_4399,N_4116);
and U4896 (N_4896,N_4477,N_4136);
and U4897 (N_4897,N_4114,N_4079);
nor U4898 (N_4898,N_4452,N_4329);
xor U4899 (N_4899,N_4256,N_4444);
nand U4900 (N_4900,N_4234,N_4298);
nand U4901 (N_4901,N_4092,N_4295);
nor U4902 (N_4902,N_4037,N_4124);
or U4903 (N_4903,N_4414,N_4122);
nand U4904 (N_4904,N_4379,N_4410);
xnor U4905 (N_4905,N_4468,N_4497);
nor U4906 (N_4906,N_4498,N_4114);
nand U4907 (N_4907,N_4104,N_4173);
and U4908 (N_4908,N_4201,N_4075);
or U4909 (N_4909,N_4069,N_4074);
or U4910 (N_4910,N_4441,N_4331);
nor U4911 (N_4911,N_4238,N_4269);
nand U4912 (N_4912,N_4234,N_4405);
and U4913 (N_4913,N_4165,N_4039);
and U4914 (N_4914,N_4153,N_4327);
and U4915 (N_4915,N_4421,N_4191);
and U4916 (N_4916,N_4257,N_4083);
or U4917 (N_4917,N_4004,N_4043);
and U4918 (N_4918,N_4269,N_4368);
nor U4919 (N_4919,N_4167,N_4071);
nor U4920 (N_4920,N_4272,N_4234);
or U4921 (N_4921,N_4304,N_4278);
and U4922 (N_4922,N_4360,N_4428);
nor U4923 (N_4923,N_4489,N_4461);
or U4924 (N_4924,N_4271,N_4149);
and U4925 (N_4925,N_4260,N_4217);
nand U4926 (N_4926,N_4128,N_4170);
and U4927 (N_4927,N_4339,N_4371);
nor U4928 (N_4928,N_4413,N_4351);
and U4929 (N_4929,N_4393,N_4272);
nand U4930 (N_4930,N_4480,N_4036);
and U4931 (N_4931,N_4276,N_4317);
and U4932 (N_4932,N_4305,N_4329);
or U4933 (N_4933,N_4443,N_4032);
and U4934 (N_4934,N_4236,N_4448);
nand U4935 (N_4935,N_4130,N_4304);
nand U4936 (N_4936,N_4236,N_4383);
or U4937 (N_4937,N_4005,N_4480);
and U4938 (N_4938,N_4352,N_4190);
nand U4939 (N_4939,N_4433,N_4101);
and U4940 (N_4940,N_4422,N_4379);
nand U4941 (N_4941,N_4464,N_4409);
or U4942 (N_4942,N_4375,N_4384);
or U4943 (N_4943,N_4045,N_4101);
xnor U4944 (N_4944,N_4099,N_4247);
or U4945 (N_4945,N_4154,N_4349);
nor U4946 (N_4946,N_4291,N_4197);
nor U4947 (N_4947,N_4219,N_4264);
and U4948 (N_4948,N_4412,N_4145);
nor U4949 (N_4949,N_4322,N_4405);
and U4950 (N_4950,N_4235,N_4369);
nand U4951 (N_4951,N_4150,N_4125);
or U4952 (N_4952,N_4475,N_4012);
or U4953 (N_4953,N_4383,N_4353);
and U4954 (N_4954,N_4251,N_4052);
and U4955 (N_4955,N_4348,N_4439);
and U4956 (N_4956,N_4131,N_4006);
and U4957 (N_4957,N_4119,N_4148);
nand U4958 (N_4958,N_4336,N_4086);
nor U4959 (N_4959,N_4068,N_4234);
and U4960 (N_4960,N_4332,N_4292);
nor U4961 (N_4961,N_4134,N_4397);
nand U4962 (N_4962,N_4400,N_4003);
or U4963 (N_4963,N_4396,N_4244);
or U4964 (N_4964,N_4454,N_4083);
nor U4965 (N_4965,N_4446,N_4442);
nand U4966 (N_4966,N_4289,N_4283);
nor U4967 (N_4967,N_4048,N_4046);
nand U4968 (N_4968,N_4092,N_4191);
or U4969 (N_4969,N_4457,N_4185);
nand U4970 (N_4970,N_4125,N_4464);
or U4971 (N_4971,N_4497,N_4064);
nor U4972 (N_4972,N_4402,N_4180);
or U4973 (N_4973,N_4066,N_4154);
nand U4974 (N_4974,N_4431,N_4149);
nor U4975 (N_4975,N_4372,N_4451);
nand U4976 (N_4976,N_4259,N_4443);
nand U4977 (N_4977,N_4491,N_4312);
and U4978 (N_4978,N_4235,N_4357);
nand U4979 (N_4979,N_4174,N_4033);
and U4980 (N_4980,N_4408,N_4292);
nand U4981 (N_4981,N_4301,N_4160);
or U4982 (N_4982,N_4165,N_4408);
or U4983 (N_4983,N_4415,N_4458);
xnor U4984 (N_4984,N_4315,N_4314);
or U4985 (N_4985,N_4308,N_4274);
nand U4986 (N_4986,N_4370,N_4017);
nor U4987 (N_4987,N_4401,N_4451);
nor U4988 (N_4988,N_4032,N_4362);
and U4989 (N_4989,N_4433,N_4000);
and U4990 (N_4990,N_4177,N_4104);
or U4991 (N_4991,N_4461,N_4253);
or U4992 (N_4992,N_4251,N_4217);
and U4993 (N_4993,N_4477,N_4188);
nand U4994 (N_4994,N_4222,N_4409);
and U4995 (N_4995,N_4244,N_4315);
and U4996 (N_4996,N_4114,N_4292);
or U4997 (N_4997,N_4086,N_4077);
or U4998 (N_4998,N_4051,N_4327);
or U4999 (N_4999,N_4486,N_4452);
or UO_0 (O_0,N_4910,N_4942);
nand UO_1 (O_1,N_4861,N_4882);
and UO_2 (O_2,N_4961,N_4676);
nor UO_3 (O_3,N_4598,N_4839);
or UO_4 (O_4,N_4774,N_4565);
nand UO_5 (O_5,N_4878,N_4706);
xnor UO_6 (O_6,N_4502,N_4743);
nand UO_7 (O_7,N_4896,N_4843);
xor UO_8 (O_8,N_4507,N_4891);
nor UO_9 (O_9,N_4504,N_4958);
xnor UO_10 (O_10,N_4576,N_4629);
nand UO_11 (O_11,N_4543,N_4756);
and UO_12 (O_12,N_4711,N_4990);
nor UO_13 (O_13,N_4523,N_4768);
nand UO_14 (O_14,N_4590,N_4541);
or UO_15 (O_15,N_4944,N_4763);
or UO_16 (O_16,N_4716,N_4638);
nor UO_17 (O_17,N_4617,N_4951);
nand UO_18 (O_18,N_4644,N_4677);
or UO_19 (O_19,N_4783,N_4694);
nor UO_20 (O_20,N_4559,N_4776);
or UO_21 (O_21,N_4745,N_4720);
or UO_22 (O_22,N_4691,N_4948);
and UO_23 (O_23,N_4815,N_4957);
and UO_24 (O_24,N_4669,N_4719);
or UO_25 (O_25,N_4715,N_4589);
nand UO_26 (O_26,N_4821,N_4905);
and UO_27 (O_27,N_4764,N_4618);
nor UO_28 (O_28,N_4608,N_4980);
nor UO_29 (O_29,N_4784,N_4655);
nand UO_30 (O_30,N_4521,N_4533);
nand UO_31 (O_31,N_4788,N_4965);
nand UO_32 (O_32,N_4793,N_4832);
nand UO_33 (O_33,N_4562,N_4828);
nand UO_34 (O_34,N_4888,N_4561);
or UO_35 (O_35,N_4983,N_4846);
nor UO_36 (O_36,N_4600,N_4702);
or UO_37 (O_37,N_4883,N_4982);
nor UO_38 (O_38,N_4831,N_4588);
nor UO_39 (O_39,N_4704,N_4989);
nor UO_40 (O_40,N_4761,N_4824);
nor UO_41 (O_41,N_4940,N_4722);
or UO_42 (O_42,N_4605,N_4673);
nor UO_43 (O_43,N_4963,N_4500);
and UO_44 (O_44,N_4640,N_4651);
and UO_45 (O_45,N_4795,N_4757);
or UO_46 (O_46,N_4852,N_4628);
and UO_47 (O_47,N_4712,N_4721);
and UO_48 (O_48,N_4515,N_4741);
or UO_49 (O_49,N_4614,N_4875);
nand UO_50 (O_50,N_4700,N_4976);
and UO_51 (O_51,N_4975,N_4789);
xor UO_52 (O_52,N_4501,N_4879);
nand UO_53 (O_53,N_4890,N_4800);
and UO_54 (O_54,N_4916,N_4857);
nor UO_55 (O_55,N_4556,N_4529);
and UO_56 (O_56,N_4863,N_4670);
and UO_57 (O_57,N_4886,N_4796);
and UO_58 (O_58,N_4946,N_4920);
and UO_59 (O_59,N_4518,N_4934);
nand UO_60 (O_60,N_4889,N_4953);
nand UO_61 (O_61,N_4892,N_4802);
and UO_62 (O_62,N_4558,N_4530);
and UO_63 (O_63,N_4850,N_4977);
and UO_64 (O_64,N_4750,N_4936);
or UO_65 (O_65,N_4578,N_4675);
nand UO_66 (O_66,N_4729,N_4632);
or UO_67 (O_67,N_4820,N_4767);
nor UO_68 (O_68,N_4667,N_4639);
or UO_69 (O_69,N_4775,N_4622);
xnor UO_70 (O_70,N_4998,N_4973);
nand UO_71 (O_71,N_4734,N_4709);
nor UO_72 (O_72,N_4952,N_4621);
nand UO_73 (O_73,N_4927,N_4563);
nand UO_74 (O_74,N_4587,N_4781);
or UO_75 (O_75,N_4897,N_4739);
nor UO_76 (O_76,N_4812,N_4705);
nor UO_77 (O_77,N_4917,N_4898);
or UO_78 (O_78,N_4935,N_4817);
nand UO_79 (O_79,N_4754,N_4791);
or UO_80 (O_80,N_4746,N_4527);
or UO_81 (O_81,N_4553,N_4580);
nor UO_82 (O_82,N_4735,N_4698);
nor UO_83 (O_83,N_4923,N_4645);
nor UO_84 (O_84,N_4868,N_4924);
and UO_85 (O_85,N_4506,N_4760);
and UO_86 (O_86,N_4713,N_4780);
or UO_87 (O_87,N_4751,N_4841);
nor UO_88 (O_88,N_4851,N_4929);
or UO_89 (O_89,N_4634,N_4664);
and UO_90 (O_90,N_4803,N_4642);
nand UO_91 (O_91,N_4593,N_4604);
nor UO_92 (O_92,N_4742,N_4571);
nand UO_93 (O_93,N_4643,N_4818);
nand UO_94 (O_94,N_4876,N_4695);
or UO_95 (O_95,N_4822,N_4960);
nand UO_96 (O_96,N_4583,N_4657);
nand UO_97 (O_97,N_4860,N_4652);
nor UO_98 (O_98,N_4845,N_4922);
nand UO_99 (O_99,N_4869,N_4591);
or UO_100 (O_100,N_4955,N_4894);
nor UO_101 (O_101,N_4992,N_4972);
nand UO_102 (O_102,N_4988,N_4524);
or UO_103 (O_103,N_4690,N_4904);
or UO_104 (O_104,N_4597,N_4925);
and UO_105 (O_105,N_4727,N_4833);
nand UO_106 (O_106,N_4542,N_4577);
nand UO_107 (O_107,N_4752,N_4686);
and UO_108 (O_108,N_4707,N_4999);
nor UO_109 (O_109,N_4732,N_4679);
nand UO_110 (O_110,N_4870,N_4648);
nor UO_111 (O_111,N_4551,N_4807);
and UO_112 (O_112,N_4726,N_4612);
or UO_113 (O_113,N_4625,N_4819);
nor UO_114 (O_114,N_4848,N_4699);
and UO_115 (O_115,N_4666,N_4725);
or UO_116 (O_116,N_4596,N_4684);
nand UO_117 (O_117,N_4792,N_4979);
nand UO_118 (O_118,N_4912,N_4616);
nand UO_119 (O_119,N_4785,N_4908);
nand UO_120 (O_120,N_4872,N_4575);
and UO_121 (O_121,N_4855,N_4615);
nand UO_122 (O_122,N_4717,N_4685);
nand UO_123 (O_123,N_4613,N_4826);
or UO_124 (O_124,N_4810,N_4835);
and UO_125 (O_125,N_4602,N_4765);
nand UO_126 (O_126,N_4997,N_4987);
or UO_127 (O_127,N_4801,N_4816);
or UO_128 (O_128,N_4755,N_4599);
nand UO_129 (O_129,N_4630,N_4748);
and UO_130 (O_130,N_4641,N_4962);
nor UO_131 (O_131,N_4656,N_4631);
nor UO_132 (O_132,N_4862,N_4730);
or UO_133 (O_133,N_4737,N_4660);
or UO_134 (O_134,N_4964,N_4692);
or UO_135 (O_135,N_4881,N_4659);
or UO_136 (O_136,N_4689,N_4526);
xor UO_137 (O_137,N_4856,N_4938);
or UO_138 (O_138,N_4967,N_4701);
nand UO_139 (O_139,N_4736,N_4688);
and UO_140 (O_140,N_4672,N_4546);
nor UO_141 (O_141,N_4681,N_4581);
and UO_142 (O_142,N_4762,N_4865);
and UO_143 (O_143,N_4528,N_4867);
nor UO_144 (O_144,N_4647,N_4753);
and UO_145 (O_145,N_4624,N_4646);
or UO_146 (O_146,N_4520,N_4805);
nand UO_147 (O_147,N_4509,N_4813);
nand UO_148 (O_148,N_4537,N_4584);
or UO_149 (O_149,N_4930,N_4594);
or UO_150 (O_150,N_4663,N_4683);
or UO_151 (O_151,N_4579,N_4510);
nor UO_152 (O_152,N_4902,N_4947);
nor UO_153 (O_153,N_4895,N_4610);
nand UO_154 (O_154,N_4971,N_4877);
nor UO_155 (O_155,N_4939,N_4758);
and UO_156 (O_156,N_4539,N_4569);
or UO_157 (O_157,N_4519,N_4635);
nor UO_158 (O_158,N_4834,N_4859);
nand UO_159 (O_159,N_4601,N_4858);
nor UO_160 (O_160,N_4728,N_4586);
nand UO_161 (O_161,N_4825,N_4738);
nor UO_162 (O_162,N_4811,N_4931);
nand UO_163 (O_163,N_4844,N_4836);
and UO_164 (O_164,N_4880,N_4668);
nor UO_165 (O_165,N_4847,N_4918);
nand UO_166 (O_166,N_4854,N_4933);
nor UO_167 (O_167,N_4654,N_4874);
xnor UO_168 (O_168,N_4724,N_4945);
and UO_169 (O_169,N_4550,N_4840);
nand UO_170 (O_170,N_4514,N_4978);
and UO_171 (O_171,N_4516,N_4970);
and UO_172 (O_172,N_4779,N_4680);
xor UO_173 (O_173,N_4928,N_4693);
nand UO_174 (O_174,N_4566,N_4603);
nand UO_175 (O_175,N_4585,N_4560);
nand UO_176 (O_176,N_4993,N_4592);
xnor UO_177 (O_177,N_4544,N_4909);
or UO_178 (O_178,N_4708,N_4564);
nor UO_179 (O_179,N_4653,N_4658);
and UO_180 (O_180,N_4773,N_4893);
xnor UO_181 (O_181,N_4532,N_4797);
and UO_182 (O_182,N_4540,N_4505);
nand UO_183 (O_183,N_4574,N_4759);
or UO_184 (O_184,N_4986,N_4853);
nand UO_185 (O_185,N_4513,N_4956);
nor UO_186 (O_186,N_4770,N_4567);
and UO_187 (O_187,N_4536,N_4919);
nor UO_188 (O_188,N_4508,N_4548);
xor UO_189 (O_189,N_4549,N_4913);
and UO_190 (O_190,N_4786,N_4678);
nand UO_191 (O_191,N_4838,N_4906);
nor UO_192 (O_192,N_4782,N_4790);
and UO_193 (O_193,N_4723,N_4899);
nor UO_194 (O_194,N_4921,N_4718);
nand UO_195 (O_195,N_4837,N_4914);
nor UO_196 (O_196,N_4557,N_4649);
nor UO_197 (O_197,N_4627,N_4950);
or UO_198 (O_198,N_4849,N_4827);
or UO_199 (O_199,N_4554,N_4573);
nand UO_200 (O_200,N_4512,N_4814);
nor UO_201 (O_201,N_4799,N_4703);
and UO_202 (O_202,N_4682,N_4984);
nor UO_203 (O_203,N_4766,N_4772);
or UO_204 (O_204,N_4864,N_4937);
nor UO_205 (O_205,N_4996,N_4661);
nor UO_206 (O_206,N_4995,N_4626);
nor UO_207 (O_207,N_4915,N_4687);
or UO_208 (O_208,N_4941,N_4787);
or UO_209 (O_209,N_4525,N_4674);
and UO_210 (O_210,N_4974,N_4830);
or UO_211 (O_211,N_4985,N_4749);
and UO_212 (O_212,N_4884,N_4620);
nor UO_213 (O_213,N_4733,N_4968);
nand UO_214 (O_214,N_4804,N_4991);
nor UO_215 (O_215,N_4954,N_4901);
nor UO_216 (O_216,N_4769,N_4606);
and UO_217 (O_217,N_4966,N_4871);
nand UO_218 (O_218,N_4623,N_4932);
or UO_219 (O_219,N_4545,N_4650);
or UO_220 (O_220,N_4531,N_4959);
nand UO_221 (O_221,N_4842,N_4911);
or UO_222 (O_222,N_4926,N_4794);
or UO_223 (O_223,N_4873,N_4777);
or UO_224 (O_224,N_4696,N_4535);
nor UO_225 (O_225,N_4697,N_4503);
or UO_226 (O_226,N_4517,N_4747);
or UO_227 (O_227,N_4636,N_4714);
nand UO_228 (O_228,N_4744,N_4903);
nor UO_229 (O_229,N_4637,N_4710);
and UO_230 (O_230,N_4522,N_4609);
nor UO_231 (O_231,N_4943,N_4595);
and UO_232 (O_232,N_4534,N_4607);
nor UO_233 (O_233,N_4823,N_4572);
or UO_234 (O_234,N_4552,N_4887);
or UO_235 (O_235,N_4885,N_4778);
nor UO_236 (O_236,N_4671,N_4829);
or UO_237 (O_237,N_4555,N_4981);
nand UO_238 (O_238,N_4633,N_4866);
nand UO_239 (O_239,N_4582,N_4740);
and UO_240 (O_240,N_4511,N_4619);
nand UO_241 (O_241,N_4662,N_4907);
and UO_242 (O_242,N_4665,N_4611);
nand UO_243 (O_243,N_4771,N_4969);
and UO_244 (O_244,N_4547,N_4949);
or UO_245 (O_245,N_4900,N_4568);
xnor UO_246 (O_246,N_4806,N_4808);
nor UO_247 (O_247,N_4570,N_4994);
and UO_248 (O_248,N_4798,N_4731);
nor UO_249 (O_249,N_4809,N_4538);
or UO_250 (O_250,N_4856,N_4916);
and UO_251 (O_251,N_4514,N_4628);
nand UO_252 (O_252,N_4859,N_4801);
nor UO_253 (O_253,N_4772,N_4510);
nor UO_254 (O_254,N_4943,N_4616);
nand UO_255 (O_255,N_4862,N_4826);
and UO_256 (O_256,N_4983,N_4833);
and UO_257 (O_257,N_4903,N_4926);
or UO_258 (O_258,N_4828,N_4730);
nor UO_259 (O_259,N_4513,N_4954);
or UO_260 (O_260,N_4797,N_4510);
and UO_261 (O_261,N_4748,N_4524);
nor UO_262 (O_262,N_4770,N_4582);
and UO_263 (O_263,N_4984,N_4636);
nor UO_264 (O_264,N_4524,N_4662);
or UO_265 (O_265,N_4771,N_4615);
or UO_266 (O_266,N_4604,N_4737);
nor UO_267 (O_267,N_4625,N_4707);
nor UO_268 (O_268,N_4745,N_4948);
and UO_269 (O_269,N_4754,N_4818);
nand UO_270 (O_270,N_4689,N_4606);
xnor UO_271 (O_271,N_4853,N_4921);
or UO_272 (O_272,N_4515,N_4560);
and UO_273 (O_273,N_4754,N_4738);
nand UO_274 (O_274,N_4549,N_4697);
or UO_275 (O_275,N_4530,N_4705);
and UO_276 (O_276,N_4812,N_4998);
xnor UO_277 (O_277,N_4876,N_4636);
or UO_278 (O_278,N_4801,N_4817);
or UO_279 (O_279,N_4666,N_4842);
nor UO_280 (O_280,N_4767,N_4722);
xnor UO_281 (O_281,N_4726,N_4731);
nand UO_282 (O_282,N_4533,N_4837);
nor UO_283 (O_283,N_4640,N_4558);
nand UO_284 (O_284,N_4809,N_4623);
nor UO_285 (O_285,N_4892,N_4794);
and UO_286 (O_286,N_4933,N_4904);
nor UO_287 (O_287,N_4798,N_4581);
and UO_288 (O_288,N_4873,N_4756);
or UO_289 (O_289,N_4686,N_4888);
or UO_290 (O_290,N_4780,N_4821);
and UO_291 (O_291,N_4990,N_4572);
or UO_292 (O_292,N_4785,N_4643);
nor UO_293 (O_293,N_4968,N_4949);
nor UO_294 (O_294,N_4711,N_4892);
nand UO_295 (O_295,N_4748,N_4805);
and UO_296 (O_296,N_4709,N_4644);
nand UO_297 (O_297,N_4883,N_4847);
nor UO_298 (O_298,N_4944,N_4888);
and UO_299 (O_299,N_4980,N_4563);
or UO_300 (O_300,N_4770,N_4577);
nand UO_301 (O_301,N_4903,N_4604);
nand UO_302 (O_302,N_4784,N_4848);
nor UO_303 (O_303,N_4816,N_4583);
or UO_304 (O_304,N_4943,N_4979);
nand UO_305 (O_305,N_4580,N_4543);
and UO_306 (O_306,N_4912,N_4690);
or UO_307 (O_307,N_4859,N_4588);
nand UO_308 (O_308,N_4870,N_4936);
and UO_309 (O_309,N_4923,N_4608);
nor UO_310 (O_310,N_4999,N_4892);
and UO_311 (O_311,N_4678,N_4672);
nand UO_312 (O_312,N_4511,N_4729);
nand UO_313 (O_313,N_4529,N_4504);
and UO_314 (O_314,N_4542,N_4995);
nand UO_315 (O_315,N_4597,N_4722);
and UO_316 (O_316,N_4639,N_4700);
and UO_317 (O_317,N_4762,N_4868);
nand UO_318 (O_318,N_4804,N_4529);
xnor UO_319 (O_319,N_4945,N_4978);
nand UO_320 (O_320,N_4788,N_4937);
xor UO_321 (O_321,N_4640,N_4993);
and UO_322 (O_322,N_4868,N_4572);
or UO_323 (O_323,N_4878,N_4912);
and UO_324 (O_324,N_4908,N_4844);
and UO_325 (O_325,N_4783,N_4946);
and UO_326 (O_326,N_4757,N_4718);
nand UO_327 (O_327,N_4903,N_4997);
and UO_328 (O_328,N_4521,N_4751);
nand UO_329 (O_329,N_4698,N_4983);
and UO_330 (O_330,N_4545,N_4961);
or UO_331 (O_331,N_4631,N_4822);
nand UO_332 (O_332,N_4564,N_4982);
or UO_333 (O_333,N_4705,N_4753);
nand UO_334 (O_334,N_4853,N_4741);
nor UO_335 (O_335,N_4765,N_4816);
nor UO_336 (O_336,N_4859,N_4881);
and UO_337 (O_337,N_4630,N_4977);
and UO_338 (O_338,N_4705,N_4622);
and UO_339 (O_339,N_4604,N_4556);
nor UO_340 (O_340,N_4791,N_4787);
or UO_341 (O_341,N_4659,N_4809);
nor UO_342 (O_342,N_4740,N_4856);
and UO_343 (O_343,N_4615,N_4533);
and UO_344 (O_344,N_4574,N_4993);
nand UO_345 (O_345,N_4568,N_4631);
and UO_346 (O_346,N_4625,N_4658);
nor UO_347 (O_347,N_4563,N_4973);
or UO_348 (O_348,N_4552,N_4744);
nand UO_349 (O_349,N_4746,N_4500);
or UO_350 (O_350,N_4616,N_4509);
nand UO_351 (O_351,N_4881,N_4549);
and UO_352 (O_352,N_4809,N_4951);
nand UO_353 (O_353,N_4516,N_4507);
nand UO_354 (O_354,N_4737,N_4745);
nand UO_355 (O_355,N_4775,N_4644);
and UO_356 (O_356,N_4985,N_4739);
or UO_357 (O_357,N_4794,N_4612);
nor UO_358 (O_358,N_4827,N_4873);
nand UO_359 (O_359,N_4534,N_4904);
nor UO_360 (O_360,N_4876,N_4875);
and UO_361 (O_361,N_4731,N_4969);
nand UO_362 (O_362,N_4869,N_4998);
nand UO_363 (O_363,N_4745,N_4777);
nor UO_364 (O_364,N_4744,N_4772);
or UO_365 (O_365,N_4668,N_4732);
and UO_366 (O_366,N_4908,N_4569);
or UO_367 (O_367,N_4554,N_4760);
nor UO_368 (O_368,N_4984,N_4822);
and UO_369 (O_369,N_4788,N_4672);
or UO_370 (O_370,N_4959,N_4951);
or UO_371 (O_371,N_4659,N_4642);
nand UO_372 (O_372,N_4563,N_4718);
or UO_373 (O_373,N_4590,N_4651);
and UO_374 (O_374,N_4842,N_4740);
or UO_375 (O_375,N_4699,N_4855);
or UO_376 (O_376,N_4805,N_4921);
and UO_377 (O_377,N_4820,N_4544);
or UO_378 (O_378,N_4775,N_4669);
nand UO_379 (O_379,N_4883,N_4513);
nand UO_380 (O_380,N_4825,N_4786);
nand UO_381 (O_381,N_4956,N_4692);
nand UO_382 (O_382,N_4500,N_4894);
nand UO_383 (O_383,N_4855,N_4585);
or UO_384 (O_384,N_4543,N_4815);
nand UO_385 (O_385,N_4671,N_4780);
nand UO_386 (O_386,N_4973,N_4735);
or UO_387 (O_387,N_4749,N_4868);
nor UO_388 (O_388,N_4659,N_4748);
nand UO_389 (O_389,N_4572,N_4517);
nand UO_390 (O_390,N_4951,N_4636);
or UO_391 (O_391,N_4820,N_4862);
or UO_392 (O_392,N_4814,N_4605);
nand UO_393 (O_393,N_4716,N_4982);
xor UO_394 (O_394,N_4670,N_4851);
and UO_395 (O_395,N_4945,N_4888);
or UO_396 (O_396,N_4999,N_4748);
nor UO_397 (O_397,N_4705,N_4700);
and UO_398 (O_398,N_4635,N_4934);
or UO_399 (O_399,N_4778,N_4769);
nand UO_400 (O_400,N_4734,N_4586);
and UO_401 (O_401,N_4764,N_4710);
and UO_402 (O_402,N_4530,N_4580);
nor UO_403 (O_403,N_4781,N_4605);
nand UO_404 (O_404,N_4515,N_4509);
nand UO_405 (O_405,N_4561,N_4710);
nand UO_406 (O_406,N_4679,N_4567);
or UO_407 (O_407,N_4851,N_4759);
or UO_408 (O_408,N_4809,N_4726);
xor UO_409 (O_409,N_4562,N_4815);
nor UO_410 (O_410,N_4838,N_4860);
xnor UO_411 (O_411,N_4638,N_4921);
nand UO_412 (O_412,N_4646,N_4823);
nand UO_413 (O_413,N_4564,N_4872);
or UO_414 (O_414,N_4611,N_4966);
nand UO_415 (O_415,N_4511,N_4615);
nor UO_416 (O_416,N_4719,N_4810);
and UO_417 (O_417,N_4987,N_4831);
and UO_418 (O_418,N_4570,N_4964);
or UO_419 (O_419,N_4557,N_4741);
and UO_420 (O_420,N_4860,N_4903);
and UO_421 (O_421,N_4967,N_4601);
and UO_422 (O_422,N_4592,N_4741);
or UO_423 (O_423,N_4580,N_4816);
and UO_424 (O_424,N_4968,N_4700);
nor UO_425 (O_425,N_4942,N_4502);
nand UO_426 (O_426,N_4878,N_4943);
nor UO_427 (O_427,N_4992,N_4509);
or UO_428 (O_428,N_4673,N_4642);
or UO_429 (O_429,N_4861,N_4698);
or UO_430 (O_430,N_4776,N_4863);
or UO_431 (O_431,N_4692,N_4543);
nor UO_432 (O_432,N_4537,N_4640);
or UO_433 (O_433,N_4645,N_4862);
or UO_434 (O_434,N_4855,N_4963);
nand UO_435 (O_435,N_4504,N_4738);
and UO_436 (O_436,N_4513,N_4540);
xnor UO_437 (O_437,N_4746,N_4899);
or UO_438 (O_438,N_4997,N_4780);
and UO_439 (O_439,N_4947,N_4951);
nand UO_440 (O_440,N_4886,N_4972);
or UO_441 (O_441,N_4566,N_4694);
nand UO_442 (O_442,N_4640,N_4769);
nor UO_443 (O_443,N_4586,N_4668);
nand UO_444 (O_444,N_4936,N_4525);
nand UO_445 (O_445,N_4839,N_4952);
nor UO_446 (O_446,N_4749,N_4946);
nor UO_447 (O_447,N_4639,N_4845);
and UO_448 (O_448,N_4947,N_4943);
and UO_449 (O_449,N_4747,N_4524);
or UO_450 (O_450,N_4977,N_4665);
and UO_451 (O_451,N_4864,N_4821);
nand UO_452 (O_452,N_4762,N_4753);
and UO_453 (O_453,N_4679,N_4641);
nand UO_454 (O_454,N_4619,N_4674);
nor UO_455 (O_455,N_4595,N_4700);
nor UO_456 (O_456,N_4708,N_4693);
nand UO_457 (O_457,N_4683,N_4997);
nand UO_458 (O_458,N_4690,N_4557);
nor UO_459 (O_459,N_4543,N_4549);
nand UO_460 (O_460,N_4721,N_4575);
and UO_461 (O_461,N_4854,N_4942);
nand UO_462 (O_462,N_4868,N_4821);
and UO_463 (O_463,N_4615,N_4845);
and UO_464 (O_464,N_4910,N_4651);
nand UO_465 (O_465,N_4645,N_4649);
nor UO_466 (O_466,N_4796,N_4658);
nand UO_467 (O_467,N_4675,N_4602);
nand UO_468 (O_468,N_4780,N_4891);
nand UO_469 (O_469,N_4586,N_4506);
nand UO_470 (O_470,N_4541,N_4852);
nor UO_471 (O_471,N_4897,N_4567);
or UO_472 (O_472,N_4626,N_4876);
or UO_473 (O_473,N_4574,N_4904);
nor UO_474 (O_474,N_4957,N_4878);
nand UO_475 (O_475,N_4598,N_4937);
nor UO_476 (O_476,N_4553,N_4729);
or UO_477 (O_477,N_4994,N_4523);
and UO_478 (O_478,N_4969,N_4876);
and UO_479 (O_479,N_4662,N_4645);
or UO_480 (O_480,N_4631,N_4925);
nor UO_481 (O_481,N_4986,N_4500);
or UO_482 (O_482,N_4832,N_4946);
xor UO_483 (O_483,N_4914,N_4686);
nor UO_484 (O_484,N_4561,N_4942);
and UO_485 (O_485,N_4627,N_4899);
nor UO_486 (O_486,N_4726,N_4823);
nor UO_487 (O_487,N_4939,N_4895);
nand UO_488 (O_488,N_4684,N_4866);
nand UO_489 (O_489,N_4622,N_4970);
nand UO_490 (O_490,N_4656,N_4524);
xnor UO_491 (O_491,N_4520,N_4865);
nor UO_492 (O_492,N_4557,N_4931);
or UO_493 (O_493,N_4632,N_4769);
and UO_494 (O_494,N_4658,N_4520);
and UO_495 (O_495,N_4555,N_4826);
nor UO_496 (O_496,N_4632,N_4981);
nand UO_497 (O_497,N_4540,N_4868);
nand UO_498 (O_498,N_4930,N_4926);
or UO_499 (O_499,N_4593,N_4742);
nor UO_500 (O_500,N_4909,N_4990);
and UO_501 (O_501,N_4527,N_4838);
nor UO_502 (O_502,N_4911,N_4615);
nand UO_503 (O_503,N_4760,N_4703);
nor UO_504 (O_504,N_4875,N_4579);
nor UO_505 (O_505,N_4625,N_4903);
and UO_506 (O_506,N_4950,N_4542);
nor UO_507 (O_507,N_4593,N_4757);
nor UO_508 (O_508,N_4588,N_4976);
nand UO_509 (O_509,N_4838,N_4694);
nand UO_510 (O_510,N_4518,N_4778);
nor UO_511 (O_511,N_4566,N_4808);
or UO_512 (O_512,N_4828,N_4835);
or UO_513 (O_513,N_4733,N_4508);
and UO_514 (O_514,N_4880,N_4588);
nor UO_515 (O_515,N_4931,N_4502);
or UO_516 (O_516,N_4776,N_4923);
or UO_517 (O_517,N_4892,N_4700);
nor UO_518 (O_518,N_4779,N_4802);
nor UO_519 (O_519,N_4568,N_4947);
nand UO_520 (O_520,N_4547,N_4820);
or UO_521 (O_521,N_4989,N_4987);
and UO_522 (O_522,N_4864,N_4647);
and UO_523 (O_523,N_4700,N_4744);
and UO_524 (O_524,N_4658,N_4602);
xor UO_525 (O_525,N_4643,N_4798);
and UO_526 (O_526,N_4678,N_4693);
and UO_527 (O_527,N_4769,N_4565);
xnor UO_528 (O_528,N_4602,N_4645);
nand UO_529 (O_529,N_4537,N_4829);
or UO_530 (O_530,N_4843,N_4544);
and UO_531 (O_531,N_4750,N_4983);
nand UO_532 (O_532,N_4737,N_4669);
or UO_533 (O_533,N_4809,N_4856);
or UO_534 (O_534,N_4988,N_4511);
or UO_535 (O_535,N_4544,N_4687);
nand UO_536 (O_536,N_4629,N_4504);
and UO_537 (O_537,N_4742,N_4781);
nor UO_538 (O_538,N_4717,N_4873);
or UO_539 (O_539,N_4541,N_4803);
and UO_540 (O_540,N_4906,N_4966);
and UO_541 (O_541,N_4530,N_4791);
nor UO_542 (O_542,N_4532,N_4772);
nor UO_543 (O_543,N_4591,N_4507);
and UO_544 (O_544,N_4802,N_4849);
nand UO_545 (O_545,N_4967,N_4846);
or UO_546 (O_546,N_4549,N_4686);
or UO_547 (O_547,N_4881,N_4988);
and UO_548 (O_548,N_4899,N_4922);
nor UO_549 (O_549,N_4790,N_4527);
nor UO_550 (O_550,N_4842,N_4582);
nor UO_551 (O_551,N_4618,N_4529);
or UO_552 (O_552,N_4577,N_4917);
nand UO_553 (O_553,N_4612,N_4824);
nor UO_554 (O_554,N_4835,N_4755);
and UO_555 (O_555,N_4696,N_4788);
nand UO_556 (O_556,N_4959,N_4645);
nor UO_557 (O_557,N_4530,N_4778);
nand UO_558 (O_558,N_4880,N_4804);
nand UO_559 (O_559,N_4933,N_4862);
nand UO_560 (O_560,N_4913,N_4975);
nand UO_561 (O_561,N_4797,N_4696);
nor UO_562 (O_562,N_4732,N_4887);
nor UO_563 (O_563,N_4789,N_4584);
nand UO_564 (O_564,N_4500,N_4593);
or UO_565 (O_565,N_4975,N_4683);
and UO_566 (O_566,N_4773,N_4582);
nor UO_567 (O_567,N_4622,N_4534);
nand UO_568 (O_568,N_4621,N_4515);
nor UO_569 (O_569,N_4714,N_4536);
nor UO_570 (O_570,N_4582,N_4704);
nor UO_571 (O_571,N_4622,N_4883);
or UO_572 (O_572,N_4963,N_4613);
nor UO_573 (O_573,N_4713,N_4925);
and UO_574 (O_574,N_4856,N_4641);
or UO_575 (O_575,N_4954,N_4856);
nand UO_576 (O_576,N_4871,N_4696);
nor UO_577 (O_577,N_4644,N_4612);
and UO_578 (O_578,N_4691,N_4656);
nand UO_579 (O_579,N_4937,N_4738);
nand UO_580 (O_580,N_4987,N_4848);
nor UO_581 (O_581,N_4904,N_4763);
or UO_582 (O_582,N_4841,N_4811);
nor UO_583 (O_583,N_4840,N_4789);
nand UO_584 (O_584,N_4974,N_4727);
nor UO_585 (O_585,N_4824,N_4826);
nand UO_586 (O_586,N_4907,N_4624);
nand UO_587 (O_587,N_4994,N_4550);
or UO_588 (O_588,N_4633,N_4992);
or UO_589 (O_589,N_4885,N_4704);
and UO_590 (O_590,N_4911,N_4938);
or UO_591 (O_591,N_4607,N_4500);
nor UO_592 (O_592,N_4558,N_4778);
nor UO_593 (O_593,N_4890,N_4609);
or UO_594 (O_594,N_4991,N_4567);
nand UO_595 (O_595,N_4907,N_4755);
nand UO_596 (O_596,N_4556,N_4894);
nor UO_597 (O_597,N_4699,N_4819);
nor UO_598 (O_598,N_4918,N_4526);
nand UO_599 (O_599,N_4610,N_4892);
nor UO_600 (O_600,N_4529,N_4554);
or UO_601 (O_601,N_4975,N_4952);
nor UO_602 (O_602,N_4918,N_4598);
xor UO_603 (O_603,N_4965,N_4799);
nor UO_604 (O_604,N_4822,N_4748);
nand UO_605 (O_605,N_4509,N_4991);
and UO_606 (O_606,N_4615,N_4939);
or UO_607 (O_607,N_4630,N_4680);
or UO_608 (O_608,N_4954,N_4543);
or UO_609 (O_609,N_4532,N_4536);
and UO_610 (O_610,N_4789,N_4765);
and UO_611 (O_611,N_4765,N_4926);
nand UO_612 (O_612,N_4781,N_4939);
or UO_613 (O_613,N_4502,N_4767);
nor UO_614 (O_614,N_4509,N_4570);
nand UO_615 (O_615,N_4984,N_4705);
nor UO_616 (O_616,N_4975,N_4597);
or UO_617 (O_617,N_4765,N_4861);
or UO_618 (O_618,N_4677,N_4834);
and UO_619 (O_619,N_4902,N_4737);
or UO_620 (O_620,N_4858,N_4561);
nor UO_621 (O_621,N_4562,N_4658);
nand UO_622 (O_622,N_4706,N_4722);
nor UO_623 (O_623,N_4658,N_4828);
or UO_624 (O_624,N_4844,N_4863);
nand UO_625 (O_625,N_4672,N_4870);
nor UO_626 (O_626,N_4638,N_4778);
nand UO_627 (O_627,N_4535,N_4879);
nand UO_628 (O_628,N_4668,N_4540);
nor UO_629 (O_629,N_4864,N_4975);
nand UO_630 (O_630,N_4900,N_4515);
nand UO_631 (O_631,N_4575,N_4590);
nor UO_632 (O_632,N_4871,N_4865);
or UO_633 (O_633,N_4703,N_4577);
nand UO_634 (O_634,N_4736,N_4855);
nand UO_635 (O_635,N_4880,N_4842);
nor UO_636 (O_636,N_4931,N_4987);
nor UO_637 (O_637,N_4782,N_4778);
and UO_638 (O_638,N_4948,N_4657);
and UO_639 (O_639,N_4663,N_4513);
nand UO_640 (O_640,N_4733,N_4685);
and UO_641 (O_641,N_4885,N_4888);
nand UO_642 (O_642,N_4698,N_4973);
and UO_643 (O_643,N_4889,N_4930);
nor UO_644 (O_644,N_4741,N_4635);
nor UO_645 (O_645,N_4839,N_4961);
and UO_646 (O_646,N_4875,N_4938);
nand UO_647 (O_647,N_4992,N_4952);
or UO_648 (O_648,N_4545,N_4601);
xor UO_649 (O_649,N_4513,N_4730);
or UO_650 (O_650,N_4763,N_4582);
and UO_651 (O_651,N_4777,N_4998);
nand UO_652 (O_652,N_4556,N_4946);
nor UO_653 (O_653,N_4607,N_4771);
nor UO_654 (O_654,N_4541,N_4666);
and UO_655 (O_655,N_4906,N_4626);
nor UO_656 (O_656,N_4615,N_4967);
nand UO_657 (O_657,N_4841,N_4736);
and UO_658 (O_658,N_4648,N_4694);
xnor UO_659 (O_659,N_4859,N_4773);
or UO_660 (O_660,N_4699,N_4676);
and UO_661 (O_661,N_4607,N_4981);
nor UO_662 (O_662,N_4814,N_4557);
or UO_663 (O_663,N_4799,N_4983);
nand UO_664 (O_664,N_4749,N_4752);
nand UO_665 (O_665,N_4755,N_4544);
and UO_666 (O_666,N_4621,N_4928);
nand UO_667 (O_667,N_4613,N_4871);
nor UO_668 (O_668,N_4958,N_4594);
or UO_669 (O_669,N_4851,N_4508);
or UO_670 (O_670,N_4768,N_4665);
nor UO_671 (O_671,N_4637,N_4946);
or UO_672 (O_672,N_4539,N_4904);
nand UO_673 (O_673,N_4878,N_4871);
nor UO_674 (O_674,N_4993,N_4542);
nand UO_675 (O_675,N_4609,N_4578);
and UO_676 (O_676,N_4947,N_4753);
and UO_677 (O_677,N_4860,N_4552);
nor UO_678 (O_678,N_4677,N_4978);
or UO_679 (O_679,N_4630,N_4548);
nand UO_680 (O_680,N_4837,N_4705);
and UO_681 (O_681,N_4885,N_4570);
xnor UO_682 (O_682,N_4661,N_4845);
and UO_683 (O_683,N_4840,N_4643);
nand UO_684 (O_684,N_4581,N_4675);
or UO_685 (O_685,N_4637,N_4628);
xnor UO_686 (O_686,N_4878,N_4734);
xor UO_687 (O_687,N_4658,N_4943);
and UO_688 (O_688,N_4662,N_4876);
nor UO_689 (O_689,N_4753,N_4982);
and UO_690 (O_690,N_4934,N_4581);
nor UO_691 (O_691,N_4969,N_4543);
nand UO_692 (O_692,N_4731,N_4896);
nand UO_693 (O_693,N_4550,N_4895);
and UO_694 (O_694,N_4659,N_4862);
and UO_695 (O_695,N_4772,N_4567);
and UO_696 (O_696,N_4620,N_4741);
or UO_697 (O_697,N_4648,N_4816);
or UO_698 (O_698,N_4545,N_4632);
and UO_699 (O_699,N_4896,N_4902);
nand UO_700 (O_700,N_4947,N_4521);
or UO_701 (O_701,N_4598,N_4858);
or UO_702 (O_702,N_4516,N_4679);
or UO_703 (O_703,N_4814,N_4843);
or UO_704 (O_704,N_4603,N_4907);
and UO_705 (O_705,N_4709,N_4702);
nor UO_706 (O_706,N_4570,N_4635);
nand UO_707 (O_707,N_4546,N_4610);
or UO_708 (O_708,N_4962,N_4649);
and UO_709 (O_709,N_4870,N_4862);
nor UO_710 (O_710,N_4980,N_4920);
nand UO_711 (O_711,N_4691,N_4563);
and UO_712 (O_712,N_4523,N_4921);
and UO_713 (O_713,N_4541,N_4572);
nor UO_714 (O_714,N_4892,N_4800);
and UO_715 (O_715,N_4560,N_4669);
and UO_716 (O_716,N_4625,N_4738);
and UO_717 (O_717,N_4683,N_4830);
and UO_718 (O_718,N_4820,N_4847);
or UO_719 (O_719,N_4734,N_4972);
nor UO_720 (O_720,N_4642,N_4552);
nand UO_721 (O_721,N_4857,N_4605);
nand UO_722 (O_722,N_4849,N_4652);
or UO_723 (O_723,N_4778,N_4681);
nor UO_724 (O_724,N_4717,N_4871);
nand UO_725 (O_725,N_4910,N_4746);
or UO_726 (O_726,N_4957,N_4864);
and UO_727 (O_727,N_4597,N_4947);
nand UO_728 (O_728,N_4971,N_4822);
nor UO_729 (O_729,N_4510,N_4809);
nand UO_730 (O_730,N_4638,N_4743);
and UO_731 (O_731,N_4678,N_4853);
and UO_732 (O_732,N_4658,N_4704);
nand UO_733 (O_733,N_4949,N_4783);
nand UO_734 (O_734,N_4857,N_4963);
nand UO_735 (O_735,N_4806,N_4776);
and UO_736 (O_736,N_4892,N_4578);
and UO_737 (O_737,N_4862,N_4618);
nand UO_738 (O_738,N_4535,N_4700);
nand UO_739 (O_739,N_4823,N_4840);
nor UO_740 (O_740,N_4807,N_4838);
and UO_741 (O_741,N_4932,N_4557);
and UO_742 (O_742,N_4985,N_4726);
nand UO_743 (O_743,N_4764,N_4583);
nand UO_744 (O_744,N_4533,N_4817);
nand UO_745 (O_745,N_4615,N_4824);
nand UO_746 (O_746,N_4567,N_4862);
nand UO_747 (O_747,N_4643,N_4573);
xnor UO_748 (O_748,N_4613,N_4901);
nand UO_749 (O_749,N_4536,N_4647);
and UO_750 (O_750,N_4569,N_4834);
nor UO_751 (O_751,N_4734,N_4541);
nor UO_752 (O_752,N_4784,N_4715);
and UO_753 (O_753,N_4883,N_4538);
and UO_754 (O_754,N_4843,N_4551);
and UO_755 (O_755,N_4695,N_4521);
nor UO_756 (O_756,N_4723,N_4524);
or UO_757 (O_757,N_4710,N_4834);
nand UO_758 (O_758,N_4996,N_4916);
and UO_759 (O_759,N_4920,N_4897);
nand UO_760 (O_760,N_4888,N_4933);
nand UO_761 (O_761,N_4866,N_4505);
or UO_762 (O_762,N_4724,N_4729);
nand UO_763 (O_763,N_4634,N_4712);
and UO_764 (O_764,N_4661,N_4750);
and UO_765 (O_765,N_4696,N_4682);
or UO_766 (O_766,N_4514,N_4944);
nand UO_767 (O_767,N_4594,N_4809);
nand UO_768 (O_768,N_4667,N_4860);
nand UO_769 (O_769,N_4647,N_4620);
and UO_770 (O_770,N_4543,N_4745);
nor UO_771 (O_771,N_4873,N_4815);
or UO_772 (O_772,N_4752,N_4817);
or UO_773 (O_773,N_4505,N_4599);
and UO_774 (O_774,N_4830,N_4721);
nor UO_775 (O_775,N_4941,N_4822);
or UO_776 (O_776,N_4617,N_4993);
xnor UO_777 (O_777,N_4536,N_4643);
nor UO_778 (O_778,N_4931,N_4566);
or UO_779 (O_779,N_4510,N_4532);
nor UO_780 (O_780,N_4620,N_4902);
or UO_781 (O_781,N_4535,N_4742);
or UO_782 (O_782,N_4924,N_4946);
or UO_783 (O_783,N_4758,N_4794);
nor UO_784 (O_784,N_4771,N_4868);
and UO_785 (O_785,N_4507,N_4802);
and UO_786 (O_786,N_4617,N_4634);
or UO_787 (O_787,N_4705,N_4808);
nand UO_788 (O_788,N_4728,N_4512);
nand UO_789 (O_789,N_4614,N_4805);
and UO_790 (O_790,N_4903,N_4832);
nor UO_791 (O_791,N_4704,N_4893);
nor UO_792 (O_792,N_4848,N_4780);
nor UO_793 (O_793,N_4714,N_4529);
or UO_794 (O_794,N_4677,N_4872);
and UO_795 (O_795,N_4677,N_4676);
or UO_796 (O_796,N_4872,N_4957);
and UO_797 (O_797,N_4842,N_4861);
and UO_798 (O_798,N_4661,N_4608);
nor UO_799 (O_799,N_4726,N_4934);
or UO_800 (O_800,N_4917,N_4583);
or UO_801 (O_801,N_4842,N_4754);
nor UO_802 (O_802,N_4698,N_4720);
or UO_803 (O_803,N_4515,N_4507);
nor UO_804 (O_804,N_4723,N_4816);
and UO_805 (O_805,N_4525,N_4798);
nand UO_806 (O_806,N_4810,N_4551);
nor UO_807 (O_807,N_4527,N_4803);
or UO_808 (O_808,N_4946,N_4735);
and UO_809 (O_809,N_4612,N_4572);
and UO_810 (O_810,N_4852,N_4691);
or UO_811 (O_811,N_4527,N_4976);
or UO_812 (O_812,N_4980,N_4528);
and UO_813 (O_813,N_4504,N_4724);
nor UO_814 (O_814,N_4630,N_4888);
nand UO_815 (O_815,N_4952,N_4614);
and UO_816 (O_816,N_4592,N_4599);
nand UO_817 (O_817,N_4893,N_4649);
nor UO_818 (O_818,N_4894,N_4711);
nand UO_819 (O_819,N_4835,N_4777);
or UO_820 (O_820,N_4951,N_4780);
and UO_821 (O_821,N_4752,N_4962);
nand UO_822 (O_822,N_4801,N_4537);
or UO_823 (O_823,N_4615,N_4707);
nand UO_824 (O_824,N_4901,N_4903);
and UO_825 (O_825,N_4671,N_4798);
or UO_826 (O_826,N_4591,N_4719);
or UO_827 (O_827,N_4575,N_4601);
or UO_828 (O_828,N_4916,N_4535);
nand UO_829 (O_829,N_4970,N_4954);
nand UO_830 (O_830,N_4880,N_4721);
and UO_831 (O_831,N_4962,N_4877);
nand UO_832 (O_832,N_4652,N_4662);
or UO_833 (O_833,N_4808,N_4667);
nand UO_834 (O_834,N_4707,N_4945);
or UO_835 (O_835,N_4669,N_4910);
xnor UO_836 (O_836,N_4631,N_4777);
nor UO_837 (O_837,N_4835,N_4510);
nand UO_838 (O_838,N_4777,N_4545);
nor UO_839 (O_839,N_4969,N_4643);
and UO_840 (O_840,N_4923,N_4945);
nor UO_841 (O_841,N_4789,N_4942);
or UO_842 (O_842,N_4911,N_4877);
nor UO_843 (O_843,N_4863,N_4565);
and UO_844 (O_844,N_4970,N_4741);
nand UO_845 (O_845,N_4925,N_4721);
or UO_846 (O_846,N_4953,N_4642);
xnor UO_847 (O_847,N_4667,N_4936);
and UO_848 (O_848,N_4552,N_4973);
nand UO_849 (O_849,N_4816,N_4724);
or UO_850 (O_850,N_4912,N_4837);
nor UO_851 (O_851,N_4877,N_4745);
xor UO_852 (O_852,N_4839,N_4908);
and UO_853 (O_853,N_4951,N_4760);
or UO_854 (O_854,N_4733,N_4847);
nor UO_855 (O_855,N_4813,N_4638);
or UO_856 (O_856,N_4768,N_4876);
xnor UO_857 (O_857,N_4598,N_4843);
and UO_858 (O_858,N_4668,N_4591);
and UO_859 (O_859,N_4520,N_4670);
and UO_860 (O_860,N_4641,N_4597);
nor UO_861 (O_861,N_4674,N_4686);
or UO_862 (O_862,N_4617,N_4734);
nand UO_863 (O_863,N_4585,N_4677);
or UO_864 (O_864,N_4521,N_4680);
nor UO_865 (O_865,N_4560,N_4651);
or UO_866 (O_866,N_4592,N_4702);
and UO_867 (O_867,N_4639,N_4868);
or UO_868 (O_868,N_4583,N_4518);
nor UO_869 (O_869,N_4746,N_4830);
nand UO_870 (O_870,N_4789,N_4565);
nand UO_871 (O_871,N_4792,N_4842);
nand UO_872 (O_872,N_4865,N_4961);
or UO_873 (O_873,N_4945,N_4619);
nor UO_874 (O_874,N_4994,N_4876);
and UO_875 (O_875,N_4531,N_4596);
and UO_876 (O_876,N_4922,N_4582);
nor UO_877 (O_877,N_4701,N_4758);
or UO_878 (O_878,N_4950,N_4797);
or UO_879 (O_879,N_4806,N_4969);
nor UO_880 (O_880,N_4601,N_4970);
or UO_881 (O_881,N_4974,N_4841);
nand UO_882 (O_882,N_4512,N_4879);
nor UO_883 (O_883,N_4835,N_4917);
and UO_884 (O_884,N_4786,N_4588);
and UO_885 (O_885,N_4701,N_4928);
or UO_886 (O_886,N_4796,N_4711);
and UO_887 (O_887,N_4944,N_4610);
and UO_888 (O_888,N_4757,N_4770);
and UO_889 (O_889,N_4591,N_4743);
and UO_890 (O_890,N_4682,N_4979);
nand UO_891 (O_891,N_4880,N_4597);
nor UO_892 (O_892,N_4692,N_4898);
nor UO_893 (O_893,N_4835,N_4989);
nor UO_894 (O_894,N_4659,N_4533);
nand UO_895 (O_895,N_4617,N_4504);
xor UO_896 (O_896,N_4654,N_4518);
nor UO_897 (O_897,N_4607,N_4965);
or UO_898 (O_898,N_4712,N_4572);
nand UO_899 (O_899,N_4867,N_4664);
or UO_900 (O_900,N_4965,N_4859);
nor UO_901 (O_901,N_4837,N_4554);
nand UO_902 (O_902,N_4699,N_4872);
and UO_903 (O_903,N_4642,N_4860);
nor UO_904 (O_904,N_4687,N_4888);
nor UO_905 (O_905,N_4686,N_4782);
nor UO_906 (O_906,N_4982,N_4979);
and UO_907 (O_907,N_4627,N_4632);
or UO_908 (O_908,N_4613,N_4920);
nand UO_909 (O_909,N_4796,N_4951);
xnor UO_910 (O_910,N_4846,N_4588);
and UO_911 (O_911,N_4942,N_4974);
nand UO_912 (O_912,N_4925,N_4628);
nor UO_913 (O_913,N_4604,N_4955);
and UO_914 (O_914,N_4726,N_4943);
nor UO_915 (O_915,N_4823,N_4608);
nor UO_916 (O_916,N_4699,N_4964);
or UO_917 (O_917,N_4732,N_4825);
nor UO_918 (O_918,N_4855,N_4564);
nand UO_919 (O_919,N_4996,N_4508);
and UO_920 (O_920,N_4825,N_4735);
and UO_921 (O_921,N_4805,N_4508);
nor UO_922 (O_922,N_4774,N_4740);
nand UO_923 (O_923,N_4845,N_4598);
nor UO_924 (O_924,N_4985,N_4921);
and UO_925 (O_925,N_4697,N_4943);
nor UO_926 (O_926,N_4953,N_4535);
and UO_927 (O_927,N_4990,N_4517);
and UO_928 (O_928,N_4965,N_4785);
or UO_929 (O_929,N_4939,N_4655);
or UO_930 (O_930,N_4706,N_4696);
or UO_931 (O_931,N_4869,N_4760);
nor UO_932 (O_932,N_4757,N_4611);
and UO_933 (O_933,N_4688,N_4554);
nor UO_934 (O_934,N_4836,N_4854);
nor UO_935 (O_935,N_4856,N_4885);
nand UO_936 (O_936,N_4768,N_4938);
nor UO_937 (O_937,N_4767,N_4548);
nand UO_938 (O_938,N_4718,N_4658);
nor UO_939 (O_939,N_4921,N_4761);
and UO_940 (O_940,N_4882,N_4511);
nor UO_941 (O_941,N_4610,N_4648);
xor UO_942 (O_942,N_4704,N_4504);
or UO_943 (O_943,N_4629,N_4954);
or UO_944 (O_944,N_4646,N_4548);
nor UO_945 (O_945,N_4927,N_4947);
or UO_946 (O_946,N_4774,N_4692);
nand UO_947 (O_947,N_4702,N_4930);
and UO_948 (O_948,N_4896,N_4500);
nor UO_949 (O_949,N_4938,N_4880);
or UO_950 (O_950,N_4510,N_4946);
nand UO_951 (O_951,N_4748,N_4672);
nand UO_952 (O_952,N_4952,N_4590);
xor UO_953 (O_953,N_4553,N_4877);
or UO_954 (O_954,N_4949,N_4709);
nand UO_955 (O_955,N_4880,N_4969);
nor UO_956 (O_956,N_4571,N_4521);
and UO_957 (O_957,N_4733,N_4758);
and UO_958 (O_958,N_4881,N_4678);
nand UO_959 (O_959,N_4569,N_4870);
nand UO_960 (O_960,N_4856,N_4893);
or UO_961 (O_961,N_4727,N_4923);
or UO_962 (O_962,N_4850,N_4573);
nand UO_963 (O_963,N_4711,N_4819);
nor UO_964 (O_964,N_4780,N_4723);
and UO_965 (O_965,N_4657,N_4685);
and UO_966 (O_966,N_4598,N_4798);
nor UO_967 (O_967,N_4641,N_4622);
or UO_968 (O_968,N_4571,N_4842);
xor UO_969 (O_969,N_4946,N_4590);
and UO_970 (O_970,N_4760,N_4615);
or UO_971 (O_971,N_4507,N_4665);
nand UO_972 (O_972,N_4857,N_4724);
or UO_973 (O_973,N_4976,N_4744);
and UO_974 (O_974,N_4961,N_4837);
and UO_975 (O_975,N_4855,N_4887);
nor UO_976 (O_976,N_4939,N_4562);
or UO_977 (O_977,N_4601,N_4727);
nand UO_978 (O_978,N_4911,N_4949);
and UO_979 (O_979,N_4653,N_4813);
or UO_980 (O_980,N_4679,N_4843);
nand UO_981 (O_981,N_4908,N_4897);
or UO_982 (O_982,N_4529,N_4659);
nor UO_983 (O_983,N_4652,N_4820);
nand UO_984 (O_984,N_4645,N_4961);
nand UO_985 (O_985,N_4759,N_4961);
nor UO_986 (O_986,N_4724,N_4878);
and UO_987 (O_987,N_4605,N_4902);
and UO_988 (O_988,N_4776,N_4699);
and UO_989 (O_989,N_4558,N_4755);
and UO_990 (O_990,N_4722,N_4830);
nor UO_991 (O_991,N_4869,N_4960);
or UO_992 (O_992,N_4598,N_4511);
or UO_993 (O_993,N_4829,N_4573);
and UO_994 (O_994,N_4803,N_4804);
or UO_995 (O_995,N_4694,N_4719);
or UO_996 (O_996,N_4521,N_4759);
and UO_997 (O_997,N_4732,N_4724);
nor UO_998 (O_998,N_4504,N_4712);
nand UO_999 (O_999,N_4833,N_4987);
endmodule