module basic_2500_25000_3000_50_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xnor U0 (N_0,In_1202,In_1014);
xor U1 (N_1,In_1735,In_29);
nor U2 (N_2,In_2297,In_1625);
or U3 (N_3,In_2180,In_1947);
nor U4 (N_4,In_480,In_576);
or U5 (N_5,In_113,In_1995);
nor U6 (N_6,In_1185,In_432);
or U7 (N_7,In_1576,In_1524);
nand U8 (N_8,In_1503,In_1969);
or U9 (N_9,In_1445,In_2095);
xnor U10 (N_10,In_1813,In_1846);
and U11 (N_11,In_57,In_2444);
or U12 (N_12,In_1169,In_1568);
nor U13 (N_13,In_141,In_1832);
xor U14 (N_14,In_1860,In_1223);
xor U15 (N_15,In_1639,In_1769);
or U16 (N_16,In_1363,In_865);
nor U17 (N_17,In_148,In_2177);
nor U18 (N_18,In_2070,In_1782);
xor U19 (N_19,In_1993,In_1716);
or U20 (N_20,In_534,In_579);
and U21 (N_21,In_1093,In_2486);
and U22 (N_22,In_1084,In_861);
and U23 (N_23,In_1573,In_239);
or U24 (N_24,In_719,In_1074);
or U25 (N_25,In_1204,In_1302);
xor U26 (N_26,In_929,In_1290);
xor U27 (N_27,In_2184,In_669);
xor U28 (N_28,In_682,In_586);
nor U29 (N_29,In_272,In_921);
nand U30 (N_30,In_288,In_2395);
nor U31 (N_31,In_257,In_250);
xnor U32 (N_32,In_961,In_144);
nand U33 (N_33,In_1795,In_2496);
or U34 (N_34,In_1622,In_552);
nand U35 (N_35,In_1234,In_2381);
and U36 (N_36,In_2198,In_85);
nand U37 (N_37,In_1222,In_131);
xnor U38 (N_38,In_1842,In_2250);
xnor U39 (N_39,In_989,In_2315);
nor U40 (N_40,In_407,In_2082);
nand U41 (N_41,In_1338,In_2153);
nand U42 (N_42,In_1551,In_1171);
and U43 (N_43,In_1188,In_493);
or U44 (N_44,In_888,In_966);
xnor U45 (N_45,In_299,In_2252);
xor U46 (N_46,In_1491,In_1684);
or U47 (N_47,In_1149,In_956);
or U48 (N_48,In_206,In_135);
and U49 (N_49,In_1066,In_1815);
and U50 (N_50,In_1968,In_847);
and U51 (N_51,In_1747,In_1816);
or U52 (N_52,In_2127,In_556);
nand U53 (N_53,In_1672,In_887);
nor U54 (N_54,In_1766,In_1225);
nand U55 (N_55,In_458,In_1138);
and U56 (N_56,In_1159,In_1714);
nor U57 (N_57,In_497,In_310);
xor U58 (N_58,In_2478,In_768);
and U59 (N_59,In_566,In_564);
xor U60 (N_60,In_1618,In_881);
and U61 (N_61,In_2441,In_2243);
nand U62 (N_62,In_2223,In_2107);
or U63 (N_63,In_1422,In_974);
and U64 (N_64,In_1603,In_1528);
or U65 (N_65,In_1796,In_1888);
or U66 (N_66,In_979,In_2222);
nand U67 (N_67,In_1167,In_1651);
nand U68 (N_68,In_1597,In_1421);
nor U69 (N_69,In_2161,In_855);
nand U70 (N_70,In_2111,In_1218);
and U71 (N_71,In_1918,In_1298);
or U72 (N_72,In_446,In_528);
or U73 (N_73,In_1304,In_952);
nor U74 (N_74,In_1897,In_1299);
nor U75 (N_75,In_1268,In_1071);
or U76 (N_76,In_212,In_190);
xnor U77 (N_77,In_987,In_173);
nor U78 (N_78,In_2339,In_725);
xnor U79 (N_79,In_2475,In_278);
nand U80 (N_80,In_474,In_2216);
and U81 (N_81,In_983,In_1498);
xor U82 (N_82,In_404,In_945);
nand U83 (N_83,In_1989,In_785);
or U84 (N_84,In_664,In_577);
or U85 (N_85,In_2455,In_1956);
and U86 (N_86,In_2356,In_2266);
or U87 (N_87,In_1067,In_1500);
xor U88 (N_88,In_228,In_1020);
or U89 (N_89,In_1770,In_147);
xnor U90 (N_90,In_23,In_409);
or U91 (N_91,In_2402,In_1615);
nand U92 (N_92,In_804,In_2069);
xor U93 (N_93,In_1056,In_2325);
or U94 (N_94,In_233,In_734);
or U95 (N_95,In_677,In_1496);
and U96 (N_96,In_210,In_1256);
or U97 (N_97,In_2330,In_1506);
and U98 (N_98,In_1613,In_1316);
nor U99 (N_99,In_428,In_2305);
xnor U100 (N_100,In_63,In_1446);
nand U101 (N_101,In_2190,In_2276);
nor U102 (N_102,In_628,In_2122);
xnor U103 (N_103,In_2316,In_529);
and U104 (N_104,In_1679,In_1254);
xor U105 (N_105,In_317,In_1411);
and U106 (N_106,In_1129,In_817);
and U107 (N_107,In_2119,In_560);
and U108 (N_108,In_764,In_2163);
xor U109 (N_109,In_1140,In_704);
nand U110 (N_110,In_1305,In_2419);
xor U111 (N_111,In_571,In_1343);
nor U112 (N_112,In_470,In_2060);
and U113 (N_113,In_2105,In_465);
nor U114 (N_114,In_905,In_2333);
xor U115 (N_115,In_2014,In_1221);
xnor U116 (N_116,In_1976,In_595);
nor U117 (N_117,In_319,In_1147);
nand U118 (N_118,In_2192,In_408);
and U119 (N_119,In_1321,In_1595);
and U120 (N_120,In_170,In_1873);
and U121 (N_121,In_256,In_2267);
or U122 (N_122,In_1749,In_2033);
and U123 (N_123,In_568,In_641);
and U124 (N_124,In_1341,In_1105);
nand U125 (N_125,In_1400,In_1023);
and U126 (N_126,In_130,In_195);
xnor U127 (N_127,In_1121,In_1201);
xnor U128 (N_128,In_2239,In_1405);
nand U129 (N_129,In_472,In_950);
and U130 (N_130,In_1228,In_1912);
and U131 (N_131,In_2350,In_187);
or U132 (N_132,In_2169,In_2071);
and U133 (N_133,In_1642,In_1541);
and U134 (N_134,In_1529,In_1035);
nand U135 (N_135,In_1864,In_1424);
or U136 (N_136,In_448,In_1374);
and U137 (N_137,In_1508,In_1726);
or U138 (N_138,In_452,In_1893);
xor U139 (N_139,In_262,In_819);
xor U140 (N_140,In_1203,In_1784);
nor U141 (N_141,In_1297,In_1010);
nand U142 (N_142,In_1178,In_638);
nor U143 (N_143,In_2370,In_588);
nand U144 (N_144,In_765,In_2152);
nand U145 (N_145,In_690,In_1307);
or U146 (N_146,In_1113,In_414);
xor U147 (N_147,In_463,In_1315);
or U148 (N_148,In_242,In_1383);
xor U149 (N_149,In_1317,In_383);
or U150 (N_150,In_2187,In_1367);
nor U151 (N_151,In_186,In_1807);
xor U152 (N_152,In_2317,In_852);
and U153 (N_153,In_467,In_582);
nor U154 (N_154,In_1898,In_623);
nand U155 (N_155,In_1678,In_812);
and U156 (N_156,In_1459,In_1200);
nor U157 (N_157,In_2128,In_1535);
or U158 (N_158,In_750,In_1328);
nand U159 (N_159,In_1854,In_1469);
and U160 (N_160,In_2135,In_980);
xnor U161 (N_161,In_589,In_1931);
xnor U162 (N_162,In_1547,In_1992);
nor U163 (N_163,In_460,In_1030);
and U164 (N_164,In_364,In_648);
nand U165 (N_165,In_535,In_977);
and U166 (N_166,In_1539,In_1017);
and U167 (N_167,In_890,In_2020);
and U168 (N_168,In_1789,In_499);
nor U169 (N_169,In_1963,In_1768);
or U170 (N_170,In_1722,In_639);
or U171 (N_171,In_732,In_26);
and U172 (N_172,In_89,In_941);
xnor U173 (N_173,In_1062,In_350);
xor U174 (N_174,In_644,In_234);
xor U175 (N_175,In_1817,In_1162);
and U176 (N_176,In_146,In_567);
nand U177 (N_177,In_326,In_959);
xor U178 (N_178,In_1665,In_166);
nor U179 (N_179,In_2299,In_2411);
nand U180 (N_180,In_316,In_1286);
and U181 (N_181,In_882,In_994);
nand U182 (N_182,In_1774,In_1476);
or U183 (N_183,In_982,In_1661);
and U184 (N_184,In_370,In_860);
nor U185 (N_185,In_2459,In_646);
and U186 (N_186,In_96,In_1802);
nor U187 (N_187,In_1249,In_2015);
nor U188 (N_188,In_1182,In_356);
and U189 (N_189,In_2327,In_680);
nor U190 (N_190,In_770,In_1991);
xnor U191 (N_191,In_1320,In_1082);
nand U192 (N_192,In_2214,In_1607);
xnor U193 (N_193,In_1765,In_5);
xor U194 (N_194,In_963,In_1578);
nor U195 (N_195,In_2258,In_1820);
nand U196 (N_196,In_502,In_1707);
and U197 (N_197,In_2043,In_308);
nor U198 (N_198,In_2462,In_1628);
and U199 (N_199,In_318,In_1692);
and U200 (N_200,In_908,In_2050);
and U201 (N_201,In_713,In_748);
nor U202 (N_202,In_2003,In_799);
and U203 (N_203,In_870,In_520);
or U204 (N_204,In_2204,In_2401);
nand U205 (N_205,In_269,In_635);
xor U206 (N_206,In_305,In_511);
or U207 (N_207,In_352,In_1194);
nand U208 (N_208,In_1455,In_2221);
and U209 (N_209,In_2264,In_1003);
and U210 (N_210,In_395,In_811);
xnor U211 (N_211,In_2200,In_999);
nor U212 (N_212,In_1423,In_2162);
nand U213 (N_213,In_265,In_1439);
and U214 (N_214,In_1612,In_51);
nor U215 (N_215,In_2413,In_1555);
and U216 (N_216,In_620,In_140);
nor U217 (N_217,In_825,In_706);
xor U218 (N_218,In_1351,In_2287);
and U219 (N_219,In_221,In_619);
nand U220 (N_220,In_1440,In_2056);
xnor U221 (N_221,In_161,In_1242);
or U222 (N_222,In_1804,In_196);
nand U223 (N_223,In_301,In_1232);
xnor U224 (N_224,In_1208,In_2271);
nor U225 (N_225,In_878,In_1039);
xor U226 (N_226,In_1882,In_2188);
xor U227 (N_227,In_2260,In_2217);
and U228 (N_228,In_1526,In_2183);
nor U229 (N_229,In_2290,In_1834);
nand U230 (N_230,In_482,In_1664);
nor U231 (N_231,In_909,In_1031);
nor U232 (N_232,In_2320,In_975);
nand U233 (N_233,In_1384,In_138);
nand U234 (N_234,In_723,In_1072);
nor U235 (N_235,In_1983,In_1790);
xnor U236 (N_236,In_542,In_36);
or U237 (N_237,In_402,In_2032);
nor U238 (N_238,In_1457,In_2285);
and U239 (N_239,In_324,In_489);
and U240 (N_240,In_289,In_1153);
xor U241 (N_241,In_151,In_124);
nand U242 (N_242,In_1621,In_583);
xnor U243 (N_243,In_1047,In_1382);
nand U244 (N_244,In_884,In_532);
and U245 (N_245,In_1803,In_1146);
nor U246 (N_246,In_2415,In_2080);
nand U247 (N_247,In_1309,In_926);
and U248 (N_248,In_2034,In_924);
nand U249 (N_249,In_767,In_2253);
xnor U250 (N_250,In_2270,In_1744);
nand U251 (N_251,In_1037,In_1142);
and U252 (N_252,In_777,In_1365);
nand U253 (N_253,In_1273,In_1542);
and U254 (N_254,In_866,In_839);
nand U255 (N_255,In_792,In_1633);
or U256 (N_256,In_2388,In_92);
xor U257 (N_257,In_1733,In_1571);
nor U258 (N_258,In_2144,In_2058);
and U259 (N_259,In_1914,In_1552);
nand U260 (N_260,In_435,In_742);
nand U261 (N_261,In_297,In_2102);
or U262 (N_262,In_181,In_2451);
nand U263 (N_263,In_1154,In_1835);
nand U264 (N_264,In_1592,In_1436);
nor U265 (N_265,In_329,In_998);
nand U266 (N_266,In_1326,In_2254);
nor U267 (N_267,In_876,In_2343);
xor U268 (N_268,In_1604,In_390);
nand U269 (N_269,In_285,In_679);
nand U270 (N_270,In_1441,In_2115);
nor U271 (N_271,In_2248,In_97);
nand U272 (N_272,In_123,In_238);
nand U273 (N_273,In_1870,In_2324);
or U274 (N_274,In_503,In_418);
nand U275 (N_275,In_443,In_2084);
xnor U276 (N_276,In_1915,In_231);
nand U277 (N_277,In_1157,In_311);
xor U278 (N_278,In_2336,In_867);
and U279 (N_279,In_1674,In_76);
or U280 (N_280,In_1981,In_1531);
or U281 (N_281,In_1636,In_2427);
or U282 (N_282,In_1549,In_649);
or U283 (N_283,In_930,In_1923);
xnor U284 (N_284,In_423,In_1151);
or U285 (N_285,In_1483,In_830);
and U286 (N_286,In_354,In_1884);
nor U287 (N_287,In_1731,In_292);
nand U288 (N_288,In_806,In_1009);
and U289 (N_289,In_385,In_507);
nor U290 (N_290,In_633,In_986);
nor U291 (N_291,In_2349,In_2372);
nand U292 (N_292,In_2430,In_728);
nand U293 (N_293,In_521,In_397);
or U294 (N_294,In_1743,In_1434);
and U295 (N_295,In_656,In_508);
nor U296 (N_296,In_1277,In_2498);
nor U297 (N_297,In_16,In_1101);
nor U298 (N_298,In_509,In_1184);
and U299 (N_299,In_1408,In_2371);
nand U300 (N_300,In_340,In_1451);
xnor U301 (N_301,In_2143,In_2129);
and U302 (N_302,In_1990,In_1094);
nand U303 (N_303,In_1065,In_720);
and U304 (N_304,In_1024,In_66);
xnor U305 (N_305,In_2054,In_377);
nand U306 (N_306,In_1401,In_0);
and U307 (N_307,In_1713,In_678);
nand U308 (N_308,In_2164,In_222);
xnor U309 (N_309,In_2345,In_949);
or U310 (N_310,In_932,In_596);
xor U311 (N_311,In_2039,In_2277);
nand U312 (N_312,In_45,In_1294);
xor U313 (N_313,In_298,In_14);
nand U314 (N_314,In_209,In_1841);
xor U315 (N_315,In_787,In_1895);
and U316 (N_316,In_111,In_759);
nand U317 (N_317,In_286,In_1510);
xnor U318 (N_318,In_653,In_1243);
and U319 (N_319,In_1904,In_2306);
xor U320 (N_320,In_2382,In_1306);
or U321 (N_321,In_1724,In_2113);
or U322 (N_322,In_199,In_2145);
nand U323 (N_323,In_1300,In_1448);
and U324 (N_324,In_1193,In_46);
and U325 (N_325,In_1984,In_2348);
or U326 (N_326,In_1695,In_545);
nor U327 (N_327,In_1754,In_55);
or U328 (N_328,In_1970,In_304);
xor U329 (N_329,In_1080,In_1544);
nor U330 (N_330,In_2340,In_2347);
nand U331 (N_331,In_2310,In_1532);
or U332 (N_332,In_661,In_1504);
or U333 (N_333,In_2137,In_1128);
nor U334 (N_334,In_240,In_450);
nand U335 (N_335,In_525,In_2093);
nor U336 (N_336,In_2213,In_133);
nor U337 (N_337,In_2472,In_2199);
nand U338 (N_338,In_33,In_1165);
nor U339 (N_339,In_769,In_1033);
nor U340 (N_340,In_1605,In_2083);
nand U341 (N_341,In_374,In_651);
nand U342 (N_342,In_2394,In_59);
and U343 (N_343,In_1737,In_25);
nor U344 (N_344,In_1189,In_1939);
nor U345 (N_345,In_1516,In_2328);
nand U346 (N_346,In_2311,In_339);
nand U347 (N_347,In_2241,In_2283);
or U348 (N_348,In_153,In_1879);
and U349 (N_349,In_1346,In_838);
nand U350 (N_350,In_516,In_1929);
nand U351 (N_351,In_673,In_1301);
nor U352 (N_352,In_1703,In_2424);
and U353 (N_353,In_2040,In_874);
and U354 (N_354,In_630,In_2458);
or U355 (N_355,In_1881,In_1572);
and U356 (N_356,In_2052,In_551);
or U357 (N_357,In_781,In_2284);
xnor U358 (N_358,In_47,In_1805);
or U359 (N_359,In_687,In_205);
nand U360 (N_360,In_968,In_1831);
nor U361 (N_361,In_2263,In_1746);
xnor U362 (N_362,In_2460,In_2046);
nand U363 (N_363,In_689,In_2425);
or U364 (N_364,In_2295,In_700);
xor U365 (N_365,In_2406,In_859);
nor U366 (N_366,In_530,In_2368);
nor U367 (N_367,In_2166,In_1442);
or U368 (N_368,In_84,In_1525);
nand U369 (N_369,In_1117,In_2175);
or U370 (N_370,In_622,In_268);
or U371 (N_371,In_58,In_976);
and U372 (N_372,In_1533,In_1191);
nor U373 (N_373,In_1686,In_684);
nand U374 (N_374,In_1959,In_83);
nand U375 (N_375,In_2236,In_2302);
or U376 (N_376,In_1347,In_1000);
nor U377 (N_377,In_1279,In_451);
xnor U378 (N_378,In_970,In_2124);
or U379 (N_379,In_1673,In_343);
xnor U380 (N_380,In_2318,In_2351);
and U381 (N_381,In_1919,In_1131);
nor U382 (N_382,In_2219,In_219);
or U383 (N_383,In_1414,In_1059);
or U384 (N_384,In_1458,In_2022);
or U385 (N_385,In_2097,In_1892);
nand U386 (N_386,In_1838,In_1291);
and U387 (N_387,In_1104,In_411);
or U388 (N_388,In_2298,In_175);
or U389 (N_389,In_718,In_2027);
nand U390 (N_390,In_1415,In_2151);
nand U391 (N_391,In_658,In_697);
nor U392 (N_392,In_565,In_1269);
xor U393 (N_393,In_2439,In_371);
nor U394 (N_394,In_834,In_441);
nand U395 (N_395,In_1567,In_614);
xor U396 (N_396,In_245,In_1785);
and U397 (N_397,In_1527,In_632);
xor U398 (N_398,In_1312,In_1876);
xnor U399 (N_399,In_2181,In_681);
nor U400 (N_400,In_2231,In_709);
nand U401 (N_401,In_406,In_864);
nand U402 (N_402,In_698,In_1112);
and U403 (N_403,In_688,In_918);
nand U404 (N_404,In_1951,In_2142);
and U405 (N_405,In_889,In_1878);
or U406 (N_406,In_366,In_1658);
and U407 (N_407,In_626,In_320);
or U408 (N_408,In_1245,In_1683);
or U409 (N_409,In_1199,In_569);
xnor U410 (N_410,In_1362,In_1404);
nor U411 (N_411,In_1935,In_543);
nor U412 (N_412,In_1289,In_1610);
nor U413 (N_413,In_456,In_88);
nand U414 (N_414,In_2265,In_727);
or U415 (N_415,In_561,In_1644);
nor U416 (N_416,In_2049,In_2047);
and U417 (N_417,In_895,In_105);
nor U418 (N_418,In_666,In_1013);
nand U419 (N_419,In_2293,In_302);
and U420 (N_420,In_121,In_1545);
and U421 (N_421,In_1760,In_2361);
or U422 (N_422,In_20,In_1478);
xor U423 (N_423,In_2450,In_156);
and U424 (N_424,In_1505,In_801);
or U425 (N_425,In_1987,In_831);
and U426 (N_426,In_1356,In_192);
or U427 (N_427,In_2326,In_2041);
or U428 (N_428,In_1352,In_1064);
or U429 (N_429,In_808,In_1641);
nor U430 (N_430,In_841,In_602);
and U431 (N_431,In_1659,In_1797);
nand U432 (N_432,In_2449,In_922);
and U433 (N_433,In_821,In_107);
nand U434 (N_434,In_657,In_1553);
nand U435 (N_435,In_1509,In_1982);
and U436 (N_436,In_1775,In_1360);
or U437 (N_437,In_2148,In_693);
and U438 (N_438,In_1358,In_805);
nand U439 (N_439,In_1034,In_143);
nor U440 (N_440,In_1851,In_869);
and U441 (N_441,In_321,In_518);
xor U442 (N_442,In_476,In_424);
xor U443 (N_443,In_1863,In_763);
xor U444 (N_444,In_1327,In_621);
nor U445 (N_445,In_1164,In_2433);
nand U446 (N_446,In_1669,In_1702);
or U447 (N_447,In_1076,In_214);
nand U448 (N_448,In_1303,In_880);
or U449 (N_449,In_2090,In_574);
nand U450 (N_450,In_1018,In_30);
nand U451 (N_451,In_984,In_1687);
xnor U452 (N_452,In_1255,In_330);
nor U453 (N_453,In_2292,In_943);
nand U454 (N_454,In_267,In_1593);
or U455 (N_455,In_2416,In_18);
xnor U456 (N_456,In_942,In_2467);
nor U457 (N_457,In_389,In_2412);
nand U458 (N_458,In_372,In_1250);
nor U459 (N_459,In_2029,In_608);
nor U460 (N_460,In_2079,In_2123);
nor U461 (N_461,In_54,In_1588);
nor U462 (N_462,In_655,In_1041);
nand U463 (N_463,In_53,In_331);
xor U464 (N_464,In_2256,In_1522);
nor U465 (N_465,In_1426,In_2136);
and U466 (N_466,In_116,In_1825);
or U467 (N_467,In_2076,In_1560);
and U468 (N_468,In_1574,In_1152);
nor U469 (N_469,In_2023,In_1889);
or U470 (N_470,In_323,In_1430);
nor U471 (N_471,In_2464,In_99);
nand U472 (N_472,In_1580,In_1109);
or U473 (N_473,In_183,In_1399);
or U474 (N_474,In_94,In_490);
nor U475 (N_475,In_2384,In_1319);
nor U476 (N_476,In_271,In_419);
xor U477 (N_477,In_382,In_388);
nor U478 (N_478,In_1172,In_826);
nor U479 (N_479,In_916,In_1403);
and U480 (N_480,In_437,In_562);
or U481 (N_481,In_1627,In_1908);
nor U482 (N_482,In_229,In_1594);
or U483 (N_483,In_363,In_2331);
or U484 (N_484,In_629,In_1718);
nor U485 (N_485,In_31,In_422);
nor U486 (N_486,In_972,In_346);
and U487 (N_487,In_716,In_627);
or U488 (N_488,In_899,In_2456);
nand U489 (N_489,In_894,In_2101);
xor U490 (N_490,In_538,In_2120);
and U491 (N_491,In_1847,In_2473);
nor U492 (N_492,In_1750,In_1468);
nand U493 (N_493,In_592,In_11);
nand U494 (N_494,In_177,In_2156);
xnor U495 (N_495,In_2037,In_501);
xor U496 (N_496,In_1417,In_1287);
and U497 (N_497,In_392,In_1481);
or U498 (N_498,In_2396,In_722);
and U499 (N_499,In_1322,In_284);
xnor U500 (N_500,In_606,In_1126);
or U501 (N_501,In_605,N_290);
nand U502 (N_502,In_1027,In_2393);
nand U503 (N_503,In_2036,In_580);
nor U504 (N_504,N_297,In_2089);
or U505 (N_505,N_115,In_1342);
nand U506 (N_506,N_246,In_1649);
nor U507 (N_507,In_739,In_2321);
and U508 (N_508,N_369,N_322);
or U509 (N_509,In_1937,In_1083);
and U510 (N_510,N_171,In_1587);
nand U511 (N_511,In_281,In_654);
or U512 (N_512,In_9,In_1652);
or U513 (N_513,In_1058,In_2383);
nor U514 (N_514,In_616,In_2346);
or U515 (N_515,N_61,In_544);
nor U516 (N_516,In_2038,In_438);
xor U517 (N_517,In_791,In_208);
or U518 (N_518,In_1958,In_1700);
nor U519 (N_519,N_373,In_1492);
nand U520 (N_520,In_934,In_634);
nor U521 (N_521,In_686,In_886);
nand U522 (N_522,In_1960,In_235);
or U523 (N_523,N_52,In_1438);
nand U524 (N_524,In_375,In_104);
xnor U525 (N_525,N_350,In_1063);
and U526 (N_526,In_1464,N_445);
nor U527 (N_527,In_559,In_1962);
and U528 (N_528,In_1032,N_384);
nand U529 (N_529,In_2159,In_236);
and U530 (N_530,In_1911,In_243);
and U531 (N_531,N_210,N_193);
xnor U532 (N_532,In_1773,In_360);
or U533 (N_533,N_28,N_162);
nor U534 (N_534,N_359,In_1479);
and U535 (N_535,In_912,In_1556);
and U536 (N_536,In_1662,In_1559);
xor U537 (N_537,In_504,In_479);
or U538 (N_538,N_425,In_872);
nor U539 (N_539,In_1463,N_264);
or U540 (N_540,In_2422,In_1739);
nor U541 (N_541,In_558,In_149);
nor U542 (N_542,N_427,In_707);
nand U543 (N_543,N_421,In_1630);
nor U544 (N_544,In_923,In_617);
and U545 (N_545,In_2085,In_1057);
nor U546 (N_546,N_1,In_1776);
xnor U547 (N_547,N_431,In_2010);
or U548 (N_548,In_1704,In_1614);
nand U549 (N_549,In_1762,In_2203);
xnor U550 (N_550,In_1028,In_32);
nand U551 (N_551,In_1462,In_2209);
or U552 (N_552,In_997,In_1311);
nand U553 (N_553,In_2471,In_786);
nor U554 (N_554,In_2028,In_244);
xor U555 (N_555,In_1709,In_1370);
or U556 (N_556,In_873,N_366);
or U557 (N_557,In_2303,In_461);
nand U558 (N_558,N_319,In_1168);
or U559 (N_559,In_902,In_1973);
nand U560 (N_560,N_14,In_2398);
nand U561 (N_561,In_447,In_1132);
or U562 (N_562,In_1231,In_1206);
or U563 (N_563,In_587,In_751);
xnor U564 (N_564,In_2245,In_992);
nor U565 (N_565,In_1158,In_1917);
xor U566 (N_566,N_367,In_376);
nand U567 (N_567,N_341,In_1753);
and U568 (N_568,In_1901,In_1418);
xor U569 (N_569,In_731,N_176);
xnor U570 (N_570,In_1477,In_512);
nand U571 (N_571,In_398,In_2308);
nand U572 (N_572,In_481,In_1853);
and U573 (N_573,N_294,In_2157);
or U574 (N_574,N_447,In_2002);
or U575 (N_575,N_5,In_379);
and U576 (N_576,In_188,In_1265);
nand U577 (N_577,In_1977,N_484);
and U578 (N_578,In_2081,In_2171);
and U579 (N_579,In_736,In_1396);
xnor U580 (N_580,In_1332,In_1934);
and U581 (N_581,In_809,In_368);
and U582 (N_582,In_1606,N_175);
nor U583 (N_583,In_965,N_168);
and U584 (N_584,In_610,N_180);
xnor U585 (N_585,N_407,In_2001);
and U586 (N_586,In_676,In_1045);
nor U587 (N_587,In_776,N_352);
and U588 (N_588,In_2319,In_2132);
nor U589 (N_589,In_836,In_1314);
xor U590 (N_590,N_111,In_612);
xnor U591 (N_591,In_1857,In_2208);
xor U592 (N_592,N_135,In_2379);
or U593 (N_593,In_1611,In_1681);
xnor U594 (N_594,In_2488,In_261);
nor U595 (N_595,In_717,In_1647);
xor U596 (N_596,In_1575,In_1619);
xor U597 (N_597,In_2117,In_1433);
nand U598 (N_598,In_1558,In_1261);
nor U599 (N_599,N_252,In_380);
or U600 (N_600,In_1238,In_2461);
or U601 (N_601,In_893,In_1213);
nor U602 (N_602,In_1,In_1029);
and U603 (N_603,In_2004,In_594);
nand U604 (N_604,In_853,In_1967);
xnor U605 (N_605,In_90,In_1209);
and U606 (N_606,In_771,In_2167);
xor U607 (N_607,In_2363,In_252);
nand U608 (N_608,N_439,N_87);
nor U609 (N_609,In_1246,In_1247);
and U610 (N_610,In_1461,In_1386);
xor U611 (N_611,In_2304,N_63);
and U612 (N_612,In_487,In_1357);
and U613 (N_613,In_1116,In_2255);
or U614 (N_614,In_1648,In_334);
or U615 (N_615,In_2149,In_484);
nand U616 (N_616,In_1953,N_460);
xnor U617 (N_617,N_17,In_1016);
and U618 (N_618,In_1262,In_691);
and U619 (N_619,In_531,In_1626);
xor U620 (N_620,N_30,N_119);
and U621 (N_621,In_2121,N_121);
nand U622 (N_622,In_797,In_488);
nor U623 (N_623,In_904,N_11);
and U624 (N_624,N_133,In_1519);
xnor U625 (N_625,In_2454,In_1177);
or U626 (N_626,N_335,In_2096);
and U627 (N_627,N_68,N_413);
or U628 (N_628,In_2019,N_476);
nor U629 (N_629,In_1450,In_158);
nor U630 (N_630,In_2249,In_69);
nor U631 (N_631,N_126,In_1339);
nand U632 (N_632,N_38,In_746);
nor U633 (N_633,In_41,N_430);
and U634 (N_634,N_327,In_2278);
or U635 (N_635,In_1467,In_824);
xor U636 (N_636,In_433,In_1608);
xnor U637 (N_637,In_2366,In_1089);
or U638 (N_638,In_2185,In_1978);
nor U639 (N_639,In_896,In_2435);
xnor U640 (N_640,In_1745,N_276);
or U641 (N_641,In_118,N_0);
nor U642 (N_642,In_119,N_55);
nor U643 (N_643,In_2007,In_1283);
and U644 (N_644,In_990,In_1771);
xnor U645 (N_645,N_240,In_1861);
nor U646 (N_646,In_248,N_403);
or U647 (N_647,In_251,In_1645);
and U648 (N_648,In_2274,N_338);
xnor U649 (N_649,In_755,In_1638);
xnor U650 (N_650,In_936,In_394);
or U651 (N_651,In_2309,In_1124);
xor U652 (N_652,In_1174,N_35);
nand U653 (N_653,In_294,In_152);
and U654 (N_654,N_262,In_1927);
or U655 (N_655,N_138,In_1125);
nand U656 (N_656,In_357,N_435);
nand U657 (N_657,In_1650,N_295);
nor U658 (N_658,N_215,In_2103);
and U659 (N_659,N_261,In_264);
or U660 (N_660,N_195,In_2008);
xor U661 (N_661,In_197,N_227);
xor U662 (N_662,N_385,In_2061);
nor U663 (N_663,N_344,In_2476);
xor U664 (N_664,In_1643,N_77);
nand U665 (N_665,In_2092,In_2296);
nor U666 (N_666,In_712,In_2426);
or U667 (N_667,In_2016,In_2094);
xor U668 (N_668,In_2334,N_239);
or U669 (N_669,In_1836,In_253);
xnor U670 (N_670,In_67,N_333);
nor U671 (N_671,N_383,In_1091);
nor U672 (N_672,In_2044,In_840);
xor U673 (N_673,In_1100,In_1756);
nand U674 (N_674,In_217,In_1330);
or U675 (N_675,N_426,In_845);
xnor U676 (N_676,In_948,In_1591);
or U677 (N_677,N_219,In_1295);
xnor U678 (N_678,In_2342,In_1444);
nand U679 (N_679,In_1053,In_1623);
nor U680 (N_680,In_1274,In_2474);
and U681 (N_681,In_1596,In_854);
or U682 (N_682,In_1215,In_486);
nand U683 (N_683,In_1848,N_471);
nand U684 (N_684,In_1398,In_1368);
xor U685 (N_685,In_546,In_607);
xor U686 (N_686,In_803,In_820);
nand U687 (N_687,In_1734,In_1600);
nor U688 (N_688,N_377,In_312);
xor U689 (N_689,In_1230,N_480);
or U690 (N_690,N_187,N_483);
nor U691 (N_691,N_161,N_78);
and U692 (N_692,In_519,In_464);
xnor U693 (N_693,In_2035,In_2259);
and U694 (N_694,In_100,In_440);
or U695 (N_695,N_91,In_2369);
nand U696 (N_696,In_2341,N_89);
xnor U697 (N_697,N_96,In_139);
nand U698 (N_698,In_1378,N_199);
and U699 (N_699,In_1830,In_1998);
xor U700 (N_700,N_389,In_892);
nand U701 (N_701,N_288,In_2240);
nand U702 (N_702,In_1660,In_1666);
and U703 (N_703,In_386,In_2055);
nand U704 (N_704,N_353,In_2457);
xor U705 (N_705,In_1260,N_32);
xor U706 (N_706,In_898,In_127);
and U707 (N_707,In_1812,In_883);
and U708 (N_708,In_498,N_250);
nor U709 (N_709,In_526,In_1335);
and U710 (N_710,N_90,In_1829);
xnor U711 (N_711,In_2206,N_108);
and U712 (N_712,In_1219,In_851);
xnor U713 (N_713,In_954,In_2048);
nand U714 (N_714,In_1921,In_1723);
or U715 (N_715,In_1845,In_1624);
or U716 (N_716,In_1198,In_1653);
nor U717 (N_717,In_749,In_1364);
xor U718 (N_718,In_1671,In_1470);
and U719 (N_719,N_420,N_27);
nand U720 (N_720,In_1263,In_232);
or U721 (N_721,In_1211,N_347);
and U722 (N_722,In_2026,In_2017);
or U723 (N_723,In_598,In_2228);
nor U724 (N_724,In_1480,In_2448);
or U725 (N_725,N_213,N_283);
nand U726 (N_726,In_2352,In_933);
xnor U727 (N_727,In_541,In_2168);
and U728 (N_728,In_2075,In_715);
xnor U729 (N_729,N_456,In_790);
or U730 (N_730,In_609,In_1757);
nand U731 (N_731,N_43,In_2446);
and U732 (N_732,In_2359,In_2495);
xnor U733 (N_733,In_345,N_296);
and U734 (N_734,In_1233,N_354);
or U735 (N_735,N_147,N_258);
and U736 (N_736,In_2499,N_475);
or U737 (N_737,N_285,In_237);
nand U738 (N_738,In_180,In_2404);
nand U739 (N_739,In_813,In_1118);
nor U740 (N_740,In_857,In_555);
nand U741 (N_741,In_2251,In_2358);
or U742 (N_742,In_1859,N_18);
or U743 (N_743,In_1195,In_2063);
or U744 (N_744,N_363,In_15);
nor U745 (N_745,In_174,In_1190);
xor U746 (N_746,In_2195,In_1849);
xor U747 (N_747,N_33,In_259);
nor U748 (N_748,In_721,N_120);
nor U749 (N_749,In_1925,N_62);
nand U750 (N_750,In_1486,In_1308);
nand U751 (N_751,In_1742,N_107);
nor U752 (N_752,In_313,In_705);
xor U753 (N_753,In_849,In_737);
nand U754 (N_754,In_24,In_584);
nand U755 (N_755,In_275,In_436);
or U756 (N_756,In_900,N_398);
nand U757 (N_757,In_2098,N_76);
or U758 (N_758,In_290,In_1902);
nand U759 (N_759,In_2353,In_1495);
nor U760 (N_760,In_2130,In_1550);
or U761 (N_761,N_123,In_585);
xor U762 (N_762,N_306,In_513);
or U763 (N_763,N_72,In_95);
xor U764 (N_764,In_471,In_2237);
nor U765 (N_765,N_42,In_49);
nor U766 (N_766,N_146,In_1429);
and U767 (N_767,In_871,In_1096);
nand U768 (N_768,In_710,In_17);
xnor U769 (N_769,N_188,In_1361);
xnor U770 (N_770,In_77,In_2197);
and U771 (N_771,In_927,In_1699);
nor U772 (N_772,In_2099,In_1964);
nor U773 (N_773,In_810,N_441);
xnor U774 (N_774,In_2453,In_1933);
nand U775 (N_775,N_124,N_149);
and U776 (N_776,N_396,In_103);
nand U777 (N_777,N_159,In_1620);
nand U778 (N_778,N_64,N_282);
nand U779 (N_779,N_36,N_293);
or U780 (N_780,In_747,In_2232);
xnor U781 (N_781,N_301,In_483);
nand U782 (N_782,In_897,N_418);
xnor U783 (N_783,N_234,In_1657);
and U784 (N_784,In_515,In_1903);
and U785 (N_785,N_411,In_1136);
nand U786 (N_786,In_754,N_182);
xor U787 (N_787,In_730,In_1292);
and U788 (N_788,In_1388,N_298);
and U789 (N_789,N_102,In_75);
nor U790 (N_790,N_79,In_1949);
or U791 (N_791,N_125,In_1920);
nor U792 (N_792,In_1811,N_179);
nand U793 (N_793,In_2172,In_1865);
xnor U794 (N_794,In_1176,In_108);
and U795 (N_795,N_356,In_702);
nand U796 (N_796,In_672,In_1932);
nor U797 (N_797,In_369,In_52);
nor U798 (N_798,In_1839,In_1452);
nor U799 (N_799,In_1663,In_1271);
nand U800 (N_800,In_744,N_200);
nand U801 (N_801,In_1248,N_424);
nor U802 (N_802,N_3,In_1454);
or U803 (N_803,In_1493,In_996);
and U804 (N_804,N_479,In_835);
and U805 (N_805,In_1554,In_211);
nand U806 (N_806,N_348,N_37);
nand U807 (N_807,In_194,N_60);
nand U808 (N_808,N_45,In_1676);
xor U809 (N_809,In_303,In_1466);
xor U810 (N_810,N_485,In_1565);
and U811 (N_811,N_81,In_2178);
and U812 (N_812,In_1940,In_1517);
nand U813 (N_813,In_1137,N_253);
or U814 (N_814,N_209,In_1792);
and U815 (N_815,In_2141,In_1585);
nor U816 (N_816,In_1534,In_1050);
or U817 (N_817,In_1668,In_10);
nand U818 (N_818,N_406,N_229);
or U819 (N_819,In_1075,N_164);
xor U820 (N_820,In_1353,In_2);
nor U821 (N_821,N_422,In_1957);
nand U822 (N_822,In_573,In_1680);
xnor U823 (N_823,In_157,In_1781);
nor U824 (N_824,N_65,In_1867);
nand U825 (N_825,In_207,In_1015);
nor U826 (N_826,In_2344,N_85);
xnor U827 (N_827,In_906,In_2150);
nor U828 (N_828,In_536,In_1108);
nand U829 (N_829,In_2329,In_421);
and U830 (N_830,In_2154,In_2059);
or U831 (N_831,In_1099,In_935);
nand U832 (N_832,In_125,In_2489);
xnor U833 (N_833,In_1971,In_74);
nand U834 (N_834,In_2077,In_4);
or U835 (N_835,N_136,N_464);
xor U836 (N_836,In_1521,N_6);
nand U837 (N_837,In_2385,In_846);
nor U838 (N_838,In_907,In_2390);
or U839 (N_839,In_2497,In_159);
and U840 (N_840,N_117,N_141);
xnor U841 (N_841,In_1473,In_2088);
xnor U842 (N_842,In_128,In_336);
and U843 (N_843,In_1098,In_249);
xor U844 (N_844,In_2288,N_236);
or U845 (N_845,In_1701,N_393);
and U846 (N_846,In_1155,In_1051);
nand U847 (N_847,In_2322,In_957);
and U848 (N_848,N_254,N_312);
nand U849 (N_849,N_249,In_1410);
xnor U850 (N_850,In_2269,N_50);
nand U851 (N_851,In_1764,N_402);
nor U852 (N_852,In_1052,In_1090);
nor U853 (N_853,In_1637,In_775);
or U854 (N_854,In_937,In_1728);
and U855 (N_855,In_1584,In_557);
and U856 (N_856,In_1334,In_1252);
xnor U857 (N_857,N_110,In_1419);
xnor U858 (N_858,In_213,N_345);
or U859 (N_859,N_470,In_1883);
nor U860 (N_860,In_784,In_1348);
nand U861 (N_861,In_1079,In_112);
or U862 (N_862,In_2337,In_1397);
and U863 (N_863,In_223,N_291);
nand U864 (N_864,In_953,In_2391);
or U865 (N_865,N_255,In_660);
nand U866 (N_866,In_624,In_3);
and U867 (N_867,In_2307,In_1691);
nand U868 (N_868,In_276,In_335);
or U869 (N_869,In_1453,In_695);
nor U870 (N_870,In_724,In_1081);
or U871 (N_871,In_1523,In_2000);
and U872 (N_872,In_1907,In_1793);
and U873 (N_873,In_517,In_1285);
nor U874 (N_874,N_34,N_139);
xor U875 (N_875,In_1345,N_364);
and U876 (N_876,In_1371,N_388);
xnor U877 (N_877,In_647,In_2155);
xnor U878 (N_878,N_183,N_19);
and U879 (N_879,In_109,In_2131);
xor U880 (N_880,In_2112,N_173);
nor U881 (N_881,N_47,In_1821);
or U882 (N_882,In_2074,In_527);
xor U883 (N_883,N_142,In_1752);
or U884 (N_884,In_459,In_2230);
or U885 (N_885,In_1740,In_2280);
xnor U886 (N_886,In_399,In_2053);
xnor U887 (N_887,N_243,In_1391);
xor U888 (N_888,In_353,In_844);
nor U889 (N_889,In_400,N_375);
xor U890 (N_890,In_349,In_1844);
nand U891 (N_891,In_920,N_399);
nor U892 (N_892,In_1788,In_971);
or U893 (N_893,N_153,In_1425);
and U894 (N_894,In_1006,In_241);
nand U895 (N_895,In_193,In_2139);
nand U896 (N_896,N_166,In_172);
nand U897 (N_897,In_1278,In_2138);
xnor U898 (N_898,In_533,In_1507);
or U899 (N_899,In_413,In_1667);
nand U900 (N_900,In_2442,In_129);
nor U901 (N_901,N_334,N_326);
or U902 (N_902,In_879,In_1284);
and U903 (N_903,In_393,In_1518);
nor U904 (N_904,In_126,In_981);
nor U905 (N_905,N_458,In_1373);
nand U906 (N_906,N_130,N_315);
nor U907 (N_907,In_163,In_1946);
nor U908 (N_908,In_86,In_150);
nor U909 (N_909,In_1706,In_1166);
or U910 (N_910,N_289,In_2005);
nor U911 (N_911,In_1955,In_2443);
and U912 (N_912,In_1272,In_1586);
nor U913 (N_913,In_401,N_268);
xor U914 (N_914,In_1996,N_332);
and U915 (N_915,In_603,N_305);
or U916 (N_916,N_207,In_938);
nand U917 (N_917,In_554,In_283);
xnor U918 (N_918,In_1985,In_2261);
xnor U919 (N_919,In_2434,In_2170);
or U920 (N_920,N_487,In_1293);
and U921 (N_921,In_1823,In_1837);
or U922 (N_922,In_903,In_1210);
nor U923 (N_923,N_203,In_202);
xor U924 (N_924,N_97,In_2281);
and U925 (N_925,In_1288,In_176);
nand U926 (N_926,In_611,In_1872);
xnor U927 (N_927,In_2410,N_372);
or U928 (N_928,In_1022,In_1943);
nand U929 (N_929,N_163,In_494);
nand U930 (N_930,N_310,N_271);
nand U931 (N_931,N_256,In_2469);
xor U932 (N_932,In_145,N_67);
or U933 (N_933,N_453,In_1994);
or U934 (N_934,In_373,In_2235);
xor U935 (N_935,In_273,N_331);
xor U936 (N_936,In_1456,N_20);
xnor U937 (N_937,In_735,In_405);
nor U938 (N_938,In_524,In_1980);
xor U939 (N_939,In_358,In_155);
and U940 (N_940,N_286,In_1337);
nor U941 (N_941,In_215,N_300);
nand U942 (N_942,In_417,In_1372);
xor U943 (N_943,N_459,In_940);
nor U944 (N_944,In_101,In_1655);
and U945 (N_945,In_2365,In_1187);
nor U946 (N_946,In_287,N_39);
and U947 (N_947,In_802,In_365);
xor U948 (N_948,N_48,In_191);
xor U949 (N_949,In_492,In_1224);
and U950 (N_950,In_915,In_1561);
nor U951 (N_951,In_1380,In_255);
and U952 (N_952,N_66,In_28);
nor U953 (N_953,In_1974,In_2432);
or U954 (N_954,In_652,N_454);
nand U955 (N_955,In_1938,In_1253);
and U956 (N_956,N_75,N_143);
xor U957 (N_957,In_1924,N_80);
xor U958 (N_958,In_2257,In_1950);
nand U959 (N_959,N_314,N_84);
xnor U960 (N_960,In_1928,N_244);
and U961 (N_961,N_51,In_1711);
and U962 (N_962,In_1721,In_1548);
nor U963 (N_963,In_201,In_993);
or U964 (N_964,N_9,In_296);
or U965 (N_965,In_2086,In_991);
or U966 (N_966,In_1227,In_663);
and U967 (N_967,In_1179,N_281);
nor U968 (N_968,In_1282,In_2247);
xnor U969 (N_969,N_225,N_54);
or U970 (N_970,In_7,In_2160);
nand U971 (N_971,In_2400,In_581);
nand U972 (N_972,In_1395,In_1712);
or U973 (N_973,N_49,In_1086);
nor U974 (N_974,N_233,In_2392);
nor U975 (N_975,In_2134,In_1186);
nor U976 (N_976,In_960,N_444);
xor U977 (N_977,In_1540,In_738);
and U978 (N_978,In_1460,In_1115);
xor U979 (N_979,In_1012,N_370);
nor U980 (N_980,In_1040,In_495);
nand U981 (N_981,In_473,N_29);
xor U982 (N_982,N_40,In_636);
or U983 (N_983,In_1824,In_50);
xor U984 (N_984,In_1906,In_2323);
nor U985 (N_985,In_73,N_160);
nand U986 (N_986,In_1494,N_194);
or U987 (N_987,In_468,In_815);
xor U988 (N_988,In_1393,In_2194);
nor U989 (N_989,In_1427,In_412);
and U990 (N_990,In_1385,In_2423);
and U991 (N_991,In_1511,In_35);
and U992 (N_992,In_1891,In_445);
xor U993 (N_993,In_444,N_127);
and U994 (N_994,In_685,In_2173);
xnor U995 (N_995,In_1390,N_329);
xor U996 (N_996,In_1780,In_1007);
nand U997 (N_997,In_593,In_1002);
nand U998 (N_998,In_1689,In_2387);
and U999 (N_999,In_549,In_2042);
nor U1000 (N_1000,In_1355,In_1377);
or U1001 (N_1001,N_735,In_1799);
or U1002 (N_1002,N_504,N_759);
nor U1003 (N_1003,In_293,N_442);
and U1004 (N_1004,N_392,N_644);
nand U1005 (N_1005,In_1161,N_643);
xnor U1006 (N_1006,In_714,In_1435);
and U1007 (N_1007,In_2376,In_2332);
and U1008 (N_1008,N_566,N_515);
nand U1009 (N_1009,N_636,N_852);
nor U1010 (N_1010,N_708,N_563);
and U1011 (N_1011,In_1044,In_553);
nor U1012 (N_1012,In_858,N_811);
nor U1013 (N_1013,N_232,N_23);
and U1014 (N_1014,In_485,In_1123);
and U1015 (N_1015,In_1207,N_73);
or U1016 (N_1016,In_740,In_1472);
and U1017 (N_1017,N_496,In_537);
or U1018 (N_1018,N_920,In_944);
or U1019 (N_1019,N_618,N_799);
and U1020 (N_1020,In_2362,N_351);
or U1021 (N_1021,In_114,In_1566);
xnor U1022 (N_1022,In_1150,N_899);
or U1023 (N_1023,In_179,N_378);
nand U1024 (N_1024,N_775,N_371);
xor U1025 (N_1025,In_2314,N_647);
xor U1026 (N_1026,N_841,N_555);
nand U1027 (N_1027,In_117,In_439);
xnor U1028 (N_1028,In_701,In_61);
xor U1029 (N_1029,In_2057,In_224);
nand U1030 (N_1030,In_184,N_581);
and U1031 (N_1031,N_813,In_1850);
nor U1032 (N_1032,N_22,In_1609);
nand U1033 (N_1033,In_2051,In_2480);
xnor U1034 (N_1034,In_2147,In_2273);
or U1035 (N_1035,N_526,N_746);
nand U1036 (N_1036,In_514,N_358);
xor U1037 (N_1037,N_877,In_2466);
nand U1038 (N_1038,N_651,N_503);
and U1039 (N_1039,In_2226,In_756);
and U1040 (N_1040,N_936,N_664);
and U1041 (N_1041,In_2364,In_795);
and U1042 (N_1042,In_1629,N_911);
xor U1043 (N_1043,N_559,In_1599);
nor U1044 (N_1044,N_21,N_957);
nand U1045 (N_1045,N_621,In_1229);
nand U1046 (N_1046,N_712,In_2490);
and U1047 (N_1047,In_1758,N_237);
nand U1048 (N_1048,In_1786,N_944);
xnor U1049 (N_1049,In_843,N_46);
or U1050 (N_1050,In_1688,In_396);
xor U1051 (N_1051,N_122,N_473);
xnor U1052 (N_1052,N_208,In_1095);
xnor U1053 (N_1053,N_238,N_630);
xor U1054 (N_1054,In_1868,N_951);
nand U1055 (N_1055,In_1379,N_678);
or U1056 (N_1056,N_886,In_455);
or U1057 (N_1057,N_603,N_145);
or U1058 (N_1058,In_829,N_280);
nor U1059 (N_1059,In_225,In_43);
nor U1060 (N_1060,In_631,In_2078);
or U1061 (N_1061,In_696,N_781);
or U1062 (N_1062,N_716,In_671);
nand U1063 (N_1063,N_963,N_865);
or U1064 (N_1064,N_639,N_681);
or U1065 (N_1065,N_349,N_706);
nand U1066 (N_1066,In_1809,In_1258);
or U1067 (N_1067,N_462,N_953);
and U1068 (N_1068,In_832,N_929);
xnor U1069 (N_1069,In_1069,N_985);
and U1070 (N_1070,In_387,In_862);
or U1071 (N_1071,In_1443,N_491);
nor U1072 (N_1072,In_1730,N_631);
nand U1073 (N_1073,N_753,In_477);
or U1074 (N_1074,In_21,In_2409);
xnor U1075 (N_1075,N_762,In_2210);
nor U1076 (N_1076,In_341,In_1499);
nor U1077 (N_1077,In_962,In_2335);
or U1078 (N_1078,In_1755,In_1049);
nor U1079 (N_1079,N_825,In_591);
xnor U1080 (N_1080,N_941,In_743);
or U1081 (N_1081,In_2482,N_216);
or U1082 (N_1082,N_7,N_763);
nand U1083 (N_1083,In_362,In_1122);
and U1084 (N_1084,N_380,N_507);
and U1085 (N_1085,In_106,N_614);
or U1086 (N_1086,In_132,N_74);
xnor U1087 (N_1087,In_1487,N_520);
or U1088 (N_1088,N_864,N_844);
nor U1089 (N_1089,In_254,In_1054);
and U1090 (N_1090,N_645,In_416);
nor U1091 (N_1091,In_1180,In_415);
nor U1092 (N_1092,N_798,N_896);
nor U1093 (N_1093,N_887,N_922);
nor U1094 (N_1094,In_1008,In_1036);
xnor U1095 (N_1095,In_575,N_854);
nor U1096 (N_1096,N_308,In_37);
nand U1097 (N_1097,N_275,N_686);
or U1098 (N_1098,N_795,N_318);
xor U1099 (N_1099,N_632,N_468);
and U1100 (N_1100,In_80,N_794);
nor U1101 (N_1101,In_522,N_637);
nor U1102 (N_1102,In_670,In_2479);
nand U1103 (N_1103,In_1412,In_665);
nor U1104 (N_1104,In_1387,In_578);
or U1105 (N_1105,N_307,In_2447);
or U1106 (N_1106,In_2182,In_988);
nor U1107 (N_1107,In_2140,N_867);
and U1108 (N_1108,In_642,In_81);
nor U1109 (N_1109,N_688,N_505);
nand U1110 (N_1110,N_498,N_940);
or U1111 (N_1111,N_816,N_982);
or U1112 (N_1112,N_436,In_662);
xnor U1113 (N_1113,In_2018,N_152);
or U1114 (N_1114,In_772,N_933);
and U1115 (N_1115,N_912,N_913);
nand U1116 (N_1116,In_2436,N_44);
xor U1117 (N_1117,N_433,N_999);
or U1118 (N_1118,In_378,In_1685);
xnor U1119 (N_1119,In_1616,N_668);
xnor U1120 (N_1120,N_569,N_873);
xor U1121 (N_1121,In_1952,N_741);
or U1122 (N_1122,In_327,N_613);
or U1123 (N_1123,In_1217,N_998);
or U1124 (N_1124,N_336,In_355);
nor U1125 (N_1125,N_128,In_1634);
and U1126 (N_1126,In_1197,N_987);
or U1127 (N_1127,In_1632,In_134);
and U1128 (N_1128,In_2114,In_625);
or U1129 (N_1129,N_455,In_2389);
xnor U1130 (N_1130,N_144,In_1376);
nand U1131 (N_1131,In_2360,N_304);
nor U1132 (N_1132,In_1717,In_1997);
nand U1133 (N_1133,N_748,In_914);
nor U1134 (N_1134,In_761,N_705);
and U1135 (N_1135,N_542,N_368);
and U1136 (N_1136,In_167,N_492);
nor U1137 (N_1137,In_547,N_376);
or U1138 (N_1138,In_778,In_22);
and U1139 (N_1139,N_437,N_457);
nor U1140 (N_1140,In_62,N_616);
nand U1141 (N_1141,N_549,N_568);
or U1142 (N_1142,N_155,In_510);
nand U1143 (N_1143,N_885,N_840);
xor U1144 (N_1144,N_792,N_342);
or U1145 (N_1145,In_762,N_374);
or U1146 (N_1146,N_397,In_947);
nand U1147 (N_1147,In_833,In_1869);
nand U1148 (N_1148,N_584,N_874);
nor U1149 (N_1149,In_1698,N_607);
xor U1150 (N_1150,In_300,N_989);
nand U1151 (N_1151,N_964,N_528);
or U1152 (N_1152,In_800,N_786);
and U1153 (N_1153,In_2165,N_962);
nor U1154 (N_1154,In_2291,In_2201);
and U1155 (N_1155,N_395,N_10);
nor U1156 (N_1156,In_2354,N_721);
or U1157 (N_1157,N_720,N_711);
nor U1158 (N_1158,In_550,N_671);
and U1159 (N_1159,N_685,In_2179);
xnor U1160 (N_1160,N_837,N_541);
nor U1161 (N_1161,N_502,In_169);
xor U1162 (N_1162,N_57,In_1130);
nand U1163 (N_1163,In_203,N_414);
xor U1164 (N_1164,In_1800,N_273);
or U1165 (N_1165,In_2202,In_2399);
and U1166 (N_1166,N_615,N_652);
xor U1167 (N_1167,In_1736,N_946);
nand U1168 (N_1168,In_1954,In_425);
nand U1169 (N_1169,N_13,In_466);
nor U1170 (N_1170,N_517,In_939);
nand U1171 (N_1171,N_585,N_25);
or U1172 (N_1172,N_465,In_1875);
nand U1173 (N_1173,In_2481,In_2193);
nor U1174 (N_1174,In_793,In_2024);
nand U1175 (N_1175,In_1512,N_177);
and U1176 (N_1176,In_2065,N_627);
or U1177 (N_1177,N_861,N_829);
nor U1178 (N_1178,N_959,N_169);
nor U1179 (N_1179,N_635,In_2477);
xor U1180 (N_1180,In_1267,In_1296);
and U1181 (N_1181,In_110,N_551);
and U1182 (N_1182,In_2301,In_220);
nand U1183 (N_1183,In_2205,In_1212);
nand U1184 (N_1184,N_608,In_1913);
nor U1185 (N_1185,In_1877,In_1801);
nand U1186 (N_1186,N_834,In_1763);
nand U1187 (N_1187,In_246,In_1005);
xnor U1188 (N_1188,In_384,N_277);
or U1189 (N_1189,In_917,N_649);
xor U1190 (N_1190,N_682,N_343);
xnor U1191 (N_1191,In_674,N_659);
or U1192 (N_1192,N_790,In_1894);
nor U1193 (N_1193,N_564,N_709);
or U1194 (N_1194,In_955,N_880);
or U1195 (N_1195,N_772,In_361);
and U1196 (N_1196,N_481,N_983);
nand U1197 (N_1197,In_1060,In_2440);
nor U1198 (N_1198,In_1720,In_91);
nor U1199 (N_1199,In_347,In_729);
xor U1200 (N_1200,N_93,N_116);
or U1201 (N_1201,In_1318,N_88);
and U1202 (N_1202,In_1537,In_1732);
and U1203 (N_1203,In_469,N_697);
or U1204 (N_1204,N_739,In_1772);
or U1205 (N_1205,In_659,In_856);
xor U1206 (N_1206,In_60,N_525);
and U1207 (N_1207,N_204,N_819);
or U1208 (N_1208,In_2191,N_224);
nand U1209 (N_1209,N_910,In_2300);
nand U1210 (N_1210,In_142,In_115);
or U1211 (N_1211,N_172,In_818);
xor U1212 (N_1212,In_263,N_698);
xor U1213 (N_1213,N_995,N_599);
xor U1214 (N_1214,N_562,In_1134);
or U1215 (N_1215,In_814,In_1324);
nor U1216 (N_1216,In_1843,N_118);
nor U1217 (N_1217,N_620,In_2118);
nand U1218 (N_1218,N_95,In_1670);
nand U1219 (N_1219,N_810,N_530);
nor U1220 (N_1220,In_1369,N_101);
and U1221 (N_1221,N_86,N_494);
nor U1222 (N_1222,N_70,N_245);
xor U1223 (N_1223,In_82,In_1402);
or U1224 (N_1224,In_277,In_270);
nor U1225 (N_1225,N_31,N_24);
nor U1226 (N_1226,In_2428,In_1777);
nand U1227 (N_1227,N_972,In_1266);
nor U1228 (N_1228,N_901,In_337);
xor U1229 (N_1229,N_961,N_648);
nand U1230 (N_1230,In_1183,N_986);
nand U1231 (N_1231,In_1791,N_846);
or U1232 (N_1232,In_315,N_871);
or U1233 (N_1233,N_629,N_248);
or U1234 (N_1234,In_1930,In_420);
nor U1235 (N_1235,N_222,In_1359);
xor U1236 (N_1236,N_284,In_1148);
xnor U1237 (N_1237,N_662,N_429);
or U1238 (N_1238,In_2438,N_672);
or U1239 (N_1239,In_279,N_903);
or U1240 (N_1240,N_391,N_958);
nand U1241 (N_1241,N_676,N_993);
nor U1242 (N_1242,N_448,In_1570);
and U1243 (N_1243,In_967,N_98);
nor U1244 (N_1244,In_2031,N_103);
or U1245 (N_1245,N_131,In_102);
nor U1246 (N_1246,In_1077,N_217);
nor U1247 (N_1247,N_828,In_1856);
nand U1248 (N_1248,In_1697,N_833);
xnor U1249 (N_1249,In_2242,N_154);
nand U1250 (N_1250,In_925,In_837);
and U1251 (N_1251,In_694,In_168);
nand U1252 (N_1252,In_703,N_779);
and U1253 (N_1253,N_658,In_1887);
nor U1254 (N_1254,In_1276,In_2125);
and U1255 (N_1255,In_572,In_1942);
nand U1256 (N_1256,In_788,N_991);
xnor U1257 (N_1257,In_1323,N_715);
or U1258 (N_1258,In_1145,N_500);
and U1259 (N_1259,N_642,In_2437);
and U1260 (N_1260,In_1581,In_783);
and U1261 (N_1261,In_1871,N_596);
nand U1262 (N_1262,N_317,N_401);
nor U1263 (N_1263,In_1021,In_454);
or U1264 (N_1264,N_657,N_780);
nor U1265 (N_1265,N_624,In_200);
xor U1266 (N_1266,N_450,In_427);
xnor U1267 (N_1267,In_2030,N_690);
nand U1268 (N_1268,N_201,In_973);
nand U1269 (N_1269,In_1501,N_184);
nand U1270 (N_1270,N_730,In_1175);
or U1271 (N_1271,In_1536,N_666);
or U1272 (N_1272,N_789,N_868);
nor U1273 (N_1273,N_325,In_120);
xor U1274 (N_1274,In_2218,In_1944);
xor U1275 (N_1275,In_1916,N_853);
nand U1276 (N_1276,N_765,In_548);
or U1277 (N_1277,N_218,In_1447);
or U1278 (N_1278,N_992,N_809);
nand U1279 (N_1279,In_667,N_755);
xor U1280 (N_1280,In_523,N_510);
xor U1281 (N_1281,N_767,N_700);
nand U1282 (N_1282,N_701,In_2233);
or U1283 (N_1283,N_287,In_1437);
nor U1284 (N_1284,In_1366,N_855);
nor U1285 (N_1285,In_1602,In_1011);
and U1286 (N_1286,In_822,In_218);
nor U1287 (N_1287,N_717,In_816);
nor U1288 (N_1288,N_930,In_1899);
or U1289 (N_1289,N_533,In_1975);
and U1290 (N_1290,In_1331,In_1173);
nand U1291 (N_1291,N_752,N_751);
nand U1292 (N_1292,N_41,N_405);
xor U1293 (N_1293,In_1336,In_2262);
nand U1294 (N_1294,N_831,N_604);
nand U1295 (N_1295,In_198,N_778);
xnor U1296 (N_1296,In_885,N_921);
xnor U1297 (N_1297,In_1413,N_728);
and U1298 (N_1298,N_737,In_2289);
xor U1299 (N_1299,In_2491,N_419);
nor U1300 (N_1300,N_894,In_500);
xnor U1301 (N_1301,In_1806,In_13);
nor U1302 (N_1302,N_134,N_856);
nand U1303 (N_1303,In_2294,In_1696);
and U1304 (N_1304,N_197,In_1577);
and U1305 (N_1305,N_206,N_954);
xnor U1306 (N_1306,In_2189,In_1241);
nand U1307 (N_1307,N_540,N_302);
and U1308 (N_1308,In_1729,In_442);
or U1309 (N_1309,In_2418,N_313);
and U1310 (N_1310,In_1497,N_805);
nand U1311 (N_1311,In_2470,N_724);
nor U1312 (N_1312,In_604,In_2158);
nor U1313 (N_1313,N_650,In_2133);
nand U1314 (N_1314,In_745,N_394);
or U1315 (N_1315,In_291,In_1874);
nand U1316 (N_1316,In_430,N_800);
and U1317 (N_1317,In_1103,N_554);
and U1318 (N_1318,In_741,N_808);
nand U1319 (N_1319,In_1280,N_736);
nand U1320 (N_1320,In_1761,In_1251);
or U1321 (N_1321,N_960,In_1110);
or U1322 (N_1322,In_189,In_1111);
nor U1323 (N_1323,In_1827,In_65);
xor U1324 (N_1324,In_1693,N_605);
nand U1325 (N_1325,In_2275,N_482);
and U1326 (N_1326,In_919,N_994);
or U1327 (N_1327,N_768,In_1675);
and U1328 (N_1328,In_798,In_2108);
nor U1329 (N_1329,N_945,In_1406);
and U1330 (N_1330,In_2109,In_1767);
nor U1331 (N_1331,N_2,In_766);
or U1332 (N_1332,N_935,N_839);
xor U1333 (N_1333,In_2374,In_431);
nor U1334 (N_1334,In_2272,N_109);
or U1335 (N_1335,In_910,N_477);
or U1336 (N_1336,N_469,In_969);
nor U1337 (N_1337,N_320,N_710);
nor U1338 (N_1338,N_112,N_83);
and U1339 (N_1339,In_1244,In_789);
xor U1340 (N_1340,N_575,In_2420);
and U1341 (N_1341,In_699,In_1890);
and U1342 (N_1342,N_758,In_1631);
nor U1343 (N_1343,In_1026,In_70);
xor U1344 (N_1344,N_266,N_966);
and U1345 (N_1345,In_1910,In_978);
nor U1346 (N_1346,In_1420,In_2268);
or U1347 (N_1347,N_723,In_1349);
nand U1348 (N_1348,N_59,In_2012);
nand U1349 (N_1349,In_2313,In_2286);
nand U1350 (N_1350,N_955,In_1858);
or U1351 (N_1351,In_780,In_295);
or U1352 (N_1352,N_704,N_744);
nor U1353 (N_1353,N_889,N_522);
nor U1354 (N_1354,N_536,In_2357);
and U1355 (N_1355,In_1085,In_1156);
xnor U1356 (N_1356,N_743,In_2176);
nand U1357 (N_1357,In_2106,N_316);
or U1358 (N_1358,In_931,In_381);
nor U1359 (N_1359,In_2468,In_613);
or U1360 (N_1360,In_282,N_132);
and U1361 (N_1361,N_488,In_2380);
or U1362 (N_1362,N_597,N_570);
or U1363 (N_1363,In_307,N_740);
nand U1364 (N_1364,In_2373,N_272);
or U1365 (N_1365,In_71,In_2126);
or U1366 (N_1366,In_995,In_1945);
or U1367 (N_1367,In_1350,N_971);
and U1368 (N_1368,In_462,In_1325);
or U1369 (N_1369,N_661,In_539);
xor U1370 (N_1370,N_745,N_512);
nand U1371 (N_1371,N_818,In_946);
and U1372 (N_1372,In_1738,N_230);
and U1373 (N_1373,In_332,In_842);
and U1374 (N_1374,In_1725,N_196);
xor U1375 (N_1375,In_597,In_2465);
and U1376 (N_1376,N_663,N_490);
nor U1377 (N_1377,In_1909,N_761);
nand U1378 (N_1378,N_952,In_1564);
nor U1379 (N_1379,N_337,N_242);
xor U1380 (N_1380,N_56,N_410);
nand U1381 (N_1381,N_835,In_1257);
nor U1382 (N_1382,In_2421,In_1926);
nand U1383 (N_1383,In_901,N_412);
nor U1384 (N_1384,N_979,In_1127);
nor U1385 (N_1385,In_426,N_891);
xor U1386 (N_1386,N_299,In_1751);
xnor U1387 (N_1387,N_472,N_390);
xnor U1388 (N_1388,In_1690,In_344);
and U1389 (N_1389,N_580,In_38);
xnor U1390 (N_1390,In_863,In_1220);
nor U1391 (N_1391,N_689,N_670);
and U1392 (N_1392,In_2174,In_757);
xor U1393 (N_1393,In_1961,In_891);
xnor U1394 (N_1394,In_1070,In_823);
nand U1395 (N_1395,In_2405,N_990);
and U1396 (N_1396,In_1814,In_1822);
nand U1397 (N_1397,In_1741,N_417);
and U1398 (N_1398,N_876,In_958);
nor U1399 (N_1399,N_524,In_1862);
or U1400 (N_1400,N_446,In_171);
nand U1401 (N_1401,In_2087,N_732);
or U1402 (N_1402,In_911,N_626);
or U1403 (N_1403,In_1646,In_1719);
or U1404 (N_1404,N_211,N_228);
nand U1405 (N_1405,In_2246,In_1484);
nor U1406 (N_1406,In_2211,N_434);
nand U1407 (N_1407,N_633,N_537);
nand U1408 (N_1408,N_573,N_968);
and U1409 (N_1409,In_48,N_919);
nor U1410 (N_1410,N_674,In_64);
xor U1411 (N_1411,In_1601,In_322);
nand U1412 (N_1412,In_668,In_1163);
xor U1413 (N_1413,In_1264,N_415);
nand U1414 (N_1414,N_654,N_836);
xor U1415 (N_1415,N_719,N_679);
and U1416 (N_1416,N_589,In_1048);
nor U1417 (N_1417,N_221,In_2445);
nand U1418 (N_1418,N_981,N_947);
and U1419 (N_1419,In_2492,In_2066);
xor U1420 (N_1420,In_434,In_1557);
xnor U1421 (N_1421,In_42,N_114);
nor U1422 (N_1422,N_16,In_2009);
or U1423 (N_1423,N_906,N_774);
or U1424 (N_1424,In_1936,N_977);
nand U1425 (N_1425,In_165,N_926);
or U1426 (N_1426,In_325,In_1181);
or U1427 (N_1427,In_650,In_1748);
nand U1428 (N_1428,N_408,N_339);
nor U1429 (N_1429,N_550,In_1579);
or U1430 (N_1430,In_2196,N_557);
and U1431 (N_1431,In_1416,In_1259);
nor U1432 (N_1432,In_1589,N_148);
and U1433 (N_1433,N_793,N_279);
xnor U1434 (N_1434,In_1281,In_1810);
nand U1435 (N_1435,N_241,N_826);
nor U1436 (N_1436,In_2186,In_2279);
nand U1437 (N_1437,In_178,N_722);
nor U1438 (N_1438,In_1582,N_578);
xor U1439 (N_1439,N_235,N_428);
nand U1440 (N_1440,In_2067,N_851);
xor U1441 (N_1441,N_309,In_590);
and U1442 (N_1442,N_924,In_496);
xnor U1443 (N_1443,N_212,N_151);
xnor U1444 (N_1444,N_848,N_838);
nor U1445 (N_1445,N_214,N_545);
and U1446 (N_1446,In_1120,N_770);
nand U1447 (N_1447,In_1640,In_2006);
nand U1448 (N_1448,In_1617,N_749);
or U1449 (N_1449,In_1375,In_753);
nor U1450 (N_1450,In_93,N_565);
xor U1451 (N_1451,N_556,In_98);
nand U1452 (N_1452,N_609,N_942);
nand U1453 (N_1453,In_1787,In_429);
and U1454 (N_1454,N_872,N_593);
or U1455 (N_1455,N_489,In_1538);
xnor U1456 (N_1456,N_263,In_807);
and U1457 (N_1457,In_391,N_895);
nand U1458 (N_1458,In_1329,N_937);
xor U1459 (N_1459,N_467,N_634);
nor U1460 (N_1460,N_669,N_346);
nor U1461 (N_1461,In_2493,In_1543);
nor U1462 (N_1462,N_622,N_561);
and U1463 (N_1463,N_386,N_888);
nor U1464 (N_1464,N_692,In_1431);
nor U1465 (N_1465,N_544,In_2227);
xnor U1466 (N_1466,N_939,In_1794);
nand U1467 (N_1467,N_105,N_361);
xnor U1468 (N_1468,N_518,In_2417);
or U1469 (N_1469,In_540,N_750);
or U1470 (N_1470,In_1677,In_2212);
and U1471 (N_1471,N_617,N_628);
or U1472 (N_1472,In_87,N_731);
nor U1473 (N_1473,N_612,In_226);
nor U1474 (N_1474,N_156,In_1583);
xor U1475 (N_1475,In_2073,In_618);
and U1476 (N_1476,N_220,N_824);
nor U1477 (N_1477,In_1407,N_897);
and U1478 (N_1478,N_756,N_99);
and U1479 (N_1479,In_1988,N_858);
nor U1480 (N_1480,N_259,In_2220);
xor U1481 (N_1481,In_12,N_904);
nor U1482 (N_1482,N_725,N_907);
xnor U1483 (N_1483,N_623,In_44);
or U1484 (N_1484,N_381,In_1381);
or U1485 (N_1485,N_269,In_1474);
nand U1486 (N_1486,In_2025,N_969);
and U1487 (N_1487,N_178,In_600);
or U1488 (N_1488,N_905,In_1235);
nand U1489 (N_1489,In_1482,In_1237);
and U1490 (N_1490,N_860,N_534);
and U1491 (N_1491,In_1160,N_619);
and U1492 (N_1492,N_543,N_665);
and U1493 (N_1493,In_1654,In_328);
nor U1494 (N_1494,N_190,N_443);
nor U1495 (N_1495,In_1569,In_453);
nand U1496 (N_1496,N_538,In_2244);
and U1497 (N_1497,In_2485,In_19);
nor U1498 (N_1498,N_832,In_868);
and U1499 (N_1499,In_1896,N_572);
nor U1500 (N_1500,N_1416,N_967);
nand U1501 (N_1501,N_1179,N_1072);
xnor U1502 (N_1502,In_683,N_1366);
nor U1503 (N_1503,In_185,In_2484);
xor U1504 (N_1504,N_1350,N_1180);
nand U1505 (N_1505,N_546,N_129);
or U1506 (N_1506,N_703,N_1228);
xor U1507 (N_1507,N_973,N_1145);
and U1508 (N_1508,N_1139,N_1092);
and U1509 (N_1509,N_1182,N_696);
and U1510 (N_1510,N_1114,N_1144);
nor U1511 (N_1511,In_1828,N_191);
or U1512 (N_1512,N_529,In_1490);
or U1513 (N_1513,N_1481,N_785);
nor U1514 (N_1514,N_1442,N_1085);
xnor U1515 (N_1515,N_1287,N_1248);
nor U1516 (N_1516,N_1399,N_1002);
xnor U1517 (N_1517,N_1117,In_782);
or U1518 (N_1518,N_1334,In_351);
xnor U1519 (N_1519,N_1346,N_1116);
and U1520 (N_1520,N_1199,N_691);
and U1521 (N_1521,N_1371,N_519);
and U1522 (N_1522,N_1146,N_847);
nor U1523 (N_1523,N_1252,N_560);
or U1524 (N_1524,N_1455,N_92);
and U1525 (N_1525,N_787,N_1317);
or U1526 (N_1526,In_1900,In_599);
nor U1527 (N_1527,N_1439,N_1293);
nand U1528 (N_1528,N_606,N_452);
xor U1529 (N_1529,N_1438,N_1183);
and U1530 (N_1530,N_1196,N_1466);
xnor U1531 (N_1531,In_2386,N_1094);
and U1532 (N_1532,In_2414,In_2463);
nand U1533 (N_1533,N_1499,N_382);
nand U1534 (N_1534,N_1376,In_1106);
nand U1535 (N_1535,N_1386,In_1139);
nor U1536 (N_1536,N_1009,In_1826);
nor U1537 (N_1537,N_1381,In_39);
xor U1538 (N_1538,In_964,In_1972);
nor U1539 (N_1539,N_1225,In_692);
nor U1540 (N_1540,N_1149,N_1299);
and U1541 (N_1541,N_1148,In_306);
or U1542 (N_1542,N_1410,N_1383);
xor U1543 (N_1543,In_1727,N_695);
xnor U1544 (N_1544,N_1165,N_1233);
nand U1545 (N_1545,N_625,N_1471);
nor U1546 (N_1546,N_1461,N_1277);
and U1547 (N_1547,N_1043,N_1056);
nor U1548 (N_1548,N_729,In_1546);
or U1549 (N_1549,N_1104,N_1478);
nor U1550 (N_1550,N_1090,N_1074);
xor U1551 (N_1551,N_1375,N_760);
nand U1552 (N_1552,In_1344,N_174);
or U1553 (N_1553,In_1798,N_1367);
nor U1554 (N_1554,In_1999,In_154);
or U1555 (N_1555,N_558,N_1087);
or U1556 (N_1556,N_1185,N_324);
nand U1557 (N_1557,N_1053,In_1141);
and U1558 (N_1558,In_2494,N_1259);
nand U1559 (N_1559,N_777,N_1400);
and U1560 (N_1560,N_1156,In_2011);
nand U1561 (N_1561,N_592,N_495);
and U1562 (N_1562,In_733,N_683);
nand U1563 (N_1563,N_1262,N_400);
and U1564 (N_1564,N_1426,In_333);
xor U1565 (N_1565,N_1017,N_1073);
or U1566 (N_1566,N_1014,N_231);
nor U1567 (N_1567,N_1060,N_845);
xnor U1568 (N_1568,N_820,N_186);
nand U1569 (N_1569,In_1562,In_1656);
and U1570 (N_1570,N_582,N_1297);
nand U1571 (N_1571,N_1428,N_1464);
xnor U1572 (N_1572,N_1028,N_1331);
xnor U1573 (N_1573,N_1407,N_1440);
xor U1574 (N_1574,N_1362,In_1635);
xnor U1575 (N_1575,N_1058,N_1200);
xor U1576 (N_1576,N_1260,In_1948);
nand U1577 (N_1577,In_643,N_1134);
nor U1578 (N_1578,N_576,N_1035);
or U1579 (N_1579,N_600,N_1475);
nor U1580 (N_1580,N_694,N_274);
xor U1581 (N_1581,N_1451,In_1143);
and U1582 (N_1582,In_1216,N_1431);
and U1583 (N_1583,N_474,N_1025);
or U1584 (N_1584,N_1081,N_1445);
or U1585 (N_1585,N_1167,In_1885);
nand U1586 (N_1586,In_1840,N_984);
and U1587 (N_1587,N_506,In_1502);
nor U1588 (N_1588,In_78,N_673);
nand U1589 (N_1589,N_463,N_713);
or U1590 (N_1590,In_2116,N_553);
or U1591 (N_1591,N_1454,N_15);
nand U1592 (N_1592,N_771,N_684);
nor U1593 (N_1593,In_1226,In_1046);
or U1594 (N_1594,N_742,N_292);
nand U1595 (N_1595,N_1305,N_1359);
xor U1596 (N_1596,N_379,In_2375);
and U1597 (N_1597,In_1905,N_1192);
or U1598 (N_1598,N_976,N_863);
xor U1599 (N_1599,N_916,In_570);
nand U1600 (N_1600,N_1347,N_1234);
nand U1601 (N_1601,N_1155,In_6);
and U1602 (N_1602,In_122,N_1110);
or U1603 (N_1603,In_2064,N_523);
and U1604 (N_1604,N_1037,N_1364);
nand U1605 (N_1605,N_1276,N_1039);
nor U1606 (N_1606,N_1004,N_1460);
nand U1607 (N_1607,N_1449,N_1107);
nor U1608 (N_1608,N_1052,N_1265);
nor U1609 (N_1609,N_1207,N_928);
nor U1610 (N_1610,N_1477,In_774);
nor U1611 (N_1611,In_2224,N_1152);
nor U1612 (N_1612,N_1422,N_303);
or U1613 (N_1613,N_1418,N_773);
xor U1614 (N_1614,In_1087,In_1239);
and U1615 (N_1615,In_79,N_1082);
and U1616 (N_1616,N_532,N_591);
nand U1617 (N_1617,N_656,N_956);
nor U1618 (N_1618,N_1304,In_2397);
nor U1619 (N_1619,In_2378,N_1308);
nor U1620 (N_1620,In_314,In_1966);
and U1621 (N_1621,N_1088,In_1449);
or U1622 (N_1622,N_69,In_2452);
or U1623 (N_1623,In_2234,N_1242);
nor U1624 (N_1624,N_1336,In_247);
xnor U1625 (N_1625,N_1288,N_577);
nor U1626 (N_1626,In_491,N_707);
or U1627 (N_1627,In_601,In_1354);
xnor U1628 (N_1628,In_2207,In_457);
nor U1629 (N_1629,In_449,N_1111);
and U1630 (N_1630,N_574,N_1036);
nand U1631 (N_1631,N_181,N_1237);
or U1632 (N_1632,N_409,N_974);
nand U1633 (N_1633,N_1291,N_882);
xor U1634 (N_1634,N_754,N_1253);
and U1635 (N_1635,N_1032,N_601);
nor U1636 (N_1636,N_1197,N_687);
xor U1637 (N_1637,N_1459,N_1313);
nand U1638 (N_1638,N_1159,In_1941);
and U1639 (N_1639,N_247,N_1121);
or U1640 (N_1640,N_1250,In_1043);
or U1641 (N_1641,N_1153,N_416);
or U1642 (N_1642,N_499,N_104);
nor U1643 (N_1643,N_823,N_1143);
nand U1644 (N_1644,N_1423,N_1322);
and U1645 (N_1645,N_1390,N_1089);
nand U1646 (N_1646,N_321,In_645);
xor U1647 (N_1647,N_1370,N_1395);
nor U1648 (N_1648,N_1099,In_1144);
nor U1649 (N_1649,N_1470,N_586);
nor U1650 (N_1650,In_2045,In_1192);
and U1651 (N_1651,N_769,N_360);
nor U1652 (N_1652,In_1489,N_1224);
or U1653 (N_1653,In_2072,In_1485);
xor U1654 (N_1654,N_1493,N_1496);
xnor U1655 (N_1655,N_1137,In_1170);
nor U1656 (N_1656,N_1098,In_2355);
nand U1657 (N_1657,N_1108,N_590);
nor U1658 (N_1658,In_1196,N_1447);
nand U1659 (N_1659,N_513,N_1329);
xnor U1660 (N_1660,N_1208,N_1452);
nor U1661 (N_1661,N_948,N_497);
xor U1662 (N_1662,N_883,N_1055);
xnor U1663 (N_1663,N_1041,N_1078);
and U1664 (N_1664,In_1038,N_1086);
xnor U1665 (N_1665,N_1205,N_1427);
and U1666 (N_1666,In_2229,N_1118);
or U1667 (N_1667,In_928,N_806);
or U1668 (N_1668,N_571,N_1138);
nor U1669 (N_1669,N_1333,N_726);
xnor U1670 (N_1670,N_521,N_1097);
nand U1671 (N_1671,N_1273,N_1103);
xor U1672 (N_1672,N_478,N_1132);
xor U1673 (N_1673,In_2408,In_1779);
or U1674 (N_1674,In_2215,N_1136);
nand U1675 (N_1675,N_1169,N_1021);
or U1676 (N_1676,N_26,N_1266);
xor U1677 (N_1677,In_1270,N_1059);
xor U1678 (N_1678,In_1471,N_1275);
and U1679 (N_1679,In_1055,N_1189);
nand U1680 (N_1680,N_511,N_1236);
or U1681 (N_1681,In_640,N_988);
xnor U1682 (N_1682,N_1217,N_1332);
nor U1683 (N_1683,N_1093,N_1355);
nor U1684 (N_1684,In_403,N_862);
or U1685 (N_1685,In_258,In_951);
and U1686 (N_1686,N_1405,N_547);
nor U1687 (N_1687,N_1436,In_410);
xnor U1688 (N_1688,N_1430,N_949);
and U1689 (N_1689,N_917,N_1338);
xor U1690 (N_1690,N_1352,N_1193);
nand U1691 (N_1691,N_1022,N_1360);
or U1692 (N_1692,N_1221,N_1077);
or U1693 (N_1693,N_357,In_2091);
nor U1694 (N_1694,N_1176,N_1298);
nor U1695 (N_1695,N_1029,N_1489);
nor U1696 (N_1696,In_828,N_1498);
nor U1697 (N_1697,N_675,N_1315);
or U1698 (N_1698,N_1079,In_230);
nor U1699 (N_1699,N_1404,N_1320);
xnor U1700 (N_1700,N_1115,N_1323);
nor U1701 (N_1701,N_1421,N_340);
or U1702 (N_1702,N_660,N_934);
or U1703 (N_1703,In_827,In_1078);
nor U1704 (N_1704,N_1330,N_113);
nor U1705 (N_1705,N_655,In_137);
xnor U1706 (N_1706,N_1484,In_760);
and U1707 (N_1707,N_970,In_1922);
and U1708 (N_1708,N_1128,N_1141);
nor U1709 (N_1709,N_1160,N_1175);
nor U1710 (N_1710,N_323,N_1419);
and U1711 (N_1711,N_1168,N_1314);
and U1712 (N_1712,N_1201,N_646);
xor U1713 (N_1713,In_637,In_182);
nor U1714 (N_1714,N_965,N_4);
nand U1715 (N_1715,In_367,N_1268);
nor U1716 (N_1716,N_527,N_1063);
or U1717 (N_1717,In_1025,N_1034);
nand U1718 (N_1718,N_791,N_1384);
or U1719 (N_1719,N_1184,N_734);
or U1720 (N_1720,N_1414,N_1391);
and U1721 (N_1721,N_1321,N_1251);
nor U1722 (N_1722,N_1006,N_782);
nor U1723 (N_1723,N_1049,N_1164);
or U1724 (N_1724,In_1710,N_812);
or U1725 (N_1725,N_1046,In_1107);
nor U1726 (N_1726,N_1444,N_158);
nor U1727 (N_1727,N_1396,N_1429);
nand U1728 (N_1728,N_1497,N_1374);
or U1729 (N_1729,In_1001,In_913);
nor U1730 (N_1730,In_56,N_1337);
nand U1731 (N_1731,N_1120,N_1349);
or U1732 (N_1732,N_802,N_1354);
or U1733 (N_1733,N_1300,In_711);
nor U1734 (N_1734,N_1363,N_1129);
nand U1735 (N_1735,N_738,N_1051);
nand U1736 (N_1736,N_508,N_365);
nor U1737 (N_1737,N_1215,N_1246);
nor U1738 (N_1738,N_1406,N_1369);
xnor U1739 (N_1739,N_1212,N_1361);
and U1740 (N_1740,N_1038,In_758);
xnor U1741 (N_1741,In_1488,N_100);
nand U1742 (N_1742,N_902,In_2377);
or U1743 (N_1743,N_932,N_514);
nor U1744 (N_1744,N_1173,N_1412);
xnor U1745 (N_1745,N_137,In_1088);
xnor U1746 (N_1746,N_493,N_1019);
and U1747 (N_1747,N_1482,N_1177);
xnor U1748 (N_1748,N_1413,N_714);
or U1749 (N_1749,N_82,N_733);
nand U1750 (N_1750,In_1819,N_1171);
and U1751 (N_1751,N_1174,N_170);
and U1752 (N_1752,N_1408,N_1420);
nand U1753 (N_1753,In_563,N_1048);
or U1754 (N_1754,In_726,N_588);
and U1755 (N_1755,N_766,N_718);
or U1756 (N_1756,In_1880,N_1487);
xnor U1757 (N_1757,In_752,In_266);
and U1758 (N_1758,N_804,N_1325);
or U1759 (N_1759,N_1147,N_1324);
or U1760 (N_1760,N_892,N_1133);
and U1761 (N_1761,N_1318,N_1202);
and U1762 (N_1762,N_1388,N_461);
and U1763 (N_1763,N_1003,N_909);
nand U1764 (N_1764,In_1042,N_950);
xnor U1765 (N_1765,N_1062,In_162);
nand U1766 (N_1766,N_1295,N_1163);
nor U1767 (N_1767,N_185,N_1379);
nor U1768 (N_1768,In_2483,N_784);
nand U1769 (N_1769,N_579,N_1340);
xnor U1770 (N_1770,N_1378,N_1424);
nor U1771 (N_1771,N_451,N_1124);
nand U1772 (N_1772,N_1240,N_1382);
xor U1773 (N_1773,N_1393,In_27);
nor U1774 (N_1774,N_875,N_1031);
nand U1775 (N_1775,N_1284,N_1229);
nand U1776 (N_1776,In_359,In_2238);
or U1777 (N_1777,N_878,In_2407);
nor U1778 (N_1778,N_1270,N_1067);
nand U1779 (N_1779,In_164,N_404);
and U1780 (N_1780,In_877,N_1227);
nand U1781 (N_1781,N_1280,In_2487);
nand U1782 (N_1782,N_1071,N_1070);
nand U1783 (N_1783,N_535,N_699);
nor U1784 (N_1784,N_1373,N_610);
nor U1785 (N_1785,N_898,N_822);
and U1786 (N_1786,N_1095,N_1294);
nor U1787 (N_1787,N_1178,N_1433);
nor U1788 (N_1788,In_1428,In_8);
nand U1789 (N_1789,N_869,N_1096);
and U1790 (N_1790,In_1705,N_827);
xnor U1791 (N_1791,N_1050,N_140);
or U1792 (N_1792,N_1342,N_1007);
nand U1793 (N_1793,In_1114,N_702);
xor U1794 (N_1794,N_975,N_595);
and U1795 (N_1795,N_1278,In_1866);
and U1796 (N_1796,N_583,N_1448);
xnor U1797 (N_1797,N_927,N_1474);
or U1798 (N_1798,In_1310,N_1011);
nor U1799 (N_1799,N_1186,In_34);
or U1800 (N_1800,N_1476,N_1279);
and U1801 (N_1801,N_1457,In_1432);
or U1802 (N_1802,N_1075,In_1833);
nor U1803 (N_1803,N_859,N_1190);
and U1804 (N_1804,In_1855,N_1286);
xnor U1805 (N_1805,N_1468,In_2367);
and U1806 (N_1806,In_1004,N_1380);
xor U1807 (N_1807,N_1387,N_205);
nor U1808 (N_1808,N_1319,N_1432);
nor U1809 (N_1809,N_267,N_843);
xor U1810 (N_1810,In_875,N_1020);
and U1811 (N_1811,N_1045,N_1102);
nand U1812 (N_1812,N_796,In_1313);
nor U1813 (N_1813,N_1301,N_165);
nand U1814 (N_1814,N_1327,In_2110);
xor U1815 (N_1815,In_1073,N_1126);
or U1816 (N_1816,N_1398,N_1030);
xnor U1817 (N_1817,N_1013,N_1341);
xnor U1818 (N_1818,N_1491,In_1759);
nand U1819 (N_1819,N_1113,N_567);
nor U1820 (N_1820,N_192,N_1109);
or U1821 (N_1821,N_1213,N_1467);
nand U1822 (N_1822,In_796,N_1219);
nand U1823 (N_1823,N_1245,In_478);
nand U1824 (N_1824,N_1024,N_1065);
xnor U1825 (N_1825,In_2225,In_1979);
xnor U1826 (N_1826,N_1027,In_1392);
or U1827 (N_1827,N_1310,N_1040);
or U1828 (N_1828,In_68,N_1122);
nand U1829 (N_1829,N_1490,In_1019);
xnor U1830 (N_1830,N_641,In_40);
or U1831 (N_1831,In_2146,N_1135);
or U1832 (N_1832,In_1340,N_693);
nand U1833 (N_1833,N_1083,N_501);
nor U1834 (N_1834,In_274,N_1033);
nor U1835 (N_1835,N_594,N_1472);
xor U1836 (N_1836,N_198,In_1135);
or U1837 (N_1837,N_1264,In_338);
nand U1838 (N_1838,N_1057,N_757);
nand U1839 (N_1839,In_2282,In_1275);
nand U1840 (N_1840,In_1986,N_1339);
xor U1841 (N_1841,N_817,N_638);
or U1842 (N_1842,N_440,In_1068);
and U1843 (N_1843,N_1326,N_1042);
nor U1844 (N_1844,N_1256,N_1204);
nand U1845 (N_1845,In_794,N_539);
and U1846 (N_1846,N_260,In_1818);
and U1847 (N_1847,N_1344,In_1061);
nor U1848 (N_1848,N_1403,N_1158);
or U1849 (N_1849,N_1417,N_1357);
nand U1850 (N_1850,N_1473,N_423);
and U1851 (N_1851,N_531,In_136);
and U1852 (N_1852,In_1389,N_1054);
nor U1853 (N_1853,N_1151,In_2431);
xor U1854 (N_1854,In_2312,N_157);
or U1855 (N_1855,N_1091,N_1008);
nor U1856 (N_1856,In_1236,N_925);
and U1857 (N_1857,N_1131,N_1209);
or U1858 (N_1858,N_1267,N_1306);
nand U1859 (N_1859,N_943,N_438);
nand U1860 (N_1860,In_2338,N_1450);
and U1861 (N_1861,In_848,In_1886);
nand U1862 (N_1862,N_1203,N_1492);
xnor U1863 (N_1863,N_1302,N_1235);
nand U1864 (N_1864,N_1232,N_1161);
and U1865 (N_1865,In_1965,N_1210);
xnor U1866 (N_1866,N_1018,N_1105);
xnor U1867 (N_1867,N_1112,N_908);
xor U1868 (N_1868,N_1150,In_1682);
nor U1869 (N_1869,N_830,In_260);
xor U1870 (N_1870,In_1465,N_1479);
nor U1871 (N_1871,N_265,In_1394);
or U1872 (N_1872,N_1191,N_1241);
nand U1873 (N_1873,N_803,N_449);
and U1874 (N_1874,N_1486,N_1000);
or U1875 (N_1875,N_1411,N_226);
nor U1876 (N_1876,N_1356,In_227);
and U1877 (N_1877,N_1206,N_432);
and U1878 (N_1878,In_773,In_1205);
or U1879 (N_1879,N_1194,In_506);
or U1880 (N_1880,N_189,N_1157);
nor U1881 (N_1881,N_814,N_842);
nand U1882 (N_1882,In_2021,N_866);
nor U1883 (N_1883,N_1365,N_1254);
and U1884 (N_1884,N_466,N_747);
nand U1885 (N_1885,N_1239,In_615);
nor U1886 (N_1886,N_1106,N_362);
or U1887 (N_1887,N_1368,N_850);
and U1888 (N_1888,N_1084,N_1140);
and U1889 (N_1889,N_1285,N_1230);
nor U1890 (N_1890,N_311,N_598);
xnor U1891 (N_1891,N_1425,N_1125);
nor U1892 (N_1892,N_1066,N_1443);
or U1893 (N_1893,N_1064,N_893);
nor U1894 (N_1894,N_1195,N_278);
and U1895 (N_1895,N_167,In_309);
xnor U1896 (N_1896,In_1092,N_1181);
nor U1897 (N_1897,N_918,N_1238);
nor U1898 (N_1898,N_776,N_1292);
or U1899 (N_1899,N_1012,N_1385);
or U1900 (N_1900,N_1290,N_1162);
and U1901 (N_1901,N_1166,In_1119);
xnor U1902 (N_1902,In_2013,N_1044);
or U1903 (N_1903,N_680,N_611);
nor U1904 (N_1904,In_72,N_1249);
nand U1905 (N_1905,N_1187,N_1076);
and U1906 (N_1906,In_1694,In_1515);
nand U1907 (N_1907,N_1345,N_330);
xnor U1908 (N_1908,N_1458,N_938);
or U1909 (N_1909,N_12,N_653);
or U1910 (N_1910,N_548,N_1453);
xor U1911 (N_1911,N_1296,N_1328);
or U1912 (N_1912,N_1001,N_1047);
and U1913 (N_1913,In_2104,N_1243);
nor U1914 (N_1914,N_257,N_1437);
and U1915 (N_1915,In_348,N_1061);
and U1916 (N_1916,N_849,N_1123);
nor U1917 (N_1917,N_997,N_1100);
nand U1918 (N_1918,In_216,N_1389);
nand U1919 (N_1919,N_1226,N_1495);
nand U1920 (N_1920,In_1214,N_1434);
and U1921 (N_1921,N_1335,N_807);
xnor U1922 (N_1922,N_1247,In_708);
nand U1923 (N_1923,N_1488,N_1446);
or U1924 (N_1924,N_1353,N_783);
nand U1925 (N_1925,N_1465,N_915);
nor U1926 (N_1926,N_270,In_1513);
and U1927 (N_1927,In_2403,N_900);
xor U1928 (N_1928,N_1343,In_204);
xnor U1929 (N_1929,In_160,N_58);
xnor U1930 (N_1930,N_788,N_797);
xnor U1931 (N_1931,In_1520,N_1401);
or U1932 (N_1932,In_1590,N_677);
or U1933 (N_1933,N_1377,N_1494);
xnor U1934 (N_1934,N_223,N_821);
or U1935 (N_1935,In_2062,In_280);
and U1936 (N_1936,N_602,N_1172);
or U1937 (N_1937,N_1272,N_1303);
nand U1938 (N_1938,In_1240,N_815);
nor U1939 (N_1939,N_1220,In_1133);
xnor U1940 (N_1940,In_1852,N_1281);
xor U1941 (N_1941,N_1469,In_505);
and U1942 (N_1942,N_667,N_1351);
and U1943 (N_1943,N_1392,N_328);
or U1944 (N_1944,N_1257,In_2100);
or U1945 (N_1945,N_1005,N_1023);
xnor U1946 (N_1946,N_727,N_857);
or U1947 (N_1947,In_850,N_923);
xor U1948 (N_1948,N_890,N_1142);
nand U1949 (N_1949,N_1218,N_1274);
nand U1950 (N_1950,N_1223,N_1188);
xor U1951 (N_1951,N_1080,N_1309);
and U1952 (N_1952,N_801,N_1068);
xor U1953 (N_1953,N_1312,N_1258);
xor U1954 (N_1954,N_1435,N_1069);
or U1955 (N_1955,N_1394,N_150);
nand U1956 (N_1956,N_870,In_1563);
nand U1957 (N_1957,N_1261,N_1211);
nand U1958 (N_1958,N_996,N_1222);
and U1959 (N_1959,In_1708,In_1530);
xnor U1960 (N_1960,N_1016,In_1808);
nand U1961 (N_1961,N_1263,N_1101);
xnor U1962 (N_1962,N_1283,N_1255);
or U1963 (N_1963,In_1102,N_1198);
nor U1964 (N_1964,N_1409,In_1097);
or U1965 (N_1965,In_985,In_1715);
nor U1966 (N_1966,In_1409,N_1154);
and U1967 (N_1967,In_1333,N_1463);
or U1968 (N_1968,N_980,N_640);
or U1969 (N_1969,N_251,N_1462);
nand U1970 (N_1970,N_1214,N_1119);
nor U1971 (N_1971,N_1372,N_1485);
nand U1972 (N_1972,N_1231,N_884);
and U1973 (N_1973,N_1127,N_1010);
or U1974 (N_1974,In_342,N_1316);
or U1975 (N_1975,N_1415,N_764);
and U1976 (N_1976,In_2429,N_1358);
nor U1977 (N_1977,N_914,N_1348);
xor U1978 (N_1978,N_355,N_53);
nand U1979 (N_1979,N_1289,N_931);
xnor U1980 (N_1980,N_1216,N_1307);
or U1981 (N_1981,N_1441,N_879);
nand U1982 (N_1982,N_1269,N_1015);
nand U1983 (N_1983,In_1514,N_1483);
nor U1984 (N_1984,N_587,In_1783);
or U1985 (N_1985,In_675,N_1170);
or U1986 (N_1986,In_1475,N_387);
nand U1987 (N_1987,N_509,N_94);
nand U1988 (N_1988,N_1244,In_2068);
or U1989 (N_1989,N_1026,In_1778);
nor U1990 (N_1990,N_552,In_1598);
xnor U1991 (N_1991,N_1456,N_1311);
nor U1992 (N_1992,In_475,N_8);
xor U1993 (N_1993,N_106,N_486);
nor U1994 (N_1994,N_516,N_881);
and U1995 (N_1995,N_1397,N_1271);
nand U1996 (N_1996,N_1282,N_1130);
or U1997 (N_1997,In_779,N_202);
and U1998 (N_1998,N_71,N_978);
nand U1999 (N_1999,N_1402,N_1480);
nand U2000 (N_2000,N_1646,N_1744);
and U2001 (N_2001,N_1791,N_1567);
nor U2002 (N_2002,N_1746,N_1750);
or U2003 (N_2003,N_1693,N_1639);
or U2004 (N_2004,N_1894,N_1900);
xnor U2005 (N_2005,N_1770,N_1829);
or U2006 (N_2006,N_1775,N_1505);
nor U2007 (N_2007,N_1534,N_1841);
nand U2008 (N_2008,N_1551,N_1546);
nor U2009 (N_2009,N_1988,N_1997);
nand U2010 (N_2010,N_1983,N_1709);
or U2011 (N_2011,N_1947,N_1718);
xor U2012 (N_2012,N_1805,N_1539);
and U2013 (N_2013,N_1656,N_1783);
xor U2014 (N_2014,N_1871,N_1712);
xnor U2015 (N_2015,N_1713,N_1765);
and U2016 (N_2016,N_1743,N_1967);
nand U2017 (N_2017,N_1984,N_1762);
or U2018 (N_2018,N_1819,N_1586);
nor U2019 (N_2019,N_1690,N_1549);
and U2020 (N_2020,N_1878,N_1961);
or U2021 (N_2021,N_1608,N_1589);
nor U2022 (N_2022,N_1563,N_1824);
nor U2023 (N_2023,N_1730,N_1973);
nand U2024 (N_2024,N_1521,N_1566);
nor U2025 (N_2025,N_1588,N_1859);
or U2026 (N_2026,N_1732,N_1647);
and U2027 (N_2027,N_1514,N_1554);
xor U2028 (N_2028,N_1526,N_1689);
or U2029 (N_2029,N_1501,N_1793);
and U2030 (N_2030,N_1842,N_1668);
nor U2031 (N_2031,N_1508,N_1923);
nand U2032 (N_2032,N_1748,N_1565);
or U2033 (N_2033,N_1834,N_1777);
or U2034 (N_2034,N_1917,N_1812);
xnor U2035 (N_2035,N_1694,N_1527);
or U2036 (N_2036,N_1616,N_1674);
nand U2037 (N_2037,N_1734,N_1627);
xnor U2038 (N_2038,N_1556,N_1665);
nand U2039 (N_2039,N_1700,N_1888);
and U2040 (N_2040,N_1768,N_1663);
nor U2041 (N_2041,N_1843,N_1632);
nand U2042 (N_2042,N_1965,N_1681);
nor U2043 (N_2043,N_1897,N_1810);
nor U2044 (N_2044,N_1679,N_1804);
or U2045 (N_2045,N_1745,N_1821);
xor U2046 (N_2046,N_1962,N_1517);
and U2047 (N_2047,N_1720,N_1981);
and U2048 (N_2048,N_1890,N_1908);
nand U2049 (N_2049,N_1999,N_1560);
or U2050 (N_2050,N_1672,N_1673);
xnor U2051 (N_2051,N_1500,N_1918);
xor U2052 (N_2052,N_1664,N_1895);
nor U2053 (N_2053,N_1938,N_1891);
or U2054 (N_2054,N_1741,N_1683);
or U2055 (N_2055,N_1598,N_1564);
or U2056 (N_2056,N_1740,N_1870);
and U2057 (N_2057,N_1574,N_1711);
nand U2058 (N_2058,N_1951,N_1789);
or U2059 (N_2059,N_1899,N_1570);
nor U2060 (N_2060,N_1807,N_1980);
nand U2061 (N_2061,N_1593,N_1503);
or U2062 (N_2062,N_1990,N_1728);
nand U2063 (N_2063,N_1725,N_1820);
or U2064 (N_2064,N_1902,N_1707);
xor U2065 (N_2065,N_1660,N_1544);
or U2066 (N_2066,N_1524,N_1912);
nor U2067 (N_2067,N_1848,N_1604);
nor U2068 (N_2068,N_1953,N_1630);
nor U2069 (N_2069,N_1957,N_1706);
nor U2070 (N_2070,N_1826,N_1607);
or U2071 (N_2071,N_1942,N_1787);
nor U2072 (N_2072,N_1628,N_1652);
nand U2073 (N_2073,N_1772,N_1766);
xnor U2074 (N_2074,N_1515,N_1946);
or U2075 (N_2075,N_1913,N_1635);
nor U2076 (N_2076,N_1619,N_1803);
nor U2077 (N_2077,N_1653,N_1576);
xnor U2078 (N_2078,N_1738,N_1520);
and U2079 (N_2079,N_1631,N_1506);
or U2080 (N_2080,N_1661,N_1833);
or U2081 (N_2081,N_1737,N_1698);
nand U2082 (N_2082,N_1531,N_1671);
nor U2083 (N_2083,N_1915,N_1816);
nor U2084 (N_2084,N_1776,N_1781);
nand U2085 (N_2085,N_1729,N_1756);
and U2086 (N_2086,N_1522,N_1782);
or U2087 (N_2087,N_1626,N_1778);
xnor U2088 (N_2088,N_1599,N_1600);
or U2089 (N_2089,N_1852,N_1795);
nand U2090 (N_2090,N_1755,N_1952);
or U2091 (N_2091,N_1922,N_1592);
and U2092 (N_2092,N_1930,N_1533);
xor U2093 (N_2093,N_1529,N_1949);
nand U2094 (N_2094,N_1623,N_1788);
nand U2095 (N_2095,N_1655,N_1977);
and U2096 (N_2096,N_1591,N_1507);
or U2097 (N_2097,N_1684,N_1525);
nand U2098 (N_2098,N_1995,N_1873);
nand U2099 (N_2099,N_1751,N_1892);
nor U2100 (N_2100,N_1864,N_1948);
nand U2101 (N_2101,N_1595,N_1644);
nand U2102 (N_2102,N_1569,N_1649);
nor U2103 (N_2103,N_1510,N_1794);
nor U2104 (N_2104,N_1889,N_1613);
xor U2105 (N_2105,N_1643,N_1699);
nand U2106 (N_2106,N_1686,N_1580);
xor U2107 (N_2107,N_1813,N_1611);
nand U2108 (N_2108,N_1722,N_1753);
or U2109 (N_2109,N_1637,N_1943);
xnor U2110 (N_2110,N_1519,N_1982);
or U2111 (N_2111,N_1759,N_1538);
nand U2112 (N_2112,N_1537,N_1928);
or U2113 (N_2113,N_1906,N_1676);
or U2114 (N_2114,N_1909,N_1861);
xor U2115 (N_2115,N_1840,N_1597);
or U2116 (N_2116,N_1638,N_1692);
xor U2117 (N_2117,N_1696,N_1811);
or U2118 (N_2118,N_1921,N_1955);
nor U2119 (N_2119,N_1670,N_1998);
nand U2120 (N_2120,N_1622,N_1513);
xnor U2121 (N_2121,N_1845,N_1979);
nor U2122 (N_2122,N_1809,N_1960);
xor U2123 (N_2123,N_1528,N_1991);
and U2124 (N_2124,N_1887,N_1761);
and U2125 (N_2125,N_1835,N_1907);
and U2126 (N_2126,N_1994,N_1937);
nand U2127 (N_2127,N_1872,N_1610);
nor U2128 (N_2128,N_1502,N_1735);
and U2129 (N_2129,N_1509,N_1971);
xor U2130 (N_2130,N_1704,N_1553);
and U2131 (N_2131,N_1799,N_1964);
nand U2132 (N_2132,N_1545,N_1881);
nand U2133 (N_2133,N_1936,N_1739);
nand U2134 (N_2134,N_1996,N_1587);
and U2135 (N_2135,N_1986,N_1710);
xnor U2136 (N_2136,N_1577,N_1987);
and U2137 (N_2137,N_1903,N_1769);
nor U2138 (N_2138,N_1877,N_1659);
xnor U2139 (N_2139,N_1924,N_1992);
or U2140 (N_2140,N_1701,N_1688);
xnor U2141 (N_2141,N_1633,N_1950);
xnor U2142 (N_2142,N_1780,N_1828);
nor U2143 (N_2143,N_1714,N_1880);
xnor U2144 (N_2144,N_1806,N_1562);
nand U2145 (N_2145,N_1849,N_1581);
nand U2146 (N_2146,N_1669,N_1944);
and U2147 (N_2147,N_1530,N_1940);
or U2148 (N_2148,N_1905,N_1721);
xnor U2149 (N_2149,N_1621,N_1797);
or U2150 (N_2150,N_1875,N_1733);
nand U2151 (N_2151,N_1682,N_1879);
or U2152 (N_2152,N_1963,N_1885);
nor U2153 (N_2153,N_1609,N_1926);
and U2154 (N_2154,N_1559,N_1540);
nand U2155 (N_2155,N_1723,N_1624);
and U2156 (N_2156,N_1650,N_1561);
or U2157 (N_2157,N_1667,N_1705);
or U2158 (N_2158,N_1516,N_1550);
nor U2159 (N_2159,N_1959,N_1792);
or U2160 (N_2160,N_1708,N_1754);
xnor U2161 (N_2161,N_1869,N_1954);
and U2162 (N_2162,N_1774,N_1945);
xor U2163 (N_2163,N_1867,N_1863);
nor U2164 (N_2164,N_1882,N_1583);
and U2165 (N_2165,N_1822,N_1974);
nand U2166 (N_2166,N_1697,N_1747);
nor U2167 (N_2167,N_1901,N_1886);
nand U2168 (N_2168,N_1585,N_1798);
nand U2169 (N_2169,N_1818,N_1830);
nand U2170 (N_2170,N_1978,N_1868);
nand U2171 (N_2171,N_1504,N_1796);
nand U2172 (N_2172,N_1853,N_1618);
xor U2173 (N_2173,N_1866,N_1985);
nand U2174 (N_2174,N_1941,N_1972);
or U2175 (N_2175,N_1839,N_1784);
xor U2176 (N_2176,N_1617,N_1658);
or U2177 (N_2177,N_1862,N_1717);
xor U2178 (N_2178,N_1636,N_1846);
or U2179 (N_2179,N_1858,N_1573);
nand U2180 (N_2180,N_1651,N_1956);
xor U2181 (N_2181,N_1851,N_1548);
or U2182 (N_2182,N_1874,N_1800);
nor U2183 (N_2183,N_1572,N_1703);
xnor U2184 (N_2184,N_1555,N_1685);
nand U2185 (N_2185,N_1929,N_1547);
and U2186 (N_2186,N_1865,N_1975);
xor U2187 (N_2187,N_1657,N_1629);
or U2188 (N_2188,N_1620,N_1677);
xor U2189 (N_2189,N_1838,N_1675);
xnor U2190 (N_2190,N_1634,N_1702);
xnor U2191 (N_2191,N_1808,N_1605);
nor U2192 (N_2192,N_1920,N_1640);
nor U2193 (N_2193,N_1823,N_1687);
nor U2194 (N_2194,N_1584,N_1582);
xor U2195 (N_2195,N_1541,N_1910);
xor U2196 (N_2196,N_1914,N_1844);
nand U2197 (N_2197,N_1736,N_1831);
or U2198 (N_2198,N_1976,N_1571);
and U2199 (N_2199,N_1535,N_1785);
xnor U2200 (N_2200,N_1898,N_1726);
and U2201 (N_2201,N_1814,N_1779);
or U2202 (N_2202,N_1856,N_1932);
nor U2203 (N_2203,N_1927,N_1645);
nand U2204 (N_2204,N_1578,N_1860);
nor U2205 (N_2205,N_1542,N_1641);
nor U2206 (N_2206,N_1802,N_1727);
or U2207 (N_2207,N_1742,N_1678);
nand U2208 (N_2208,N_1773,N_1933);
xor U2209 (N_2209,N_1764,N_1969);
xor U2210 (N_2210,N_1614,N_1966);
or U2211 (N_2211,N_1536,N_1786);
and U2212 (N_2212,N_1771,N_1857);
nand U2213 (N_2213,N_1716,N_1523);
or U2214 (N_2214,N_1854,N_1575);
xnor U2215 (N_2215,N_1817,N_1603);
xor U2216 (N_2216,N_1931,N_1836);
or U2217 (N_2217,N_1602,N_1579);
nand U2218 (N_2218,N_1758,N_1847);
xor U2219 (N_2219,N_1654,N_1752);
and U2220 (N_2220,N_1518,N_1893);
nor U2221 (N_2221,N_1731,N_1642);
and U2222 (N_2222,N_1557,N_1904);
and U2223 (N_2223,N_1648,N_1680);
nor U2224 (N_2224,N_1939,N_1695);
and U2225 (N_2225,N_1715,N_1968);
nand U2226 (N_2226,N_1876,N_1724);
or U2227 (N_2227,N_1993,N_1543);
xor U2228 (N_2228,N_1925,N_1790);
xnor U2229 (N_2229,N_1850,N_1615);
nor U2230 (N_2230,N_1911,N_1590);
nor U2231 (N_2231,N_1749,N_1825);
nor U2232 (N_2232,N_1662,N_1837);
and U2233 (N_2233,N_1883,N_1532);
nor U2234 (N_2234,N_1512,N_1601);
xnor U2235 (N_2235,N_1757,N_1855);
or U2236 (N_2236,N_1827,N_1989);
xor U2237 (N_2237,N_1596,N_1815);
and U2238 (N_2238,N_1691,N_1916);
and U2239 (N_2239,N_1884,N_1958);
and U2240 (N_2240,N_1558,N_1970);
or U2241 (N_2241,N_1612,N_1919);
and U2242 (N_2242,N_1552,N_1594);
xor U2243 (N_2243,N_1760,N_1801);
xnor U2244 (N_2244,N_1568,N_1606);
or U2245 (N_2245,N_1935,N_1832);
or U2246 (N_2246,N_1719,N_1511);
xor U2247 (N_2247,N_1666,N_1767);
nand U2248 (N_2248,N_1934,N_1625);
and U2249 (N_2249,N_1763,N_1896);
or U2250 (N_2250,N_1815,N_1717);
or U2251 (N_2251,N_1578,N_1640);
nand U2252 (N_2252,N_1745,N_1511);
or U2253 (N_2253,N_1735,N_1592);
and U2254 (N_2254,N_1515,N_1804);
and U2255 (N_2255,N_1534,N_1505);
nand U2256 (N_2256,N_1903,N_1507);
and U2257 (N_2257,N_1702,N_1569);
nand U2258 (N_2258,N_1550,N_1991);
nor U2259 (N_2259,N_1982,N_1618);
nor U2260 (N_2260,N_1949,N_1830);
and U2261 (N_2261,N_1975,N_1681);
nand U2262 (N_2262,N_1864,N_1839);
nand U2263 (N_2263,N_1661,N_1873);
or U2264 (N_2264,N_1676,N_1962);
or U2265 (N_2265,N_1887,N_1649);
nand U2266 (N_2266,N_1927,N_1628);
or U2267 (N_2267,N_1584,N_1945);
xor U2268 (N_2268,N_1609,N_1741);
nand U2269 (N_2269,N_1565,N_1735);
nor U2270 (N_2270,N_1709,N_1677);
nor U2271 (N_2271,N_1869,N_1661);
or U2272 (N_2272,N_1618,N_1631);
nor U2273 (N_2273,N_1835,N_1749);
xor U2274 (N_2274,N_1875,N_1793);
or U2275 (N_2275,N_1504,N_1613);
xor U2276 (N_2276,N_1609,N_1525);
xnor U2277 (N_2277,N_1829,N_1629);
or U2278 (N_2278,N_1541,N_1615);
xnor U2279 (N_2279,N_1833,N_1925);
nand U2280 (N_2280,N_1626,N_1737);
nor U2281 (N_2281,N_1526,N_1931);
and U2282 (N_2282,N_1781,N_1600);
nand U2283 (N_2283,N_1754,N_1680);
or U2284 (N_2284,N_1727,N_1511);
or U2285 (N_2285,N_1606,N_1710);
xnor U2286 (N_2286,N_1828,N_1697);
or U2287 (N_2287,N_1759,N_1841);
nand U2288 (N_2288,N_1914,N_1741);
nor U2289 (N_2289,N_1785,N_1880);
nor U2290 (N_2290,N_1507,N_1601);
nor U2291 (N_2291,N_1833,N_1589);
or U2292 (N_2292,N_1771,N_1759);
and U2293 (N_2293,N_1542,N_1611);
nor U2294 (N_2294,N_1527,N_1896);
nor U2295 (N_2295,N_1685,N_1736);
nor U2296 (N_2296,N_1551,N_1854);
xor U2297 (N_2297,N_1888,N_1857);
nand U2298 (N_2298,N_1906,N_1698);
and U2299 (N_2299,N_1600,N_1938);
or U2300 (N_2300,N_1679,N_1632);
xor U2301 (N_2301,N_1731,N_1959);
nand U2302 (N_2302,N_1774,N_1514);
nor U2303 (N_2303,N_1957,N_1510);
nor U2304 (N_2304,N_1670,N_1900);
nand U2305 (N_2305,N_1589,N_1791);
and U2306 (N_2306,N_1941,N_1696);
and U2307 (N_2307,N_1816,N_1634);
nand U2308 (N_2308,N_1608,N_1930);
and U2309 (N_2309,N_1943,N_1696);
nand U2310 (N_2310,N_1865,N_1741);
nand U2311 (N_2311,N_1613,N_1707);
and U2312 (N_2312,N_1827,N_1501);
xor U2313 (N_2313,N_1983,N_1704);
or U2314 (N_2314,N_1903,N_1659);
nand U2315 (N_2315,N_1501,N_1567);
nor U2316 (N_2316,N_1762,N_1806);
or U2317 (N_2317,N_1906,N_1583);
nand U2318 (N_2318,N_1945,N_1984);
nand U2319 (N_2319,N_1884,N_1763);
nand U2320 (N_2320,N_1837,N_1835);
xor U2321 (N_2321,N_1625,N_1830);
xnor U2322 (N_2322,N_1807,N_1515);
xnor U2323 (N_2323,N_1953,N_1742);
nand U2324 (N_2324,N_1958,N_1582);
and U2325 (N_2325,N_1692,N_1527);
or U2326 (N_2326,N_1875,N_1525);
nand U2327 (N_2327,N_1524,N_1573);
nand U2328 (N_2328,N_1709,N_1952);
nor U2329 (N_2329,N_1996,N_1670);
xor U2330 (N_2330,N_1539,N_1625);
nand U2331 (N_2331,N_1841,N_1906);
nor U2332 (N_2332,N_1803,N_1717);
or U2333 (N_2333,N_1550,N_1763);
xnor U2334 (N_2334,N_1771,N_1716);
and U2335 (N_2335,N_1635,N_1792);
nand U2336 (N_2336,N_1683,N_1849);
nor U2337 (N_2337,N_1747,N_1941);
or U2338 (N_2338,N_1767,N_1789);
and U2339 (N_2339,N_1563,N_1922);
xnor U2340 (N_2340,N_1705,N_1693);
xnor U2341 (N_2341,N_1670,N_1853);
and U2342 (N_2342,N_1645,N_1855);
nor U2343 (N_2343,N_1551,N_1743);
and U2344 (N_2344,N_1778,N_1681);
nor U2345 (N_2345,N_1518,N_1691);
nor U2346 (N_2346,N_1991,N_1657);
or U2347 (N_2347,N_1883,N_1593);
and U2348 (N_2348,N_1618,N_1652);
nor U2349 (N_2349,N_1629,N_1702);
and U2350 (N_2350,N_1911,N_1712);
and U2351 (N_2351,N_1560,N_1687);
nor U2352 (N_2352,N_1522,N_1598);
nand U2353 (N_2353,N_1598,N_1766);
nor U2354 (N_2354,N_1792,N_1957);
nand U2355 (N_2355,N_1724,N_1839);
and U2356 (N_2356,N_1545,N_1956);
nand U2357 (N_2357,N_1678,N_1608);
xor U2358 (N_2358,N_1522,N_1664);
and U2359 (N_2359,N_1651,N_1995);
nor U2360 (N_2360,N_1614,N_1624);
nor U2361 (N_2361,N_1553,N_1614);
or U2362 (N_2362,N_1847,N_1860);
xnor U2363 (N_2363,N_1975,N_1605);
nor U2364 (N_2364,N_1567,N_1955);
xor U2365 (N_2365,N_1948,N_1915);
nand U2366 (N_2366,N_1750,N_1827);
xor U2367 (N_2367,N_1532,N_1593);
nand U2368 (N_2368,N_1586,N_1656);
nand U2369 (N_2369,N_1749,N_1634);
or U2370 (N_2370,N_1777,N_1876);
nand U2371 (N_2371,N_1949,N_1706);
xor U2372 (N_2372,N_1515,N_1738);
and U2373 (N_2373,N_1884,N_1892);
xor U2374 (N_2374,N_1596,N_1603);
xnor U2375 (N_2375,N_1908,N_1681);
or U2376 (N_2376,N_1825,N_1551);
nor U2377 (N_2377,N_1772,N_1654);
or U2378 (N_2378,N_1519,N_1958);
xor U2379 (N_2379,N_1724,N_1624);
nand U2380 (N_2380,N_1588,N_1984);
and U2381 (N_2381,N_1683,N_1980);
nand U2382 (N_2382,N_1708,N_1668);
nor U2383 (N_2383,N_1885,N_1933);
nor U2384 (N_2384,N_1767,N_1630);
nor U2385 (N_2385,N_1893,N_1612);
nor U2386 (N_2386,N_1932,N_1985);
nand U2387 (N_2387,N_1750,N_1581);
nor U2388 (N_2388,N_1644,N_1622);
nor U2389 (N_2389,N_1683,N_1834);
and U2390 (N_2390,N_1510,N_1516);
nand U2391 (N_2391,N_1597,N_1952);
or U2392 (N_2392,N_1846,N_1816);
or U2393 (N_2393,N_1634,N_1840);
nor U2394 (N_2394,N_1700,N_1697);
or U2395 (N_2395,N_1725,N_1559);
and U2396 (N_2396,N_1640,N_1607);
nand U2397 (N_2397,N_1968,N_1629);
or U2398 (N_2398,N_1797,N_1990);
nand U2399 (N_2399,N_1816,N_1639);
nor U2400 (N_2400,N_1811,N_1989);
or U2401 (N_2401,N_1731,N_1663);
nand U2402 (N_2402,N_1943,N_1509);
and U2403 (N_2403,N_1976,N_1903);
and U2404 (N_2404,N_1987,N_1651);
nand U2405 (N_2405,N_1650,N_1769);
xor U2406 (N_2406,N_1726,N_1821);
nor U2407 (N_2407,N_1707,N_1791);
xnor U2408 (N_2408,N_1946,N_1533);
and U2409 (N_2409,N_1632,N_1865);
or U2410 (N_2410,N_1845,N_1662);
nor U2411 (N_2411,N_1704,N_1711);
xnor U2412 (N_2412,N_1746,N_1727);
nand U2413 (N_2413,N_1585,N_1730);
nor U2414 (N_2414,N_1906,N_1621);
nor U2415 (N_2415,N_1662,N_1537);
or U2416 (N_2416,N_1810,N_1996);
and U2417 (N_2417,N_1549,N_1718);
xnor U2418 (N_2418,N_1897,N_1958);
xor U2419 (N_2419,N_1958,N_1881);
nand U2420 (N_2420,N_1639,N_1738);
xnor U2421 (N_2421,N_1581,N_1874);
or U2422 (N_2422,N_1706,N_1608);
or U2423 (N_2423,N_1640,N_1694);
or U2424 (N_2424,N_1539,N_1530);
or U2425 (N_2425,N_1736,N_1636);
xnor U2426 (N_2426,N_1597,N_1634);
or U2427 (N_2427,N_1643,N_1980);
xnor U2428 (N_2428,N_1698,N_1696);
nand U2429 (N_2429,N_1971,N_1731);
or U2430 (N_2430,N_1644,N_1742);
and U2431 (N_2431,N_1808,N_1737);
nand U2432 (N_2432,N_1914,N_1626);
or U2433 (N_2433,N_1715,N_1927);
or U2434 (N_2434,N_1713,N_1934);
or U2435 (N_2435,N_1668,N_1534);
nand U2436 (N_2436,N_1526,N_1547);
or U2437 (N_2437,N_1747,N_1585);
or U2438 (N_2438,N_1906,N_1519);
xnor U2439 (N_2439,N_1973,N_1987);
xnor U2440 (N_2440,N_1695,N_1628);
xnor U2441 (N_2441,N_1981,N_1808);
or U2442 (N_2442,N_1561,N_1608);
nor U2443 (N_2443,N_1719,N_1988);
nand U2444 (N_2444,N_1948,N_1819);
or U2445 (N_2445,N_1949,N_1548);
or U2446 (N_2446,N_1611,N_1514);
or U2447 (N_2447,N_1876,N_1942);
xor U2448 (N_2448,N_1577,N_1806);
or U2449 (N_2449,N_1626,N_1645);
and U2450 (N_2450,N_1506,N_1600);
or U2451 (N_2451,N_1637,N_1833);
nor U2452 (N_2452,N_1801,N_1509);
nand U2453 (N_2453,N_1978,N_1710);
nor U2454 (N_2454,N_1505,N_1509);
nor U2455 (N_2455,N_1754,N_1827);
nand U2456 (N_2456,N_1678,N_1699);
nand U2457 (N_2457,N_1990,N_1971);
xnor U2458 (N_2458,N_1575,N_1540);
nor U2459 (N_2459,N_1585,N_1675);
or U2460 (N_2460,N_1613,N_1693);
or U2461 (N_2461,N_1906,N_1757);
or U2462 (N_2462,N_1903,N_1994);
xor U2463 (N_2463,N_1519,N_1661);
and U2464 (N_2464,N_1595,N_1692);
and U2465 (N_2465,N_1658,N_1879);
nor U2466 (N_2466,N_1963,N_1794);
or U2467 (N_2467,N_1621,N_1726);
xnor U2468 (N_2468,N_1710,N_1596);
and U2469 (N_2469,N_1590,N_1967);
xor U2470 (N_2470,N_1880,N_1749);
xor U2471 (N_2471,N_1639,N_1891);
nand U2472 (N_2472,N_1581,N_1556);
and U2473 (N_2473,N_1534,N_1504);
nor U2474 (N_2474,N_1535,N_1952);
nor U2475 (N_2475,N_1506,N_1668);
or U2476 (N_2476,N_1693,N_1907);
nor U2477 (N_2477,N_1729,N_1792);
or U2478 (N_2478,N_1634,N_1716);
and U2479 (N_2479,N_1548,N_1514);
and U2480 (N_2480,N_1693,N_1804);
xor U2481 (N_2481,N_1759,N_1655);
nor U2482 (N_2482,N_1671,N_1640);
or U2483 (N_2483,N_1885,N_1888);
and U2484 (N_2484,N_1888,N_1869);
nor U2485 (N_2485,N_1590,N_1616);
or U2486 (N_2486,N_1525,N_1549);
xnor U2487 (N_2487,N_1929,N_1926);
xnor U2488 (N_2488,N_1551,N_1649);
xor U2489 (N_2489,N_1787,N_1648);
or U2490 (N_2490,N_1838,N_1981);
and U2491 (N_2491,N_1658,N_1631);
nor U2492 (N_2492,N_1658,N_1818);
or U2493 (N_2493,N_1896,N_1816);
and U2494 (N_2494,N_1848,N_1609);
nor U2495 (N_2495,N_1795,N_1728);
or U2496 (N_2496,N_1611,N_1668);
xor U2497 (N_2497,N_1882,N_1694);
or U2498 (N_2498,N_1689,N_1522);
nand U2499 (N_2499,N_1997,N_1719);
or U2500 (N_2500,N_2151,N_2415);
xor U2501 (N_2501,N_2334,N_2159);
nor U2502 (N_2502,N_2399,N_2410);
nand U2503 (N_2503,N_2173,N_2047);
and U2504 (N_2504,N_2488,N_2146);
nor U2505 (N_2505,N_2437,N_2093);
xnor U2506 (N_2506,N_2029,N_2434);
or U2507 (N_2507,N_2493,N_2270);
nand U2508 (N_2508,N_2492,N_2196);
xor U2509 (N_2509,N_2221,N_2172);
nor U2510 (N_2510,N_2001,N_2244);
nand U2511 (N_2511,N_2157,N_2327);
nand U2512 (N_2512,N_2165,N_2286);
and U2513 (N_2513,N_2379,N_2238);
and U2514 (N_2514,N_2461,N_2080);
nand U2515 (N_2515,N_2186,N_2102);
nand U2516 (N_2516,N_2245,N_2273);
nand U2517 (N_2517,N_2212,N_2442);
xor U2518 (N_2518,N_2272,N_2048);
nor U2519 (N_2519,N_2130,N_2494);
or U2520 (N_2520,N_2193,N_2224);
and U2521 (N_2521,N_2315,N_2027);
nand U2522 (N_2522,N_2333,N_2064);
and U2523 (N_2523,N_2141,N_2483);
and U2524 (N_2524,N_2388,N_2112);
or U2525 (N_2525,N_2233,N_2061);
and U2526 (N_2526,N_2430,N_2370);
nand U2527 (N_2527,N_2435,N_2291);
xor U2528 (N_2528,N_2252,N_2121);
and U2529 (N_2529,N_2046,N_2055);
nand U2530 (N_2530,N_2153,N_2177);
xnor U2531 (N_2531,N_2418,N_2246);
nor U2532 (N_2532,N_2076,N_2427);
nor U2533 (N_2533,N_2038,N_2409);
xnor U2534 (N_2534,N_2373,N_2429);
and U2535 (N_2535,N_2470,N_2145);
or U2536 (N_2536,N_2087,N_2105);
nand U2537 (N_2537,N_2411,N_2417);
and U2538 (N_2538,N_2036,N_2302);
xor U2539 (N_2539,N_2469,N_2353);
xor U2540 (N_2540,N_2445,N_2421);
or U2541 (N_2541,N_2416,N_2419);
nand U2542 (N_2542,N_2197,N_2241);
or U2543 (N_2543,N_2015,N_2452);
and U2544 (N_2544,N_2480,N_2387);
xor U2545 (N_2545,N_2187,N_2219);
nand U2546 (N_2546,N_2365,N_2009);
nor U2547 (N_2547,N_2086,N_2360);
nand U2548 (N_2548,N_2479,N_2440);
xnor U2549 (N_2549,N_2220,N_2462);
and U2550 (N_2550,N_2344,N_2215);
nand U2551 (N_2551,N_2201,N_2489);
and U2552 (N_2552,N_2084,N_2362);
nor U2553 (N_2553,N_2366,N_2401);
nand U2554 (N_2554,N_2089,N_2279);
nand U2555 (N_2555,N_2391,N_2303);
and U2556 (N_2556,N_2178,N_2184);
or U2557 (N_2557,N_2211,N_2176);
or U2558 (N_2558,N_2345,N_2495);
xor U2559 (N_2559,N_2283,N_2405);
or U2560 (N_2560,N_2295,N_2318);
nor U2561 (N_2561,N_2192,N_2464);
xor U2562 (N_2562,N_2074,N_2234);
xor U2563 (N_2563,N_2132,N_2348);
or U2564 (N_2564,N_2065,N_2250);
xor U2565 (N_2565,N_2395,N_2383);
xnor U2566 (N_2566,N_2031,N_2347);
nand U2567 (N_2567,N_2406,N_2376);
nand U2568 (N_2568,N_2191,N_2280);
nor U2569 (N_2569,N_2218,N_2206);
xor U2570 (N_2570,N_2354,N_2448);
and U2571 (N_2571,N_2491,N_2322);
nand U2572 (N_2572,N_2033,N_2476);
nor U2573 (N_2573,N_2320,N_2021);
xnor U2574 (N_2574,N_2499,N_2271);
nor U2575 (N_2575,N_2482,N_2095);
xnor U2576 (N_2576,N_2335,N_2122);
nand U2577 (N_2577,N_2123,N_2228);
or U2578 (N_2578,N_2020,N_2116);
xor U2579 (N_2579,N_2040,N_2386);
or U2580 (N_2580,N_2203,N_2382);
nand U2581 (N_2581,N_2068,N_2100);
xnor U2582 (N_2582,N_2057,N_2003);
or U2583 (N_2583,N_2077,N_2359);
nand U2584 (N_2584,N_2161,N_2456);
xor U2585 (N_2585,N_2441,N_2477);
xnor U2586 (N_2586,N_2230,N_2090);
and U2587 (N_2587,N_2231,N_2164);
nor U2588 (N_2588,N_2439,N_2496);
xor U2589 (N_2589,N_2413,N_2371);
xor U2590 (N_2590,N_2056,N_2285);
nor U2591 (N_2591,N_2200,N_2357);
xnor U2592 (N_2592,N_2258,N_2147);
nand U2593 (N_2593,N_2372,N_2222);
and U2594 (N_2594,N_2180,N_2138);
xnor U2595 (N_2595,N_2490,N_2396);
nor U2596 (N_2596,N_2288,N_2171);
nand U2597 (N_2597,N_2075,N_2097);
xor U2598 (N_2598,N_2447,N_2332);
or U2599 (N_2599,N_2152,N_2329);
or U2600 (N_2600,N_2170,N_2078);
nand U2601 (N_2601,N_2127,N_2367);
nor U2602 (N_2602,N_2264,N_2085);
nand U2603 (N_2603,N_2485,N_2301);
or U2604 (N_2604,N_2254,N_2341);
nor U2605 (N_2605,N_2240,N_2390);
xnor U2606 (N_2606,N_2298,N_2094);
nand U2607 (N_2607,N_2443,N_2158);
xnor U2608 (N_2608,N_2316,N_2169);
and U2609 (N_2609,N_2135,N_2330);
nor U2610 (N_2610,N_2028,N_2162);
nand U2611 (N_2611,N_2239,N_2008);
nand U2612 (N_2612,N_2126,N_2392);
and U2613 (N_2613,N_2174,N_2109);
nor U2614 (N_2614,N_2314,N_2167);
xnor U2615 (N_2615,N_2004,N_2181);
nand U2616 (N_2616,N_2251,N_2012);
and U2617 (N_2617,N_2136,N_2481);
xor U2618 (N_2618,N_2284,N_2025);
xor U2619 (N_2619,N_2111,N_2398);
xor U2620 (N_2620,N_2281,N_2039);
nor U2621 (N_2621,N_2384,N_2227);
or U2622 (N_2622,N_2317,N_2467);
and U2623 (N_2623,N_2118,N_2260);
and U2624 (N_2624,N_2050,N_2324);
and U2625 (N_2625,N_2142,N_2185);
nor U2626 (N_2626,N_2129,N_2081);
or U2627 (N_2627,N_2451,N_2319);
or U2628 (N_2628,N_2338,N_2044);
and U2629 (N_2629,N_2007,N_2101);
xor U2630 (N_2630,N_2179,N_2275);
or U2631 (N_2631,N_2304,N_2342);
and U2632 (N_2632,N_2454,N_2140);
or U2633 (N_2633,N_2358,N_2300);
nand U2634 (N_2634,N_2474,N_2407);
or U2635 (N_2635,N_2099,N_2088);
xor U2636 (N_2636,N_2000,N_2313);
or U2637 (N_2637,N_2189,N_2160);
and U2638 (N_2638,N_2067,N_2062);
and U2639 (N_2639,N_2190,N_2060);
and U2640 (N_2640,N_2011,N_2265);
nor U2641 (N_2641,N_2223,N_2328);
nand U2642 (N_2642,N_2144,N_2389);
or U2643 (N_2643,N_2325,N_2226);
and U2644 (N_2644,N_2378,N_2471);
and U2645 (N_2645,N_2455,N_2049);
or U2646 (N_2646,N_2175,N_2486);
nand U2647 (N_2647,N_2069,N_2030);
xnor U2648 (N_2648,N_2487,N_2019);
nand U2649 (N_2649,N_2072,N_2278);
nor U2650 (N_2650,N_2091,N_2349);
or U2651 (N_2651,N_2213,N_2119);
and U2652 (N_2652,N_2182,N_2249);
or U2653 (N_2653,N_2287,N_2433);
or U2654 (N_2654,N_2356,N_2051);
xnor U2655 (N_2655,N_2183,N_2351);
nor U2656 (N_2656,N_2497,N_2262);
and U2657 (N_2657,N_2117,N_2210);
nor U2658 (N_2658,N_2242,N_2267);
and U2659 (N_2659,N_2473,N_2243);
xor U2660 (N_2660,N_2308,N_2374);
nand U2661 (N_2661,N_2498,N_2259);
or U2662 (N_2662,N_2014,N_2071);
or U2663 (N_2663,N_2198,N_2294);
nor U2664 (N_2664,N_2305,N_2079);
and U2665 (N_2665,N_2216,N_2394);
nor U2666 (N_2666,N_2150,N_2400);
and U2667 (N_2667,N_2034,N_2043);
xnor U2668 (N_2668,N_2045,N_2110);
xnor U2669 (N_2669,N_2310,N_2208);
and U2670 (N_2670,N_2247,N_2053);
nor U2671 (N_2671,N_2339,N_2229);
nand U2672 (N_2672,N_2195,N_2148);
xor U2673 (N_2673,N_2042,N_2380);
or U2674 (N_2674,N_2214,N_2326);
xor U2675 (N_2675,N_2484,N_2266);
and U2676 (N_2676,N_2052,N_2309);
nand U2677 (N_2677,N_2468,N_2299);
or U2678 (N_2678,N_2312,N_2472);
and U2679 (N_2679,N_2236,N_2006);
nand U2680 (N_2680,N_2307,N_2232);
nor U2681 (N_2681,N_2114,N_2368);
nor U2682 (N_2682,N_2292,N_2449);
or U2683 (N_2683,N_2016,N_2125);
or U2684 (N_2684,N_2022,N_2438);
xor U2685 (N_2685,N_2024,N_2154);
nor U2686 (N_2686,N_2155,N_2414);
xnor U2687 (N_2687,N_2202,N_2010);
nor U2688 (N_2688,N_2453,N_2096);
or U2689 (N_2689,N_2336,N_2018);
or U2690 (N_2690,N_2041,N_2289);
and U2691 (N_2691,N_2054,N_2460);
nand U2692 (N_2692,N_2428,N_2321);
and U2693 (N_2693,N_2137,N_2194);
xnor U2694 (N_2694,N_2005,N_2013);
or U2695 (N_2695,N_2276,N_2035);
nand U2696 (N_2696,N_2032,N_2343);
or U2697 (N_2697,N_2363,N_2478);
and U2698 (N_2698,N_2459,N_2066);
nand U2699 (N_2699,N_2207,N_2364);
xor U2700 (N_2700,N_2163,N_2058);
xor U2701 (N_2701,N_2282,N_2073);
and U2702 (N_2702,N_2149,N_2465);
and U2703 (N_2703,N_2475,N_2457);
and U2704 (N_2704,N_2156,N_2422);
xor U2705 (N_2705,N_2323,N_2420);
nor U2706 (N_2706,N_2337,N_2402);
nor U2707 (N_2707,N_2466,N_2277);
or U2708 (N_2708,N_2458,N_2037);
nand U2709 (N_2709,N_2404,N_2352);
and U2710 (N_2710,N_2306,N_2355);
xnor U2711 (N_2711,N_2103,N_2120);
nor U2712 (N_2712,N_2293,N_2235);
or U2713 (N_2713,N_2346,N_2115);
and U2714 (N_2714,N_2063,N_2431);
xor U2715 (N_2715,N_2253,N_2403);
nand U2716 (N_2716,N_2269,N_2268);
nand U2717 (N_2717,N_2381,N_2026);
or U2718 (N_2718,N_2426,N_2436);
nand U2719 (N_2719,N_2199,N_2393);
nor U2720 (N_2720,N_2423,N_2257);
nor U2721 (N_2721,N_2092,N_2340);
or U2722 (N_2722,N_2205,N_2385);
xor U2723 (N_2723,N_2424,N_2023);
or U2724 (N_2724,N_2425,N_2059);
xor U2725 (N_2725,N_2261,N_2331);
and U2726 (N_2726,N_2104,N_2108);
and U2727 (N_2727,N_2113,N_2133);
xor U2728 (N_2728,N_2412,N_2397);
or U2729 (N_2729,N_2255,N_2017);
xnor U2730 (N_2730,N_2375,N_2143);
nor U2731 (N_2731,N_2432,N_2188);
or U2732 (N_2732,N_2450,N_2209);
nand U2733 (N_2733,N_2311,N_2408);
nor U2734 (N_2734,N_2248,N_2131);
nand U2735 (N_2735,N_2070,N_2290);
xnor U2736 (N_2736,N_2082,N_2274);
nor U2737 (N_2737,N_2444,N_2166);
xor U2738 (N_2738,N_2134,N_2217);
and U2739 (N_2739,N_2446,N_2083);
nand U2740 (N_2740,N_2107,N_2463);
xor U2741 (N_2741,N_2369,N_2350);
nor U2742 (N_2742,N_2124,N_2168);
nor U2743 (N_2743,N_2204,N_2297);
nand U2744 (N_2744,N_2263,N_2098);
and U2745 (N_2745,N_2128,N_2361);
and U2746 (N_2746,N_2256,N_2377);
and U2747 (N_2747,N_2237,N_2139);
nor U2748 (N_2748,N_2002,N_2296);
nor U2749 (N_2749,N_2225,N_2106);
nand U2750 (N_2750,N_2276,N_2214);
or U2751 (N_2751,N_2378,N_2012);
and U2752 (N_2752,N_2149,N_2255);
xor U2753 (N_2753,N_2347,N_2147);
nand U2754 (N_2754,N_2223,N_2048);
xor U2755 (N_2755,N_2079,N_2009);
xor U2756 (N_2756,N_2068,N_2067);
nand U2757 (N_2757,N_2012,N_2350);
nor U2758 (N_2758,N_2209,N_2443);
nand U2759 (N_2759,N_2047,N_2312);
or U2760 (N_2760,N_2195,N_2480);
nor U2761 (N_2761,N_2003,N_2406);
or U2762 (N_2762,N_2169,N_2000);
or U2763 (N_2763,N_2003,N_2121);
nor U2764 (N_2764,N_2038,N_2347);
xnor U2765 (N_2765,N_2045,N_2123);
nand U2766 (N_2766,N_2100,N_2458);
xor U2767 (N_2767,N_2109,N_2172);
and U2768 (N_2768,N_2494,N_2197);
nand U2769 (N_2769,N_2391,N_2306);
nand U2770 (N_2770,N_2286,N_2216);
nor U2771 (N_2771,N_2367,N_2194);
nand U2772 (N_2772,N_2462,N_2295);
xor U2773 (N_2773,N_2238,N_2059);
or U2774 (N_2774,N_2399,N_2495);
and U2775 (N_2775,N_2293,N_2157);
and U2776 (N_2776,N_2353,N_2101);
or U2777 (N_2777,N_2405,N_2461);
nand U2778 (N_2778,N_2064,N_2262);
or U2779 (N_2779,N_2355,N_2316);
nand U2780 (N_2780,N_2305,N_2421);
nor U2781 (N_2781,N_2385,N_2366);
xor U2782 (N_2782,N_2418,N_2471);
and U2783 (N_2783,N_2220,N_2001);
nor U2784 (N_2784,N_2093,N_2233);
and U2785 (N_2785,N_2371,N_2233);
nor U2786 (N_2786,N_2308,N_2072);
nand U2787 (N_2787,N_2265,N_2186);
nand U2788 (N_2788,N_2235,N_2435);
or U2789 (N_2789,N_2285,N_2497);
or U2790 (N_2790,N_2364,N_2169);
xnor U2791 (N_2791,N_2442,N_2481);
or U2792 (N_2792,N_2451,N_2195);
xor U2793 (N_2793,N_2198,N_2436);
nand U2794 (N_2794,N_2458,N_2173);
nor U2795 (N_2795,N_2307,N_2323);
and U2796 (N_2796,N_2349,N_2280);
and U2797 (N_2797,N_2177,N_2038);
nand U2798 (N_2798,N_2356,N_2375);
nand U2799 (N_2799,N_2396,N_2436);
xor U2800 (N_2800,N_2420,N_2135);
or U2801 (N_2801,N_2039,N_2151);
or U2802 (N_2802,N_2075,N_2492);
nand U2803 (N_2803,N_2395,N_2296);
nor U2804 (N_2804,N_2065,N_2331);
xnor U2805 (N_2805,N_2190,N_2428);
and U2806 (N_2806,N_2465,N_2243);
or U2807 (N_2807,N_2492,N_2366);
and U2808 (N_2808,N_2484,N_2094);
nor U2809 (N_2809,N_2238,N_2482);
xnor U2810 (N_2810,N_2165,N_2323);
and U2811 (N_2811,N_2169,N_2068);
nor U2812 (N_2812,N_2397,N_2443);
and U2813 (N_2813,N_2338,N_2231);
nand U2814 (N_2814,N_2161,N_2337);
nand U2815 (N_2815,N_2345,N_2109);
or U2816 (N_2816,N_2352,N_2466);
nand U2817 (N_2817,N_2303,N_2360);
and U2818 (N_2818,N_2017,N_2002);
or U2819 (N_2819,N_2305,N_2460);
nand U2820 (N_2820,N_2147,N_2096);
xnor U2821 (N_2821,N_2145,N_2111);
xnor U2822 (N_2822,N_2410,N_2456);
and U2823 (N_2823,N_2342,N_2207);
or U2824 (N_2824,N_2363,N_2394);
nor U2825 (N_2825,N_2307,N_2479);
and U2826 (N_2826,N_2178,N_2036);
nand U2827 (N_2827,N_2289,N_2356);
xnor U2828 (N_2828,N_2027,N_2280);
or U2829 (N_2829,N_2135,N_2092);
nand U2830 (N_2830,N_2229,N_2499);
xnor U2831 (N_2831,N_2365,N_2439);
nand U2832 (N_2832,N_2191,N_2039);
and U2833 (N_2833,N_2253,N_2443);
nor U2834 (N_2834,N_2366,N_2046);
nor U2835 (N_2835,N_2427,N_2205);
or U2836 (N_2836,N_2281,N_2229);
and U2837 (N_2837,N_2498,N_2324);
xnor U2838 (N_2838,N_2411,N_2374);
xnor U2839 (N_2839,N_2187,N_2358);
and U2840 (N_2840,N_2137,N_2114);
nor U2841 (N_2841,N_2369,N_2332);
xnor U2842 (N_2842,N_2286,N_2462);
and U2843 (N_2843,N_2137,N_2321);
xor U2844 (N_2844,N_2434,N_2103);
or U2845 (N_2845,N_2212,N_2358);
and U2846 (N_2846,N_2001,N_2391);
and U2847 (N_2847,N_2418,N_2247);
nand U2848 (N_2848,N_2013,N_2123);
and U2849 (N_2849,N_2181,N_2416);
or U2850 (N_2850,N_2170,N_2229);
and U2851 (N_2851,N_2414,N_2165);
and U2852 (N_2852,N_2456,N_2185);
nor U2853 (N_2853,N_2240,N_2020);
nand U2854 (N_2854,N_2442,N_2072);
or U2855 (N_2855,N_2422,N_2163);
and U2856 (N_2856,N_2411,N_2396);
xnor U2857 (N_2857,N_2039,N_2292);
and U2858 (N_2858,N_2082,N_2120);
and U2859 (N_2859,N_2115,N_2483);
nor U2860 (N_2860,N_2211,N_2461);
xnor U2861 (N_2861,N_2305,N_2273);
and U2862 (N_2862,N_2276,N_2406);
xor U2863 (N_2863,N_2447,N_2193);
xor U2864 (N_2864,N_2297,N_2181);
nor U2865 (N_2865,N_2268,N_2096);
nor U2866 (N_2866,N_2013,N_2194);
nand U2867 (N_2867,N_2120,N_2365);
nand U2868 (N_2868,N_2133,N_2063);
and U2869 (N_2869,N_2128,N_2066);
or U2870 (N_2870,N_2358,N_2469);
xor U2871 (N_2871,N_2254,N_2479);
or U2872 (N_2872,N_2341,N_2064);
or U2873 (N_2873,N_2113,N_2312);
and U2874 (N_2874,N_2301,N_2169);
and U2875 (N_2875,N_2497,N_2348);
nand U2876 (N_2876,N_2333,N_2189);
xor U2877 (N_2877,N_2285,N_2157);
nand U2878 (N_2878,N_2003,N_2179);
xor U2879 (N_2879,N_2003,N_2014);
nand U2880 (N_2880,N_2074,N_2076);
and U2881 (N_2881,N_2276,N_2241);
nor U2882 (N_2882,N_2425,N_2007);
and U2883 (N_2883,N_2123,N_2442);
and U2884 (N_2884,N_2118,N_2045);
or U2885 (N_2885,N_2431,N_2252);
nor U2886 (N_2886,N_2181,N_2249);
or U2887 (N_2887,N_2342,N_2458);
nor U2888 (N_2888,N_2023,N_2158);
and U2889 (N_2889,N_2499,N_2354);
or U2890 (N_2890,N_2161,N_2311);
or U2891 (N_2891,N_2038,N_2000);
nor U2892 (N_2892,N_2230,N_2236);
xnor U2893 (N_2893,N_2228,N_2186);
nor U2894 (N_2894,N_2001,N_2165);
nor U2895 (N_2895,N_2117,N_2165);
xnor U2896 (N_2896,N_2080,N_2277);
xor U2897 (N_2897,N_2481,N_2246);
nand U2898 (N_2898,N_2140,N_2008);
nor U2899 (N_2899,N_2134,N_2093);
and U2900 (N_2900,N_2051,N_2013);
nand U2901 (N_2901,N_2341,N_2054);
xnor U2902 (N_2902,N_2288,N_2424);
nand U2903 (N_2903,N_2063,N_2128);
and U2904 (N_2904,N_2213,N_2091);
or U2905 (N_2905,N_2475,N_2263);
nand U2906 (N_2906,N_2094,N_2266);
and U2907 (N_2907,N_2294,N_2173);
and U2908 (N_2908,N_2065,N_2388);
xnor U2909 (N_2909,N_2309,N_2213);
nand U2910 (N_2910,N_2449,N_2458);
nand U2911 (N_2911,N_2385,N_2195);
nand U2912 (N_2912,N_2328,N_2137);
nor U2913 (N_2913,N_2314,N_2408);
nand U2914 (N_2914,N_2021,N_2030);
nor U2915 (N_2915,N_2253,N_2398);
nor U2916 (N_2916,N_2390,N_2025);
nand U2917 (N_2917,N_2080,N_2315);
nand U2918 (N_2918,N_2324,N_2478);
or U2919 (N_2919,N_2155,N_2487);
or U2920 (N_2920,N_2250,N_2318);
and U2921 (N_2921,N_2274,N_2010);
xnor U2922 (N_2922,N_2431,N_2185);
nor U2923 (N_2923,N_2075,N_2113);
nor U2924 (N_2924,N_2316,N_2429);
nand U2925 (N_2925,N_2164,N_2257);
nand U2926 (N_2926,N_2279,N_2400);
xnor U2927 (N_2927,N_2364,N_2379);
xnor U2928 (N_2928,N_2097,N_2093);
and U2929 (N_2929,N_2412,N_2015);
or U2930 (N_2930,N_2032,N_2096);
nor U2931 (N_2931,N_2323,N_2099);
xnor U2932 (N_2932,N_2052,N_2022);
or U2933 (N_2933,N_2063,N_2232);
xor U2934 (N_2934,N_2316,N_2300);
and U2935 (N_2935,N_2052,N_2256);
or U2936 (N_2936,N_2052,N_2000);
xnor U2937 (N_2937,N_2357,N_2361);
or U2938 (N_2938,N_2240,N_2343);
nor U2939 (N_2939,N_2327,N_2341);
and U2940 (N_2940,N_2490,N_2157);
or U2941 (N_2941,N_2155,N_2126);
or U2942 (N_2942,N_2382,N_2046);
xnor U2943 (N_2943,N_2323,N_2210);
or U2944 (N_2944,N_2354,N_2335);
nor U2945 (N_2945,N_2125,N_2450);
xor U2946 (N_2946,N_2429,N_2351);
nand U2947 (N_2947,N_2017,N_2408);
nand U2948 (N_2948,N_2416,N_2467);
and U2949 (N_2949,N_2349,N_2036);
nor U2950 (N_2950,N_2090,N_2159);
or U2951 (N_2951,N_2193,N_2115);
xnor U2952 (N_2952,N_2308,N_2022);
and U2953 (N_2953,N_2147,N_2405);
xnor U2954 (N_2954,N_2301,N_2167);
nor U2955 (N_2955,N_2025,N_2079);
nor U2956 (N_2956,N_2460,N_2446);
nand U2957 (N_2957,N_2078,N_2251);
xnor U2958 (N_2958,N_2167,N_2416);
xor U2959 (N_2959,N_2144,N_2385);
xnor U2960 (N_2960,N_2205,N_2369);
xor U2961 (N_2961,N_2432,N_2083);
nor U2962 (N_2962,N_2041,N_2171);
and U2963 (N_2963,N_2003,N_2112);
nor U2964 (N_2964,N_2129,N_2490);
nor U2965 (N_2965,N_2499,N_2086);
nor U2966 (N_2966,N_2063,N_2417);
and U2967 (N_2967,N_2329,N_2189);
nor U2968 (N_2968,N_2053,N_2166);
or U2969 (N_2969,N_2481,N_2334);
nand U2970 (N_2970,N_2159,N_2361);
nand U2971 (N_2971,N_2346,N_2458);
or U2972 (N_2972,N_2416,N_2484);
and U2973 (N_2973,N_2328,N_2478);
xor U2974 (N_2974,N_2232,N_2162);
xor U2975 (N_2975,N_2289,N_2432);
nor U2976 (N_2976,N_2265,N_2120);
nor U2977 (N_2977,N_2284,N_2170);
and U2978 (N_2978,N_2352,N_2302);
or U2979 (N_2979,N_2283,N_2073);
and U2980 (N_2980,N_2383,N_2441);
xnor U2981 (N_2981,N_2403,N_2436);
nand U2982 (N_2982,N_2183,N_2398);
nor U2983 (N_2983,N_2333,N_2389);
or U2984 (N_2984,N_2145,N_2332);
nor U2985 (N_2985,N_2471,N_2486);
or U2986 (N_2986,N_2302,N_2265);
or U2987 (N_2987,N_2461,N_2468);
nand U2988 (N_2988,N_2245,N_2264);
and U2989 (N_2989,N_2289,N_2209);
nand U2990 (N_2990,N_2496,N_2148);
nor U2991 (N_2991,N_2031,N_2275);
or U2992 (N_2992,N_2286,N_2032);
nor U2993 (N_2993,N_2010,N_2432);
nand U2994 (N_2994,N_2131,N_2430);
or U2995 (N_2995,N_2187,N_2357);
xor U2996 (N_2996,N_2075,N_2017);
nor U2997 (N_2997,N_2302,N_2495);
nand U2998 (N_2998,N_2276,N_2360);
xnor U2999 (N_2999,N_2351,N_2069);
and U3000 (N_3000,N_2504,N_2603);
nand U3001 (N_3001,N_2904,N_2980);
xor U3002 (N_3002,N_2695,N_2615);
or U3003 (N_3003,N_2543,N_2688);
nor U3004 (N_3004,N_2701,N_2941);
and U3005 (N_3005,N_2671,N_2654);
and U3006 (N_3006,N_2714,N_2763);
or U3007 (N_3007,N_2638,N_2925);
or U3008 (N_3008,N_2785,N_2847);
or U3009 (N_3009,N_2508,N_2815);
or U3010 (N_3010,N_2720,N_2711);
xnor U3011 (N_3011,N_2857,N_2844);
and U3012 (N_3012,N_2580,N_2996);
nor U3013 (N_3013,N_2790,N_2716);
xnor U3014 (N_3014,N_2723,N_2624);
nor U3015 (N_3015,N_2923,N_2893);
xnor U3016 (N_3016,N_2617,N_2949);
nor U3017 (N_3017,N_2816,N_2717);
xor U3018 (N_3018,N_2601,N_2787);
xor U3019 (N_3019,N_2590,N_2878);
xnor U3020 (N_3020,N_2674,N_2541);
and U3021 (N_3021,N_2849,N_2999);
xor U3022 (N_3022,N_2957,N_2839);
nand U3023 (N_3023,N_2606,N_2780);
and U3024 (N_3024,N_2843,N_2776);
nand U3025 (N_3025,N_2599,N_2709);
or U3026 (N_3026,N_2691,N_2639);
nand U3027 (N_3027,N_2917,N_2680);
xnor U3028 (N_3028,N_2517,N_2683);
and U3029 (N_3029,N_2833,N_2838);
or U3030 (N_3030,N_2666,N_2636);
nand U3031 (N_3031,N_2708,N_2991);
or U3032 (N_3032,N_2511,N_2745);
nand U3033 (N_3033,N_2876,N_2575);
nor U3034 (N_3034,N_2736,N_2643);
nor U3035 (N_3035,N_2842,N_2576);
nor U3036 (N_3036,N_2867,N_2952);
and U3037 (N_3037,N_2529,N_2903);
nand U3038 (N_3038,N_2871,N_2907);
and U3039 (N_3039,N_2530,N_2573);
or U3040 (N_3040,N_2733,N_2966);
nand U3041 (N_3041,N_2538,N_2805);
or U3042 (N_3042,N_2918,N_2731);
and U3043 (N_3043,N_2678,N_2783);
xnor U3044 (N_3044,N_2846,N_2692);
and U3045 (N_3045,N_2932,N_2775);
or U3046 (N_3046,N_2747,N_2571);
xnor U3047 (N_3047,N_2858,N_2649);
xnor U3048 (N_3048,N_2964,N_2682);
nand U3049 (N_3049,N_2946,N_2569);
and U3050 (N_3050,N_2620,N_2902);
nand U3051 (N_3051,N_2528,N_2597);
and U3052 (N_3052,N_2670,N_2760);
nand U3053 (N_3053,N_2725,N_2684);
or U3054 (N_3054,N_2799,N_2697);
xnor U3055 (N_3055,N_2753,N_2728);
nor U3056 (N_3056,N_2631,N_2548);
nand U3057 (N_3057,N_2718,N_2859);
nor U3058 (N_3058,N_2770,N_2761);
and U3059 (N_3059,N_2500,N_2598);
nor U3060 (N_3060,N_2628,N_2744);
or U3061 (N_3061,N_2627,N_2924);
nand U3062 (N_3062,N_2641,N_2979);
xor U3063 (N_3063,N_2762,N_2502);
or U3064 (N_3064,N_2935,N_2927);
and U3065 (N_3065,N_2607,N_2807);
nand U3066 (N_3066,N_2983,N_2901);
or U3067 (N_3067,N_2749,N_2881);
nor U3068 (N_3068,N_2735,N_2604);
and U3069 (N_3069,N_2765,N_2911);
nand U3070 (N_3070,N_2591,N_2592);
nand U3071 (N_3071,N_2612,N_2668);
and U3072 (N_3072,N_2687,N_2919);
or U3073 (N_3073,N_2795,N_2945);
and U3074 (N_3074,N_2686,N_2921);
xnor U3075 (N_3075,N_2653,N_2806);
or U3076 (N_3076,N_2885,N_2933);
or U3077 (N_3077,N_2809,N_2880);
or U3078 (N_3078,N_2756,N_2811);
or U3079 (N_3079,N_2755,N_2507);
and U3080 (N_3080,N_2644,N_2694);
or U3081 (N_3081,N_2832,N_2836);
or U3082 (N_3082,N_2552,N_2655);
or U3083 (N_3083,N_2936,N_2888);
nor U3084 (N_3084,N_2581,N_2732);
or U3085 (N_3085,N_2845,N_2953);
or U3086 (N_3086,N_2984,N_2647);
and U3087 (N_3087,N_2712,N_2937);
or U3088 (N_3088,N_2704,N_2928);
nor U3089 (N_3089,N_2681,N_2820);
xnor U3090 (N_3090,N_2740,N_2989);
or U3091 (N_3091,N_2633,N_2873);
xnor U3092 (N_3092,N_2588,N_2967);
and U3093 (N_3093,N_2690,N_2501);
nor U3094 (N_3094,N_2729,N_2738);
and U3095 (N_3095,N_2512,N_2719);
and U3096 (N_3096,N_2974,N_2951);
and U3097 (N_3097,N_2840,N_2677);
nor U3098 (N_3098,N_2658,N_2519);
and U3099 (N_3099,N_2825,N_2884);
nor U3100 (N_3100,N_2862,N_2819);
nand U3101 (N_3101,N_2531,N_2894);
xnor U3102 (N_3102,N_2960,N_2710);
or U3103 (N_3103,N_2778,N_2613);
and U3104 (N_3104,N_2782,N_2988);
and U3105 (N_3105,N_2594,N_2887);
xor U3106 (N_3106,N_2535,N_2546);
and U3107 (N_3107,N_2922,N_2864);
or U3108 (N_3108,N_2514,N_2585);
nor U3109 (N_3109,N_2856,N_2982);
nand U3110 (N_3110,N_2852,N_2558);
or U3111 (N_3111,N_2900,N_2913);
nor U3112 (N_3112,N_2771,N_2899);
nor U3113 (N_3113,N_2727,N_2797);
nand U3114 (N_3114,N_2827,N_2956);
nand U3115 (N_3115,N_2520,N_2975);
or U3116 (N_3116,N_2540,N_2772);
nand U3117 (N_3117,N_2889,N_2834);
xor U3118 (N_3118,N_2616,N_2985);
xor U3119 (N_3119,N_2970,N_2545);
and U3120 (N_3120,N_2905,N_2800);
and U3121 (N_3121,N_2623,N_2987);
xor U3122 (N_3122,N_2971,N_2931);
nand U3123 (N_3123,N_2605,N_2525);
xnor U3124 (N_3124,N_2958,N_2882);
nand U3125 (N_3125,N_2976,N_2555);
or U3126 (N_3126,N_2930,N_2835);
xnor U3127 (N_3127,N_2568,N_2837);
xor U3128 (N_3128,N_2669,N_2865);
xor U3129 (N_3129,N_2963,N_2685);
and U3130 (N_3130,N_2635,N_2934);
xor U3131 (N_3131,N_2897,N_2640);
xor U3132 (N_3132,N_2828,N_2866);
xor U3133 (N_3133,N_2944,N_2777);
nor U3134 (N_3134,N_2767,N_2860);
nand U3135 (N_3135,N_2879,N_2503);
xnor U3136 (N_3136,N_2977,N_2657);
nand U3137 (N_3137,N_2564,N_2877);
nand U3138 (N_3138,N_2853,N_2516);
or U3139 (N_3139,N_2579,N_2943);
or U3140 (N_3140,N_2673,N_2527);
xnor U3141 (N_3141,N_2774,N_2572);
or U3142 (N_3142,N_2892,N_2562);
and U3143 (N_3143,N_2886,N_2618);
xnor U3144 (N_3144,N_2915,N_2992);
or U3145 (N_3145,N_2786,N_2537);
or U3146 (N_3146,N_2830,N_2608);
and U3147 (N_3147,N_2506,N_2600);
nand U3148 (N_3148,N_2713,N_2582);
or U3149 (N_3149,N_2533,N_2758);
nor U3150 (N_3150,N_2978,N_2542);
nor U3151 (N_3151,N_2817,N_2706);
or U3152 (N_3152,N_2757,N_2962);
or U3153 (N_3153,N_2869,N_2891);
and U3154 (N_3154,N_2823,N_2651);
nor U3155 (N_3155,N_2619,N_2947);
xnor U3156 (N_3156,N_2750,N_2629);
nor U3157 (N_3157,N_2645,N_2549);
and U3158 (N_3158,N_2648,N_2773);
and U3159 (N_3159,N_2812,N_2621);
nor U3160 (N_3160,N_2589,N_2965);
or U3161 (N_3161,N_2521,N_2997);
and U3162 (N_3162,N_2539,N_2524);
nand U3163 (N_3163,N_2950,N_2981);
nand U3164 (N_3164,N_2577,N_2788);
and U3165 (N_3165,N_2560,N_2698);
or U3166 (N_3166,N_2672,N_2929);
or U3167 (N_3167,N_2986,N_2587);
nand U3168 (N_3168,N_2565,N_2870);
or U3169 (N_3169,N_2522,N_2802);
nand U3170 (N_3170,N_2909,N_2920);
nor U3171 (N_3171,N_2781,N_2754);
nand U3172 (N_3172,N_2707,N_2662);
and U3173 (N_3173,N_2509,N_2526);
xnor U3174 (N_3174,N_2779,N_2743);
nor U3175 (N_3175,N_2872,N_2973);
nand U3176 (N_3176,N_2896,N_2665);
nand U3177 (N_3177,N_2764,N_2926);
or U3178 (N_3178,N_2699,N_2939);
nand U3179 (N_3179,N_2742,N_2954);
and U3180 (N_3180,N_2563,N_2803);
or U3181 (N_3181,N_2863,N_2570);
or U3182 (N_3182,N_2792,N_2826);
nor U3183 (N_3183,N_2890,N_2968);
and U3184 (N_3184,N_2700,N_2663);
or U3185 (N_3185,N_2741,N_2822);
or U3186 (N_3186,N_2689,N_2659);
or U3187 (N_3187,N_2515,N_2730);
nor U3188 (N_3188,N_2650,N_2768);
nand U3189 (N_3189,N_2523,N_2550);
xor U3190 (N_3190,N_2664,N_2895);
nand U3191 (N_3191,N_2726,N_2796);
nand U3192 (N_3192,N_2505,N_2534);
and U3193 (N_3193,N_2721,N_2660);
and U3194 (N_3194,N_2804,N_2547);
or U3195 (N_3195,N_2912,N_2855);
or U3196 (N_3196,N_2995,N_2990);
or U3197 (N_3197,N_2578,N_2583);
xor U3198 (N_3198,N_2818,N_2910);
and U3199 (N_3199,N_2906,N_2574);
nor U3200 (N_3200,N_2532,N_2661);
nand U3201 (N_3201,N_2993,N_2829);
xnor U3202 (N_3202,N_2868,N_2908);
nand U3203 (N_3203,N_2609,N_2544);
nand U3204 (N_3204,N_2848,N_2602);
or U3205 (N_3205,N_2551,N_2994);
xnor U3206 (N_3206,N_2794,N_2814);
and U3207 (N_3207,N_2898,N_2566);
xnor U3208 (N_3208,N_2518,N_2722);
nand U3209 (N_3209,N_2789,N_2675);
nand U3210 (N_3210,N_2808,N_2676);
or U3211 (N_3211,N_2630,N_2705);
nor U3212 (N_3212,N_2969,N_2998);
xnor U3213 (N_3213,N_2959,N_2938);
nor U3214 (N_3214,N_2637,N_2593);
and U3215 (N_3215,N_2751,N_2611);
and U3216 (N_3216,N_2567,N_2824);
nand U3217 (N_3217,N_2784,N_2737);
xnor U3218 (N_3218,N_2614,N_2916);
nor U3219 (N_3219,N_2801,N_2854);
nor U3220 (N_3220,N_2940,N_2556);
xnor U3221 (N_3221,N_2955,N_2702);
and U3222 (N_3222,N_2584,N_2942);
nand U3223 (N_3223,N_2793,N_2739);
or U3224 (N_3224,N_2610,N_2632);
and U3225 (N_3225,N_2850,N_2703);
nor U3226 (N_3226,N_2748,N_2759);
nor U3227 (N_3227,N_2961,N_2667);
nor U3228 (N_3228,N_2646,N_2510);
nand U3229 (N_3229,N_2724,N_2972);
and U3230 (N_3230,N_2746,N_2693);
and U3231 (N_3231,N_2513,N_2586);
nor U3232 (N_3232,N_2841,N_2553);
or U3233 (N_3233,N_2561,N_2596);
nand U3234 (N_3234,N_2874,N_2821);
nand U3235 (N_3235,N_2696,N_2791);
and U3236 (N_3236,N_2914,N_2766);
xor U3237 (N_3237,N_2813,N_2536);
xor U3238 (N_3238,N_2622,N_2769);
nor U3239 (N_3239,N_2559,N_2851);
xnor U3240 (N_3240,N_2595,N_2734);
nor U3241 (N_3241,N_2948,N_2634);
and U3242 (N_3242,N_2554,N_2715);
nor U3243 (N_3243,N_2861,N_2656);
nand U3244 (N_3244,N_2883,N_2831);
nor U3245 (N_3245,N_2752,N_2626);
xor U3246 (N_3246,N_2798,N_2875);
or U3247 (N_3247,N_2679,N_2625);
nor U3248 (N_3248,N_2810,N_2652);
and U3249 (N_3249,N_2642,N_2557);
nor U3250 (N_3250,N_2780,N_2549);
or U3251 (N_3251,N_2962,N_2582);
nand U3252 (N_3252,N_2730,N_2768);
and U3253 (N_3253,N_2890,N_2891);
nand U3254 (N_3254,N_2688,N_2714);
nand U3255 (N_3255,N_2855,N_2535);
xnor U3256 (N_3256,N_2824,N_2605);
nor U3257 (N_3257,N_2633,N_2915);
nand U3258 (N_3258,N_2595,N_2654);
or U3259 (N_3259,N_2528,N_2636);
and U3260 (N_3260,N_2714,N_2535);
and U3261 (N_3261,N_2746,N_2999);
xor U3262 (N_3262,N_2500,N_2829);
or U3263 (N_3263,N_2612,N_2727);
nor U3264 (N_3264,N_2714,N_2760);
nor U3265 (N_3265,N_2624,N_2798);
xnor U3266 (N_3266,N_2755,N_2752);
xnor U3267 (N_3267,N_2973,N_2894);
and U3268 (N_3268,N_2974,N_2541);
nor U3269 (N_3269,N_2565,N_2852);
or U3270 (N_3270,N_2653,N_2553);
nand U3271 (N_3271,N_2644,N_2714);
nand U3272 (N_3272,N_2743,N_2653);
or U3273 (N_3273,N_2523,N_2641);
or U3274 (N_3274,N_2931,N_2784);
and U3275 (N_3275,N_2665,N_2611);
or U3276 (N_3276,N_2839,N_2670);
and U3277 (N_3277,N_2683,N_2963);
xnor U3278 (N_3278,N_2905,N_2852);
and U3279 (N_3279,N_2551,N_2561);
nor U3280 (N_3280,N_2720,N_2843);
xor U3281 (N_3281,N_2613,N_2532);
and U3282 (N_3282,N_2508,N_2948);
and U3283 (N_3283,N_2550,N_2804);
xnor U3284 (N_3284,N_2758,N_2915);
nand U3285 (N_3285,N_2746,N_2857);
and U3286 (N_3286,N_2730,N_2613);
nand U3287 (N_3287,N_2504,N_2818);
xor U3288 (N_3288,N_2924,N_2730);
xor U3289 (N_3289,N_2909,N_2581);
nor U3290 (N_3290,N_2509,N_2673);
xnor U3291 (N_3291,N_2634,N_2960);
or U3292 (N_3292,N_2822,N_2770);
or U3293 (N_3293,N_2718,N_2917);
nand U3294 (N_3294,N_2799,N_2767);
and U3295 (N_3295,N_2680,N_2973);
nand U3296 (N_3296,N_2951,N_2579);
and U3297 (N_3297,N_2570,N_2834);
nand U3298 (N_3298,N_2599,N_2741);
xnor U3299 (N_3299,N_2997,N_2508);
nor U3300 (N_3300,N_2829,N_2518);
or U3301 (N_3301,N_2751,N_2911);
nand U3302 (N_3302,N_2945,N_2964);
and U3303 (N_3303,N_2707,N_2518);
or U3304 (N_3304,N_2794,N_2972);
nor U3305 (N_3305,N_2544,N_2726);
nor U3306 (N_3306,N_2655,N_2574);
xnor U3307 (N_3307,N_2520,N_2617);
and U3308 (N_3308,N_2796,N_2958);
or U3309 (N_3309,N_2673,N_2528);
and U3310 (N_3310,N_2500,N_2896);
or U3311 (N_3311,N_2935,N_2967);
nor U3312 (N_3312,N_2607,N_2949);
nand U3313 (N_3313,N_2886,N_2690);
xnor U3314 (N_3314,N_2646,N_2920);
nor U3315 (N_3315,N_2634,N_2919);
or U3316 (N_3316,N_2518,N_2960);
xor U3317 (N_3317,N_2851,N_2792);
and U3318 (N_3318,N_2861,N_2531);
or U3319 (N_3319,N_2972,N_2504);
and U3320 (N_3320,N_2671,N_2845);
xor U3321 (N_3321,N_2931,N_2788);
nand U3322 (N_3322,N_2854,N_2803);
and U3323 (N_3323,N_2763,N_2932);
nand U3324 (N_3324,N_2900,N_2725);
or U3325 (N_3325,N_2969,N_2865);
xor U3326 (N_3326,N_2775,N_2783);
xnor U3327 (N_3327,N_2866,N_2593);
nand U3328 (N_3328,N_2865,N_2970);
nand U3329 (N_3329,N_2784,N_2805);
nand U3330 (N_3330,N_2646,N_2719);
nand U3331 (N_3331,N_2616,N_2915);
nand U3332 (N_3332,N_2924,N_2563);
and U3333 (N_3333,N_2500,N_2798);
nand U3334 (N_3334,N_2645,N_2809);
xor U3335 (N_3335,N_2820,N_2701);
nor U3336 (N_3336,N_2589,N_2503);
and U3337 (N_3337,N_2847,N_2906);
xor U3338 (N_3338,N_2601,N_2682);
or U3339 (N_3339,N_2736,N_2563);
or U3340 (N_3340,N_2917,N_2710);
or U3341 (N_3341,N_2580,N_2745);
nor U3342 (N_3342,N_2532,N_2758);
xnor U3343 (N_3343,N_2928,N_2647);
or U3344 (N_3344,N_2854,N_2500);
xnor U3345 (N_3345,N_2976,N_2666);
nand U3346 (N_3346,N_2724,N_2692);
and U3347 (N_3347,N_2563,N_2669);
nor U3348 (N_3348,N_2590,N_2834);
nand U3349 (N_3349,N_2672,N_2643);
and U3350 (N_3350,N_2550,N_2912);
and U3351 (N_3351,N_2684,N_2829);
or U3352 (N_3352,N_2899,N_2768);
nor U3353 (N_3353,N_2816,N_2852);
xor U3354 (N_3354,N_2651,N_2848);
nand U3355 (N_3355,N_2520,N_2759);
or U3356 (N_3356,N_2831,N_2704);
and U3357 (N_3357,N_2616,N_2813);
nand U3358 (N_3358,N_2912,N_2789);
nor U3359 (N_3359,N_2563,N_2730);
nor U3360 (N_3360,N_2904,N_2971);
and U3361 (N_3361,N_2815,N_2840);
nor U3362 (N_3362,N_2696,N_2930);
nand U3363 (N_3363,N_2539,N_2573);
nor U3364 (N_3364,N_2598,N_2811);
nor U3365 (N_3365,N_2765,N_2846);
or U3366 (N_3366,N_2513,N_2987);
and U3367 (N_3367,N_2790,N_2705);
xor U3368 (N_3368,N_2903,N_2835);
xor U3369 (N_3369,N_2598,N_2764);
nor U3370 (N_3370,N_2896,N_2686);
and U3371 (N_3371,N_2828,N_2770);
or U3372 (N_3372,N_2861,N_2738);
nor U3373 (N_3373,N_2909,N_2534);
nor U3374 (N_3374,N_2530,N_2809);
nand U3375 (N_3375,N_2883,N_2874);
nor U3376 (N_3376,N_2809,N_2520);
nor U3377 (N_3377,N_2598,N_2871);
nor U3378 (N_3378,N_2995,N_2767);
and U3379 (N_3379,N_2655,N_2511);
and U3380 (N_3380,N_2517,N_2759);
nand U3381 (N_3381,N_2755,N_2657);
and U3382 (N_3382,N_2872,N_2805);
and U3383 (N_3383,N_2717,N_2938);
and U3384 (N_3384,N_2581,N_2858);
and U3385 (N_3385,N_2811,N_2824);
nor U3386 (N_3386,N_2604,N_2768);
xor U3387 (N_3387,N_2636,N_2660);
nand U3388 (N_3388,N_2966,N_2858);
xnor U3389 (N_3389,N_2784,N_2535);
nor U3390 (N_3390,N_2952,N_2629);
nor U3391 (N_3391,N_2595,N_2582);
and U3392 (N_3392,N_2957,N_2944);
nand U3393 (N_3393,N_2869,N_2920);
nor U3394 (N_3394,N_2661,N_2837);
and U3395 (N_3395,N_2528,N_2838);
nand U3396 (N_3396,N_2516,N_2988);
nand U3397 (N_3397,N_2877,N_2692);
xnor U3398 (N_3398,N_2798,N_2789);
or U3399 (N_3399,N_2574,N_2963);
and U3400 (N_3400,N_2898,N_2872);
and U3401 (N_3401,N_2500,N_2879);
and U3402 (N_3402,N_2548,N_2771);
or U3403 (N_3403,N_2511,N_2843);
or U3404 (N_3404,N_2843,N_2854);
nand U3405 (N_3405,N_2622,N_2627);
and U3406 (N_3406,N_2821,N_2845);
nor U3407 (N_3407,N_2656,N_2545);
xnor U3408 (N_3408,N_2745,N_2531);
nor U3409 (N_3409,N_2501,N_2551);
nor U3410 (N_3410,N_2787,N_2933);
xnor U3411 (N_3411,N_2800,N_2743);
or U3412 (N_3412,N_2988,N_2713);
xor U3413 (N_3413,N_2698,N_2888);
nor U3414 (N_3414,N_2738,N_2997);
and U3415 (N_3415,N_2803,N_2864);
and U3416 (N_3416,N_2557,N_2880);
nor U3417 (N_3417,N_2778,N_2640);
xor U3418 (N_3418,N_2544,N_2692);
or U3419 (N_3419,N_2881,N_2504);
xor U3420 (N_3420,N_2885,N_2753);
or U3421 (N_3421,N_2525,N_2833);
nand U3422 (N_3422,N_2847,N_2536);
nand U3423 (N_3423,N_2726,N_2674);
nand U3424 (N_3424,N_2831,N_2691);
nand U3425 (N_3425,N_2778,N_2518);
nand U3426 (N_3426,N_2651,N_2582);
nand U3427 (N_3427,N_2763,N_2880);
nand U3428 (N_3428,N_2740,N_2806);
nor U3429 (N_3429,N_2597,N_2856);
nand U3430 (N_3430,N_2577,N_2650);
nor U3431 (N_3431,N_2642,N_2881);
or U3432 (N_3432,N_2554,N_2811);
nor U3433 (N_3433,N_2682,N_2642);
nand U3434 (N_3434,N_2778,N_2905);
nor U3435 (N_3435,N_2910,N_2887);
xnor U3436 (N_3436,N_2640,N_2771);
nand U3437 (N_3437,N_2816,N_2573);
nor U3438 (N_3438,N_2744,N_2736);
and U3439 (N_3439,N_2617,N_2682);
xor U3440 (N_3440,N_2591,N_2656);
and U3441 (N_3441,N_2689,N_2853);
nand U3442 (N_3442,N_2801,N_2567);
nor U3443 (N_3443,N_2832,N_2733);
nor U3444 (N_3444,N_2720,N_2583);
xor U3445 (N_3445,N_2658,N_2930);
nor U3446 (N_3446,N_2528,N_2839);
nand U3447 (N_3447,N_2615,N_2515);
xnor U3448 (N_3448,N_2623,N_2669);
or U3449 (N_3449,N_2560,N_2780);
nor U3450 (N_3450,N_2538,N_2914);
nor U3451 (N_3451,N_2841,N_2699);
and U3452 (N_3452,N_2636,N_2575);
nor U3453 (N_3453,N_2857,N_2779);
and U3454 (N_3454,N_2696,N_2803);
or U3455 (N_3455,N_2810,N_2558);
or U3456 (N_3456,N_2772,N_2992);
or U3457 (N_3457,N_2597,N_2710);
xnor U3458 (N_3458,N_2628,N_2962);
nand U3459 (N_3459,N_2951,N_2962);
or U3460 (N_3460,N_2629,N_2850);
or U3461 (N_3461,N_2867,N_2827);
xnor U3462 (N_3462,N_2547,N_2919);
and U3463 (N_3463,N_2815,N_2908);
and U3464 (N_3464,N_2633,N_2935);
and U3465 (N_3465,N_2787,N_2736);
and U3466 (N_3466,N_2990,N_2674);
xor U3467 (N_3467,N_2732,N_2555);
xor U3468 (N_3468,N_2502,N_2563);
and U3469 (N_3469,N_2628,N_2643);
nand U3470 (N_3470,N_2629,N_2944);
nand U3471 (N_3471,N_2796,N_2696);
and U3472 (N_3472,N_2642,N_2993);
or U3473 (N_3473,N_2880,N_2711);
or U3474 (N_3474,N_2777,N_2981);
and U3475 (N_3475,N_2556,N_2736);
nand U3476 (N_3476,N_2824,N_2701);
or U3477 (N_3477,N_2675,N_2727);
nand U3478 (N_3478,N_2950,N_2567);
or U3479 (N_3479,N_2736,N_2981);
nand U3480 (N_3480,N_2653,N_2988);
and U3481 (N_3481,N_2900,N_2689);
and U3482 (N_3482,N_2845,N_2735);
nand U3483 (N_3483,N_2890,N_2951);
and U3484 (N_3484,N_2773,N_2607);
nand U3485 (N_3485,N_2973,N_2713);
and U3486 (N_3486,N_2602,N_2517);
or U3487 (N_3487,N_2750,N_2709);
nor U3488 (N_3488,N_2777,N_2627);
nand U3489 (N_3489,N_2711,N_2816);
and U3490 (N_3490,N_2733,N_2554);
or U3491 (N_3491,N_2800,N_2952);
nand U3492 (N_3492,N_2717,N_2690);
and U3493 (N_3493,N_2649,N_2872);
and U3494 (N_3494,N_2539,N_2867);
and U3495 (N_3495,N_2610,N_2985);
nor U3496 (N_3496,N_2668,N_2979);
xnor U3497 (N_3497,N_2560,N_2749);
nor U3498 (N_3498,N_2626,N_2525);
or U3499 (N_3499,N_2829,N_2832);
or U3500 (N_3500,N_3025,N_3274);
nand U3501 (N_3501,N_3017,N_3233);
nand U3502 (N_3502,N_3270,N_3458);
xor U3503 (N_3503,N_3123,N_3186);
nand U3504 (N_3504,N_3333,N_3417);
nor U3505 (N_3505,N_3452,N_3448);
and U3506 (N_3506,N_3325,N_3214);
xor U3507 (N_3507,N_3153,N_3120);
and U3508 (N_3508,N_3354,N_3093);
nand U3509 (N_3509,N_3007,N_3192);
or U3510 (N_3510,N_3100,N_3241);
or U3511 (N_3511,N_3237,N_3356);
nor U3512 (N_3512,N_3175,N_3201);
nor U3513 (N_3513,N_3204,N_3286);
nor U3514 (N_3514,N_3482,N_3173);
nand U3515 (N_3515,N_3311,N_3495);
or U3516 (N_3516,N_3283,N_3171);
nand U3517 (N_3517,N_3329,N_3215);
and U3518 (N_3518,N_3338,N_3413);
or U3519 (N_3519,N_3009,N_3132);
nor U3520 (N_3520,N_3264,N_3036);
nand U3521 (N_3521,N_3468,N_3184);
xnor U3522 (N_3522,N_3365,N_3076);
nand U3523 (N_3523,N_3483,N_3141);
nand U3524 (N_3524,N_3383,N_3353);
nor U3525 (N_3525,N_3396,N_3190);
nor U3526 (N_3526,N_3053,N_3169);
or U3527 (N_3527,N_3364,N_3322);
and U3528 (N_3528,N_3045,N_3013);
nand U3529 (N_3529,N_3326,N_3112);
nand U3530 (N_3530,N_3081,N_3402);
nand U3531 (N_3531,N_3213,N_3397);
or U3532 (N_3532,N_3263,N_3341);
nand U3533 (N_3533,N_3472,N_3023);
and U3534 (N_3534,N_3390,N_3499);
xnor U3535 (N_3535,N_3208,N_3029);
nand U3536 (N_3536,N_3166,N_3267);
xnor U3537 (N_3537,N_3209,N_3463);
nor U3538 (N_3538,N_3371,N_3447);
xor U3539 (N_3539,N_3096,N_3276);
or U3540 (N_3540,N_3490,N_3005);
or U3541 (N_3541,N_3321,N_3350);
nand U3542 (N_3542,N_3497,N_3442);
nor U3543 (N_3543,N_3031,N_3072);
nor U3544 (N_3544,N_3145,N_3282);
nor U3545 (N_3545,N_3470,N_3052);
or U3546 (N_3546,N_3334,N_3489);
and U3547 (N_3547,N_3296,N_3420);
nand U3548 (N_3548,N_3273,N_3125);
or U3549 (N_3549,N_3484,N_3080);
xor U3550 (N_3550,N_3393,N_3091);
and U3551 (N_3551,N_3077,N_3000);
nor U3552 (N_3552,N_3070,N_3040);
nor U3553 (N_3553,N_3252,N_3224);
nand U3554 (N_3554,N_3436,N_3256);
nor U3555 (N_3555,N_3275,N_3126);
xnor U3556 (N_3556,N_3466,N_3340);
or U3557 (N_3557,N_3099,N_3083);
and U3558 (N_3558,N_3240,N_3058);
xor U3559 (N_3559,N_3084,N_3082);
xor U3560 (N_3560,N_3375,N_3183);
xnor U3561 (N_3561,N_3370,N_3459);
and U3562 (N_3562,N_3071,N_3360);
nor U3563 (N_3563,N_3016,N_3136);
xnor U3564 (N_3564,N_3376,N_3246);
nand U3565 (N_3565,N_3272,N_3288);
nor U3566 (N_3566,N_3069,N_3254);
and U3567 (N_3567,N_3403,N_3431);
nand U3568 (N_3568,N_3199,N_3422);
xnor U3569 (N_3569,N_3328,N_3225);
xnor U3570 (N_3570,N_3444,N_3122);
nand U3571 (N_3571,N_3331,N_3379);
nand U3572 (N_3572,N_3172,N_3075);
and U3573 (N_3573,N_3293,N_3137);
or U3574 (N_3574,N_3027,N_3011);
and U3575 (N_3575,N_3302,N_3419);
xnor U3576 (N_3576,N_3150,N_3382);
or U3577 (N_3577,N_3211,N_3299);
nand U3578 (N_3578,N_3079,N_3266);
nor U3579 (N_3579,N_3102,N_3094);
nor U3580 (N_3580,N_3163,N_3074);
or U3581 (N_3581,N_3400,N_3314);
or U3582 (N_3582,N_3337,N_3368);
and U3583 (N_3583,N_3312,N_3012);
nand U3584 (N_3584,N_3301,N_3015);
or U3585 (N_3585,N_3164,N_3279);
nand U3586 (N_3586,N_3129,N_3307);
nor U3587 (N_3587,N_3243,N_3244);
and U3588 (N_3588,N_3180,N_3048);
or U3589 (N_3589,N_3151,N_3496);
or U3590 (N_3590,N_3265,N_3221);
nor U3591 (N_3591,N_3441,N_3154);
or U3592 (N_3592,N_3097,N_3373);
nand U3593 (N_3593,N_3462,N_3219);
nand U3594 (N_3594,N_3366,N_3453);
and U3595 (N_3595,N_3471,N_3239);
xor U3596 (N_3596,N_3090,N_3167);
nand U3597 (N_3597,N_3140,N_3234);
or U3598 (N_3598,N_3253,N_3037);
nand U3599 (N_3599,N_3238,N_3477);
nor U3600 (N_3600,N_3106,N_3491);
and U3601 (N_3601,N_3412,N_3161);
and U3602 (N_3602,N_3101,N_3024);
and U3603 (N_3603,N_3144,N_3158);
xnor U3604 (N_3604,N_3454,N_3380);
or U3605 (N_3605,N_3255,N_3050);
and U3606 (N_3606,N_3271,N_3259);
nor U3607 (N_3607,N_3345,N_3139);
xnor U3608 (N_3608,N_3210,N_3377);
and U3609 (N_3609,N_3168,N_3087);
xor U3610 (N_3610,N_3235,N_3010);
or U3611 (N_3611,N_3105,N_3443);
and U3612 (N_3612,N_3474,N_3033);
nor U3613 (N_3613,N_3086,N_3218);
xor U3614 (N_3614,N_3438,N_3202);
xnor U3615 (N_3615,N_3044,N_3404);
or U3616 (N_3616,N_3284,N_3498);
and U3617 (N_3617,N_3116,N_3188);
xor U3618 (N_3618,N_3135,N_3232);
or U3619 (N_3619,N_3295,N_3064);
xnor U3620 (N_3620,N_3460,N_3392);
nor U3621 (N_3621,N_3156,N_3281);
nand U3622 (N_3622,N_3449,N_3378);
or U3623 (N_3623,N_3309,N_3138);
xnor U3624 (N_3624,N_3313,N_3065);
nor U3625 (N_3625,N_3230,N_3361);
xor U3626 (N_3626,N_3303,N_3111);
or U3627 (N_3627,N_3424,N_3191);
nand U3628 (N_3628,N_3160,N_3318);
xnor U3629 (N_3629,N_3001,N_3268);
xnor U3630 (N_3630,N_3056,N_3467);
and U3631 (N_3631,N_3432,N_3063);
xor U3632 (N_3632,N_3465,N_3359);
nand U3633 (N_3633,N_3133,N_3428);
xnor U3634 (N_3634,N_3294,N_3363);
or U3635 (N_3635,N_3369,N_3030);
and U3636 (N_3636,N_3385,N_3226);
nand U3637 (N_3637,N_3475,N_3389);
nor U3638 (N_3638,N_3049,N_3236);
nor U3639 (N_3639,N_3060,N_3486);
xor U3640 (N_3640,N_3195,N_3223);
nor U3641 (N_3641,N_3391,N_3405);
nand U3642 (N_3642,N_3217,N_3026);
nand U3643 (N_3643,N_3189,N_3054);
nand U3644 (N_3644,N_3018,N_3316);
or U3645 (N_3645,N_3034,N_3127);
or U3646 (N_3646,N_3117,N_3249);
xnor U3647 (N_3647,N_3014,N_3348);
nor U3648 (N_3648,N_3410,N_3411);
nor U3649 (N_3649,N_3261,N_3386);
xnor U3650 (N_3650,N_3019,N_3388);
nand U3651 (N_3651,N_3062,N_3197);
nand U3652 (N_3652,N_3165,N_3146);
xnor U3653 (N_3653,N_3229,N_3245);
and U3654 (N_3654,N_3124,N_3032);
xor U3655 (N_3655,N_3046,N_3148);
or U3656 (N_3656,N_3004,N_3194);
or U3657 (N_3657,N_3352,N_3319);
xnor U3658 (N_3658,N_3399,N_3178);
nor U3659 (N_3659,N_3473,N_3055);
nor U3660 (N_3660,N_3078,N_3297);
nand U3661 (N_3661,N_3061,N_3258);
nand U3662 (N_3662,N_3176,N_3152);
or U3663 (N_3663,N_3203,N_3398);
xnor U3664 (N_3664,N_3437,N_3181);
nor U3665 (N_3665,N_3439,N_3315);
or U3666 (N_3666,N_3035,N_3287);
and U3667 (N_3667,N_3022,N_3242);
or U3668 (N_3668,N_3006,N_3095);
or U3669 (N_3669,N_3142,N_3248);
nor U3670 (N_3670,N_3343,N_3205);
nor U3671 (N_3671,N_3308,N_3415);
or U3672 (N_3672,N_3357,N_3098);
or U3673 (N_3673,N_3469,N_3277);
or U3674 (N_3674,N_3231,N_3433);
xnor U3675 (N_3675,N_3162,N_3485);
or U3676 (N_3676,N_3119,N_3028);
nand U3677 (N_3677,N_3409,N_3440);
or U3678 (N_3678,N_3347,N_3488);
xnor U3679 (N_3679,N_3220,N_3320);
nor U3680 (N_3680,N_3250,N_3446);
nand U3681 (N_3681,N_3157,N_3107);
or U3682 (N_3682,N_3342,N_3159);
and U3683 (N_3683,N_3479,N_3193);
or U3684 (N_3684,N_3324,N_3306);
or U3685 (N_3685,N_3073,N_3198);
nor U3686 (N_3686,N_3381,N_3110);
and U3687 (N_3687,N_3323,N_3174);
nor U3688 (N_3688,N_3108,N_3332);
nand U3689 (N_3689,N_3427,N_3425);
or U3690 (N_3690,N_3304,N_3416);
and U3691 (N_3691,N_3290,N_3351);
nand U3692 (N_3692,N_3008,N_3057);
and U3693 (N_3693,N_3051,N_3260);
nand U3694 (N_3694,N_3021,N_3131);
xor U3695 (N_3695,N_3104,N_3450);
or U3696 (N_3696,N_3109,N_3251);
and U3697 (N_3697,N_3113,N_3280);
or U3698 (N_3698,N_3430,N_3434);
or U3699 (N_3699,N_3121,N_3085);
or U3700 (N_3700,N_3003,N_3187);
nand U3701 (N_3701,N_3374,N_3336);
nand U3702 (N_3702,N_3339,N_3196);
nor U3703 (N_3703,N_3464,N_3041);
xnor U3704 (N_3704,N_3043,N_3414);
or U3705 (N_3705,N_3092,N_3384);
nor U3706 (N_3706,N_3421,N_3401);
or U3707 (N_3707,N_3118,N_3227);
and U3708 (N_3708,N_3222,N_3408);
xor U3709 (N_3709,N_3066,N_3426);
xor U3710 (N_3710,N_3406,N_3456);
xnor U3711 (N_3711,N_3372,N_3039);
xnor U3712 (N_3712,N_3269,N_3327);
and U3713 (N_3713,N_3206,N_3114);
nor U3714 (N_3714,N_3278,N_3247);
nor U3715 (N_3715,N_3185,N_3300);
xor U3716 (N_3716,N_3346,N_3262);
xor U3717 (N_3717,N_3335,N_3291);
xnor U3718 (N_3718,N_3494,N_3394);
nand U3719 (N_3719,N_3423,N_3115);
nor U3720 (N_3720,N_3289,N_3493);
nor U3721 (N_3721,N_3445,N_3429);
xnor U3722 (N_3722,N_3047,N_3042);
or U3723 (N_3723,N_3310,N_3182);
xnor U3724 (N_3724,N_3305,N_3395);
nor U3725 (N_3725,N_3207,N_3200);
xor U3726 (N_3726,N_3367,N_3317);
or U3727 (N_3727,N_3088,N_3147);
and U3728 (N_3728,N_3068,N_3038);
and U3729 (N_3729,N_3387,N_3002);
nand U3730 (N_3730,N_3355,N_3179);
xnor U3731 (N_3731,N_3358,N_3487);
xnor U3732 (N_3732,N_3130,N_3103);
nor U3733 (N_3733,N_3461,N_3418);
or U3734 (N_3734,N_3457,N_3344);
nor U3735 (N_3735,N_3149,N_3089);
nor U3736 (N_3736,N_3476,N_3481);
nor U3737 (N_3737,N_3298,N_3407);
nand U3738 (N_3738,N_3059,N_3134);
nor U3739 (N_3739,N_3285,N_3451);
nor U3740 (N_3740,N_3170,N_3455);
or U3741 (N_3741,N_3128,N_3330);
xnor U3742 (N_3742,N_3155,N_3292);
nor U3743 (N_3743,N_3020,N_3216);
nand U3744 (N_3744,N_3257,N_3212);
nand U3745 (N_3745,N_3349,N_3177);
nor U3746 (N_3746,N_3143,N_3067);
nor U3747 (N_3747,N_3492,N_3480);
nand U3748 (N_3748,N_3228,N_3362);
xor U3749 (N_3749,N_3478,N_3435);
nand U3750 (N_3750,N_3039,N_3330);
nor U3751 (N_3751,N_3277,N_3370);
nor U3752 (N_3752,N_3145,N_3122);
nor U3753 (N_3753,N_3397,N_3091);
xnor U3754 (N_3754,N_3063,N_3142);
nand U3755 (N_3755,N_3166,N_3118);
xor U3756 (N_3756,N_3284,N_3338);
xnor U3757 (N_3757,N_3327,N_3449);
and U3758 (N_3758,N_3215,N_3412);
xor U3759 (N_3759,N_3107,N_3399);
nor U3760 (N_3760,N_3210,N_3400);
and U3761 (N_3761,N_3094,N_3367);
xnor U3762 (N_3762,N_3257,N_3439);
nor U3763 (N_3763,N_3073,N_3351);
nor U3764 (N_3764,N_3417,N_3409);
or U3765 (N_3765,N_3121,N_3367);
xnor U3766 (N_3766,N_3201,N_3474);
nand U3767 (N_3767,N_3076,N_3481);
nor U3768 (N_3768,N_3420,N_3451);
nor U3769 (N_3769,N_3070,N_3440);
nor U3770 (N_3770,N_3059,N_3365);
xor U3771 (N_3771,N_3201,N_3104);
and U3772 (N_3772,N_3071,N_3244);
xnor U3773 (N_3773,N_3106,N_3287);
or U3774 (N_3774,N_3267,N_3377);
nand U3775 (N_3775,N_3216,N_3068);
or U3776 (N_3776,N_3042,N_3081);
and U3777 (N_3777,N_3455,N_3160);
or U3778 (N_3778,N_3262,N_3137);
nor U3779 (N_3779,N_3115,N_3419);
xnor U3780 (N_3780,N_3233,N_3027);
or U3781 (N_3781,N_3492,N_3251);
or U3782 (N_3782,N_3401,N_3191);
or U3783 (N_3783,N_3495,N_3365);
nor U3784 (N_3784,N_3145,N_3227);
xor U3785 (N_3785,N_3078,N_3412);
and U3786 (N_3786,N_3221,N_3375);
nor U3787 (N_3787,N_3058,N_3497);
nor U3788 (N_3788,N_3371,N_3240);
xor U3789 (N_3789,N_3088,N_3000);
xnor U3790 (N_3790,N_3210,N_3229);
nand U3791 (N_3791,N_3249,N_3464);
nor U3792 (N_3792,N_3333,N_3460);
nor U3793 (N_3793,N_3410,N_3348);
nand U3794 (N_3794,N_3235,N_3206);
or U3795 (N_3795,N_3226,N_3269);
or U3796 (N_3796,N_3011,N_3364);
nor U3797 (N_3797,N_3163,N_3353);
nand U3798 (N_3798,N_3391,N_3438);
nand U3799 (N_3799,N_3317,N_3102);
nor U3800 (N_3800,N_3220,N_3465);
xor U3801 (N_3801,N_3430,N_3301);
or U3802 (N_3802,N_3309,N_3411);
or U3803 (N_3803,N_3031,N_3041);
or U3804 (N_3804,N_3468,N_3085);
nor U3805 (N_3805,N_3493,N_3201);
xnor U3806 (N_3806,N_3310,N_3139);
and U3807 (N_3807,N_3102,N_3148);
or U3808 (N_3808,N_3139,N_3321);
xor U3809 (N_3809,N_3349,N_3364);
xnor U3810 (N_3810,N_3249,N_3010);
nor U3811 (N_3811,N_3279,N_3168);
or U3812 (N_3812,N_3417,N_3204);
xor U3813 (N_3813,N_3409,N_3426);
or U3814 (N_3814,N_3373,N_3272);
nand U3815 (N_3815,N_3483,N_3148);
xnor U3816 (N_3816,N_3276,N_3071);
or U3817 (N_3817,N_3148,N_3336);
xor U3818 (N_3818,N_3410,N_3210);
and U3819 (N_3819,N_3259,N_3047);
nand U3820 (N_3820,N_3032,N_3130);
nor U3821 (N_3821,N_3160,N_3458);
xnor U3822 (N_3822,N_3007,N_3479);
and U3823 (N_3823,N_3248,N_3298);
xor U3824 (N_3824,N_3219,N_3031);
xnor U3825 (N_3825,N_3325,N_3441);
xnor U3826 (N_3826,N_3287,N_3065);
and U3827 (N_3827,N_3353,N_3454);
nand U3828 (N_3828,N_3206,N_3394);
or U3829 (N_3829,N_3188,N_3239);
and U3830 (N_3830,N_3464,N_3010);
nor U3831 (N_3831,N_3333,N_3437);
nand U3832 (N_3832,N_3226,N_3180);
nor U3833 (N_3833,N_3024,N_3034);
nor U3834 (N_3834,N_3080,N_3395);
and U3835 (N_3835,N_3097,N_3350);
or U3836 (N_3836,N_3328,N_3164);
nand U3837 (N_3837,N_3146,N_3324);
nor U3838 (N_3838,N_3344,N_3473);
and U3839 (N_3839,N_3044,N_3345);
nor U3840 (N_3840,N_3473,N_3386);
nand U3841 (N_3841,N_3490,N_3182);
xnor U3842 (N_3842,N_3444,N_3259);
xor U3843 (N_3843,N_3436,N_3053);
and U3844 (N_3844,N_3139,N_3129);
xnor U3845 (N_3845,N_3021,N_3479);
nand U3846 (N_3846,N_3376,N_3163);
nand U3847 (N_3847,N_3168,N_3016);
and U3848 (N_3848,N_3023,N_3284);
or U3849 (N_3849,N_3116,N_3386);
and U3850 (N_3850,N_3162,N_3199);
nor U3851 (N_3851,N_3366,N_3372);
and U3852 (N_3852,N_3434,N_3174);
or U3853 (N_3853,N_3255,N_3243);
nor U3854 (N_3854,N_3153,N_3400);
or U3855 (N_3855,N_3134,N_3148);
xor U3856 (N_3856,N_3332,N_3111);
nor U3857 (N_3857,N_3207,N_3402);
or U3858 (N_3858,N_3376,N_3060);
nor U3859 (N_3859,N_3329,N_3316);
nor U3860 (N_3860,N_3086,N_3232);
nor U3861 (N_3861,N_3313,N_3320);
and U3862 (N_3862,N_3448,N_3490);
nor U3863 (N_3863,N_3111,N_3393);
xnor U3864 (N_3864,N_3184,N_3033);
nor U3865 (N_3865,N_3366,N_3036);
xor U3866 (N_3866,N_3024,N_3482);
xor U3867 (N_3867,N_3331,N_3332);
and U3868 (N_3868,N_3496,N_3229);
xor U3869 (N_3869,N_3006,N_3245);
nor U3870 (N_3870,N_3325,N_3270);
nor U3871 (N_3871,N_3174,N_3142);
and U3872 (N_3872,N_3135,N_3244);
nand U3873 (N_3873,N_3095,N_3130);
xor U3874 (N_3874,N_3325,N_3066);
or U3875 (N_3875,N_3207,N_3239);
nand U3876 (N_3876,N_3173,N_3409);
or U3877 (N_3877,N_3077,N_3457);
nand U3878 (N_3878,N_3315,N_3499);
xor U3879 (N_3879,N_3376,N_3379);
or U3880 (N_3880,N_3322,N_3361);
nor U3881 (N_3881,N_3086,N_3491);
xor U3882 (N_3882,N_3186,N_3371);
xnor U3883 (N_3883,N_3342,N_3423);
xnor U3884 (N_3884,N_3415,N_3419);
or U3885 (N_3885,N_3427,N_3484);
or U3886 (N_3886,N_3247,N_3065);
or U3887 (N_3887,N_3441,N_3388);
xnor U3888 (N_3888,N_3425,N_3261);
and U3889 (N_3889,N_3006,N_3048);
or U3890 (N_3890,N_3046,N_3190);
nor U3891 (N_3891,N_3155,N_3362);
nand U3892 (N_3892,N_3096,N_3272);
and U3893 (N_3893,N_3275,N_3343);
and U3894 (N_3894,N_3385,N_3408);
nand U3895 (N_3895,N_3493,N_3257);
xor U3896 (N_3896,N_3331,N_3429);
or U3897 (N_3897,N_3082,N_3222);
and U3898 (N_3898,N_3323,N_3232);
xnor U3899 (N_3899,N_3082,N_3319);
or U3900 (N_3900,N_3263,N_3336);
nand U3901 (N_3901,N_3409,N_3287);
and U3902 (N_3902,N_3031,N_3367);
or U3903 (N_3903,N_3049,N_3111);
nor U3904 (N_3904,N_3279,N_3145);
and U3905 (N_3905,N_3353,N_3447);
nand U3906 (N_3906,N_3416,N_3309);
xor U3907 (N_3907,N_3272,N_3061);
nor U3908 (N_3908,N_3491,N_3040);
or U3909 (N_3909,N_3000,N_3264);
nor U3910 (N_3910,N_3348,N_3361);
and U3911 (N_3911,N_3142,N_3440);
nor U3912 (N_3912,N_3118,N_3434);
nor U3913 (N_3913,N_3182,N_3168);
or U3914 (N_3914,N_3442,N_3096);
or U3915 (N_3915,N_3392,N_3455);
or U3916 (N_3916,N_3126,N_3407);
and U3917 (N_3917,N_3385,N_3186);
and U3918 (N_3918,N_3154,N_3274);
nor U3919 (N_3919,N_3314,N_3376);
xnor U3920 (N_3920,N_3367,N_3049);
xnor U3921 (N_3921,N_3017,N_3327);
nand U3922 (N_3922,N_3470,N_3422);
nand U3923 (N_3923,N_3095,N_3431);
or U3924 (N_3924,N_3083,N_3291);
xnor U3925 (N_3925,N_3469,N_3323);
nand U3926 (N_3926,N_3456,N_3179);
and U3927 (N_3927,N_3030,N_3201);
nor U3928 (N_3928,N_3458,N_3065);
xnor U3929 (N_3929,N_3110,N_3355);
xnor U3930 (N_3930,N_3219,N_3133);
or U3931 (N_3931,N_3126,N_3150);
nand U3932 (N_3932,N_3479,N_3294);
and U3933 (N_3933,N_3383,N_3491);
or U3934 (N_3934,N_3460,N_3048);
and U3935 (N_3935,N_3438,N_3485);
nand U3936 (N_3936,N_3290,N_3342);
xnor U3937 (N_3937,N_3194,N_3271);
nand U3938 (N_3938,N_3011,N_3073);
nor U3939 (N_3939,N_3009,N_3221);
and U3940 (N_3940,N_3320,N_3180);
or U3941 (N_3941,N_3494,N_3401);
nand U3942 (N_3942,N_3474,N_3303);
or U3943 (N_3943,N_3159,N_3497);
and U3944 (N_3944,N_3153,N_3469);
nor U3945 (N_3945,N_3046,N_3138);
and U3946 (N_3946,N_3289,N_3271);
nor U3947 (N_3947,N_3058,N_3337);
nor U3948 (N_3948,N_3255,N_3456);
xor U3949 (N_3949,N_3175,N_3103);
and U3950 (N_3950,N_3240,N_3156);
nor U3951 (N_3951,N_3175,N_3034);
nand U3952 (N_3952,N_3008,N_3428);
or U3953 (N_3953,N_3415,N_3460);
or U3954 (N_3954,N_3485,N_3403);
nand U3955 (N_3955,N_3143,N_3344);
xnor U3956 (N_3956,N_3311,N_3371);
or U3957 (N_3957,N_3118,N_3248);
xnor U3958 (N_3958,N_3465,N_3090);
nor U3959 (N_3959,N_3029,N_3062);
or U3960 (N_3960,N_3378,N_3256);
or U3961 (N_3961,N_3384,N_3016);
nor U3962 (N_3962,N_3225,N_3050);
nor U3963 (N_3963,N_3379,N_3162);
nor U3964 (N_3964,N_3089,N_3138);
xnor U3965 (N_3965,N_3353,N_3171);
nand U3966 (N_3966,N_3308,N_3049);
or U3967 (N_3967,N_3457,N_3066);
or U3968 (N_3968,N_3099,N_3102);
nor U3969 (N_3969,N_3441,N_3464);
or U3970 (N_3970,N_3461,N_3075);
and U3971 (N_3971,N_3181,N_3051);
and U3972 (N_3972,N_3091,N_3322);
and U3973 (N_3973,N_3330,N_3111);
and U3974 (N_3974,N_3074,N_3309);
and U3975 (N_3975,N_3041,N_3153);
nand U3976 (N_3976,N_3191,N_3149);
nand U3977 (N_3977,N_3368,N_3358);
and U3978 (N_3978,N_3295,N_3008);
or U3979 (N_3979,N_3390,N_3429);
xnor U3980 (N_3980,N_3447,N_3412);
xnor U3981 (N_3981,N_3473,N_3070);
nor U3982 (N_3982,N_3128,N_3021);
and U3983 (N_3983,N_3102,N_3379);
xor U3984 (N_3984,N_3024,N_3433);
nand U3985 (N_3985,N_3275,N_3097);
xor U3986 (N_3986,N_3428,N_3296);
xnor U3987 (N_3987,N_3171,N_3112);
nand U3988 (N_3988,N_3420,N_3403);
or U3989 (N_3989,N_3462,N_3428);
nand U3990 (N_3990,N_3179,N_3419);
nand U3991 (N_3991,N_3382,N_3088);
or U3992 (N_3992,N_3085,N_3499);
xor U3993 (N_3993,N_3268,N_3404);
and U3994 (N_3994,N_3203,N_3130);
or U3995 (N_3995,N_3285,N_3288);
or U3996 (N_3996,N_3302,N_3290);
xor U3997 (N_3997,N_3292,N_3267);
or U3998 (N_3998,N_3213,N_3349);
xor U3999 (N_3999,N_3157,N_3396);
xnor U4000 (N_4000,N_3766,N_3843);
xor U4001 (N_4001,N_3706,N_3791);
or U4002 (N_4002,N_3880,N_3730);
and U4003 (N_4003,N_3670,N_3871);
nand U4004 (N_4004,N_3907,N_3870);
or U4005 (N_4005,N_3586,N_3527);
xnor U4006 (N_4006,N_3583,N_3787);
or U4007 (N_4007,N_3926,N_3979);
xor U4008 (N_4008,N_3633,N_3933);
or U4009 (N_4009,N_3585,N_3705);
nor U4010 (N_4010,N_3686,N_3785);
nand U4011 (N_4011,N_3923,N_3515);
nand U4012 (N_4012,N_3577,N_3797);
and U4013 (N_4013,N_3507,N_3689);
xor U4014 (N_4014,N_3734,N_3779);
or U4015 (N_4015,N_3827,N_3680);
nor U4016 (N_4016,N_3549,N_3852);
or U4017 (N_4017,N_3988,N_3716);
xnor U4018 (N_4018,N_3816,N_3719);
and U4019 (N_4019,N_3729,N_3920);
nor U4020 (N_4020,N_3715,N_3864);
nor U4021 (N_4021,N_3838,N_3620);
nor U4022 (N_4022,N_3755,N_3641);
xnor U4023 (N_4023,N_3846,N_3899);
nand U4024 (N_4024,N_3690,N_3801);
nor U4025 (N_4025,N_3661,N_3989);
and U4026 (N_4026,N_3713,N_3834);
xnor U4027 (N_4027,N_3731,N_3921);
nor U4028 (N_4028,N_3688,N_3974);
nor U4029 (N_4029,N_3879,N_3819);
xnor U4030 (N_4030,N_3558,N_3998);
xnor U4031 (N_4031,N_3721,N_3659);
xor U4032 (N_4032,N_3683,N_3516);
xnor U4033 (N_4033,N_3518,N_3556);
or U4034 (N_4034,N_3836,N_3963);
and U4035 (N_4035,N_3636,N_3997);
nor U4036 (N_4036,N_3931,N_3991);
nor U4037 (N_4037,N_3622,N_3693);
and U4038 (N_4038,N_3543,N_3678);
nand U4039 (N_4039,N_3874,N_3614);
nand U4040 (N_4040,N_3775,N_3742);
nor U4041 (N_4041,N_3948,N_3635);
or U4042 (N_4042,N_3526,N_3833);
nand U4043 (N_4043,N_3668,N_3523);
xor U4044 (N_4044,N_3859,N_3664);
nand U4045 (N_4045,N_3889,N_3563);
nor U4046 (N_4046,N_3517,N_3919);
xnor U4047 (N_4047,N_3888,N_3799);
xor U4048 (N_4048,N_3818,N_3831);
nand U4049 (N_4049,N_3732,N_3821);
and U4050 (N_4050,N_3545,N_3908);
nand U4051 (N_4051,N_3590,N_3944);
nand U4052 (N_4052,N_3939,N_3582);
nand U4053 (N_4053,N_3519,N_3924);
nand U4054 (N_4054,N_3798,N_3762);
xnor U4055 (N_4055,N_3863,N_3739);
and U4056 (N_4056,N_3576,N_3560);
nand U4057 (N_4057,N_3937,N_3538);
or U4058 (N_4058,N_3595,N_3749);
nand U4059 (N_4059,N_3505,N_3840);
or U4060 (N_4060,N_3929,N_3587);
or U4061 (N_4061,N_3682,N_3610);
nand U4062 (N_4062,N_3566,N_3504);
or U4063 (N_4063,N_3905,N_3599);
xnor U4064 (N_4064,N_3783,N_3769);
or U4065 (N_4065,N_3649,N_3972);
xnor U4066 (N_4066,N_3913,N_3892);
xor U4067 (N_4067,N_3665,N_3945);
or U4068 (N_4068,N_3709,N_3890);
nand U4069 (N_4069,N_3814,N_3660);
or U4070 (N_4070,N_3841,N_3579);
nand U4071 (N_4071,N_3760,N_3868);
nor U4072 (N_4072,N_3946,N_3956);
nand U4073 (N_4073,N_3758,N_3860);
nand U4074 (N_4074,N_3973,N_3652);
and U4075 (N_4075,N_3906,N_3904);
or U4076 (N_4076,N_3826,N_3932);
nand U4077 (N_4077,N_3949,N_3565);
nand U4078 (N_4078,N_3609,N_3621);
or U4079 (N_4079,N_3681,N_3789);
or U4080 (N_4080,N_3741,N_3695);
xnor U4081 (N_4081,N_3679,N_3663);
nand U4082 (N_4082,N_3521,N_3725);
nor U4083 (N_4083,N_3938,N_3829);
or U4084 (N_4084,N_3568,N_3772);
xor U4085 (N_4085,N_3915,N_3588);
nor U4086 (N_4086,N_3650,N_3809);
xnor U4087 (N_4087,N_3562,N_3986);
nand U4088 (N_4088,N_3786,N_3625);
or U4089 (N_4089,N_3965,N_3942);
nand U4090 (N_4090,N_3858,N_3528);
nand U4091 (N_4091,N_3959,N_3940);
nor U4092 (N_4092,N_3631,N_3862);
nand U4093 (N_4093,N_3765,N_3856);
nand U4094 (N_4094,N_3896,N_3849);
xnor U4095 (N_4095,N_3736,N_3756);
nand U4096 (N_4096,N_3669,N_3574);
nand U4097 (N_4097,N_3780,N_3916);
or U4098 (N_4098,N_3532,N_3615);
nor U4099 (N_4099,N_3509,N_3687);
or U4100 (N_4100,N_3651,N_3629);
nand U4101 (N_4101,N_3624,N_3943);
and U4102 (N_4102,N_3600,N_3975);
nor U4103 (N_4103,N_3544,N_3684);
xnor U4104 (N_4104,N_3767,N_3807);
and U4105 (N_4105,N_3551,N_3601);
xnor U4106 (N_4106,N_3676,N_3643);
xor U4107 (N_4107,N_3744,N_3570);
nand U4108 (N_4108,N_3591,N_3995);
xnor U4109 (N_4109,N_3983,N_3522);
or U4110 (N_4110,N_3993,N_3984);
and U4111 (N_4111,N_3540,N_3738);
nor U4112 (N_4112,N_3722,N_3724);
and U4113 (N_4113,N_3881,N_3764);
nor U4114 (N_4114,N_3808,N_3753);
xnor U4115 (N_4115,N_3746,N_3968);
and U4116 (N_4116,N_3961,N_3637);
and U4117 (N_4117,N_3578,N_3674);
nand U4118 (N_4118,N_3817,N_3593);
or U4119 (N_4119,N_3820,N_3876);
nand U4120 (N_4120,N_3812,N_3966);
nand U4121 (N_4121,N_3743,N_3605);
nand U4122 (N_4122,N_3805,N_3553);
xor U4123 (N_4123,N_3964,N_3781);
xnor U4124 (N_4124,N_3550,N_3960);
xnor U4125 (N_4125,N_3694,N_3941);
nor U4126 (N_4126,N_3733,N_3604);
or U4127 (N_4127,N_3757,N_3999);
nand U4128 (N_4128,N_3928,N_3717);
nand U4129 (N_4129,N_3912,N_3955);
nor U4130 (N_4130,N_3514,N_3763);
or U4131 (N_4131,N_3703,N_3697);
or U4132 (N_4132,N_3878,N_3866);
or U4133 (N_4133,N_3950,N_3842);
nand U4134 (N_4134,N_3559,N_3897);
nor U4135 (N_4135,N_3525,N_3754);
or U4136 (N_4136,N_3875,N_3934);
nor U4137 (N_4137,N_3745,N_3813);
or U4138 (N_4138,N_3692,N_3784);
xnor U4139 (N_4139,N_3996,N_3770);
nor U4140 (N_4140,N_3911,N_3554);
nand U4141 (N_4141,N_3580,N_3796);
xor U4142 (N_4142,N_3804,N_3644);
or U4143 (N_4143,N_3704,N_3894);
and U4144 (N_4144,N_3608,N_3909);
nor U4145 (N_4145,N_3882,N_3639);
nand U4146 (N_4146,N_3853,N_3634);
nand U4147 (N_4147,N_3822,N_3778);
xor U4148 (N_4148,N_3501,N_3655);
or U4149 (N_4149,N_3985,N_3832);
xnor U4150 (N_4150,N_3656,N_3930);
nand U4151 (N_4151,N_3830,N_3638);
or U4152 (N_4152,N_3978,N_3511);
xnor U4153 (N_4153,N_3954,N_3869);
nand U4154 (N_4154,N_3802,N_3837);
or U4155 (N_4155,N_3803,N_3536);
xnor U4156 (N_4156,N_3728,N_3951);
and U4157 (N_4157,N_3740,N_3542);
nor U4158 (N_4158,N_3546,N_3512);
xor U4159 (N_4159,N_3750,N_3500);
and U4160 (N_4160,N_3782,N_3606);
nand U4161 (N_4161,N_3596,N_3994);
and U4162 (N_4162,N_3701,N_3971);
nor U4163 (N_4163,N_3761,N_3794);
nor U4164 (N_4164,N_3602,N_3903);
nand U4165 (N_4165,N_3675,N_3710);
nor U4166 (N_4166,N_3751,N_3877);
or U4167 (N_4167,N_3584,N_3917);
and U4168 (N_4168,N_3886,N_3564);
or U4169 (N_4169,N_3530,N_3673);
xnor U4170 (N_4170,N_3884,N_3845);
xor U4171 (N_4171,N_3508,N_3571);
nor U4172 (N_4172,N_3976,N_3748);
xnor U4173 (N_4173,N_3777,N_3502);
nand U4174 (N_4174,N_3541,N_3967);
nor U4175 (N_4175,N_3539,N_3616);
or U4176 (N_4176,N_3691,N_3700);
nand U4177 (N_4177,N_3922,N_3828);
and U4178 (N_4178,N_3806,N_3685);
nand U4179 (N_4179,N_3646,N_3914);
and U4180 (N_4180,N_3752,N_3552);
nor U4181 (N_4181,N_3824,N_3788);
nand U4182 (N_4182,N_3657,N_3531);
or U4183 (N_4183,N_3815,N_3698);
nor U4184 (N_4184,N_3711,N_3712);
xnor U4185 (N_4185,N_3953,N_3795);
xor U4186 (N_4186,N_3537,N_3793);
or U4187 (N_4187,N_3533,N_3572);
and U4188 (N_4188,N_3720,N_3589);
and U4189 (N_4189,N_3901,N_3918);
xnor U4190 (N_4190,N_3503,N_3768);
or U4191 (N_4191,N_3895,N_3873);
or U4192 (N_4192,N_3969,N_3970);
xor U4193 (N_4193,N_3548,N_3534);
nand U4194 (N_4194,N_3623,N_3759);
or U4195 (N_4195,N_3861,N_3823);
nor U4196 (N_4196,N_3855,N_3800);
and U4197 (N_4197,N_3524,N_3927);
nand U4198 (N_4198,N_3723,N_3677);
or U4199 (N_4199,N_3613,N_3573);
nand U4200 (N_4200,N_3575,N_3883);
and U4201 (N_4201,N_3628,N_3667);
nor U4202 (N_4202,N_3598,N_3936);
and U4203 (N_4203,N_3603,N_3555);
and U4204 (N_4204,N_3718,N_3776);
xor U4205 (N_4205,N_3850,N_3569);
xor U4206 (N_4206,N_3594,N_3654);
and U4207 (N_4207,N_3699,N_3672);
and U4208 (N_4208,N_3708,N_3825);
nor U4209 (N_4209,N_3547,N_3990);
nand U4210 (N_4210,N_3726,N_3611);
nor U4211 (N_4211,N_3520,N_3612);
nor U4212 (N_4212,N_3848,N_3773);
xor U4213 (N_4213,N_3957,N_3771);
nand U4214 (N_4214,N_3992,N_3925);
xor U4215 (N_4215,N_3617,N_3958);
xor U4216 (N_4216,N_3630,N_3696);
nor U4217 (N_4217,N_3727,N_3510);
nor U4218 (N_4218,N_3645,N_3902);
nand U4219 (N_4219,N_3702,N_3653);
nand U4220 (N_4220,N_3658,N_3535);
or U4221 (N_4221,N_3872,N_3947);
or U4222 (N_4222,N_3607,N_3632);
xor U4223 (N_4223,N_3671,N_3592);
or U4224 (N_4224,N_3952,N_3774);
and U4225 (N_4225,N_3640,N_3557);
nand U4226 (N_4226,N_3735,N_3662);
nand U4227 (N_4227,N_3935,N_3910);
and U4228 (N_4228,N_3981,N_3987);
or U4229 (N_4229,N_3865,N_3887);
xor U4230 (N_4230,N_3857,N_3648);
or U4231 (N_4231,N_3737,N_3891);
nor U4232 (N_4232,N_3561,N_3529);
or U4233 (N_4233,N_3893,N_3618);
nand U4234 (N_4234,N_3867,N_3790);
or U4235 (N_4235,N_3885,N_3581);
or U4236 (N_4236,N_3647,N_3980);
nand U4237 (N_4237,N_3962,N_3810);
nand U4238 (N_4238,N_3666,N_3839);
or U4239 (N_4239,N_3619,N_3835);
nor U4240 (N_4240,N_3714,N_3626);
and U4241 (N_4241,N_3707,N_3900);
xnor U4242 (N_4242,N_3811,N_3747);
xnor U4243 (N_4243,N_3982,N_3597);
or U4244 (N_4244,N_3567,N_3513);
xnor U4245 (N_4245,N_3844,N_3847);
xnor U4246 (N_4246,N_3898,N_3851);
or U4247 (N_4247,N_3642,N_3854);
nand U4248 (N_4248,N_3506,N_3792);
and U4249 (N_4249,N_3977,N_3627);
xor U4250 (N_4250,N_3842,N_3810);
or U4251 (N_4251,N_3992,N_3577);
or U4252 (N_4252,N_3843,N_3813);
nand U4253 (N_4253,N_3961,N_3628);
nor U4254 (N_4254,N_3740,N_3930);
xnor U4255 (N_4255,N_3873,N_3721);
xnor U4256 (N_4256,N_3547,N_3899);
nor U4257 (N_4257,N_3981,N_3880);
or U4258 (N_4258,N_3925,N_3760);
xor U4259 (N_4259,N_3761,N_3585);
or U4260 (N_4260,N_3998,N_3528);
and U4261 (N_4261,N_3816,N_3844);
nand U4262 (N_4262,N_3679,N_3610);
nor U4263 (N_4263,N_3816,N_3726);
or U4264 (N_4264,N_3505,N_3590);
nand U4265 (N_4265,N_3799,N_3959);
or U4266 (N_4266,N_3991,N_3745);
and U4267 (N_4267,N_3798,N_3509);
or U4268 (N_4268,N_3792,N_3615);
and U4269 (N_4269,N_3681,N_3865);
nand U4270 (N_4270,N_3736,N_3975);
or U4271 (N_4271,N_3804,N_3932);
nand U4272 (N_4272,N_3502,N_3676);
and U4273 (N_4273,N_3522,N_3659);
and U4274 (N_4274,N_3631,N_3762);
nor U4275 (N_4275,N_3556,N_3516);
nand U4276 (N_4276,N_3883,N_3630);
xnor U4277 (N_4277,N_3843,N_3912);
nor U4278 (N_4278,N_3506,N_3984);
or U4279 (N_4279,N_3797,N_3538);
and U4280 (N_4280,N_3724,N_3665);
xor U4281 (N_4281,N_3597,N_3860);
or U4282 (N_4282,N_3789,N_3720);
or U4283 (N_4283,N_3919,N_3841);
nand U4284 (N_4284,N_3880,N_3536);
xor U4285 (N_4285,N_3724,N_3700);
nand U4286 (N_4286,N_3548,N_3522);
or U4287 (N_4287,N_3822,N_3800);
nor U4288 (N_4288,N_3817,N_3563);
nand U4289 (N_4289,N_3626,N_3624);
or U4290 (N_4290,N_3537,N_3822);
xnor U4291 (N_4291,N_3541,N_3943);
nand U4292 (N_4292,N_3726,N_3980);
xnor U4293 (N_4293,N_3863,N_3603);
and U4294 (N_4294,N_3548,N_3877);
xnor U4295 (N_4295,N_3994,N_3549);
and U4296 (N_4296,N_3820,N_3568);
or U4297 (N_4297,N_3853,N_3897);
nor U4298 (N_4298,N_3537,N_3788);
and U4299 (N_4299,N_3795,N_3938);
or U4300 (N_4300,N_3567,N_3969);
nor U4301 (N_4301,N_3909,N_3777);
and U4302 (N_4302,N_3732,N_3943);
xor U4303 (N_4303,N_3603,N_3675);
nor U4304 (N_4304,N_3923,N_3502);
xor U4305 (N_4305,N_3826,N_3931);
and U4306 (N_4306,N_3857,N_3891);
and U4307 (N_4307,N_3538,N_3537);
xnor U4308 (N_4308,N_3563,N_3581);
nor U4309 (N_4309,N_3738,N_3999);
and U4310 (N_4310,N_3523,N_3966);
and U4311 (N_4311,N_3864,N_3838);
nand U4312 (N_4312,N_3652,N_3750);
xnor U4313 (N_4313,N_3587,N_3562);
and U4314 (N_4314,N_3946,N_3696);
xor U4315 (N_4315,N_3967,N_3621);
xor U4316 (N_4316,N_3816,N_3802);
xnor U4317 (N_4317,N_3791,N_3609);
nand U4318 (N_4318,N_3575,N_3548);
nand U4319 (N_4319,N_3614,N_3907);
or U4320 (N_4320,N_3565,N_3786);
nor U4321 (N_4321,N_3972,N_3543);
nand U4322 (N_4322,N_3541,N_3584);
nand U4323 (N_4323,N_3818,N_3861);
xor U4324 (N_4324,N_3561,N_3891);
and U4325 (N_4325,N_3902,N_3724);
and U4326 (N_4326,N_3554,N_3667);
nor U4327 (N_4327,N_3637,N_3784);
or U4328 (N_4328,N_3610,N_3884);
and U4329 (N_4329,N_3928,N_3624);
xor U4330 (N_4330,N_3723,N_3542);
nand U4331 (N_4331,N_3585,N_3622);
nor U4332 (N_4332,N_3736,N_3632);
and U4333 (N_4333,N_3540,N_3679);
or U4334 (N_4334,N_3664,N_3740);
or U4335 (N_4335,N_3728,N_3664);
or U4336 (N_4336,N_3531,N_3501);
xor U4337 (N_4337,N_3975,N_3908);
nand U4338 (N_4338,N_3960,N_3728);
or U4339 (N_4339,N_3877,N_3520);
xor U4340 (N_4340,N_3646,N_3875);
nand U4341 (N_4341,N_3569,N_3869);
xnor U4342 (N_4342,N_3575,N_3634);
xor U4343 (N_4343,N_3677,N_3785);
or U4344 (N_4344,N_3508,N_3898);
or U4345 (N_4345,N_3522,N_3521);
xnor U4346 (N_4346,N_3787,N_3908);
nor U4347 (N_4347,N_3627,N_3819);
nand U4348 (N_4348,N_3817,N_3542);
nand U4349 (N_4349,N_3900,N_3774);
or U4350 (N_4350,N_3619,N_3695);
xnor U4351 (N_4351,N_3696,N_3787);
and U4352 (N_4352,N_3934,N_3779);
xnor U4353 (N_4353,N_3852,N_3943);
and U4354 (N_4354,N_3619,N_3601);
nor U4355 (N_4355,N_3512,N_3784);
xnor U4356 (N_4356,N_3938,N_3607);
and U4357 (N_4357,N_3542,N_3978);
nand U4358 (N_4358,N_3847,N_3828);
nor U4359 (N_4359,N_3779,N_3889);
and U4360 (N_4360,N_3646,N_3690);
xor U4361 (N_4361,N_3878,N_3890);
nand U4362 (N_4362,N_3797,N_3894);
nand U4363 (N_4363,N_3794,N_3610);
nand U4364 (N_4364,N_3808,N_3827);
and U4365 (N_4365,N_3962,N_3618);
xnor U4366 (N_4366,N_3968,N_3635);
or U4367 (N_4367,N_3712,N_3916);
or U4368 (N_4368,N_3908,N_3709);
and U4369 (N_4369,N_3808,N_3635);
and U4370 (N_4370,N_3765,N_3852);
nor U4371 (N_4371,N_3700,N_3637);
or U4372 (N_4372,N_3921,N_3894);
xor U4373 (N_4373,N_3752,N_3614);
nand U4374 (N_4374,N_3939,N_3815);
xnor U4375 (N_4375,N_3948,N_3998);
nor U4376 (N_4376,N_3632,N_3603);
or U4377 (N_4377,N_3797,N_3576);
and U4378 (N_4378,N_3667,N_3825);
nand U4379 (N_4379,N_3734,N_3608);
xnor U4380 (N_4380,N_3526,N_3600);
nor U4381 (N_4381,N_3763,N_3937);
xor U4382 (N_4382,N_3740,N_3586);
nand U4383 (N_4383,N_3829,N_3645);
xor U4384 (N_4384,N_3703,N_3787);
and U4385 (N_4385,N_3692,N_3755);
and U4386 (N_4386,N_3934,N_3970);
and U4387 (N_4387,N_3745,N_3761);
nor U4388 (N_4388,N_3978,N_3621);
xnor U4389 (N_4389,N_3776,N_3707);
xor U4390 (N_4390,N_3688,N_3718);
nand U4391 (N_4391,N_3526,N_3683);
and U4392 (N_4392,N_3888,N_3877);
nand U4393 (N_4393,N_3870,N_3616);
nand U4394 (N_4394,N_3856,N_3542);
nor U4395 (N_4395,N_3668,N_3656);
nor U4396 (N_4396,N_3733,N_3967);
or U4397 (N_4397,N_3546,N_3602);
nand U4398 (N_4398,N_3779,N_3663);
nand U4399 (N_4399,N_3893,N_3855);
xor U4400 (N_4400,N_3544,N_3833);
xnor U4401 (N_4401,N_3712,N_3702);
xor U4402 (N_4402,N_3959,N_3994);
or U4403 (N_4403,N_3792,N_3513);
xnor U4404 (N_4404,N_3947,N_3789);
and U4405 (N_4405,N_3745,N_3543);
or U4406 (N_4406,N_3981,N_3800);
nor U4407 (N_4407,N_3811,N_3973);
xnor U4408 (N_4408,N_3888,N_3807);
and U4409 (N_4409,N_3932,N_3859);
nor U4410 (N_4410,N_3571,N_3611);
nor U4411 (N_4411,N_3908,N_3649);
nand U4412 (N_4412,N_3701,N_3995);
or U4413 (N_4413,N_3905,N_3811);
and U4414 (N_4414,N_3620,N_3805);
xor U4415 (N_4415,N_3918,N_3894);
nand U4416 (N_4416,N_3868,N_3865);
nor U4417 (N_4417,N_3915,N_3928);
xor U4418 (N_4418,N_3664,N_3618);
or U4419 (N_4419,N_3927,N_3816);
xnor U4420 (N_4420,N_3600,N_3817);
nor U4421 (N_4421,N_3885,N_3703);
and U4422 (N_4422,N_3694,N_3690);
nand U4423 (N_4423,N_3718,N_3915);
and U4424 (N_4424,N_3977,N_3725);
nand U4425 (N_4425,N_3868,N_3606);
nand U4426 (N_4426,N_3580,N_3864);
nor U4427 (N_4427,N_3578,N_3586);
and U4428 (N_4428,N_3547,N_3562);
nor U4429 (N_4429,N_3780,N_3559);
or U4430 (N_4430,N_3987,N_3851);
nor U4431 (N_4431,N_3658,N_3778);
xor U4432 (N_4432,N_3774,N_3980);
and U4433 (N_4433,N_3971,N_3673);
and U4434 (N_4434,N_3764,N_3865);
and U4435 (N_4435,N_3786,N_3793);
nand U4436 (N_4436,N_3844,N_3671);
nor U4437 (N_4437,N_3641,N_3758);
xor U4438 (N_4438,N_3608,N_3538);
nor U4439 (N_4439,N_3761,N_3868);
nor U4440 (N_4440,N_3917,N_3984);
nor U4441 (N_4441,N_3882,N_3815);
and U4442 (N_4442,N_3756,N_3734);
xor U4443 (N_4443,N_3755,N_3592);
or U4444 (N_4444,N_3865,N_3971);
and U4445 (N_4445,N_3743,N_3574);
nand U4446 (N_4446,N_3501,N_3639);
nand U4447 (N_4447,N_3851,N_3610);
or U4448 (N_4448,N_3841,N_3715);
nor U4449 (N_4449,N_3693,N_3656);
xor U4450 (N_4450,N_3811,N_3603);
and U4451 (N_4451,N_3680,N_3755);
and U4452 (N_4452,N_3754,N_3694);
nand U4453 (N_4453,N_3578,N_3679);
and U4454 (N_4454,N_3893,N_3820);
xnor U4455 (N_4455,N_3915,N_3688);
or U4456 (N_4456,N_3599,N_3745);
nand U4457 (N_4457,N_3887,N_3584);
xnor U4458 (N_4458,N_3973,N_3657);
xnor U4459 (N_4459,N_3783,N_3811);
nor U4460 (N_4460,N_3646,N_3818);
nand U4461 (N_4461,N_3874,N_3621);
nand U4462 (N_4462,N_3937,N_3932);
nand U4463 (N_4463,N_3787,N_3865);
xor U4464 (N_4464,N_3771,N_3657);
xor U4465 (N_4465,N_3854,N_3954);
nor U4466 (N_4466,N_3502,N_3876);
or U4467 (N_4467,N_3584,N_3952);
and U4468 (N_4468,N_3592,N_3902);
nand U4469 (N_4469,N_3728,N_3864);
nor U4470 (N_4470,N_3805,N_3974);
xor U4471 (N_4471,N_3516,N_3655);
nand U4472 (N_4472,N_3895,N_3991);
and U4473 (N_4473,N_3926,N_3572);
xnor U4474 (N_4474,N_3764,N_3879);
xnor U4475 (N_4475,N_3534,N_3862);
nor U4476 (N_4476,N_3643,N_3925);
xor U4477 (N_4477,N_3639,N_3631);
nor U4478 (N_4478,N_3597,N_3813);
nand U4479 (N_4479,N_3611,N_3517);
xnor U4480 (N_4480,N_3808,N_3559);
xnor U4481 (N_4481,N_3893,N_3697);
or U4482 (N_4482,N_3709,N_3912);
xnor U4483 (N_4483,N_3778,N_3808);
nor U4484 (N_4484,N_3987,N_3782);
nand U4485 (N_4485,N_3821,N_3522);
xor U4486 (N_4486,N_3684,N_3697);
nor U4487 (N_4487,N_3822,N_3644);
nand U4488 (N_4488,N_3924,N_3884);
nand U4489 (N_4489,N_3724,N_3752);
or U4490 (N_4490,N_3971,N_3939);
nor U4491 (N_4491,N_3839,N_3809);
or U4492 (N_4492,N_3892,N_3981);
or U4493 (N_4493,N_3754,N_3580);
nor U4494 (N_4494,N_3537,N_3646);
nor U4495 (N_4495,N_3993,N_3904);
or U4496 (N_4496,N_3742,N_3749);
and U4497 (N_4497,N_3878,N_3824);
and U4498 (N_4498,N_3701,N_3622);
xnor U4499 (N_4499,N_3706,N_3749);
and U4500 (N_4500,N_4135,N_4285);
nor U4501 (N_4501,N_4361,N_4388);
and U4502 (N_4502,N_4342,N_4360);
and U4503 (N_4503,N_4468,N_4432);
nand U4504 (N_4504,N_4470,N_4258);
nor U4505 (N_4505,N_4460,N_4349);
nand U4506 (N_4506,N_4306,N_4448);
nor U4507 (N_4507,N_4020,N_4050);
nor U4508 (N_4508,N_4359,N_4469);
nor U4509 (N_4509,N_4440,N_4387);
and U4510 (N_4510,N_4352,N_4145);
or U4511 (N_4511,N_4398,N_4243);
xnor U4512 (N_4512,N_4056,N_4236);
nor U4513 (N_4513,N_4175,N_4066);
or U4514 (N_4514,N_4199,N_4430);
and U4515 (N_4515,N_4491,N_4231);
nor U4516 (N_4516,N_4402,N_4362);
xnor U4517 (N_4517,N_4194,N_4278);
or U4518 (N_4518,N_4429,N_4416);
or U4519 (N_4519,N_4094,N_4311);
or U4520 (N_4520,N_4249,N_4302);
nor U4521 (N_4521,N_4414,N_4033);
and U4522 (N_4522,N_4325,N_4040);
nand U4523 (N_4523,N_4304,N_4444);
xnor U4524 (N_4524,N_4275,N_4161);
nand U4525 (N_4525,N_4277,N_4484);
nand U4526 (N_4526,N_4413,N_4452);
xor U4527 (N_4527,N_4228,N_4259);
or U4528 (N_4528,N_4169,N_4167);
or U4529 (N_4529,N_4417,N_4380);
xnor U4530 (N_4530,N_4187,N_4477);
and U4531 (N_4531,N_4442,N_4262);
nor U4532 (N_4532,N_4492,N_4490);
xnor U4533 (N_4533,N_4334,N_4282);
nand U4534 (N_4534,N_4412,N_4377);
and U4535 (N_4535,N_4127,N_4105);
or U4536 (N_4536,N_4441,N_4292);
xor U4537 (N_4537,N_4357,N_4439);
xnor U4538 (N_4538,N_4345,N_4177);
nor U4539 (N_4539,N_4181,N_4091);
nor U4540 (N_4540,N_4021,N_4158);
nor U4541 (N_4541,N_4042,N_4088);
and U4542 (N_4542,N_4084,N_4198);
nor U4543 (N_4543,N_4039,N_4001);
or U4544 (N_4544,N_4497,N_4443);
xor U4545 (N_4545,N_4202,N_4142);
nand U4546 (N_4546,N_4384,N_4205);
or U4547 (N_4547,N_4261,N_4293);
or U4548 (N_4548,N_4059,N_4230);
and U4549 (N_4549,N_4272,N_4340);
and U4550 (N_4550,N_4227,N_4101);
and U4551 (N_4551,N_4346,N_4068);
xor U4552 (N_4552,N_4025,N_4263);
and U4553 (N_4553,N_4485,N_4086);
and U4554 (N_4554,N_4465,N_4240);
nor U4555 (N_4555,N_4095,N_4499);
nand U4556 (N_4556,N_4211,N_4179);
xor U4557 (N_4557,N_4218,N_4012);
or U4558 (N_4558,N_4244,N_4295);
nand U4559 (N_4559,N_4073,N_4449);
nor U4560 (N_4560,N_4341,N_4270);
and U4561 (N_4561,N_4148,N_4036);
and U4562 (N_4562,N_4496,N_4234);
xnor U4563 (N_4563,N_4216,N_4106);
xor U4564 (N_4564,N_4407,N_4140);
nor U4565 (N_4565,N_4297,N_4048);
nor U4566 (N_4566,N_4172,N_4269);
and U4567 (N_4567,N_4393,N_4152);
or U4568 (N_4568,N_4321,N_4260);
xor U4569 (N_4569,N_4305,N_4403);
and U4570 (N_4570,N_4112,N_4283);
nand U4571 (N_4571,N_4118,N_4296);
nand U4572 (N_4572,N_4327,N_4072);
nor U4573 (N_4573,N_4410,N_4002);
xnor U4574 (N_4574,N_4298,N_4107);
xor U4575 (N_4575,N_4222,N_4008);
nand U4576 (N_4576,N_4022,N_4239);
xor U4577 (N_4577,N_4146,N_4397);
and U4578 (N_4578,N_4336,N_4281);
or U4579 (N_4579,N_4354,N_4369);
or U4580 (N_4580,N_4482,N_4134);
and U4581 (N_4581,N_4189,N_4015);
nand U4582 (N_4582,N_4424,N_4071);
and U4583 (N_4583,N_4375,N_4013);
or U4584 (N_4584,N_4195,N_4157);
nor U4585 (N_4585,N_4391,N_4217);
and U4586 (N_4586,N_4274,N_4489);
xor U4587 (N_4587,N_4248,N_4338);
nand U4588 (N_4588,N_4447,N_4303);
nor U4589 (N_4589,N_4209,N_4326);
or U4590 (N_4590,N_4390,N_4166);
nand U4591 (N_4591,N_4097,N_4320);
nor U4592 (N_4592,N_4486,N_4203);
nor U4593 (N_4593,N_4319,N_4017);
or U4594 (N_4594,N_4079,N_4007);
or U4595 (N_4595,N_4365,N_4103);
or U4596 (N_4596,N_4294,N_4456);
xor U4597 (N_4597,N_4016,N_4450);
and U4598 (N_4598,N_4138,N_4253);
and U4599 (N_4599,N_4433,N_4206);
or U4600 (N_4600,N_4437,N_4459);
or U4601 (N_4601,N_4406,N_4241);
nor U4602 (N_4602,N_4180,N_4356);
nand U4603 (N_4603,N_4351,N_4368);
or U4604 (N_4604,N_4032,N_4207);
and U4605 (N_4605,N_4358,N_4291);
nand U4606 (N_4606,N_4472,N_4220);
or U4607 (N_4607,N_4264,N_4348);
nor U4608 (N_4608,N_4215,N_4266);
nor U4609 (N_4609,N_4196,N_4041);
nand U4610 (N_4610,N_4401,N_4102);
xnor U4611 (N_4611,N_4493,N_4367);
or U4612 (N_4612,N_4461,N_4399);
nand U4613 (N_4613,N_4045,N_4344);
xnor U4614 (N_4614,N_4419,N_4164);
xor U4615 (N_4615,N_4256,N_4431);
nor U4616 (N_4616,N_4333,N_4197);
nor U4617 (N_4617,N_4004,N_4251);
or U4618 (N_4618,N_4034,N_4474);
nor U4619 (N_4619,N_4287,N_4463);
and U4620 (N_4620,N_4223,N_4063);
or U4621 (N_4621,N_4471,N_4064);
xnor U4622 (N_4622,N_4159,N_4254);
nor U4623 (N_4623,N_4347,N_4316);
nand U4624 (N_4624,N_4090,N_4109);
xor U4625 (N_4625,N_4343,N_4317);
or U4626 (N_4626,N_4149,N_4422);
nand U4627 (N_4627,N_4435,N_4370);
or U4628 (N_4628,N_4130,N_4323);
nor U4629 (N_4629,N_4427,N_4183);
or U4630 (N_4630,N_4372,N_4160);
xor U4631 (N_4631,N_4268,N_4481);
nand U4632 (N_4632,N_4114,N_4003);
and U4633 (N_4633,N_4237,N_4191);
or U4634 (N_4634,N_4132,N_4210);
xnor U4635 (N_4635,N_4280,N_4185);
xor U4636 (N_4636,N_4353,N_4495);
nand U4637 (N_4637,N_4136,N_4462);
or U4638 (N_4638,N_4364,N_4383);
nand U4639 (N_4639,N_4310,N_4480);
xnor U4640 (N_4640,N_4080,N_4190);
or U4641 (N_4641,N_4168,N_4252);
nand U4642 (N_4642,N_4005,N_4156);
xor U4643 (N_4643,N_4178,N_4043);
and U4644 (N_4644,N_4478,N_4286);
and U4645 (N_4645,N_4395,N_4426);
nor U4646 (N_4646,N_4479,N_4379);
and U4647 (N_4647,N_4255,N_4250);
xor U4648 (N_4648,N_4028,N_4133);
nor U4649 (N_4649,N_4014,N_4494);
or U4650 (N_4650,N_4301,N_4279);
nand U4651 (N_4651,N_4246,N_4212);
xor U4652 (N_4652,N_4300,N_4137);
or U4653 (N_4653,N_4330,N_4221);
and U4654 (N_4654,N_4093,N_4290);
nand U4655 (N_4655,N_4049,N_4058);
xnor U4656 (N_4656,N_4044,N_4061);
nand U4657 (N_4657,N_4089,N_4163);
or U4658 (N_4658,N_4047,N_4242);
or U4659 (N_4659,N_4081,N_4055);
and U4660 (N_4660,N_4193,N_4052);
nand U4661 (N_4661,N_4077,N_4308);
nor U4662 (N_4662,N_4315,N_4087);
or U4663 (N_4663,N_4322,N_4229);
nand U4664 (N_4664,N_4313,N_4184);
nand U4665 (N_4665,N_4420,N_4129);
xnor U4666 (N_4666,N_4085,N_4092);
and U4667 (N_4667,N_4117,N_4035);
and U4668 (N_4668,N_4010,N_4144);
nor U4669 (N_4669,N_4385,N_4476);
nand U4670 (N_4670,N_4267,N_4192);
nor U4671 (N_4671,N_4464,N_4067);
nand U4672 (N_4672,N_4386,N_4428);
or U4673 (N_4673,N_4075,N_4488);
xnor U4674 (N_4674,N_4188,N_4309);
nor U4675 (N_4675,N_4404,N_4155);
xor U4676 (N_4676,N_4143,N_4366);
and U4677 (N_4677,N_4423,N_4128);
nand U4678 (N_4678,N_4312,N_4247);
nand U4679 (N_4679,N_4186,N_4408);
and U4680 (N_4680,N_4100,N_4139);
nor U4681 (N_4681,N_4200,N_4062);
nand U4682 (N_4682,N_4418,N_4376);
xnor U4683 (N_4683,N_4070,N_4078);
or U4684 (N_4684,N_4031,N_4154);
xnor U4685 (N_4685,N_4284,N_4389);
and U4686 (N_4686,N_4457,N_4337);
xnor U4687 (N_4687,N_4265,N_4053);
nor U4688 (N_4688,N_4467,N_4453);
nand U4689 (N_4689,N_4069,N_4475);
xor U4690 (N_4690,N_4276,N_4057);
and U4691 (N_4691,N_4454,N_4458);
nand U4692 (N_4692,N_4498,N_4288);
nor U4693 (N_4693,N_4037,N_4483);
nor U4694 (N_4694,N_4332,N_4065);
nand U4695 (N_4695,N_4124,N_4394);
nor U4696 (N_4696,N_4214,N_4434);
or U4697 (N_4697,N_4331,N_4208);
and U4698 (N_4698,N_4108,N_4026);
or U4699 (N_4699,N_4224,N_4436);
or U4700 (N_4700,N_4019,N_4099);
nor U4701 (N_4701,N_4307,N_4378);
or U4702 (N_4702,N_4382,N_4355);
xnor U4703 (N_4703,N_4150,N_4176);
nand U4704 (N_4704,N_4335,N_4174);
nand U4705 (N_4705,N_4451,N_4018);
or U4706 (N_4706,N_4121,N_4038);
nor U4707 (N_4707,N_4235,N_4473);
xnor U4708 (N_4708,N_4120,N_4411);
nand U4709 (N_4709,N_4400,N_4363);
xor U4710 (N_4710,N_4030,N_4487);
nor U4711 (N_4711,N_4415,N_4225);
nor U4712 (N_4712,N_4153,N_4373);
xor U4713 (N_4713,N_4060,N_4374);
and U4714 (N_4714,N_4076,N_4054);
and U4715 (N_4715,N_4409,N_4233);
nand U4716 (N_4716,N_4219,N_4111);
nor U4717 (N_4717,N_4392,N_4238);
xor U4718 (N_4718,N_4029,N_4011);
nor U4719 (N_4719,N_4289,N_4381);
and U4720 (N_4720,N_4455,N_4350);
nor U4721 (N_4721,N_4110,N_4271);
nand U4722 (N_4722,N_4204,N_4115);
or U4723 (N_4723,N_4147,N_4083);
or U4724 (N_4724,N_4466,N_4098);
and U4725 (N_4725,N_4104,N_4445);
xnor U4726 (N_4726,N_4141,N_4329);
nor U4727 (N_4727,N_4116,N_4182);
xnor U4728 (N_4728,N_4405,N_4339);
nor U4729 (N_4729,N_4328,N_4046);
and U4730 (N_4730,N_4299,N_4226);
nor U4731 (N_4731,N_4396,N_4123);
and U4732 (N_4732,N_4113,N_4446);
nor U4733 (N_4733,N_4082,N_4170);
and U4734 (N_4734,N_4213,N_4324);
nand U4735 (N_4735,N_4126,N_4151);
or U4736 (N_4736,N_4257,N_4000);
or U4737 (N_4737,N_4027,N_4122);
nor U4738 (N_4738,N_4051,N_4162);
xnor U4739 (N_4739,N_4096,N_4074);
or U4740 (N_4740,N_4245,N_4438);
or U4741 (N_4741,N_4201,N_4131);
xnor U4742 (N_4742,N_4165,N_4009);
and U4743 (N_4743,N_4425,N_4273);
xor U4744 (N_4744,N_4421,N_4371);
and U4745 (N_4745,N_4023,N_4171);
nand U4746 (N_4746,N_4318,N_4173);
xor U4747 (N_4747,N_4125,N_4314);
xor U4748 (N_4748,N_4119,N_4006);
or U4749 (N_4749,N_4232,N_4024);
or U4750 (N_4750,N_4032,N_4235);
xor U4751 (N_4751,N_4479,N_4110);
xor U4752 (N_4752,N_4385,N_4224);
nor U4753 (N_4753,N_4295,N_4171);
and U4754 (N_4754,N_4276,N_4419);
nor U4755 (N_4755,N_4096,N_4387);
nor U4756 (N_4756,N_4416,N_4495);
or U4757 (N_4757,N_4434,N_4160);
or U4758 (N_4758,N_4275,N_4064);
nand U4759 (N_4759,N_4097,N_4266);
and U4760 (N_4760,N_4042,N_4258);
xnor U4761 (N_4761,N_4297,N_4306);
nor U4762 (N_4762,N_4166,N_4090);
or U4763 (N_4763,N_4070,N_4286);
or U4764 (N_4764,N_4333,N_4379);
and U4765 (N_4765,N_4235,N_4096);
xor U4766 (N_4766,N_4185,N_4465);
nand U4767 (N_4767,N_4121,N_4005);
and U4768 (N_4768,N_4458,N_4065);
xnor U4769 (N_4769,N_4458,N_4267);
nor U4770 (N_4770,N_4306,N_4345);
nor U4771 (N_4771,N_4250,N_4423);
nor U4772 (N_4772,N_4200,N_4360);
xor U4773 (N_4773,N_4032,N_4344);
and U4774 (N_4774,N_4193,N_4493);
and U4775 (N_4775,N_4284,N_4062);
xor U4776 (N_4776,N_4143,N_4378);
nor U4777 (N_4777,N_4033,N_4093);
xnor U4778 (N_4778,N_4362,N_4412);
nand U4779 (N_4779,N_4035,N_4059);
and U4780 (N_4780,N_4326,N_4216);
or U4781 (N_4781,N_4250,N_4102);
xnor U4782 (N_4782,N_4315,N_4272);
nor U4783 (N_4783,N_4004,N_4169);
nor U4784 (N_4784,N_4306,N_4299);
nor U4785 (N_4785,N_4268,N_4204);
nor U4786 (N_4786,N_4079,N_4251);
and U4787 (N_4787,N_4034,N_4299);
xnor U4788 (N_4788,N_4001,N_4215);
and U4789 (N_4789,N_4161,N_4023);
xnor U4790 (N_4790,N_4179,N_4334);
xnor U4791 (N_4791,N_4169,N_4218);
or U4792 (N_4792,N_4239,N_4469);
xor U4793 (N_4793,N_4438,N_4347);
or U4794 (N_4794,N_4036,N_4301);
and U4795 (N_4795,N_4307,N_4182);
and U4796 (N_4796,N_4077,N_4285);
and U4797 (N_4797,N_4020,N_4279);
nor U4798 (N_4798,N_4263,N_4058);
xnor U4799 (N_4799,N_4147,N_4041);
or U4800 (N_4800,N_4404,N_4330);
or U4801 (N_4801,N_4367,N_4351);
or U4802 (N_4802,N_4455,N_4289);
nor U4803 (N_4803,N_4455,N_4277);
xnor U4804 (N_4804,N_4422,N_4482);
xnor U4805 (N_4805,N_4089,N_4023);
or U4806 (N_4806,N_4431,N_4162);
nor U4807 (N_4807,N_4086,N_4132);
xnor U4808 (N_4808,N_4229,N_4112);
or U4809 (N_4809,N_4326,N_4158);
and U4810 (N_4810,N_4445,N_4100);
nand U4811 (N_4811,N_4221,N_4463);
or U4812 (N_4812,N_4049,N_4234);
and U4813 (N_4813,N_4312,N_4206);
or U4814 (N_4814,N_4490,N_4194);
or U4815 (N_4815,N_4496,N_4488);
and U4816 (N_4816,N_4194,N_4485);
xor U4817 (N_4817,N_4154,N_4321);
xor U4818 (N_4818,N_4361,N_4382);
or U4819 (N_4819,N_4234,N_4382);
or U4820 (N_4820,N_4097,N_4110);
nor U4821 (N_4821,N_4188,N_4290);
or U4822 (N_4822,N_4412,N_4099);
nand U4823 (N_4823,N_4360,N_4408);
nor U4824 (N_4824,N_4193,N_4341);
nor U4825 (N_4825,N_4471,N_4101);
nand U4826 (N_4826,N_4425,N_4185);
and U4827 (N_4827,N_4300,N_4167);
xnor U4828 (N_4828,N_4131,N_4262);
or U4829 (N_4829,N_4067,N_4368);
or U4830 (N_4830,N_4148,N_4089);
nor U4831 (N_4831,N_4035,N_4160);
or U4832 (N_4832,N_4378,N_4473);
and U4833 (N_4833,N_4349,N_4050);
nand U4834 (N_4834,N_4263,N_4323);
nand U4835 (N_4835,N_4301,N_4168);
nor U4836 (N_4836,N_4119,N_4045);
nor U4837 (N_4837,N_4237,N_4124);
and U4838 (N_4838,N_4417,N_4309);
and U4839 (N_4839,N_4154,N_4186);
xnor U4840 (N_4840,N_4000,N_4326);
or U4841 (N_4841,N_4128,N_4411);
and U4842 (N_4842,N_4041,N_4234);
nor U4843 (N_4843,N_4466,N_4219);
xor U4844 (N_4844,N_4339,N_4440);
nor U4845 (N_4845,N_4372,N_4214);
nand U4846 (N_4846,N_4341,N_4004);
and U4847 (N_4847,N_4483,N_4077);
or U4848 (N_4848,N_4388,N_4269);
or U4849 (N_4849,N_4425,N_4261);
and U4850 (N_4850,N_4470,N_4133);
nor U4851 (N_4851,N_4436,N_4160);
or U4852 (N_4852,N_4252,N_4454);
xor U4853 (N_4853,N_4298,N_4087);
nor U4854 (N_4854,N_4477,N_4341);
and U4855 (N_4855,N_4426,N_4085);
and U4856 (N_4856,N_4207,N_4474);
or U4857 (N_4857,N_4485,N_4397);
and U4858 (N_4858,N_4452,N_4065);
xor U4859 (N_4859,N_4322,N_4301);
nor U4860 (N_4860,N_4445,N_4474);
nand U4861 (N_4861,N_4366,N_4363);
xnor U4862 (N_4862,N_4103,N_4106);
or U4863 (N_4863,N_4055,N_4477);
and U4864 (N_4864,N_4409,N_4206);
and U4865 (N_4865,N_4412,N_4342);
xnor U4866 (N_4866,N_4381,N_4386);
or U4867 (N_4867,N_4394,N_4011);
xnor U4868 (N_4868,N_4455,N_4326);
nor U4869 (N_4869,N_4156,N_4033);
and U4870 (N_4870,N_4106,N_4449);
xor U4871 (N_4871,N_4188,N_4232);
nand U4872 (N_4872,N_4055,N_4436);
xor U4873 (N_4873,N_4025,N_4417);
or U4874 (N_4874,N_4251,N_4378);
nor U4875 (N_4875,N_4182,N_4478);
and U4876 (N_4876,N_4046,N_4225);
and U4877 (N_4877,N_4202,N_4133);
or U4878 (N_4878,N_4297,N_4332);
or U4879 (N_4879,N_4173,N_4004);
and U4880 (N_4880,N_4121,N_4447);
nor U4881 (N_4881,N_4302,N_4319);
nand U4882 (N_4882,N_4385,N_4275);
xor U4883 (N_4883,N_4225,N_4371);
and U4884 (N_4884,N_4108,N_4082);
nor U4885 (N_4885,N_4157,N_4355);
xnor U4886 (N_4886,N_4334,N_4443);
or U4887 (N_4887,N_4059,N_4076);
nor U4888 (N_4888,N_4282,N_4125);
nand U4889 (N_4889,N_4245,N_4369);
or U4890 (N_4890,N_4164,N_4268);
and U4891 (N_4891,N_4471,N_4202);
nand U4892 (N_4892,N_4055,N_4137);
xor U4893 (N_4893,N_4396,N_4227);
or U4894 (N_4894,N_4353,N_4169);
nand U4895 (N_4895,N_4325,N_4138);
nand U4896 (N_4896,N_4078,N_4277);
xnor U4897 (N_4897,N_4099,N_4158);
nand U4898 (N_4898,N_4498,N_4454);
and U4899 (N_4899,N_4127,N_4473);
or U4900 (N_4900,N_4220,N_4099);
xnor U4901 (N_4901,N_4170,N_4151);
nor U4902 (N_4902,N_4148,N_4340);
nand U4903 (N_4903,N_4325,N_4341);
nor U4904 (N_4904,N_4425,N_4281);
nor U4905 (N_4905,N_4302,N_4445);
or U4906 (N_4906,N_4076,N_4237);
or U4907 (N_4907,N_4066,N_4019);
or U4908 (N_4908,N_4454,N_4017);
nand U4909 (N_4909,N_4460,N_4031);
and U4910 (N_4910,N_4165,N_4149);
and U4911 (N_4911,N_4462,N_4315);
nor U4912 (N_4912,N_4375,N_4450);
nor U4913 (N_4913,N_4428,N_4321);
xnor U4914 (N_4914,N_4375,N_4444);
nor U4915 (N_4915,N_4045,N_4312);
or U4916 (N_4916,N_4096,N_4320);
or U4917 (N_4917,N_4003,N_4411);
nor U4918 (N_4918,N_4096,N_4134);
or U4919 (N_4919,N_4280,N_4129);
or U4920 (N_4920,N_4166,N_4267);
nand U4921 (N_4921,N_4296,N_4043);
nor U4922 (N_4922,N_4388,N_4025);
nand U4923 (N_4923,N_4402,N_4476);
and U4924 (N_4924,N_4428,N_4245);
and U4925 (N_4925,N_4103,N_4141);
nand U4926 (N_4926,N_4112,N_4012);
xor U4927 (N_4927,N_4496,N_4463);
and U4928 (N_4928,N_4476,N_4434);
or U4929 (N_4929,N_4487,N_4397);
xor U4930 (N_4930,N_4425,N_4196);
xor U4931 (N_4931,N_4218,N_4398);
nor U4932 (N_4932,N_4040,N_4012);
nand U4933 (N_4933,N_4348,N_4265);
and U4934 (N_4934,N_4011,N_4079);
nor U4935 (N_4935,N_4332,N_4416);
xnor U4936 (N_4936,N_4436,N_4263);
xnor U4937 (N_4937,N_4178,N_4284);
and U4938 (N_4938,N_4002,N_4185);
and U4939 (N_4939,N_4261,N_4018);
and U4940 (N_4940,N_4025,N_4446);
and U4941 (N_4941,N_4141,N_4231);
and U4942 (N_4942,N_4260,N_4488);
nand U4943 (N_4943,N_4094,N_4445);
or U4944 (N_4944,N_4164,N_4155);
nand U4945 (N_4945,N_4014,N_4351);
xnor U4946 (N_4946,N_4430,N_4338);
or U4947 (N_4947,N_4425,N_4122);
nand U4948 (N_4948,N_4060,N_4083);
and U4949 (N_4949,N_4094,N_4081);
xnor U4950 (N_4950,N_4201,N_4164);
xor U4951 (N_4951,N_4247,N_4100);
xor U4952 (N_4952,N_4469,N_4299);
nor U4953 (N_4953,N_4087,N_4192);
or U4954 (N_4954,N_4435,N_4394);
xnor U4955 (N_4955,N_4059,N_4345);
nand U4956 (N_4956,N_4152,N_4274);
and U4957 (N_4957,N_4130,N_4271);
nand U4958 (N_4958,N_4270,N_4373);
nand U4959 (N_4959,N_4252,N_4143);
xor U4960 (N_4960,N_4354,N_4173);
xnor U4961 (N_4961,N_4477,N_4282);
xnor U4962 (N_4962,N_4454,N_4079);
or U4963 (N_4963,N_4462,N_4014);
xor U4964 (N_4964,N_4198,N_4301);
nor U4965 (N_4965,N_4421,N_4416);
nand U4966 (N_4966,N_4346,N_4120);
nor U4967 (N_4967,N_4275,N_4162);
or U4968 (N_4968,N_4161,N_4056);
xor U4969 (N_4969,N_4460,N_4227);
or U4970 (N_4970,N_4308,N_4391);
nand U4971 (N_4971,N_4298,N_4247);
and U4972 (N_4972,N_4462,N_4472);
xor U4973 (N_4973,N_4449,N_4212);
or U4974 (N_4974,N_4282,N_4031);
and U4975 (N_4975,N_4476,N_4140);
xor U4976 (N_4976,N_4365,N_4176);
or U4977 (N_4977,N_4043,N_4308);
or U4978 (N_4978,N_4282,N_4295);
nand U4979 (N_4979,N_4171,N_4183);
and U4980 (N_4980,N_4400,N_4145);
nor U4981 (N_4981,N_4195,N_4200);
nand U4982 (N_4982,N_4468,N_4461);
nor U4983 (N_4983,N_4096,N_4284);
and U4984 (N_4984,N_4129,N_4454);
nor U4985 (N_4985,N_4407,N_4436);
xnor U4986 (N_4986,N_4406,N_4288);
nand U4987 (N_4987,N_4050,N_4298);
nor U4988 (N_4988,N_4269,N_4412);
nand U4989 (N_4989,N_4391,N_4300);
and U4990 (N_4990,N_4330,N_4271);
nand U4991 (N_4991,N_4229,N_4436);
nand U4992 (N_4992,N_4264,N_4116);
nand U4993 (N_4993,N_4252,N_4056);
xnor U4994 (N_4994,N_4322,N_4015);
nand U4995 (N_4995,N_4338,N_4014);
and U4996 (N_4996,N_4367,N_4119);
or U4997 (N_4997,N_4009,N_4408);
nor U4998 (N_4998,N_4369,N_4319);
and U4999 (N_4999,N_4306,N_4244);
xor U5000 (N_5000,N_4609,N_4707);
nor U5001 (N_5001,N_4839,N_4690);
xnor U5002 (N_5002,N_4850,N_4944);
nor U5003 (N_5003,N_4894,N_4951);
nand U5004 (N_5004,N_4519,N_4513);
and U5005 (N_5005,N_4774,N_4835);
nor U5006 (N_5006,N_4514,N_4813);
xnor U5007 (N_5007,N_4714,N_4970);
or U5008 (N_5008,N_4916,N_4784);
nor U5009 (N_5009,N_4711,N_4565);
nor U5010 (N_5010,N_4875,N_4673);
and U5011 (N_5011,N_4636,N_4789);
xnor U5012 (N_5012,N_4740,N_4718);
nand U5013 (N_5013,N_4820,N_4729);
and U5014 (N_5014,N_4666,N_4543);
nand U5015 (N_5015,N_4917,N_4960);
and U5016 (N_5016,N_4770,N_4624);
and U5017 (N_5017,N_4931,N_4908);
and U5018 (N_5018,N_4903,N_4566);
xor U5019 (N_5019,N_4956,N_4606);
nor U5020 (N_5020,N_4777,N_4874);
or U5021 (N_5021,N_4795,N_4897);
nand U5022 (N_5022,N_4744,N_4504);
nor U5023 (N_5023,N_4571,N_4989);
and U5024 (N_5024,N_4832,N_4676);
or U5025 (N_5025,N_4709,N_4845);
or U5026 (N_5026,N_4937,N_4564);
xor U5027 (N_5027,N_4940,N_4807);
or U5028 (N_5028,N_4708,N_4867);
and U5029 (N_5029,N_4806,N_4568);
nand U5030 (N_5030,N_4500,N_4539);
nand U5031 (N_5031,N_4846,N_4618);
and U5032 (N_5032,N_4720,N_4596);
and U5033 (N_5033,N_4507,N_4642);
nand U5034 (N_5034,N_4523,N_4857);
nor U5035 (N_5035,N_4927,N_4930);
nand U5036 (N_5036,N_4630,N_4688);
or U5037 (N_5037,N_4621,N_4724);
xnor U5038 (N_5038,N_4805,N_4809);
or U5039 (N_5039,N_4595,N_4751);
nand U5040 (N_5040,N_4728,N_4785);
xor U5041 (N_5041,N_4652,N_4992);
nand U5042 (N_5042,N_4984,N_4852);
nor U5043 (N_5043,N_4985,N_4858);
nor U5044 (N_5044,N_4623,N_4753);
nand U5045 (N_5045,N_4815,N_4684);
xnor U5046 (N_5046,N_4675,N_4547);
and U5047 (N_5047,N_4581,N_4589);
and U5048 (N_5048,N_4727,N_4996);
nor U5049 (N_5049,N_4518,N_4665);
nor U5050 (N_5050,N_4671,N_4638);
nor U5051 (N_5051,N_4554,N_4509);
nor U5052 (N_5052,N_4735,N_4861);
and U5053 (N_5053,N_4731,N_4631);
xnor U5054 (N_5054,N_4923,N_4537);
nor U5055 (N_5055,N_4948,N_4963);
nand U5056 (N_5056,N_4526,N_4814);
nor U5057 (N_5057,N_4669,N_4981);
and U5058 (N_5058,N_4515,N_4936);
or U5059 (N_5059,N_4767,N_4559);
and U5060 (N_5060,N_4869,N_4639);
and U5061 (N_5061,N_4921,N_4644);
nor U5062 (N_5062,N_4502,N_4549);
nand U5063 (N_5063,N_4569,N_4841);
xnor U5064 (N_5064,N_4578,N_4531);
or U5065 (N_5065,N_4836,N_4590);
xor U5066 (N_5066,N_4763,N_4953);
nor U5067 (N_5067,N_4612,N_4692);
nand U5068 (N_5068,N_4683,N_4743);
or U5069 (N_5069,N_4752,N_4717);
nor U5070 (N_5070,N_4762,N_4732);
nor U5071 (N_5071,N_4971,N_4754);
nand U5072 (N_5072,N_4677,N_4958);
or U5073 (N_5073,N_4594,N_4660);
xnor U5074 (N_5074,N_4983,N_4540);
nand U5075 (N_5075,N_4713,N_4508);
nand U5076 (N_5076,N_4640,N_4796);
xnor U5077 (N_5077,N_4959,N_4831);
and U5078 (N_5078,N_4964,N_4776);
or U5079 (N_5079,N_4653,N_4616);
nor U5080 (N_5080,N_4705,N_4878);
xnor U5081 (N_5081,N_4524,N_4693);
nor U5082 (N_5082,N_4561,N_4965);
nor U5083 (N_5083,N_4755,N_4912);
nand U5084 (N_5084,N_4888,N_4901);
nand U5085 (N_5085,N_4579,N_4804);
or U5086 (N_5086,N_4607,N_4911);
and U5087 (N_5087,N_4574,N_4702);
or U5088 (N_5088,N_4925,N_4935);
xor U5089 (N_5089,N_4674,N_4800);
xor U5090 (N_5090,N_4918,N_4773);
and U5091 (N_5091,N_4748,N_4881);
nor U5092 (N_5092,N_4745,N_4979);
nand U5093 (N_5093,N_4641,N_4906);
nand U5094 (N_5094,N_4952,N_4860);
or U5095 (N_5095,N_4961,N_4527);
nor U5096 (N_5096,N_4704,N_4847);
and U5097 (N_5097,N_4764,N_4957);
or U5098 (N_5098,N_4866,N_4900);
nor U5099 (N_5099,N_4876,N_4859);
nor U5100 (N_5100,N_4601,N_4975);
nor U5101 (N_5101,N_4591,N_4721);
xnor U5102 (N_5102,N_4782,N_4628);
and U5103 (N_5103,N_4863,N_4864);
xnor U5104 (N_5104,N_4670,N_4598);
and U5105 (N_5105,N_4833,N_4822);
nand U5106 (N_5106,N_4871,N_4988);
or U5107 (N_5107,N_4781,N_4608);
or U5108 (N_5108,N_4637,N_4620);
nand U5109 (N_5109,N_4698,N_4715);
and U5110 (N_5110,N_4824,N_4538);
nand U5111 (N_5111,N_4757,N_4525);
nand U5112 (N_5112,N_4768,N_4560);
nand U5113 (N_5113,N_4534,N_4694);
and U5114 (N_5114,N_4946,N_4703);
xnor U5115 (N_5115,N_4950,N_4928);
xnor U5116 (N_5116,N_4577,N_4759);
nor U5117 (N_5117,N_4633,N_4741);
or U5118 (N_5118,N_4627,N_4974);
nand U5119 (N_5119,N_4765,N_4837);
and U5120 (N_5120,N_4778,N_4879);
and U5121 (N_5121,N_4862,N_4873);
and U5122 (N_5122,N_4650,N_4766);
and U5123 (N_5123,N_4798,N_4772);
or U5124 (N_5124,N_4583,N_4934);
or U5125 (N_5125,N_4919,N_4615);
nand U5126 (N_5126,N_4885,N_4746);
nand U5127 (N_5127,N_4629,N_4649);
nor U5128 (N_5128,N_4887,N_4883);
or U5129 (N_5129,N_4730,N_4659);
nand U5130 (N_5130,N_4699,N_4818);
nand U5131 (N_5131,N_4853,N_4501);
and U5132 (N_5132,N_4736,N_4611);
nor U5133 (N_5133,N_4510,N_4987);
xnor U5134 (N_5134,N_4605,N_4910);
xnor U5135 (N_5135,N_4613,N_4647);
nor U5136 (N_5136,N_4710,N_4546);
nand U5137 (N_5137,N_4749,N_4733);
and U5138 (N_5138,N_4760,N_4695);
or U5139 (N_5139,N_4954,N_4780);
and U5140 (N_5140,N_4821,N_4791);
and U5141 (N_5141,N_4582,N_4542);
nor U5142 (N_5142,N_4976,N_4816);
and U5143 (N_5143,N_4891,N_4779);
and U5144 (N_5144,N_4899,N_4902);
nand U5145 (N_5145,N_4962,N_4812);
or U5146 (N_5146,N_4856,N_4758);
or U5147 (N_5147,N_4977,N_4726);
or U5148 (N_5148,N_4828,N_4572);
nor U5149 (N_5149,N_4563,N_4663);
and U5150 (N_5150,N_4716,N_4994);
or U5151 (N_5151,N_4843,N_4972);
xor U5152 (N_5152,N_4680,N_4679);
nand U5153 (N_5153,N_4775,N_4553);
or U5154 (N_5154,N_4520,N_4756);
xor U5155 (N_5155,N_4686,N_4827);
and U5156 (N_5156,N_4998,N_4512);
and U5157 (N_5157,N_4980,N_4622);
and U5158 (N_5158,N_4678,N_4750);
xor U5159 (N_5159,N_4942,N_4747);
xnor U5160 (N_5160,N_4943,N_4761);
nor U5161 (N_5161,N_4592,N_4528);
or U5162 (N_5162,N_4913,N_4722);
or U5163 (N_5163,N_4969,N_4632);
xor U5164 (N_5164,N_4895,N_4511);
nor U5165 (N_5165,N_4551,N_4562);
and U5166 (N_5166,N_4924,N_4570);
and U5167 (N_5167,N_4602,N_4681);
nor U5168 (N_5168,N_4982,N_4575);
xor U5169 (N_5169,N_4790,N_4898);
xor U5170 (N_5170,N_4799,N_4604);
or U5171 (N_5171,N_4588,N_4738);
or U5172 (N_5172,N_4771,N_4868);
nand U5173 (N_5173,N_4643,N_4792);
nand U5174 (N_5174,N_4522,N_4685);
nor U5175 (N_5175,N_4848,N_4955);
nand U5176 (N_5176,N_4658,N_4548);
or U5177 (N_5177,N_4558,N_4610);
xor U5178 (N_5178,N_4997,N_4990);
nor U5179 (N_5179,N_4645,N_4646);
and U5180 (N_5180,N_4825,N_4600);
nand U5181 (N_5181,N_4668,N_4712);
xnor U5182 (N_5182,N_4801,N_4929);
and U5183 (N_5183,N_4597,N_4995);
or U5184 (N_5184,N_4783,N_4978);
xor U5185 (N_5185,N_4909,N_4719);
nor U5186 (N_5186,N_4786,N_4840);
or U5187 (N_5187,N_4947,N_4967);
and U5188 (N_5188,N_4614,N_4915);
nor U5189 (N_5189,N_4672,N_4593);
nor U5190 (N_5190,N_4541,N_4886);
nand U5191 (N_5191,N_4986,N_4580);
and U5192 (N_5192,N_4793,N_4905);
or U5193 (N_5193,N_4661,N_4877);
or U5194 (N_5194,N_4973,N_4505);
nand U5195 (N_5195,N_4892,N_4794);
xnor U5196 (N_5196,N_4872,N_4657);
nor U5197 (N_5197,N_4844,N_4556);
xor U5198 (N_5198,N_4890,N_4889);
xnor U5199 (N_5199,N_4904,N_4576);
or U5200 (N_5200,N_4907,N_4634);
nor U5201 (N_5201,N_4654,N_4966);
xor U5202 (N_5202,N_4584,N_4701);
or U5203 (N_5203,N_4855,N_4819);
nand U5204 (N_5204,N_4769,N_4922);
nor U5205 (N_5205,N_4920,N_4991);
nand U5206 (N_5206,N_4626,N_4817);
xor U5207 (N_5207,N_4550,N_4968);
nor U5208 (N_5208,N_4896,N_4842);
nor U5209 (N_5209,N_4557,N_4586);
and U5210 (N_5210,N_4545,N_4737);
xor U5211 (N_5211,N_4742,N_4797);
or U5212 (N_5212,N_4585,N_4939);
or U5213 (N_5213,N_4503,N_4734);
nor U5214 (N_5214,N_4849,N_4826);
nor U5215 (N_5215,N_4723,N_4725);
xor U5216 (N_5216,N_4893,N_4926);
nand U5217 (N_5217,N_4999,N_4697);
or U5218 (N_5218,N_4656,N_4803);
nor U5219 (N_5219,N_4625,N_4506);
and U5220 (N_5220,N_4619,N_4808);
xor U5221 (N_5221,N_4664,N_4532);
or U5222 (N_5222,N_4882,N_4830);
nand U5223 (N_5223,N_4938,N_4706);
nor U5224 (N_5224,N_4536,N_4567);
xor U5225 (N_5225,N_4838,N_4802);
or U5226 (N_5226,N_4635,N_4949);
nand U5227 (N_5227,N_4599,N_4914);
nor U5228 (N_5228,N_4823,N_4667);
and U5229 (N_5229,N_4811,N_4648);
nand U5230 (N_5230,N_4993,N_4662);
and U5231 (N_5231,N_4517,N_4555);
and U5232 (N_5232,N_4535,N_4603);
or U5233 (N_5233,N_4941,N_4854);
xnor U5234 (N_5234,N_4530,N_4552);
nor U5235 (N_5235,N_4700,N_4682);
and U5236 (N_5236,N_4691,N_4651);
nor U5237 (N_5237,N_4945,N_4529);
or U5238 (N_5238,N_4788,N_4787);
nand U5239 (N_5239,N_4587,N_4573);
nand U5240 (N_5240,N_4617,N_4829);
nand U5241 (N_5241,N_4933,N_4655);
xnor U5242 (N_5242,N_4932,N_4689);
xor U5243 (N_5243,N_4880,N_4516);
xnor U5244 (N_5244,N_4544,N_4870);
nand U5245 (N_5245,N_4884,N_4521);
xor U5246 (N_5246,N_4687,N_4533);
xor U5247 (N_5247,N_4739,N_4696);
and U5248 (N_5248,N_4851,N_4865);
nand U5249 (N_5249,N_4810,N_4834);
nand U5250 (N_5250,N_4903,N_4668);
nand U5251 (N_5251,N_4694,N_4922);
nand U5252 (N_5252,N_4941,N_4887);
nand U5253 (N_5253,N_4782,N_4633);
nand U5254 (N_5254,N_4911,N_4805);
and U5255 (N_5255,N_4508,N_4591);
nand U5256 (N_5256,N_4718,N_4926);
nand U5257 (N_5257,N_4877,N_4680);
nor U5258 (N_5258,N_4622,N_4656);
nand U5259 (N_5259,N_4668,N_4792);
and U5260 (N_5260,N_4810,N_4524);
or U5261 (N_5261,N_4993,N_4881);
and U5262 (N_5262,N_4536,N_4629);
nand U5263 (N_5263,N_4807,N_4903);
xor U5264 (N_5264,N_4610,N_4704);
nor U5265 (N_5265,N_4546,N_4871);
xor U5266 (N_5266,N_4919,N_4519);
xnor U5267 (N_5267,N_4598,N_4982);
or U5268 (N_5268,N_4730,N_4614);
nand U5269 (N_5269,N_4927,N_4639);
nor U5270 (N_5270,N_4946,N_4989);
xnor U5271 (N_5271,N_4841,N_4968);
nor U5272 (N_5272,N_4511,N_4846);
or U5273 (N_5273,N_4910,N_4768);
or U5274 (N_5274,N_4694,N_4614);
nand U5275 (N_5275,N_4617,N_4722);
nor U5276 (N_5276,N_4891,N_4940);
or U5277 (N_5277,N_4896,N_4853);
nor U5278 (N_5278,N_4713,N_4532);
or U5279 (N_5279,N_4658,N_4868);
nand U5280 (N_5280,N_4671,N_4995);
nand U5281 (N_5281,N_4824,N_4634);
and U5282 (N_5282,N_4933,N_4954);
nor U5283 (N_5283,N_4692,N_4958);
and U5284 (N_5284,N_4603,N_4924);
nor U5285 (N_5285,N_4594,N_4996);
xnor U5286 (N_5286,N_4673,N_4547);
or U5287 (N_5287,N_4565,N_4999);
nand U5288 (N_5288,N_4761,N_4590);
xor U5289 (N_5289,N_4831,N_4943);
nand U5290 (N_5290,N_4816,N_4940);
nand U5291 (N_5291,N_4820,N_4700);
nand U5292 (N_5292,N_4525,N_4586);
or U5293 (N_5293,N_4905,N_4671);
and U5294 (N_5294,N_4526,N_4797);
nand U5295 (N_5295,N_4956,N_4968);
nor U5296 (N_5296,N_4603,N_4750);
nand U5297 (N_5297,N_4751,N_4764);
nand U5298 (N_5298,N_4506,N_4646);
and U5299 (N_5299,N_4847,N_4900);
or U5300 (N_5300,N_4877,N_4879);
nor U5301 (N_5301,N_4532,N_4650);
xnor U5302 (N_5302,N_4666,N_4778);
xor U5303 (N_5303,N_4636,N_4765);
or U5304 (N_5304,N_4946,N_4824);
nand U5305 (N_5305,N_4727,N_4772);
xor U5306 (N_5306,N_4728,N_4902);
xor U5307 (N_5307,N_4584,N_4560);
nor U5308 (N_5308,N_4869,N_4803);
xnor U5309 (N_5309,N_4646,N_4538);
xor U5310 (N_5310,N_4738,N_4772);
and U5311 (N_5311,N_4977,N_4815);
nand U5312 (N_5312,N_4906,N_4575);
xor U5313 (N_5313,N_4666,N_4824);
xor U5314 (N_5314,N_4562,N_4590);
xnor U5315 (N_5315,N_4773,N_4663);
or U5316 (N_5316,N_4679,N_4829);
or U5317 (N_5317,N_4558,N_4611);
nand U5318 (N_5318,N_4612,N_4823);
nand U5319 (N_5319,N_4948,N_4524);
nor U5320 (N_5320,N_4884,N_4722);
nor U5321 (N_5321,N_4626,N_4747);
nand U5322 (N_5322,N_4570,N_4976);
nand U5323 (N_5323,N_4980,N_4516);
nor U5324 (N_5324,N_4932,N_4853);
and U5325 (N_5325,N_4723,N_4785);
xnor U5326 (N_5326,N_4597,N_4556);
nand U5327 (N_5327,N_4993,N_4847);
and U5328 (N_5328,N_4565,N_4988);
xnor U5329 (N_5329,N_4704,N_4977);
or U5330 (N_5330,N_4795,N_4934);
nand U5331 (N_5331,N_4702,N_4648);
nor U5332 (N_5332,N_4818,N_4633);
xor U5333 (N_5333,N_4731,N_4873);
xnor U5334 (N_5334,N_4768,N_4944);
nand U5335 (N_5335,N_4886,N_4949);
or U5336 (N_5336,N_4538,N_4942);
and U5337 (N_5337,N_4909,N_4537);
nor U5338 (N_5338,N_4910,N_4871);
xor U5339 (N_5339,N_4685,N_4589);
nor U5340 (N_5340,N_4642,N_4544);
or U5341 (N_5341,N_4853,N_4636);
nor U5342 (N_5342,N_4810,N_4531);
xor U5343 (N_5343,N_4898,N_4674);
and U5344 (N_5344,N_4864,N_4838);
or U5345 (N_5345,N_4982,N_4835);
or U5346 (N_5346,N_4815,N_4818);
nor U5347 (N_5347,N_4595,N_4787);
nor U5348 (N_5348,N_4806,N_4874);
or U5349 (N_5349,N_4768,N_4958);
nand U5350 (N_5350,N_4549,N_4607);
nor U5351 (N_5351,N_4788,N_4585);
or U5352 (N_5352,N_4688,N_4563);
nand U5353 (N_5353,N_4844,N_4933);
nand U5354 (N_5354,N_4881,N_4779);
nor U5355 (N_5355,N_4508,N_4604);
and U5356 (N_5356,N_4870,N_4706);
nor U5357 (N_5357,N_4942,N_4874);
and U5358 (N_5358,N_4716,N_4878);
nor U5359 (N_5359,N_4969,N_4667);
nand U5360 (N_5360,N_4892,N_4844);
xnor U5361 (N_5361,N_4749,N_4948);
and U5362 (N_5362,N_4949,N_4851);
or U5363 (N_5363,N_4502,N_4991);
and U5364 (N_5364,N_4670,N_4519);
and U5365 (N_5365,N_4748,N_4986);
nor U5366 (N_5366,N_4801,N_4770);
nor U5367 (N_5367,N_4959,N_4981);
nand U5368 (N_5368,N_4866,N_4938);
nor U5369 (N_5369,N_4897,N_4919);
nor U5370 (N_5370,N_4755,N_4651);
or U5371 (N_5371,N_4604,N_4692);
and U5372 (N_5372,N_4991,N_4603);
nor U5373 (N_5373,N_4639,N_4805);
xnor U5374 (N_5374,N_4621,N_4646);
nor U5375 (N_5375,N_4945,N_4543);
or U5376 (N_5376,N_4942,N_4813);
and U5377 (N_5377,N_4762,N_4967);
nand U5378 (N_5378,N_4701,N_4734);
and U5379 (N_5379,N_4747,N_4896);
nor U5380 (N_5380,N_4759,N_4562);
nand U5381 (N_5381,N_4682,N_4880);
xnor U5382 (N_5382,N_4512,N_4857);
nand U5383 (N_5383,N_4967,N_4567);
xnor U5384 (N_5384,N_4613,N_4588);
nor U5385 (N_5385,N_4756,N_4996);
or U5386 (N_5386,N_4529,N_4783);
xnor U5387 (N_5387,N_4573,N_4836);
xor U5388 (N_5388,N_4980,N_4775);
nor U5389 (N_5389,N_4601,N_4537);
nor U5390 (N_5390,N_4630,N_4534);
nor U5391 (N_5391,N_4930,N_4680);
or U5392 (N_5392,N_4535,N_4801);
nor U5393 (N_5393,N_4689,N_4772);
nor U5394 (N_5394,N_4513,N_4670);
nand U5395 (N_5395,N_4524,N_4847);
and U5396 (N_5396,N_4802,N_4577);
or U5397 (N_5397,N_4782,N_4947);
nand U5398 (N_5398,N_4732,N_4741);
nor U5399 (N_5399,N_4763,N_4813);
xor U5400 (N_5400,N_4807,N_4649);
nor U5401 (N_5401,N_4824,N_4749);
nor U5402 (N_5402,N_4883,N_4684);
and U5403 (N_5403,N_4647,N_4745);
and U5404 (N_5404,N_4543,N_4727);
xor U5405 (N_5405,N_4971,N_4515);
nor U5406 (N_5406,N_4918,N_4700);
or U5407 (N_5407,N_4553,N_4923);
nor U5408 (N_5408,N_4824,N_4516);
xor U5409 (N_5409,N_4822,N_4841);
nor U5410 (N_5410,N_4951,N_4785);
nor U5411 (N_5411,N_4925,N_4554);
xor U5412 (N_5412,N_4571,N_4795);
xor U5413 (N_5413,N_4969,N_4581);
nand U5414 (N_5414,N_4847,N_4971);
and U5415 (N_5415,N_4908,N_4779);
or U5416 (N_5416,N_4897,N_4780);
nor U5417 (N_5417,N_4694,N_4569);
nor U5418 (N_5418,N_4711,N_4569);
nor U5419 (N_5419,N_4519,N_4683);
xnor U5420 (N_5420,N_4811,N_4649);
nand U5421 (N_5421,N_4574,N_4971);
nand U5422 (N_5422,N_4568,N_4559);
nand U5423 (N_5423,N_4718,N_4603);
and U5424 (N_5424,N_4705,N_4620);
nor U5425 (N_5425,N_4979,N_4811);
or U5426 (N_5426,N_4745,N_4732);
nor U5427 (N_5427,N_4826,N_4998);
nor U5428 (N_5428,N_4979,N_4616);
xnor U5429 (N_5429,N_4696,N_4996);
nand U5430 (N_5430,N_4984,N_4859);
nor U5431 (N_5431,N_4968,N_4792);
and U5432 (N_5432,N_4678,N_4680);
nor U5433 (N_5433,N_4624,N_4839);
nor U5434 (N_5434,N_4839,N_4859);
nand U5435 (N_5435,N_4964,N_4719);
xnor U5436 (N_5436,N_4539,N_4771);
xor U5437 (N_5437,N_4868,N_4949);
nand U5438 (N_5438,N_4550,N_4903);
nand U5439 (N_5439,N_4647,N_4616);
or U5440 (N_5440,N_4660,N_4541);
xnor U5441 (N_5441,N_4945,N_4670);
nor U5442 (N_5442,N_4700,N_4644);
xnor U5443 (N_5443,N_4690,N_4937);
xnor U5444 (N_5444,N_4925,N_4719);
and U5445 (N_5445,N_4877,N_4671);
nand U5446 (N_5446,N_4637,N_4611);
xnor U5447 (N_5447,N_4609,N_4555);
or U5448 (N_5448,N_4984,N_4960);
or U5449 (N_5449,N_4608,N_4670);
xnor U5450 (N_5450,N_4926,N_4928);
and U5451 (N_5451,N_4922,N_4868);
xnor U5452 (N_5452,N_4545,N_4987);
nor U5453 (N_5453,N_4780,N_4977);
nand U5454 (N_5454,N_4731,N_4521);
or U5455 (N_5455,N_4809,N_4699);
nand U5456 (N_5456,N_4713,N_4859);
nand U5457 (N_5457,N_4509,N_4922);
or U5458 (N_5458,N_4784,N_4631);
and U5459 (N_5459,N_4856,N_4785);
nand U5460 (N_5460,N_4754,N_4810);
xnor U5461 (N_5461,N_4523,N_4624);
and U5462 (N_5462,N_4532,N_4810);
and U5463 (N_5463,N_4648,N_4587);
nor U5464 (N_5464,N_4548,N_4999);
nand U5465 (N_5465,N_4540,N_4750);
and U5466 (N_5466,N_4611,N_4983);
and U5467 (N_5467,N_4636,N_4656);
xor U5468 (N_5468,N_4605,N_4522);
xor U5469 (N_5469,N_4697,N_4982);
or U5470 (N_5470,N_4530,N_4976);
nor U5471 (N_5471,N_4590,N_4641);
and U5472 (N_5472,N_4682,N_4503);
nor U5473 (N_5473,N_4886,N_4866);
nand U5474 (N_5474,N_4573,N_4618);
or U5475 (N_5475,N_4860,N_4871);
xor U5476 (N_5476,N_4641,N_4873);
and U5477 (N_5477,N_4986,N_4645);
or U5478 (N_5478,N_4793,N_4966);
and U5479 (N_5479,N_4546,N_4941);
and U5480 (N_5480,N_4808,N_4937);
nor U5481 (N_5481,N_4824,N_4761);
nand U5482 (N_5482,N_4529,N_4992);
or U5483 (N_5483,N_4695,N_4723);
and U5484 (N_5484,N_4671,N_4826);
and U5485 (N_5485,N_4783,N_4627);
xor U5486 (N_5486,N_4740,N_4562);
nor U5487 (N_5487,N_4515,N_4622);
and U5488 (N_5488,N_4884,N_4547);
nand U5489 (N_5489,N_4897,N_4762);
nand U5490 (N_5490,N_4978,N_4708);
and U5491 (N_5491,N_4532,N_4949);
nand U5492 (N_5492,N_4642,N_4775);
nand U5493 (N_5493,N_4940,N_4990);
xor U5494 (N_5494,N_4943,N_4848);
xnor U5495 (N_5495,N_4807,N_4708);
nor U5496 (N_5496,N_4753,N_4814);
nor U5497 (N_5497,N_4521,N_4970);
nand U5498 (N_5498,N_4634,N_4729);
or U5499 (N_5499,N_4525,N_4661);
and U5500 (N_5500,N_5465,N_5041);
and U5501 (N_5501,N_5298,N_5056);
nor U5502 (N_5502,N_5384,N_5281);
or U5503 (N_5503,N_5233,N_5129);
nor U5504 (N_5504,N_5499,N_5314);
nor U5505 (N_5505,N_5348,N_5291);
nand U5506 (N_5506,N_5393,N_5242);
nor U5507 (N_5507,N_5138,N_5166);
nand U5508 (N_5508,N_5328,N_5402);
nand U5509 (N_5509,N_5164,N_5349);
nor U5510 (N_5510,N_5480,N_5126);
nand U5511 (N_5511,N_5079,N_5034);
xnor U5512 (N_5512,N_5165,N_5052);
or U5513 (N_5513,N_5346,N_5046);
and U5514 (N_5514,N_5142,N_5150);
xor U5515 (N_5515,N_5243,N_5236);
or U5516 (N_5516,N_5359,N_5389);
or U5517 (N_5517,N_5305,N_5204);
or U5518 (N_5518,N_5321,N_5273);
nand U5519 (N_5519,N_5221,N_5313);
xor U5520 (N_5520,N_5344,N_5326);
nor U5521 (N_5521,N_5331,N_5479);
and U5522 (N_5522,N_5064,N_5379);
nand U5523 (N_5523,N_5247,N_5350);
nand U5524 (N_5524,N_5159,N_5018);
and U5525 (N_5525,N_5148,N_5325);
or U5526 (N_5526,N_5154,N_5469);
nor U5527 (N_5527,N_5397,N_5157);
and U5528 (N_5528,N_5054,N_5032);
xnor U5529 (N_5529,N_5297,N_5187);
xor U5530 (N_5530,N_5422,N_5059);
or U5531 (N_5531,N_5391,N_5078);
nor U5532 (N_5532,N_5370,N_5076);
xnor U5533 (N_5533,N_5374,N_5180);
or U5534 (N_5534,N_5049,N_5169);
xnor U5535 (N_5535,N_5474,N_5105);
nand U5536 (N_5536,N_5423,N_5051);
and U5537 (N_5537,N_5140,N_5039);
xnor U5538 (N_5538,N_5323,N_5063);
nand U5539 (N_5539,N_5453,N_5436);
nand U5540 (N_5540,N_5010,N_5275);
or U5541 (N_5541,N_5403,N_5152);
nor U5542 (N_5542,N_5109,N_5451);
or U5543 (N_5543,N_5200,N_5489);
nor U5544 (N_5544,N_5383,N_5256);
or U5545 (N_5545,N_5335,N_5048);
or U5546 (N_5546,N_5405,N_5123);
or U5547 (N_5547,N_5173,N_5044);
and U5548 (N_5548,N_5011,N_5211);
and U5549 (N_5549,N_5171,N_5360);
nand U5550 (N_5550,N_5246,N_5031);
xor U5551 (N_5551,N_5339,N_5382);
and U5552 (N_5552,N_5446,N_5108);
xnor U5553 (N_5553,N_5407,N_5410);
nand U5554 (N_5554,N_5124,N_5083);
or U5555 (N_5555,N_5425,N_5160);
nor U5556 (N_5556,N_5186,N_5133);
nand U5557 (N_5557,N_5250,N_5197);
nor U5558 (N_5558,N_5327,N_5177);
nor U5559 (N_5559,N_5312,N_5294);
or U5560 (N_5560,N_5145,N_5342);
xor U5561 (N_5561,N_5361,N_5132);
and U5562 (N_5562,N_5122,N_5372);
and U5563 (N_5563,N_5225,N_5182);
nand U5564 (N_5564,N_5332,N_5042);
and U5565 (N_5565,N_5222,N_5110);
nor U5566 (N_5566,N_5174,N_5306);
nor U5567 (N_5567,N_5213,N_5475);
xnor U5568 (N_5568,N_5387,N_5006);
xnor U5569 (N_5569,N_5458,N_5426);
or U5570 (N_5570,N_5002,N_5189);
or U5571 (N_5571,N_5094,N_5424);
or U5572 (N_5572,N_5070,N_5366);
nand U5573 (N_5573,N_5215,N_5288);
nor U5574 (N_5574,N_5185,N_5438);
nor U5575 (N_5575,N_5230,N_5477);
nand U5576 (N_5576,N_5459,N_5014);
xnor U5577 (N_5577,N_5362,N_5483);
or U5578 (N_5578,N_5434,N_5183);
or U5579 (N_5579,N_5053,N_5428);
nor U5580 (N_5580,N_5228,N_5271);
nor U5581 (N_5581,N_5111,N_5482);
nor U5582 (N_5582,N_5058,N_5263);
nand U5583 (N_5583,N_5322,N_5115);
or U5584 (N_5584,N_5069,N_5158);
and U5585 (N_5585,N_5091,N_5395);
and U5586 (N_5586,N_5319,N_5285);
nor U5587 (N_5587,N_5343,N_5151);
xor U5588 (N_5588,N_5130,N_5341);
nand U5589 (N_5589,N_5210,N_5352);
and U5590 (N_5590,N_5258,N_5062);
and U5591 (N_5591,N_5196,N_5466);
and U5592 (N_5592,N_5369,N_5264);
and U5593 (N_5593,N_5439,N_5303);
xnor U5594 (N_5594,N_5337,N_5102);
nand U5595 (N_5595,N_5179,N_5199);
nor U5596 (N_5596,N_5068,N_5038);
or U5597 (N_5597,N_5050,N_5205);
xor U5598 (N_5598,N_5260,N_5286);
xnor U5599 (N_5599,N_5030,N_5016);
xor U5600 (N_5600,N_5401,N_5497);
and U5601 (N_5601,N_5252,N_5367);
and U5602 (N_5602,N_5121,N_5498);
nand U5603 (N_5603,N_5376,N_5420);
nand U5604 (N_5604,N_5487,N_5476);
and U5605 (N_5605,N_5363,N_5447);
xor U5606 (N_5606,N_5441,N_5461);
nand U5607 (N_5607,N_5101,N_5089);
and U5608 (N_5608,N_5100,N_5357);
and U5609 (N_5609,N_5047,N_5355);
nand U5610 (N_5610,N_5134,N_5368);
or U5611 (N_5611,N_5188,N_5184);
or U5612 (N_5612,N_5096,N_5345);
nor U5613 (N_5613,N_5333,N_5464);
or U5614 (N_5614,N_5104,N_5000);
and U5615 (N_5615,N_5320,N_5287);
xnor U5616 (N_5616,N_5201,N_5119);
nand U5617 (N_5617,N_5156,N_5280);
nor U5618 (N_5618,N_5057,N_5040);
nand U5619 (N_5619,N_5061,N_5442);
or U5620 (N_5620,N_5206,N_5232);
nor U5621 (N_5621,N_5013,N_5025);
xnor U5622 (N_5622,N_5417,N_5304);
or U5623 (N_5623,N_5347,N_5136);
nor U5624 (N_5624,N_5409,N_5399);
nand U5625 (N_5625,N_5444,N_5473);
nand U5626 (N_5626,N_5467,N_5373);
nand U5627 (N_5627,N_5127,N_5279);
and U5628 (N_5628,N_5147,N_5429);
xor U5629 (N_5629,N_5270,N_5463);
and U5630 (N_5630,N_5027,N_5455);
or U5631 (N_5631,N_5494,N_5231);
nand U5632 (N_5632,N_5162,N_5435);
or U5633 (N_5633,N_5026,N_5440);
nand U5634 (N_5634,N_5009,N_5324);
or U5635 (N_5635,N_5135,N_5392);
nand U5636 (N_5636,N_5308,N_5021);
and U5637 (N_5637,N_5309,N_5385);
xor U5638 (N_5638,N_5194,N_5012);
and U5639 (N_5639,N_5364,N_5244);
xnor U5640 (N_5640,N_5255,N_5223);
nand U5641 (N_5641,N_5261,N_5282);
nor U5642 (N_5642,N_5125,N_5388);
nor U5643 (N_5643,N_5290,N_5353);
and U5644 (N_5644,N_5300,N_5212);
and U5645 (N_5645,N_5356,N_5492);
xor U5646 (N_5646,N_5266,N_5045);
nor U5647 (N_5647,N_5024,N_5433);
nand U5648 (N_5648,N_5419,N_5413);
xor U5649 (N_5649,N_5106,N_5099);
nand U5650 (N_5650,N_5262,N_5155);
nor U5651 (N_5651,N_5216,N_5118);
and U5652 (N_5652,N_5239,N_5296);
xnor U5653 (N_5653,N_5253,N_5354);
or U5654 (N_5654,N_5168,N_5098);
or U5655 (N_5655,N_5128,N_5175);
or U5656 (N_5656,N_5408,N_5495);
nand U5657 (N_5657,N_5249,N_5329);
nand U5658 (N_5658,N_5033,N_5386);
and U5659 (N_5659,N_5017,N_5077);
or U5660 (N_5660,N_5161,N_5085);
or U5661 (N_5661,N_5195,N_5295);
nand U5662 (N_5662,N_5431,N_5176);
xnor U5663 (N_5663,N_5153,N_5112);
and U5664 (N_5664,N_5421,N_5146);
nor U5665 (N_5665,N_5193,N_5336);
nor U5666 (N_5666,N_5198,N_5245);
and U5667 (N_5667,N_5457,N_5005);
or U5668 (N_5668,N_5143,N_5224);
or U5669 (N_5669,N_5137,N_5003);
nor U5670 (N_5670,N_5449,N_5358);
or U5671 (N_5671,N_5090,N_5283);
or U5672 (N_5672,N_5229,N_5317);
nor U5673 (N_5673,N_5276,N_5235);
nand U5674 (N_5674,N_5073,N_5008);
xor U5675 (N_5675,N_5277,N_5214);
and U5676 (N_5676,N_5496,N_5103);
or U5677 (N_5677,N_5470,N_5398);
and U5678 (N_5678,N_5170,N_5227);
and U5679 (N_5679,N_5084,N_5378);
nor U5680 (N_5680,N_5238,N_5330);
nor U5681 (N_5681,N_5037,N_5390);
nor U5682 (N_5682,N_5074,N_5114);
nor U5683 (N_5683,N_5415,N_5484);
nand U5684 (N_5684,N_5460,N_5412);
or U5685 (N_5685,N_5203,N_5338);
and U5686 (N_5686,N_5116,N_5293);
nand U5687 (N_5687,N_5097,N_5268);
or U5688 (N_5688,N_5377,N_5269);
and U5689 (N_5689,N_5452,N_5490);
or U5690 (N_5690,N_5471,N_5139);
and U5691 (N_5691,N_5141,N_5481);
nor U5692 (N_5692,N_5302,N_5080);
xnor U5693 (N_5693,N_5207,N_5240);
or U5694 (N_5694,N_5088,N_5043);
or U5695 (N_5695,N_5394,N_5416);
and U5696 (N_5696,N_5448,N_5491);
nand U5697 (N_5697,N_5066,N_5334);
nor U5698 (N_5698,N_5248,N_5172);
nand U5699 (N_5699,N_5117,N_5086);
xor U5700 (N_5700,N_5120,N_5144);
and U5701 (N_5701,N_5015,N_5251);
nand U5702 (N_5702,N_5167,N_5226);
nand U5703 (N_5703,N_5237,N_5486);
xnor U5704 (N_5704,N_5055,N_5404);
nor U5705 (N_5705,N_5178,N_5208);
and U5706 (N_5706,N_5082,N_5406);
nor U5707 (N_5707,N_5488,N_5340);
xnor U5708 (N_5708,N_5414,N_5190);
and U5709 (N_5709,N_5004,N_5093);
or U5710 (N_5710,N_5272,N_5241);
xor U5711 (N_5711,N_5278,N_5450);
and U5712 (N_5712,N_5075,N_5478);
nor U5713 (N_5713,N_5071,N_5462);
xor U5714 (N_5714,N_5060,N_5219);
or U5715 (N_5715,N_5072,N_5191);
nor U5716 (N_5716,N_5380,N_5259);
nand U5717 (N_5717,N_5456,N_5351);
and U5718 (N_5718,N_5289,N_5485);
nor U5719 (N_5719,N_5468,N_5022);
and U5720 (N_5720,N_5472,N_5218);
or U5721 (N_5721,N_5029,N_5437);
xnor U5722 (N_5722,N_5131,N_5181);
xor U5723 (N_5723,N_5149,N_5375);
nand U5724 (N_5724,N_5254,N_5371);
or U5725 (N_5725,N_5315,N_5365);
xor U5726 (N_5726,N_5007,N_5310);
xor U5727 (N_5727,N_5316,N_5234);
nand U5728 (N_5728,N_5311,N_5209);
nand U5729 (N_5729,N_5163,N_5019);
xor U5730 (N_5730,N_5411,N_5020);
or U5731 (N_5731,N_5023,N_5081);
nor U5732 (N_5732,N_5318,N_5454);
or U5733 (N_5733,N_5493,N_5092);
xnor U5734 (N_5734,N_5001,N_5432);
nor U5735 (N_5735,N_5265,N_5267);
nor U5736 (N_5736,N_5427,N_5107);
nand U5737 (N_5737,N_5220,N_5396);
or U5738 (N_5738,N_5257,N_5400);
and U5739 (N_5739,N_5430,N_5445);
nor U5740 (N_5740,N_5381,N_5095);
and U5741 (N_5741,N_5307,N_5028);
xnor U5742 (N_5742,N_5202,N_5065);
nor U5743 (N_5743,N_5299,N_5443);
xor U5744 (N_5744,N_5274,N_5036);
or U5745 (N_5745,N_5292,N_5301);
nand U5746 (N_5746,N_5418,N_5087);
or U5747 (N_5747,N_5192,N_5217);
nand U5748 (N_5748,N_5113,N_5067);
nand U5749 (N_5749,N_5035,N_5284);
and U5750 (N_5750,N_5318,N_5366);
or U5751 (N_5751,N_5276,N_5306);
nand U5752 (N_5752,N_5292,N_5275);
nor U5753 (N_5753,N_5498,N_5260);
xor U5754 (N_5754,N_5362,N_5467);
or U5755 (N_5755,N_5101,N_5352);
or U5756 (N_5756,N_5057,N_5328);
nand U5757 (N_5757,N_5065,N_5184);
and U5758 (N_5758,N_5300,N_5178);
and U5759 (N_5759,N_5248,N_5183);
xnor U5760 (N_5760,N_5048,N_5427);
or U5761 (N_5761,N_5115,N_5039);
or U5762 (N_5762,N_5295,N_5076);
nor U5763 (N_5763,N_5246,N_5425);
xor U5764 (N_5764,N_5238,N_5444);
nand U5765 (N_5765,N_5432,N_5400);
or U5766 (N_5766,N_5210,N_5286);
nor U5767 (N_5767,N_5452,N_5055);
xnor U5768 (N_5768,N_5251,N_5413);
or U5769 (N_5769,N_5017,N_5251);
or U5770 (N_5770,N_5067,N_5056);
xor U5771 (N_5771,N_5398,N_5154);
or U5772 (N_5772,N_5326,N_5062);
nor U5773 (N_5773,N_5267,N_5396);
xnor U5774 (N_5774,N_5348,N_5350);
and U5775 (N_5775,N_5151,N_5156);
nand U5776 (N_5776,N_5260,N_5323);
nand U5777 (N_5777,N_5118,N_5231);
xnor U5778 (N_5778,N_5256,N_5245);
and U5779 (N_5779,N_5247,N_5415);
nor U5780 (N_5780,N_5315,N_5328);
nor U5781 (N_5781,N_5440,N_5163);
nand U5782 (N_5782,N_5131,N_5376);
nor U5783 (N_5783,N_5189,N_5214);
or U5784 (N_5784,N_5421,N_5044);
and U5785 (N_5785,N_5403,N_5223);
or U5786 (N_5786,N_5052,N_5022);
nand U5787 (N_5787,N_5092,N_5492);
xnor U5788 (N_5788,N_5470,N_5206);
nor U5789 (N_5789,N_5163,N_5005);
xor U5790 (N_5790,N_5096,N_5397);
nand U5791 (N_5791,N_5207,N_5238);
or U5792 (N_5792,N_5123,N_5429);
and U5793 (N_5793,N_5156,N_5218);
or U5794 (N_5794,N_5028,N_5360);
nand U5795 (N_5795,N_5484,N_5308);
and U5796 (N_5796,N_5451,N_5301);
and U5797 (N_5797,N_5125,N_5157);
or U5798 (N_5798,N_5282,N_5270);
nand U5799 (N_5799,N_5295,N_5261);
and U5800 (N_5800,N_5004,N_5451);
nand U5801 (N_5801,N_5132,N_5190);
and U5802 (N_5802,N_5231,N_5219);
and U5803 (N_5803,N_5041,N_5092);
xor U5804 (N_5804,N_5376,N_5466);
xor U5805 (N_5805,N_5088,N_5113);
or U5806 (N_5806,N_5190,N_5191);
xor U5807 (N_5807,N_5036,N_5065);
xnor U5808 (N_5808,N_5469,N_5394);
xor U5809 (N_5809,N_5296,N_5253);
nor U5810 (N_5810,N_5145,N_5207);
nand U5811 (N_5811,N_5203,N_5185);
nor U5812 (N_5812,N_5284,N_5198);
or U5813 (N_5813,N_5317,N_5164);
nor U5814 (N_5814,N_5426,N_5475);
xnor U5815 (N_5815,N_5172,N_5317);
nand U5816 (N_5816,N_5119,N_5328);
nand U5817 (N_5817,N_5251,N_5296);
and U5818 (N_5818,N_5394,N_5231);
nand U5819 (N_5819,N_5469,N_5376);
nor U5820 (N_5820,N_5101,N_5282);
nor U5821 (N_5821,N_5314,N_5079);
nor U5822 (N_5822,N_5328,N_5003);
and U5823 (N_5823,N_5181,N_5430);
or U5824 (N_5824,N_5137,N_5155);
or U5825 (N_5825,N_5074,N_5400);
xnor U5826 (N_5826,N_5182,N_5409);
xnor U5827 (N_5827,N_5463,N_5082);
nand U5828 (N_5828,N_5161,N_5200);
nand U5829 (N_5829,N_5425,N_5441);
xor U5830 (N_5830,N_5359,N_5395);
nor U5831 (N_5831,N_5424,N_5206);
or U5832 (N_5832,N_5293,N_5030);
nand U5833 (N_5833,N_5228,N_5448);
xnor U5834 (N_5834,N_5055,N_5188);
nor U5835 (N_5835,N_5166,N_5296);
nor U5836 (N_5836,N_5390,N_5220);
xnor U5837 (N_5837,N_5236,N_5079);
xnor U5838 (N_5838,N_5469,N_5245);
or U5839 (N_5839,N_5164,N_5214);
nor U5840 (N_5840,N_5110,N_5089);
nand U5841 (N_5841,N_5381,N_5139);
xor U5842 (N_5842,N_5030,N_5476);
or U5843 (N_5843,N_5149,N_5115);
xnor U5844 (N_5844,N_5307,N_5378);
and U5845 (N_5845,N_5015,N_5441);
nand U5846 (N_5846,N_5419,N_5304);
nand U5847 (N_5847,N_5093,N_5474);
nor U5848 (N_5848,N_5290,N_5089);
or U5849 (N_5849,N_5058,N_5014);
nand U5850 (N_5850,N_5321,N_5408);
nand U5851 (N_5851,N_5475,N_5284);
or U5852 (N_5852,N_5452,N_5156);
nor U5853 (N_5853,N_5261,N_5321);
nor U5854 (N_5854,N_5188,N_5224);
and U5855 (N_5855,N_5227,N_5128);
xnor U5856 (N_5856,N_5386,N_5312);
nand U5857 (N_5857,N_5448,N_5068);
nor U5858 (N_5858,N_5024,N_5190);
nand U5859 (N_5859,N_5087,N_5415);
nor U5860 (N_5860,N_5445,N_5106);
nor U5861 (N_5861,N_5436,N_5443);
xor U5862 (N_5862,N_5118,N_5381);
and U5863 (N_5863,N_5124,N_5005);
nand U5864 (N_5864,N_5414,N_5469);
and U5865 (N_5865,N_5112,N_5450);
nand U5866 (N_5866,N_5448,N_5411);
and U5867 (N_5867,N_5182,N_5281);
nor U5868 (N_5868,N_5471,N_5434);
xor U5869 (N_5869,N_5451,N_5390);
nand U5870 (N_5870,N_5182,N_5239);
or U5871 (N_5871,N_5095,N_5342);
or U5872 (N_5872,N_5356,N_5182);
nor U5873 (N_5873,N_5004,N_5013);
nor U5874 (N_5874,N_5425,N_5384);
nand U5875 (N_5875,N_5304,N_5255);
and U5876 (N_5876,N_5169,N_5477);
nor U5877 (N_5877,N_5369,N_5245);
xor U5878 (N_5878,N_5368,N_5383);
xnor U5879 (N_5879,N_5067,N_5391);
and U5880 (N_5880,N_5046,N_5090);
nor U5881 (N_5881,N_5282,N_5366);
or U5882 (N_5882,N_5409,N_5189);
or U5883 (N_5883,N_5241,N_5345);
nand U5884 (N_5884,N_5050,N_5126);
or U5885 (N_5885,N_5274,N_5409);
or U5886 (N_5886,N_5246,N_5389);
xnor U5887 (N_5887,N_5257,N_5260);
and U5888 (N_5888,N_5472,N_5433);
xnor U5889 (N_5889,N_5379,N_5496);
nor U5890 (N_5890,N_5303,N_5107);
or U5891 (N_5891,N_5081,N_5403);
or U5892 (N_5892,N_5451,N_5132);
and U5893 (N_5893,N_5199,N_5488);
or U5894 (N_5894,N_5480,N_5098);
nand U5895 (N_5895,N_5253,N_5083);
nand U5896 (N_5896,N_5488,N_5441);
nand U5897 (N_5897,N_5013,N_5419);
and U5898 (N_5898,N_5490,N_5377);
nand U5899 (N_5899,N_5305,N_5422);
and U5900 (N_5900,N_5131,N_5300);
nor U5901 (N_5901,N_5108,N_5207);
xnor U5902 (N_5902,N_5340,N_5363);
xnor U5903 (N_5903,N_5008,N_5284);
or U5904 (N_5904,N_5228,N_5280);
and U5905 (N_5905,N_5064,N_5021);
xnor U5906 (N_5906,N_5318,N_5277);
or U5907 (N_5907,N_5382,N_5013);
and U5908 (N_5908,N_5075,N_5428);
and U5909 (N_5909,N_5228,N_5327);
nor U5910 (N_5910,N_5194,N_5227);
nand U5911 (N_5911,N_5112,N_5036);
nor U5912 (N_5912,N_5175,N_5419);
nor U5913 (N_5913,N_5091,N_5368);
and U5914 (N_5914,N_5209,N_5486);
and U5915 (N_5915,N_5371,N_5187);
or U5916 (N_5916,N_5437,N_5486);
xnor U5917 (N_5917,N_5266,N_5228);
nor U5918 (N_5918,N_5432,N_5023);
and U5919 (N_5919,N_5140,N_5156);
or U5920 (N_5920,N_5247,N_5429);
nand U5921 (N_5921,N_5072,N_5013);
and U5922 (N_5922,N_5077,N_5243);
xor U5923 (N_5923,N_5376,N_5015);
xor U5924 (N_5924,N_5412,N_5383);
or U5925 (N_5925,N_5107,N_5374);
nor U5926 (N_5926,N_5168,N_5061);
and U5927 (N_5927,N_5356,N_5117);
and U5928 (N_5928,N_5077,N_5468);
and U5929 (N_5929,N_5318,N_5393);
or U5930 (N_5930,N_5492,N_5362);
nand U5931 (N_5931,N_5468,N_5125);
nand U5932 (N_5932,N_5206,N_5138);
xnor U5933 (N_5933,N_5086,N_5328);
xnor U5934 (N_5934,N_5258,N_5019);
nand U5935 (N_5935,N_5224,N_5108);
and U5936 (N_5936,N_5401,N_5173);
xor U5937 (N_5937,N_5224,N_5411);
and U5938 (N_5938,N_5395,N_5348);
nor U5939 (N_5939,N_5471,N_5293);
and U5940 (N_5940,N_5256,N_5375);
xor U5941 (N_5941,N_5026,N_5034);
or U5942 (N_5942,N_5033,N_5292);
xnor U5943 (N_5943,N_5327,N_5414);
and U5944 (N_5944,N_5350,N_5013);
and U5945 (N_5945,N_5076,N_5129);
xnor U5946 (N_5946,N_5479,N_5131);
xor U5947 (N_5947,N_5178,N_5045);
xnor U5948 (N_5948,N_5426,N_5355);
xor U5949 (N_5949,N_5203,N_5283);
nand U5950 (N_5950,N_5189,N_5444);
nor U5951 (N_5951,N_5118,N_5317);
nand U5952 (N_5952,N_5147,N_5156);
or U5953 (N_5953,N_5142,N_5175);
nor U5954 (N_5954,N_5446,N_5471);
or U5955 (N_5955,N_5035,N_5432);
nand U5956 (N_5956,N_5091,N_5099);
nand U5957 (N_5957,N_5448,N_5263);
or U5958 (N_5958,N_5287,N_5232);
and U5959 (N_5959,N_5025,N_5364);
and U5960 (N_5960,N_5134,N_5174);
and U5961 (N_5961,N_5322,N_5373);
and U5962 (N_5962,N_5108,N_5299);
xnor U5963 (N_5963,N_5132,N_5037);
xnor U5964 (N_5964,N_5313,N_5475);
xor U5965 (N_5965,N_5413,N_5039);
xor U5966 (N_5966,N_5048,N_5213);
xnor U5967 (N_5967,N_5375,N_5470);
and U5968 (N_5968,N_5051,N_5369);
nand U5969 (N_5969,N_5001,N_5373);
and U5970 (N_5970,N_5177,N_5261);
nor U5971 (N_5971,N_5089,N_5107);
and U5972 (N_5972,N_5008,N_5161);
nand U5973 (N_5973,N_5242,N_5316);
nor U5974 (N_5974,N_5425,N_5332);
and U5975 (N_5975,N_5465,N_5068);
xnor U5976 (N_5976,N_5160,N_5384);
nand U5977 (N_5977,N_5096,N_5182);
and U5978 (N_5978,N_5307,N_5435);
xor U5979 (N_5979,N_5469,N_5053);
and U5980 (N_5980,N_5124,N_5069);
nor U5981 (N_5981,N_5491,N_5249);
or U5982 (N_5982,N_5269,N_5064);
xnor U5983 (N_5983,N_5377,N_5392);
nor U5984 (N_5984,N_5197,N_5127);
xor U5985 (N_5985,N_5268,N_5220);
and U5986 (N_5986,N_5149,N_5159);
nor U5987 (N_5987,N_5045,N_5152);
xnor U5988 (N_5988,N_5215,N_5136);
xor U5989 (N_5989,N_5367,N_5278);
and U5990 (N_5990,N_5231,N_5040);
nand U5991 (N_5991,N_5437,N_5493);
nand U5992 (N_5992,N_5336,N_5054);
nand U5993 (N_5993,N_5137,N_5170);
nand U5994 (N_5994,N_5222,N_5144);
nor U5995 (N_5995,N_5048,N_5031);
and U5996 (N_5996,N_5454,N_5177);
nor U5997 (N_5997,N_5445,N_5380);
xor U5998 (N_5998,N_5499,N_5136);
and U5999 (N_5999,N_5173,N_5108);
nand U6000 (N_6000,N_5609,N_5697);
xor U6001 (N_6001,N_5894,N_5585);
and U6002 (N_6002,N_5951,N_5691);
xnor U6003 (N_6003,N_5536,N_5578);
or U6004 (N_6004,N_5808,N_5945);
nor U6005 (N_6005,N_5984,N_5912);
nor U6006 (N_6006,N_5759,N_5590);
nand U6007 (N_6007,N_5998,N_5929);
nand U6008 (N_6008,N_5553,N_5933);
xor U6009 (N_6009,N_5952,N_5742);
xnor U6010 (N_6010,N_5638,N_5762);
and U6011 (N_6011,N_5500,N_5707);
nor U6012 (N_6012,N_5508,N_5613);
or U6013 (N_6013,N_5727,N_5730);
and U6014 (N_6014,N_5736,N_5703);
xnor U6015 (N_6015,N_5812,N_5988);
or U6016 (N_6016,N_5565,N_5985);
or U6017 (N_6017,N_5934,N_5857);
and U6018 (N_6018,N_5893,N_5954);
nand U6019 (N_6019,N_5708,N_5778);
xor U6020 (N_6020,N_5949,N_5623);
or U6021 (N_6021,N_5872,N_5769);
xnor U6022 (N_6022,N_5610,N_5917);
xnor U6023 (N_6023,N_5689,N_5982);
xnor U6024 (N_6024,N_5624,N_5715);
and U6025 (N_6025,N_5836,N_5851);
or U6026 (N_6026,N_5930,N_5546);
nor U6027 (N_6027,N_5598,N_5550);
and U6028 (N_6028,N_5688,N_5973);
nand U6029 (N_6029,N_5704,N_5781);
and U6030 (N_6030,N_5579,N_5895);
and U6031 (N_6031,N_5815,N_5597);
nor U6032 (N_6032,N_5916,N_5844);
and U6033 (N_6033,N_5826,N_5757);
nor U6034 (N_6034,N_5841,N_5821);
and U6035 (N_6035,N_5687,N_5650);
or U6036 (N_6036,N_5504,N_5679);
nand U6037 (N_6037,N_5753,N_5532);
nand U6038 (N_6038,N_5557,N_5659);
and U6039 (N_6039,N_5601,N_5832);
nand U6040 (N_6040,N_5915,N_5563);
nor U6041 (N_6041,N_5962,N_5806);
xnor U6042 (N_6042,N_5822,N_5709);
nor U6043 (N_6043,N_5547,N_5847);
nor U6044 (N_6044,N_5725,N_5670);
and U6045 (N_6045,N_5586,N_5920);
or U6046 (N_6046,N_5771,N_5594);
and U6047 (N_6047,N_5502,N_5790);
nand U6048 (N_6048,N_5849,N_5554);
nand U6049 (N_6049,N_5767,N_5901);
or U6050 (N_6050,N_5943,N_5927);
and U6051 (N_6051,N_5651,N_5657);
xor U6052 (N_6052,N_5775,N_5791);
and U6053 (N_6053,N_5873,N_5542);
nand U6054 (N_6054,N_5556,N_5612);
nand U6055 (N_6055,N_5776,N_5726);
and U6056 (N_6056,N_5939,N_5800);
or U6057 (N_6057,N_5568,N_5674);
xor U6058 (N_6058,N_5859,N_5591);
nand U6059 (N_6059,N_5950,N_5676);
xor U6060 (N_6060,N_5783,N_5947);
nor U6061 (N_6061,N_5887,N_5886);
xor U6062 (N_6062,N_5575,N_5641);
xnor U6063 (N_6063,N_5528,N_5986);
and U6064 (N_6064,N_5580,N_5903);
and U6065 (N_6065,N_5908,N_5979);
and U6066 (N_6066,N_5897,N_5593);
xnor U6067 (N_6067,N_5911,N_5747);
xor U6068 (N_6068,N_5740,N_5605);
and U6069 (N_6069,N_5902,N_5566);
and U6070 (N_6070,N_5827,N_5518);
nor U6071 (N_6071,N_5526,N_5634);
or U6072 (N_6072,N_5660,N_5989);
and U6073 (N_6073,N_5662,N_5675);
or U6074 (N_6074,N_5581,N_5572);
or U6075 (N_6075,N_5999,N_5924);
xnor U6076 (N_6076,N_5639,N_5968);
xor U6077 (N_6077,N_5932,N_5900);
or U6078 (N_6078,N_5522,N_5758);
nand U6079 (N_6079,N_5507,N_5621);
xnor U6080 (N_6080,N_5538,N_5842);
nand U6081 (N_6081,N_5990,N_5737);
or U6082 (N_6082,N_5738,N_5834);
nor U6083 (N_6083,N_5548,N_5652);
or U6084 (N_6084,N_5602,N_5862);
or U6085 (N_6085,N_5763,N_5666);
nor U6086 (N_6086,N_5829,N_5777);
or U6087 (N_6087,N_5785,N_5882);
and U6088 (N_6088,N_5848,N_5571);
nor U6089 (N_6089,N_5818,N_5523);
and U6090 (N_6090,N_5506,N_5835);
nor U6091 (N_6091,N_5701,N_5549);
nand U6092 (N_6092,N_5972,N_5625);
and U6093 (N_6093,N_5875,N_5993);
nand U6094 (N_6094,N_5514,N_5997);
and U6095 (N_6095,N_5607,N_5694);
or U6096 (N_6096,N_5653,N_5587);
and U6097 (N_6097,N_5680,N_5513);
or U6098 (N_6098,N_5828,N_5569);
xor U6099 (N_6099,N_5798,N_5584);
nand U6100 (N_6100,N_5837,N_5723);
nor U6101 (N_6101,N_5987,N_5525);
and U6102 (N_6102,N_5672,N_5671);
or U6103 (N_6103,N_5696,N_5626);
xor U6104 (N_6104,N_5544,N_5501);
xor U6105 (N_6105,N_5729,N_5959);
or U6106 (N_6106,N_5642,N_5739);
and U6107 (N_6107,N_5863,N_5527);
nor U6108 (N_6108,N_5702,N_5773);
and U6109 (N_6109,N_5813,N_5884);
xor U6110 (N_6110,N_5846,N_5649);
nor U6111 (N_6111,N_5640,N_5632);
nand U6112 (N_6112,N_5937,N_5936);
or U6113 (N_6113,N_5899,N_5965);
nor U6114 (N_6114,N_5957,N_5940);
xor U6115 (N_6115,N_5868,N_5796);
nor U6116 (N_6116,N_5520,N_5716);
nor U6117 (N_6117,N_5713,N_5840);
xnor U6118 (N_6118,N_5684,N_5787);
xnor U6119 (N_6119,N_5706,N_5870);
or U6120 (N_6120,N_5963,N_5735);
and U6121 (N_6121,N_5719,N_5668);
xnor U6122 (N_6122,N_5925,N_5619);
nor U6123 (N_6123,N_5823,N_5647);
nand U6124 (N_6124,N_5533,N_5661);
and U6125 (N_6125,N_5881,N_5922);
and U6126 (N_6126,N_5732,N_5627);
nand U6127 (N_6127,N_5971,N_5620);
xnor U6128 (N_6128,N_5637,N_5938);
nand U6129 (N_6129,N_5717,N_5958);
nor U6130 (N_6130,N_5734,N_5606);
nor U6131 (N_6131,N_5695,N_5779);
nand U6132 (N_6132,N_5693,N_5817);
nand U6133 (N_6133,N_5874,N_5573);
nor U6134 (N_6134,N_5786,N_5615);
nand U6135 (N_6135,N_5750,N_5764);
nor U6136 (N_6136,N_5807,N_5978);
nor U6137 (N_6137,N_5975,N_5733);
nor U6138 (N_6138,N_5622,N_5545);
nor U6139 (N_6139,N_5770,N_5761);
and U6140 (N_6140,N_5850,N_5673);
and U6141 (N_6141,N_5705,N_5561);
xnor U6142 (N_6142,N_5755,N_5539);
and U6143 (N_6143,N_5816,N_5918);
xnor U6144 (N_6144,N_5914,N_5690);
or U6145 (N_6145,N_5512,N_5611);
and U6146 (N_6146,N_5754,N_5720);
xor U6147 (N_6147,N_5805,N_5570);
xnor U6148 (N_6148,N_5804,N_5983);
and U6149 (N_6149,N_5780,N_5710);
or U6150 (N_6150,N_5752,N_5852);
or U6151 (N_6151,N_5946,N_5782);
and U6152 (N_6152,N_5698,N_5935);
or U6153 (N_6153,N_5839,N_5564);
nand U6154 (N_6154,N_5955,N_5923);
or U6155 (N_6155,N_5644,N_5596);
xor U6156 (N_6156,N_5948,N_5751);
or U6157 (N_6157,N_5654,N_5854);
nand U6158 (N_6158,N_5756,N_5524);
xnor U6159 (N_6159,N_5853,N_5664);
and U6160 (N_6160,N_5746,N_5744);
nor U6161 (N_6161,N_5560,N_5503);
xor U6162 (N_6162,N_5636,N_5714);
nand U6163 (N_6163,N_5692,N_5718);
xnor U6164 (N_6164,N_5995,N_5741);
or U6165 (N_6165,N_5885,N_5802);
or U6166 (N_6166,N_5898,N_5825);
and U6167 (N_6167,N_5509,N_5877);
xnor U6168 (N_6168,N_5810,N_5505);
nand U6169 (N_6169,N_5977,N_5921);
and U6170 (N_6170,N_5981,N_5833);
nor U6171 (N_6171,N_5931,N_5685);
and U6172 (N_6172,N_5860,N_5941);
and U6173 (N_6173,N_5592,N_5967);
xor U6174 (N_6174,N_5552,N_5803);
nand U6175 (N_6175,N_5669,N_5712);
nand U6176 (N_6176,N_5976,N_5633);
or U6177 (N_6177,N_5876,N_5681);
and U6178 (N_6178,N_5992,N_5656);
or U6179 (N_6179,N_5559,N_5558);
or U6180 (N_6180,N_5996,N_5913);
nand U6181 (N_6181,N_5879,N_5551);
nand U6182 (N_6182,N_5910,N_5699);
nand U6183 (N_6183,N_5534,N_5583);
nand U6184 (N_6184,N_5838,N_5960);
xor U6185 (N_6185,N_5529,N_5909);
nor U6186 (N_6186,N_5510,N_5892);
nand U6187 (N_6187,N_5760,N_5831);
nand U6188 (N_6188,N_5582,N_5700);
nand U6189 (N_6189,N_5801,N_5711);
or U6190 (N_6190,N_5631,N_5797);
nor U6191 (N_6191,N_5974,N_5942);
and U6192 (N_6192,N_5743,N_5956);
or U6193 (N_6193,N_5728,N_5515);
nor U6194 (N_6194,N_5517,N_5969);
nor U6195 (N_6195,N_5600,N_5749);
and U6196 (N_6196,N_5907,N_5646);
and U6197 (N_6197,N_5814,N_5964);
xor U6198 (N_6198,N_5855,N_5889);
or U6199 (N_6199,N_5511,N_5731);
and U6200 (N_6200,N_5867,N_5896);
xor U6201 (N_6201,N_5537,N_5677);
or U6202 (N_6202,N_5686,N_5530);
or U6203 (N_6203,N_5864,N_5628);
and U6204 (N_6204,N_5721,N_5604);
nor U6205 (N_6205,N_5722,N_5926);
and U6206 (N_6206,N_5667,N_5768);
nor U6207 (N_6207,N_5635,N_5878);
or U6208 (N_6208,N_5562,N_5928);
nor U6209 (N_6209,N_5890,N_5792);
or U6210 (N_6210,N_5603,N_5799);
nand U6211 (N_6211,N_5830,N_5643);
and U6212 (N_6212,N_5577,N_5519);
nor U6213 (N_6213,N_5789,N_5766);
nand U6214 (N_6214,N_5888,N_5811);
nor U6215 (N_6215,N_5793,N_5745);
or U6216 (N_6216,N_5535,N_5991);
and U6217 (N_6217,N_5516,N_5906);
nor U6218 (N_6218,N_5865,N_5629);
and U6219 (N_6219,N_5599,N_5574);
xor U6220 (N_6220,N_5961,N_5683);
or U6221 (N_6221,N_5774,N_5891);
and U6222 (N_6222,N_5856,N_5678);
and U6223 (N_6223,N_5843,N_5589);
xor U6224 (N_6224,N_5788,N_5645);
nor U6225 (N_6225,N_5630,N_5880);
nand U6226 (N_6226,N_5648,N_5858);
xnor U6227 (N_6227,N_5845,N_5618);
nor U6228 (N_6228,N_5905,N_5617);
or U6229 (N_6229,N_5614,N_5665);
xnor U6230 (N_6230,N_5595,N_5919);
xnor U6231 (N_6231,N_5944,N_5724);
or U6232 (N_6232,N_5861,N_5994);
nor U6233 (N_6233,N_5824,N_5794);
nor U6234 (N_6234,N_5531,N_5966);
nor U6235 (N_6235,N_5795,N_5820);
nor U6236 (N_6236,N_5970,N_5576);
xor U6237 (N_6237,N_5541,N_5871);
xnor U6238 (N_6238,N_5819,N_5980);
xor U6239 (N_6239,N_5608,N_5748);
or U6240 (N_6240,N_5655,N_5616);
xor U6241 (N_6241,N_5772,N_5658);
and U6242 (N_6242,N_5543,N_5588);
nand U6243 (N_6243,N_5953,N_5540);
nand U6244 (N_6244,N_5682,N_5663);
nand U6245 (N_6245,N_5521,N_5904);
and U6246 (N_6246,N_5555,N_5567);
xor U6247 (N_6247,N_5765,N_5883);
nor U6248 (N_6248,N_5866,N_5869);
xnor U6249 (N_6249,N_5784,N_5809);
xor U6250 (N_6250,N_5901,N_5574);
xor U6251 (N_6251,N_5519,N_5585);
xor U6252 (N_6252,N_5999,N_5604);
xor U6253 (N_6253,N_5616,N_5856);
and U6254 (N_6254,N_5944,N_5671);
nor U6255 (N_6255,N_5841,N_5550);
xor U6256 (N_6256,N_5650,N_5594);
or U6257 (N_6257,N_5739,N_5912);
nand U6258 (N_6258,N_5699,N_5681);
xor U6259 (N_6259,N_5504,N_5768);
or U6260 (N_6260,N_5681,N_5927);
nor U6261 (N_6261,N_5655,N_5931);
and U6262 (N_6262,N_5561,N_5921);
or U6263 (N_6263,N_5524,N_5660);
nor U6264 (N_6264,N_5723,N_5924);
or U6265 (N_6265,N_5812,N_5561);
nor U6266 (N_6266,N_5650,N_5798);
nor U6267 (N_6267,N_5866,N_5625);
and U6268 (N_6268,N_5658,N_5889);
xnor U6269 (N_6269,N_5695,N_5783);
or U6270 (N_6270,N_5992,N_5534);
and U6271 (N_6271,N_5935,N_5707);
xnor U6272 (N_6272,N_5711,N_5559);
or U6273 (N_6273,N_5643,N_5882);
and U6274 (N_6274,N_5566,N_5568);
nand U6275 (N_6275,N_5665,N_5610);
nor U6276 (N_6276,N_5777,N_5522);
nand U6277 (N_6277,N_5591,N_5979);
nand U6278 (N_6278,N_5938,N_5605);
nor U6279 (N_6279,N_5540,N_5712);
or U6280 (N_6280,N_5596,N_5641);
and U6281 (N_6281,N_5855,N_5688);
nor U6282 (N_6282,N_5863,N_5978);
nand U6283 (N_6283,N_5839,N_5830);
nor U6284 (N_6284,N_5633,N_5559);
xor U6285 (N_6285,N_5938,N_5542);
nand U6286 (N_6286,N_5992,N_5722);
xnor U6287 (N_6287,N_5510,N_5783);
nor U6288 (N_6288,N_5596,N_5725);
xor U6289 (N_6289,N_5688,N_5859);
nor U6290 (N_6290,N_5871,N_5695);
xor U6291 (N_6291,N_5727,N_5689);
and U6292 (N_6292,N_5705,N_5691);
xnor U6293 (N_6293,N_5672,N_5522);
or U6294 (N_6294,N_5554,N_5504);
nand U6295 (N_6295,N_5927,N_5622);
nor U6296 (N_6296,N_5715,N_5511);
or U6297 (N_6297,N_5967,N_5590);
xnor U6298 (N_6298,N_5802,N_5908);
or U6299 (N_6299,N_5868,N_5550);
nor U6300 (N_6300,N_5775,N_5645);
nor U6301 (N_6301,N_5670,N_5881);
xnor U6302 (N_6302,N_5539,N_5877);
nor U6303 (N_6303,N_5698,N_5557);
and U6304 (N_6304,N_5618,N_5652);
nand U6305 (N_6305,N_5830,N_5789);
or U6306 (N_6306,N_5953,N_5945);
nor U6307 (N_6307,N_5677,N_5600);
xor U6308 (N_6308,N_5849,N_5838);
or U6309 (N_6309,N_5603,N_5942);
nor U6310 (N_6310,N_5559,N_5580);
or U6311 (N_6311,N_5814,N_5552);
xnor U6312 (N_6312,N_5817,N_5734);
nand U6313 (N_6313,N_5596,N_5551);
xor U6314 (N_6314,N_5738,N_5642);
nor U6315 (N_6315,N_5762,N_5614);
xnor U6316 (N_6316,N_5530,N_5512);
nor U6317 (N_6317,N_5584,N_5825);
xnor U6318 (N_6318,N_5981,N_5877);
and U6319 (N_6319,N_5614,N_5803);
and U6320 (N_6320,N_5595,N_5880);
nor U6321 (N_6321,N_5731,N_5723);
xor U6322 (N_6322,N_5838,N_5702);
or U6323 (N_6323,N_5929,N_5957);
and U6324 (N_6324,N_5964,N_5567);
xnor U6325 (N_6325,N_5563,N_5862);
xor U6326 (N_6326,N_5704,N_5780);
xnor U6327 (N_6327,N_5968,N_5663);
xnor U6328 (N_6328,N_5809,N_5958);
nor U6329 (N_6329,N_5827,N_5884);
xnor U6330 (N_6330,N_5988,N_5886);
xor U6331 (N_6331,N_5646,N_5556);
nand U6332 (N_6332,N_5959,N_5767);
and U6333 (N_6333,N_5731,N_5552);
xnor U6334 (N_6334,N_5990,N_5510);
and U6335 (N_6335,N_5557,N_5893);
xor U6336 (N_6336,N_5904,N_5606);
and U6337 (N_6337,N_5797,N_5515);
and U6338 (N_6338,N_5961,N_5696);
or U6339 (N_6339,N_5939,N_5761);
nor U6340 (N_6340,N_5693,N_5800);
nand U6341 (N_6341,N_5535,N_5565);
nor U6342 (N_6342,N_5534,N_5868);
nand U6343 (N_6343,N_5697,N_5844);
and U6344 (N_6344,N_5639,N_5528);
or U6345 (N_6345,N_5938,N_5850);
or U6346 (N_6346,N_5554,N_5923);
xor U6347 (N_6347,N_5978,N_5631);
and U6348 (N_6348,N_5831,N_5645);
xor U6349 (N_6349,N_5775,N_5622);
or U6350 (N_6350,N_5522,N_5741);
and U6351 (N_6351,N_5927,N_5653);
nand U6352 (N_6352,N_5989,N_5636);
or U6353 (N_6353,N_5775,N_5868);
xnor U6354 (N_6354,N_5630,N_5732);
or U6355 (N_6355,N_5918,N_5535);
or U6356 (N_6356,N_5709,N_5585);
nand U6357 (N_6357,N_5805,N_5840);
nand U6358 (N_6358,N_5779,N_5784);
nor U6359 (N_6359,N_5753,N_5755);
nor U6360 (N_6360,N_5789,N_5605);
nor U6361 (N_6361,N_5715,N_5527);
nand U6362 (N_6362,N_5795,N_5663);
or U6363 (N_6363,N_5715,N_5873);
or U6364 (N_6364,N_5871,N_5743);
nor U6365 (N_6365,N_5755,N_5700);
xnor U6366 (N_6366,N_5798,N_5837);
nor U6367 (N_6367,N_5846,N_5885);
nand U6368 (N_6368,N_5630,N_5925);
xnor U6369 (N_6369,N_5902,N_5793);
nand U6370 (N_6370,N_5705,N_5584);
and U6371 (N_6371,N_5857,N_5803);
or U6372 (N_6372,N_5862,N_5508);
nor U6373 (N_6373,N_5824,N_5653);
xnor U6374 (N_6374,N_5877,N_5852);
and U6375 (N_6375,N_5699,N_5769);
and U6376 (N_6376,N_5606,N_5942);
nor U6377 (N_6377,N_5786,N_5753);
or U6378 (N_6378,N_5504,N_5543);
or U6379 (N_6379,N_5921,N_5628);
or U6380 (N_6380,N_5780,N_5769);
nor U6381 (N_6381,N_5586,N_5540);
nor U6382 (N_6382,N_5546,N_5625);
or U6383 (N_6383,N_5614,N_5684);
nor U6384 (N_6384,N_5894,N_5619);
nor U6385 (N_6385,N_5511,N_5846);
xor U6386 (N_6386,N_5840,N_5592);
xnor U6387 (N_6387,N_5518,N_5659);
or U6388 (N_6388,N_5614,N_5692);
nand U6389 (N_6389,N_5940,N_5938);
and U6390 (N_6390,N_5982,N_5705);
nor U6391 (N_6391,N_5917,N_5532);
xor U6392 (N_6392,N_5952,N_5955);
xor U6393 (N_6393,N_5917,N_5576);
nor U6394 (N_6394,N_5726,N_5841);
or U6395 (N_6395,N_5654,N_5563);
or U6396 (N_6396,N_5733,N_5840);
nand U6397 (N_6397,N_5760,N_5536);
or U6398 (N_6398,N_5600,N_5697);
nor U6399 (N_6399,N_5572,N_5871);
nor U6400 (N_6400,N_5547,N_5542);
nand U6401 (N_6401,N_5750,N_5844);
or U6402 (N_6402,N_5919,N_5731);
and U6403 (N_6403,N_5641,N_5633);
xnor U6404 (N_6404,N_5902,N_5933);
or U6405 (N_6405,N_5866,N_5911);
xnor U6406 (N_6406,N_5791,N_5718);
and U6407 (N_6407,N_5658,N_5914);
nor U6408 (N_6408,N_5960,N_5814);
and U6409 (N_6409,N_5785,N_5553);
and U6410 (N_6410,N_5708,N_5727);
and U6411 (N_6411,N_5755,N_5828);
nand U6412 (N_6412,N_5694,N_5902);
nor U6413 (N_6413,N_5500,N_5961);
or U6414 (N_6414,N_5557,N_5657);
xnor U6415 (N_6415,N_5637,N_5644);
nand U6416 (N_6416,N_5927,N_5585);
nor U6417 (N_6417,N_5751,N_5684);
nor U6418 (N_6418,N_5583,N_5573);
or U6419 (N_6419,N_5604,N_5743);
nand U6420 (N_6420,N_5587,N_5505);
or U6421 (N_6421,N_5535,N_5795);
and U6422 (N_6422,N_5966,N_5747);
or U6423 (N_6423,N_5783,N_5714);
xnor U6424 (N_6424,N_5837,N_5603);
xnor U6425 (N_6425,N_5629,N_5973);
nand U6426 (N_6426,N_5900,N_5528);
nor U6427 (N_6427,N_5645,N_5872);
nand U6428 (N_6428,N_5568,N_5877);
nand U6429 (N_6429,N_5728,N_5977);
nand U6430 (N_6430,N_5643,N_5583);
nor U6431 (N_6431,N_5809,N_5811);
xor U6432 (N_6432,N_5815,N_5818);
or U6433 (N_6433,N_5803,N_5659);
nand U6434 (N_6434,N_5570,N_5542);
nor U6435 (N_6435,N_5854,N_5996);
or U6436 (N_6436,N_5939,N_5555);
and U6437 (N_6437,N_5517,N_5848);
xnor U6438 (N_6438,N_5738,N_5748);
or U6439 (N_6439,N_5887,N_5730);
and U6440 (N_6440,N_5909,N_5809);
or U6441 (N_6441,N_5957,N_5802);
xnor U6442 (N_6442,N_5785,N_5970);
xor U6443 (N_6443,N_5884,N_5846);
or U6444 (N_6444,N_5717,N_5929);
xor U6445 (N_6445,N_5970,N_5524);
nand U6446 (N_6446,N_5845,N_5598);
nor U6447 (N_6447,N_5919,N_5715);
xnor U6448 (N_6448,N_5800,N_5742);
xnor U6449 (N_6449,N_5574,N_5667);
xor U6450 (N_6450,N_5944,N_5773);
and U6451 (N_6451,N_5597,N_5776);
nor U6452 (N_6452,N_5960,N_5859);
and U6453 (N_6453,N_5950,N_5654);
nand U6454 (N_6454,N_5760,N_5751);
and U6455 (N_6455,N_5580,N_5578);
and U6456 (N_6456,N_5613,N_5989);
nor U6457 (N_6457,N_5567,N_5641);
and U6458 (N_6458,N_5780,N_5933);
xnor U6459 (N_6459,N_5696,N_5687);
or U6460 (N_6460,N_5886,N_5783);
xor U6461 (N_6461,N_5641,N_5729);
xnor U6462 (N_6462,N_5839,N_5921);
and U6463 (N_6463,N_5653,N_5869);
xnor U6464 (N_6464,N_5874,N_5862);
and U6465 (N_6465,N_5509,N_5644);
or U6466 (N_6466,N_5523,N_5764);
nor U6467 (N_6467,N_5587,N_5571);
nor U6468 (N_6468,N_5588,N_5969);
xnor U6469 (N_6469,N_5976,N_5980);
nand U6470 (N_6470,N_5642,N_5568);
and U6471 (N_6471,N_5814,N_5898);
and U6472 (N_6472,N_5803,N_5991);
or U6473 (N_6473,N_5597,N_5535);
nand U6474 (N_6474,N_5622,N_5582);
nand U6475 (N_6475,N_5707,N_5664);
nor U6476 (N_6476,N_5573,N_5737);
nor U6477 (N_6477,N_5564,N_5836);
xnor U6478 (N_6478,N_5515,N_5662);
and U6479 (N_6479,N_5553,N_5736);
xor U6480 (N_6480,N_5986,N_5515);
nor U6481 (N_6481,N_5681,N_5625);
or U6482 (N_6482,N_5900,N_5940);
and U6483 (N_6483,N_5703,N_5546);
nand U6484 (N_6484,N_5970,N_5735);
nor U6485 (N_6485,N_5774,N_5565);
or U6486 (N_6486,N_5874,N_5645);
or U6487 (N_6487,N_5967,N_5516);
or U6488 (N_6488,N_5664,N_5553);
nor U6489 (N_6489,N_5553,N_5849);
nand U6490 (N_6490,N_5972,N_5850);
xor U6491 (N_6491,N_5962,N_5646);
nand U6492 (N_6492,N_5559,N_5894);
or U6493 (N_6493,N_5704,N_5751);
nor U6494 (N_6494,N_5683,N_5838);
and U6495 (N_6495,N_5721,N_5518);
nor U6496 (N_6496,N_5517,N_5534);
nor U6497 (N_6497,N_5654,N_5532);
nand U6498 (N_6498,N_5539,N_5708);
and U6499 (N_6499,N_5536,N_5714);
nor U6500 (N_6500,N_6188,N_6324);
nand U6501 (N_6501,N_6235,N_6282);
or U6502 (N_6502,N_6312,N_6387);
nand U6503 (N_6503,N_6109,N_6300);
or U6504 (N_6504,N_6278,N_6068);
xor U6505 (N_6505,N_6449,N_6301);
xor U6506 (N_6506,N_6355,N_6447);
nand U6507 (N_6507,N_6118,N_6227);
or U6508 (N_6508,N_6457,N_6377);
nor U6509 (N_6509,N_6178,N_6340);
xnor U6510 (N_6510,N_6439,N_6407);
xor U6511 (N_6511,N_6041,N_6175);
nand U6512 (N_6512,N_6067,N_6198);
or U6513 (N_6513,N_6002,N_6470);
nor U6514 (N_6514,N_6362,N_6464);
or U6515 (N_6515,N_6414,N_6336);
or U6516 (N_6516,N_6452,N_6455);
xnor U6517 (N_6517,N_6090,N_6213);
xor U6518 (N_6518,N_6215,N_6158);
xor U6519 (N_6519,N_6219,N_6016);
xor U6520 (N_6520,N_6234,N_6098);
xor U6521 (N_6521,N_6023,N_6124);
xnor U6522 (N_6522,N_6165,N_6454);
xnor U6523 (N_6523,N_6145,N_6202);
nand U6524 (N_6524,N_6030,N_6402);
xnor U6525 (N_6525,N_6057,N_6400);
xnor U6526 (N_6526,N_6038,N_6256);
and U6527 (N_6527,N_6248,N_6209);
or U6528 (N_6528,N_6021,N_6321);
or U6529 (N_6529,N_6149,N_6232);
xor U6530 (N_6530,N_6420,N_6385);
nand U6531 (N_6531,N_6058,N_6037);
and U6532 (N_6532,N_6172,N_6448);
nand U6533 (N_6533,N_6259,N_6076);
and U6534 (N_6534,N_6056,N_6252);
nand U6535 (N_6535,N_6040,N_6095);
and U6536 (N_6536,N_6116,N_6373);
xor U6537 (N_6537,N_6401,N_6126);
or U6538 (N_6538,N_6157,N_6043);
and U6539 (N_6539,N_6024,N_6280);
and U6540 (N_6540,N_6254,N_6463);
and U6541 (N_6541,N_6263,N_6257);
nand U6542 (N_6542,N_6378,N_6242);
nor U6543 (N_6543,N_6123,N_6120);
nor U6544 (N_6544,N_6368,N_6425);
nor U6545 (N_6545,N_6361,N_6383);
or U6546 (N_6546,N_6372,N_6065);
nor U6547 (N_6547,N_6154,N_6322);
xor U6548 (N_6548,N_6140,N_6394);
nor U6549 (N_6549,N_6071,N_6250);
nor U6550 (N_6550,N_6207,N_6005);
or U6551 (N_6551,N_6147,N_6131);
xnor U6552 (N_6552,N_6319,N_6445);
nor U6553 (N_6553,N_6335,N_6450);
nand U6554 (N_6554,N_6033,N_6003);
nor U6555 (N_6555,N_6429,N_6471);
nand U6556 (N_6556,N_6416,N_6332);
nand U6557 (N_6557,N_6089,N_6411);
xor U6558 (N_6558,N_6081,N_6281);
xor U6559 (N_6559,N_6036,N_6063);
nand U6560 (N_6560,N_6150,N_6477);
nor U6561 (N_6561,N_6034,N_6093);
and U6562 (N_6562,N_6121,N_6231);
nand U6563 (N_6563,N_6054,N_6186);
nor U6564 (N_6564,N_6070,N_6004);
xor U6565 (N_6565,N_6212,N_6313);
and U6566 (N_6566,N_6496,N_6384);
and U6567 (N_6567,N_6039,N_6433);
xnor U6568 (N_6568,N_6430,N_6266);
xnor U6569 (N_6569,N_6277,N_6148);
and U6570 (N_6570,N_6084,N_6099);
nor U6571 (N_6571,N_6436,N_6261);
and U6572 (N_6572,N_6276,N_6304);
xor U6573 (N_6573,N_6217,N_6097);
and U6574 (N_6574,N_6087,N_6489);
nor U6575 (N_6575,N_6382,N_6046);
nand U6576 (N_6576,N_6224,N_6230);
nand U6577 (N_6577,N_6458,N_6102);
and U6578 (N_6578,N_6258,N_6006);
xor U6579 (N_6579,N_6139,N_6001);
or U6580 (N_6580,N_6194,N_6347);
nand U6581 (N_6581,N_6299,N_6160);
nand U6582 (N_6582,N_6395,N_6125);
xor U6583 (N_6583,N_6191,N_6115);
xnor U6584 (N_6584,N_6474,N_6018);
or U6585 (N_6585,N_6141,N_6424);
xnor U6586 (N_6586,N_6268,N_6246);
and U6587 (N_6587,N_6152,N_6182);
nand U6588 (N_6588,N_6262,N_6376);
xnor U6589 (N_6589,N_6438,N_6408);
and U6590 (N_6590,N_6079,N_6122);
and U6591 (N_6591,N_6468,N_6333);
and U6592 (N_6592,N_6302,N_6222);
and U6593 (N_6593,N_6074,N_6443);
or U6594 (N_6594,N_6486,N_6161);
nor U6595 (N_6595,N_6228,N_6275);
or U6596 (N_6596,N_6075,N_6360);
xnor U6597 (N_6597,N_6290,N_6239);
or U6598 (N_6598,N_6206,N_6350);
nand U6599 (N_6599,N_6069,N_6047);
nand U6600 (N_6600,N_6127,N_6293);
nand U6601 (N_6601,N_6472,N_6326);
and U6602 (N_6602,N_6328,N_6014);
nor U6603 (N_6603,N_6226,N_6241);
or U6604 (N_6604,N_6491,N_6142);
and U6605 (N_6605,N_6417,N_6091);
or U6606 (N_6606,N_6110,N_6174);
or U6607 (N_6607,N_6391,N_6351);
xnor U6608 (N_6608,N_6478,N_6442);
xnor U6609 (N_6609,N_6484,N_6113);
or U6610 (N_6610,N_6044,N_6331);
or U6611 (N_6611,N_6229,N_6273);
and U6612 (N_6612,N_6461,N_6208);
nor U6613 (N_6613,N_6143,N_6088);
or U6614 (N_6614,N_6077,N_6279);
nor U6615 (N_6615,N_6473,N_6151);
and U6616 (N_6616,N_6444,N_6431);
xor U6617 (N_6617,N_6380,N_6469);
nand U6618 (N_6618,N_6171,N_6138);
xor U6619 (N_6619,N_6316,N_6195);
or U6620 (N_6620,N_6035,N_6105);
xnor U6621 (N_6621,N_6103,N_6356);
and U6622 (N_6622,N_6497,N_6104);
or U6623 (N_6623,N_6406,N_6237);
xor U6624 (N_6624,N_6218,N_6050);
and U6625 (N_6625,N_6000,N_6495);
or U6626 (N_6626,N_6374,N_6342);
xnor U6627 (N_6627,N_6137,N_6423);
nand U6628 (N_6628,N_6240,N_6045);
and U6629 (N_6629,N_6216,N_6183);
nand U6630 (N_6630,N_6390,N_6305);
nor U6631 (N_6631,N_6185,N_6462);
xor U6632 (N_6632,N_6418,N_6236);
and U6633 (N_6633,N_6184,N_6119);
and U6634 (N_6634,N_6082,N_6187);
xor U6635 (N_6635,N_6337,N_6386);
xnor U6636 (N_6636,N_6288,N_6012);
and U6637 (N_6637,N_6271,N_6265);
or U6638 (N_6638,N_6189,N_6323);
nand U6639 (N_6639,N_6490,N_6397);
nor U6640 (N_6640,N_6211,N_6086);
and U6641 (N_6641,N_6169,N_6479);
xor U6642 (N_6642,N_6010,N_6365);
or U6643 (N_6643,N_6199,N_6349);
nand U6644 (N_6644,N_6136,N_6192);
or U6645 (N_6645,N_6247,N_6107);
and U6646 (N_6646,N_6308,N_6357);
nand U6647 (N_6647,N_6201,N_6481);
nor U6648 (N_6648,N_6432,N_6163);
and U6649 (N_6649,N_6399,N_6015);
and U6650 (N_6650,N_6428,N_6475);
nor U6651 (N_6651,N_6128,N_6393);
and U6652 (N_6652,N_6285,N_6132);
nand U6653 (N_6653,N_6060,N_6112);
and U6654 (N_6654,N_6334,N_6467);
xnor U6655 (N_6655,N_6251,N_6498);
or U6656 (N_6656,N_6066,N_6409);
or U6657 (N_6657,N_6204,N_6249);
xnor U6658 (N_6658,N_6117,N_6085);
nor U6659 (N_6659,N_6108,N_6064);
nand U6660 (N_6660,N_6164,N_6270);
xor U6661 (N_6661,N_6162,N_6482);
nor U6662 (N_6662,N_6341,N_6286);
or U6663 (N_6663,N_6398,N_6283);
xor U6664 (N_6664,N_6028,N_6094);
or U6665 (N_6665,N_6348,N_6106);
nor U6666 (N_6666,N_6296,N_6181);
or U6667 (N_6667,N_6072,N_6287);
nand U6668 (N_6668,N_6413,N_6101);
or U6669 (N_6669,N_6027,N_6415);
nand U6670 (N_6670,N_6059,N_6049);
nor U6671 (N_6671,N_6346,N_6388);
xnor U6672 (N_6672,N_6111,N_6200);
xnor U6673 (N_6673,N_6100,N_6274);
xor U6674 (N_6674,N_6245,N_6255);
nand U6675 (N_6675,N_6007,N_6303);
nor U6676 (N_6676,N_6327,N_6210);
xor U6677 (N_6677,N_6440,N_6359);
nand U6678 (N_6678,N_6170,N_6114);
nand U6679 (N_6679,N_6493,N_6166);
nand U6680 (N_6680,N_6476,N_6221);
nor U6681 (N_6681,N_6310,N_6453);
xor U6682 (N_6682,N_6367,N_6465);
and U6683 (N_6683,N_6381,N_6267);
nand U6684 (N_6684,N_6205,N_6329);
or U6685 (N_6685,N_6193,N_6480);
and U6686 (N_6686,N_6180,N_6244);
or U6687 (N_6687,N_6403,N_6214);
nand U6688 (N_6688,N_6344,N_6260);
and U6689 (N_6689,N_6153,N_6092);
and U6690 (N_6690,N_6155,N_6253);
nor U6691 (N_6691,N_6019,N_6499);
or U6692 (N_6692,N_6048,N_6318);
nand U6693 (N_6693,N_6325,N_6146);
or U6694 (N_6694,N_6156,N_6022);
and U6695 (N_6695,N_6061,N_6422);
nor U6696 (N_6696,N_6456,N_6190);
and U6697 (N_6697,N_6284,N_6083);
nand U6698 (N_6698,N_6062,N_6306);
xor U6699 (N_6699,N_6494,N_6130);
nor U6700 (N_6700,N_6441,N_6042);
nand U6701 (N_6701,N_6358,N_6295);
or U6702 (N_6702,N_6460,N_6233);
nand U6703 (N_6703,N_6029,N_6421);
nand U6704 (N_6704,N_6352,N_6291);
nor U6705 (N_6705,N_6426,N_6177);
xor U6706 (N_6706,N_6315,N_6055);
xnor U6707 (N_6707,N_6375,N_6353);
nor U6708 (N_6708,N_6392,N_6412);
xnor U6709 (N_6709,N_6289,N_6176);
and U6710 (N_6710,N_6404,N_6223);
xor U6711 (N_6711,N_6338,N_6080);
xor U6712 (N_6712,N_6051,N_6298);
or U6713 (N_6713,N_6173,N_6488);
xnor U6714 (N_6714,N_6487,N_6032);
and U6715 (N_6715,N_6446,N_6320);
xnor U6716 (N_6716,N_6379,N_6129);
nand U6717 (N_6717,N_6330,N_6317);
nor U6718 (N_6718,N_6405,N_6159);
nor U6719 (N_6719,N_6369,N_6179);
nand U6720 (N_6720,N_6011,N_6485);
xor U6721 (N_6721,N_6026,N_6017);
nor U6722 (N_6722,N_6292,N_6144);
or U6723 (N_6723,N_6366,N_6466);
nor U6724 (N_6724,N_6309,N_6363);
and U6725 (N_6725,N_6135,N_6167);
xor U6726 (N_6726,N_6196,N_6389);
xor U6727 (N_6727,N_6031,N_6197);
xnor U6728 (N_6728,N_6297,N_6419);
and U6729 (N_6729,N_6294,N_6009);
xor U6730 (N_6730,N_6053,N_6243);
nor U6731 (N_6731,N_6370,N_6434);
and U6732 (N_6732,N_6134,N_6364);
and U6733 (N_6733,N_6269,N_6343);
or U6734 (N_6734,N_6238,N_6052);
xnor U6735 (N_6735,N_6483,N_6314);
nand U6736 (N_6736,N_6264,N_6492);
or U6737 (N_6737,N_6020,N_6025);
nor U6738 (N_6738,N_6339,N_6345);
nor U6739 (N_6739,N_6371,N_6220);
nor U6740 (N_6740,N_6203,N_6410);
and U6741 (N_6741,N_6078,N_6272);
nand U6742 (N_6742,N_6354,N_6451);
nand U6743 (N_6743,N_6307,N_6437);
nor U6744 (N_6744,N_6435,N_6396);
nor U6745 (N_6745,N_6427,N_6096);
nor U6746 (N_6746,N_6008,N_6168);
nand U6747 (N_6747,N_6013,N_6073);
xnor U6748 (N_6748,N_6225,N_6459);
xor U6749 (N_6749,N_6311,N_6133);
or U6750 (N_6750,N_6002,N_6204);
and U6751 (N_6751,N_6326,N_6482);
xor U6752 (N_6752,N_6063,N_6089);
or U6753 (N_6753,N_6147,N_6058);
nor U6754 (N_6754,N_6047,N_6089);
or U6755 (N_6755,N_6268,N_6097);
nand U6756 (N_6756,N_6044,N_6374);
nor U6757 (N_6757,N_6256,N_6418);
nand U6758 (N_6758,N_6256,N_6184);
nand U6759 (N_6759,N_6396,N_6012);
xnor U6760 (N_6760,N_6443,N_6296);
nand U6761 (N_6761,N_6248,N_6337);
nand U6762 (N_6762,N_6413,N_6095);
xnor U6763 (N_6763,N_6303,N_6184);
or U6764 (N_6764,N_6219,N_6235);
xor U6765 (N_6765,N_6035,N_6080);
nor U6766 (N_6766,N_6116,N_6024);
or U6767 (N_6767,N_6088,N_6044);
nand U6768 (N_6768,N_6074,N_6427);
nand U6769 (N_6769,N_6445,N_6469);
and U6770 (N_6770,N_6164,N_6319);
and U6771 (N_6771,N_6271,N_6069);
xnor U6772 (N_6772,N_6400,N_6258);
and U6773 (N_6773,N_6497,N_6369);
or U6774 (N_6774,N_6481,N_6305);
or U6775 (N_6775,N_6312,N_6147);
xnor U6776 (N_6776,N_6316,N_6194);
nand U6777 (N_6777,N_6231,N_6148);
xnor U6778 (N_6778,N_6361,N_6407);
nand U6779 (N_6779,N_6370,N_6493);
or U6780 (N_6780,N_6221,N_6238);
nand U6781 (N_6781,N_6477,N_6430);
nand U6782 (N_6782,N_6263,N_6076);
nor U6783 (N_6783,N_6079,N_6191);
nor U6784 (N_6784,N_6379,N_6429);
xor U6785 (N_6785,N_6427,N_6335);
nand U6786 (N_6786,N_6404,N_6376);
xnor U6787 (N_6787,N_6239,N_6068);
or U6788 (N_6788,N_6162,N_6477);
xnor U6789 (N_6789,N_6354,N_6125);
nand U6790 (N_6790,N_6015,N_6322);
or U6791 (N_6791,N_6486,N_6405);
xor U6792 (N_6792,N_6311,N_6290);
xor U6793 (N_6793,N_6069,N_6383);
nor U6794 (N_6794,N_6269,N_6440);
xor U6795 (N_6795,N_6205,N_6085);
and U6796 (N_6796,N_6148,N_6134);
nand U6797 (N_6797,N_6395,N_6234);
and U6798 (N_6798,N_6449,N_6036);
xor U6799 (N_6799,N_6327,N_6168);
or U6800 (N_6800,N_6347,N_6152);
nor U6801 (N_6801,N_6233,N_6020);
nand U6802 (N_6802,N_6014,N_6057);
nand U6803 (N_6803,N_6023,N_6468);
or U6804 (N_6804,N_6380,N_6087);
xnor U6805 (N_6805,N_6346,N_6058);
nor U6806 (N_6806,N_6427,N_6133);
and U6807 (N_6807,N_6010,N_6064);
xor U6808 (N_6808,N_6285,N_6015);
nor U6809 (N_6809,N_6068,N_6303);
nand U6810 (N_6810,N_6156,N_6390);
and U6811 (N_6811,N_6370,N_6180);
or U6812 (N_6812,N_6379,N_6230);
or U6813 (N_6813,N_6086,N_6336);
xnor U6814 (N_6814,N_6008,N_6485);
nor U6815 (N_6815,N_6115,N_6092);
and U6816 (N_6816,N_6462,N_6001);
nand U6817 (N_6817,N_6224,N_6089);
or U6818 (N_6818,N_6154,N_6186);
nand U6819 (N_6819,N_6065,N_6091);
or U6820 (N_6820,N_6275,N_6485);
or U6821 (N_6821,N_6097,N_6482);
or U6822 (N_6822,N_6161,N_6309);
and U6823 (N_6823,N_6130,N_6024);
and U6824 (N_6824,N_6166,N_6012);
nand U6825 (N_6825,N_6115,N_6418);
nor U6826 (N_6826,N_6165,N_6172);
and U6827 (N_6827,N_6372,N_6278);
xnor U6828 (N_6828,N_6382,N_6080);
nand U6829 (N_6829,N_6035,N_6376);
nor U6830 (N_6830,N_6351,N_6024);
or U6831 (N_6831,N_6048,N_6162);
and U6832 (N_6832,N_6457,N_6019);
nor U6833 (N_6833,N_6227,N_6247);
xnor U6834 (N_6834,N_6180,N_6397);
or U6835 (N_6835,N_6448,N_6356);
nand U6836 (N_6836,N_6330,N_6123);
and U6837 (N_6837,N_6304,N_6278);
and U6838 (N_6838,N_6214,N_6212);
xnor U6839 (N_6839,N_6364,N_6439);
xor U6840 (N_6840,N_6263,N_6380);
nor U6841 (N_6841,N_6035,N_6455);
xor U6842 (N_6842,N_6127,N_6053);
nand U6843 (N_6843,N_6233,N_6018);
nand U6844 (N_6844,N_6056,N_6035);
and U6845 (N_6845,N_6379,N_6261);
xor U6846 (N_6846,N_6135,N_6040);
or U6847 (N_6847,N_6203,N_6186);
and U6848 (N_6848,N_6275,N_6012);
and U6849 (N_6849,N_6242,N_6201);
and U6850 (N_6850,N_6421,N_6360);
nor U6851 (N_6851,N_6485,N_6390);
and U6852 (N_6852,N_6042,N_6108);
nand U6853 (N_6853,N_6335,N_6008);
or U6854 (N_6854,N_6369,N_6351);
nand U6855 (N_6855,N_6082,N_6005);
xnor U6856 (N_6856,N_6098,N_6279);
nand U6857 (N_6857,N_6237,N_6483);
or U6858 (N_6858,N_6228,N_6199);
nand U6859 (N_6859,N_6021,N_6306);
nand U6860 (N_6860,N_6084,N_6483);
nor U6861 (N_6861,N_6316,N_6319);
nand U6862 (N_6862,N_6372,N_6487);
xor U6863 (N_6863,N_6484,N_6058);
and U6864 (N_6864,N_6224,N_6088);
or U6865 (N_6865,N_6489,N_6020);
and U6866 (N_6866,N_6161,N_6332);
nand U6867 (N_6867,N_6378,N_6117);
nor U6868 (N_6868,N_6268,N_6466);
xor U6869 (N_6869,N_6445,N_6461);
or U6870 (N_6870,N_6390,N_6097);
xnor U6871 (N_6871,N_6306,N_6274);
nand U6872 (N_6872,N_6038,N_6193);
or U6873 (N_6873,N_6307,N_6231);
and U6874 (N_6874,N_6027,N_6262);
nor U6875 (N_6875,N_6464,N_6120);
and U6876 (N_6876,N_6093,N_6105);
xnor U6877 (N_6877,N_6109,N_6456);
and U6878 (N_6878,N_6403,N_6441);
nand U6879 (N_6879,N_6353,N_6093);
or U6880 (N_6880,N_6400,N_6312);
nor U6881 (N_6881,N_6280,N_6402);
nor U6882 (N_6882,N_6060,N_6125);
and U6883 (N_6883,N_6036,N_6305);
and U6884 (N_6884,N_6051,N_6179);
and U6885 (N_6885,N_6418,N_6436);
nor U6886 (N_6886,N_6157,N_6354);
or U6887 (N_6887,N_6481,N_6283);
nand U6888 (N_6888,N_6170,N_6341);
nand U6889 (N_6889,N_6444,N_6388);
nor U6890 (N_6890,N_6224,N_6357);
xnor U6891 (N_6891,N_6276,N_6233);
xnor U6892 (N_6892,N_6434,N_6248);
xor U6893 (N_6893,N_6251,N_6385);
xor U6894 (N_6894,N_6477,N_6341);
nand U6895 (N_6895,N_6426,N_6347);
or U6896 (N_6896,N_6461,N_6287);
nand U6897 (N_6897,N_6078,N_6239);
nor U6898 (N_6898,N_6499,N_6423);
or U6899 (N_6899,N_6467,N_6356);
or U6900 (N_6900,N_6232,N_6386);
and U6901 (N_6901,N_6368,N_6344);
nor U6902 (N_6902,N_6200,N_6103);
nor U6903 (N_6903,N_6116,N_6489);
nor U6904 (N_6904,N_6094,N_6242);
xnor U6905 (N_6905,N_6472,N_6094);
nand U6906 (N_6906,N_6374,N_6151);
and U6907 (N_6907,N_6152,N_6444);
xor U6908 (N_6908,N_6437,N_6444);
nor U6909 (N_6909,N_6167,N_6482);
nor U6910 (N_6910,N_6088,N_6202);
nand U6911 (N_6911,N_6065,N_6137);
and U6912 (N_6912,N_6341,N_6208);
nand U6913 (N_6913,N_6329,N_6348);
xor U6914 (N_6914,N_6165,N_6375);
nand U6915 (N_6915,N_6147,N_6219);
nand U6916 (N_6916,N_6074,N_6161);
and U6917 (N_6917,N_6025,N_6449);
nor U6918 (N_6918,N_6321,N_6264);
xnor U6919 (N_6919,N_6084,N_6297);
and U6920 (N_6920,N_6410,N_6065);
and U6921 (N_6921,N_6081,N_6280);
nor U6922 (N_6922,N_6449,N_6458);
nand U6923 (N_6923,N_6388,N_6013);
xnor U6924 (N_6924,N_6012,N_6434);
or U6925 (N_6925,N_6241,N_6261);
nand U6926 (N_6926,N_6240,N_6074);
and U6927 (N_6927,N_6276,N_6391);
nand U6928 (N_6928,N_6366,N_6204);
xor U6929 (N_6929,N_6355,N_6499);
xor U6930 (N_6930,N_6299,N_6294);
xor U6931 (N_6931,N_6246,N_6086);
nand U6932 (N_6932,N_6246,N_6124);
and U6933 (N_6933,N_6333,N_6170);
or U6934 (N_6934,N_6106,N_6308);
nand U6935 (N_6935,N_6139,N_6094);
or U6936 (N_6936,N_6212,N_6070);
nand U6937 (N_6937,N_6020,N_6164);
nor U6938 (N_6938,N_6065,N_6425);
and U6939 (N_6939,N_6122,N_6089);
nor U6940 (N_6940,N_6489,N_6117);
or U6941 (N_6941,N_6223,N_6002);
nand U6942 (N_6942,N_6299,N_6247);
xor U6943 (N_6943,N_6016,N_6200);
and U6944 (N_6944,N_6361,N_6437);
nor U6945 (N_6945,N_6115,N_6270);
or U6946 (N_6946,N_6415,N_6135);
nand U6947 (N_6947,N_6229,N_6215);
nand U6948 (N_6948,N_6142,N_6461);
nand U6949 (N_6949,N_6057,N_6137);
and U6950 (N_6950,N_6281,N_6203);
xnor U6951 (N_6951,N_6412,N_6376);
nor U6952 (N_6952,N_6273,N_6046);
nor U6953 (N_6953,N_6427,N_6497);
or U6954 (N_6954,N_6431,N_6163);
or U6955 (N_6955,N_6369,N_6184);
xnor U6956 (N_6956,N_6216,N_6022);
or U6957 (N_6957,N_6378,N_6290);
and U6958 (N_6958,N_6060,N_6199);
nand U6959 (N_6959,N_6187,N_6115);
nand U6960 (N_6960,N_6112,N_6426);
and U6961 (N_6961,N_6368,N_6342);
nand U6962 (N_6962,N_6200,N_6214);
and U6963 (N_6963,N_6314,N_6221);
nor U6964 (N_6964,N_6466,N_6216);
and U6965 (N_6965,N_6486,N_6340);
xnor U6966 (N_6966,N_6011,N_6439);
xor U6967 (N_6967,N_6321,N_6014);
nor U6968 (N_6968,N_6330,N_6024);
or U6969 (N_6969,N_6383,N_6378);
or U6970 (N_6970,N_6169,N_6295);
nand U6971 (N_6971,N_6167,N_6211);
or U6972 (N_6972,N_6458,N_6349);
xnor U6973 (N_6973,N_6129,N_6048);
xor U6974 (N_6974,N_6429,N_6387);
nor U6975 (N_6975,N_6421,N_6168);
xnor U6976 (N_6976,N_6217,N_6450);
and U6977 (N_6977,N_6301,N_6267);
or U6978 (N_6978,N_6037,N_6186);
nor U6979 (N_6979,N_6050,N_6267);
nor U6980 (N_6980,N_6270,N_6289);
nor U6981 (N_6981,N_6286,N_6132);
and U6982 (N_6982,N_6475,N_6427);
nand U6983 (N_6983,N_6416,N_6386);
nor U6984 (N_6984,N_6083,N_6206);
nor U6985 (N_6985,N_6007,N_6251);
or U6986 (N_6986,N_6449,N_6099);
nor U6987 (N_6987,N_6326,N_6140);
xor U6988 (N_6988,N_6061,N_6233);
and U6989 (N_6989,N_6498,N_6308);
and U6990 (N_6990,N_6126,N_6054);
or U6991 (N_6991,N_6456,N_6443);
nand U6992 (N_6992,N_6469,N_6240);
xor U6993 (N_6993,N_6299,N_6491);
and U6994 (N_6994,N_6393,N_6209);
nand U6995 (N_6995,N_6282,N_6214);
and U6996 (N_6996,N_6463,N_6016);
xnor U6997 (N_6997,N_6462,N_6457);
and U6998 (N_6998,N_6189,N_6146);
or U6999 (N_6999,N_6036,N_6388);
nor U7000 (N_7000,N_6608,N_6607);
xnor U7001 (N_7001,N_6948,N_6742);
or U7002 (N_7002,N_6823,N_6939);
and U7003 (N_7003,N_6717,N_6578);
and U7004 (N_7004,N_6525,N_6516);
xnor U7005 (N_7005,N_6807,N_6985);
and U7006 (N_7006,N_6633,N_6621);
or U7007 (N_7007,N_6983,N_6693);
nor U7008 (N_7008,N_6880,N_6727);
nand U7009 (N_7009,N_6886,N_6547);
nand U7010 (N_7010,N_6788,N_6755);
xor U7011 (N_7011,N_6573,N_6800);
nand U7012 (N_7012,N_6836,N_6820);
nand U7013 (N_7013,N_6617,N_6912);
or U7014 (N_7014,N_6714,N_6585);
and U7015 (N_7015,N_6690,N_6883);
nor U7016 (N_7016,N_6802,N_6684);
xor U7017 (N_7017,N_6692,N_6670);
xnor U7018 (N_7018,N_6978,N_6879);
nor U7019 (N_7019,N_6555,N_6704);
xnor U7020 (N_7020,N_6591,N_6511);
nor U7021 (N_7021,N_6720,N_6686);
and U7022 (N_7022,N_6731,N_6520);
and U7023 (N_7023,N_6922,N_6631);
xor U7024 (N_7024,N_6762,N_6783);
xnor U7025 (N_7025,N_6812,N_6616);
nand U7026 (N_7026,N_6658,N_6507);
nand U7027 (N_7027,N_6865,N_6746);
nand U7028 (N_7028,N_6977,N_6989);
nor U7029 (N_7029,N_6514,N_6626);
xnor U7030 (N_7030,N_6903,N_6535);
nor U7031 (N_7031,N_6971,N_6504);
nand U7032 (N_7032,N_6743,N_6850);
nor U7033 (N_7033,N_6795,N_6840);
nand U7034 (N_7034,N_6534,N_6794);
nand U7035 (N_7035,N_6574,N_6605);
nand U7036 (N_7036,N_6868,N_6662);
nand U7037 (N_7037,N_6990,N_6554);
or U7038 (N_7038,N_6984,N_6908);
nor U7039 (N_7039,N_6716,N_6906);
xor U7040 (N_7040,N_6529,N_6766);
or U7041 (N_7041,N_6646,N_6805);
nand U7042 (N_7042,N_6775,N_6705);
nand U7043 (N_7043,N_6596,N_6570);
nor U7044 (N_7044,N_6799,N_6628);
nand U7045 (N_7045,N_6680,N_6828);
nand U7046 (N_7046,N_6907,N_6759);
nor U7047 (N_7047,N_6604,N_6881);
xnor U7048 (N_7048,N_6672,N_6556);
or U7049 (N_7049,N_6689,N_6998);
xnor U7050 (N_7050,N_6651,N_6835);
or U7051 (N_7051,N_6991,N_6910);
nor U7052 (N_7052,N_6764,N_6959);
nor U7053 (N_7053,N_6975,N_6715);
or U7054 (N_7054,N_6953,N_6933);
or U7055 (N_7055,N_6760,N_6640);
xnor U7056 (N_7056,N_6546,N_6653);
and U7057 (N_7057,N_6683,N_6569);
nand U7058 (N_7058,N_6947,N_6709);
nand U7059 (N_7059,N_6885,N_6756);
or U7060 (N_7060,N_6703,N_6864);
xor U7061 (N_7061,N_6895,N_6695);
or U7062 (N_7062,N_6815,N_6931);
nor U7063 (N_7063,N_6965,N_6994);
xnor U7064 (N_7064,N_6987,N_6801);
nand U7065 (N_7065,N_6976,N_6667);
or U7066 (N_7066,N_6675,N_6980);
or U7067 (N_7067,N_6758,N_6669);
and U7068 (N_7068,N_6521,N_6563);
nor U7069 (N_7069,N_6593,N_6635);
xnor U7070 (N_7070,N_6698,N_6612);
nand U7071 (N_7071,N_6736,N_6753);
and U7072 (N_7072,N_6747,N_6664);
xor U7073 (N_7073,N_6847,N_6866);
or U7074 (N_7074,N_6510,N_6924);
or U7075 (N_7075,N_6797,N_6825);
or U7076 (N_7076,N_6873,N_6738);
xnor U7077 (N_7077,N_6996,N_6702);
and U7078 (N_7078,N_6706,N_6560);
nor U7079 (N_7079,N_6963,N_6900);
or U7080 (N_7080,N_6919,N_6502);
or U7081 (N_7081,N_6988,N_6721);
xor U7082 (N_7082,N_6579,N_6543);
nor U7083 (N_7083,N_6995,N_6826);
nand U7084 (N_7084,N_6832,N_6875);
or U7085 (N_7085,N_6584,N_6606);
or U7086 (N_7086,N_6551,N_6614);
or U7087 (N_7087,N_6734,N_6613);
or U7088 (N_7088,N_6981,N_6598);
nor U7089 (N_7089,N_6558,N_6733);
nor U7090 (N_7090,N_6905,N_6878);
xnor U7091 (N_7091,N_6597,N_6940);
or U7092 (N_7092,N_6932,N_6539);
nor U7093 (N_7093,N_6874,N_6609);
xor U7094 (N_7094,N_6831,N_6972);
and U7095 (N_7095,N_6500,N_6629);
and U7096 (N_7096,N_6806,N_6618);
nor U7097 (N_7097,N_6517,N_6789);
or U7098 (N_7098,N_6851,N_6522);
and U7099 (N_7099,N_6557,N_6538);
nand U7100 (N_7100,N_6509,N_6857);
and U7101 (N_7101,N_6532,N_6652);
nand U7102 (N_7102,N_6942,N_6796);
xor U7103 (N_7103,N_6821,N_6561);
and U7104 (N_7104,N_6929,N_6843);
or U7105 (N_7105,N_6997,N_6819);
or U7106 (N_7106,N_6785,N_6968);
or U7107 (N_7107,N_6540,N_6632);
or U7108 (N_7108,N_6700,N_6917);
or U7109 (N_7109,N_6622,N_6610);
nor U7110 (N_7110,N_6542,N_6958);
and U7111 (N_7111,N_6877,N_6926);
and U7112 (N_7112,N_6528,N_6505);
xnor U7113 (N_7113,N_6711,N_6870);
nand U7114 (N_7114,N_6587,N_6624);
xnor U7115 (N_7115,N_6562,N_6956);
and U7116 (N_7116,N_6691,N_6888);
or U7117 (N_7117,N_6803,N_6636);
and U7118 (N_7118,N_6941,N_6519);
or U7119 (N_7119,N_6603,N_6712);
and U7120 (N_7120,N_6630,N_6623);
nor U7121 (N_7121,N_6583,N_6536);
or U7122 (N_7122,N_6688,N_6678);
or U7123 (N_7123,N_6944,N_6909);
nand U7124 (N_7124,N_6589,N_6838);
nor U7125 (N_7125,N_6523,N_6566);
or U7126 (N_7126,N_6592,N_6769);
nand U7127 (N_7127,N_6818,N_6575);
xor U7128 (N_7128,N_6642,N_6544);
and U7129 (N_7129,N_6781,N_6936);
nand U7130 (N_7130,N_6810,N_6829);
nand U7131 (N_7131,N_6656,N_6641);
or U7132 (N_7132,N_6827,N_6845);
and U7133 (N_7133,N_6920,N_6708);
or U7134 (N_7134,N_6601,N_6730);
nor U7135 (N_7135,N_6619,N_6580);
xor U7136 (N_7136,N_6595,N_6871);
and U7137 (N_7137,N_6779,N_6923);
xnor U7138 (N_7138,N_6999,N_6732);
or U7139 (N_7139,N_6729,N_6679);
or U7140 (N_7140,N_6659,N_6767);
xnor U7141 (N_7141,N_6896,N_6786);
xor U7142 (N_7142,N_6676,N_6884);
nor U7143 (N_7143,N_6841,N_6804);
and U7144 (N_7144,N_6790,N_6916);
nor U7145 (N_7145,N_6637,N_6848);
nand U7146 (N_7146,N_6665,N_6699);
nor U7147 (N_7147,N_6813,N_6735);
or U7148 (N_7148,N_6754,N_6969);
and U7149 (N_7149,N_6982,N_6643);
nor U7150 (N_7150,N_6882,N_6792);
nand U7151 (N_7151,N_6710,N_6625);
nor U7152 (N_7152,N_6954,N_6930);
nand U7153 (N_7153,N_6663,N_6780);
and U7154 (N_7154,N_6966,N_6674);
nor U7155 (N_7155,N_6979,N_6834);
and U7156 (N_7156,N_6576,N_6787);
nor U7157 (N_7157,N_6816,N_6645);
nor U7158 (N_7158,N_6824,N_6768);
nand U7159 (N_7159,N_6599,N_6899);
nor U7160 (N_7160,N_6513,N_6728);
nand U7161 (N_7161,N_6718,N_6950);
and U7162 (N_7162,N_6541,N_6553);
nand U7163 (N_7163,N_6568,N_6524);
nand U7164 (N_7164,N_6904,N_6748);
or U7165 (N_7165,N_6955,N_6697);
or U7166 (N_7166,N_6889,N_6654);
or U7167 (N_7167,N_6918,N_6952);
nor U7168 (N_7168,N_6822,N_6817);
nor U7169 (N_7169,N_6973,N_6713);
nand U7170 (N_7170,N_6921,N_6945);
nor U7171 (N_7171,N_6961,N_6724);
and U7172 (N_7172,N_6844,N_6739);
nand U7173 (N_7173,N_6894,N_6830);
xnor U7174 (N_7174,N_6696,N_6594);
and U7175 (N_7175,N_6545,N_6677);
xor U7176 (N_7176,N_6837,N_6937);
xor U7177 (N_7177,N_6668,N_6661);
xnor U7178 (N_7178,N_6914,N_6935);
or U7179 (N_7179,N_6811,N_6750);
and U7180 (N_7180,N_6639,N_6853);
nand U7181 (N_7181,N_6701,N_6681);
xnor U7182 (N_7182,N_6745,N_6620);
and U7183 (N_7183,N_6992,N_6970);
xnor U7184 (N_7184,N_6986,N_6993);
xor U7185 (N_7185,N_6778,N_6773);
and U7186 (N_7186,N_6809,N_6655);
or U7187 (N_7187,N_6862,N_6559);
nand U7188 (N_7188,N_6749,N_6531);
nor U7189 (N_7189,N_6856,N_6765);
and U7190 (N_7190,N_6564,N_6673);
and U7191 (N_7191,N_6915,N_6627);
xor U7192 (N_7192,N_6565,N_6657);
or U7193 (N_7193,N_6671,N_6590);
xnor U7194 (N_7194,N_6776,N_6549);
xor U7195 (N_7195,N_6707,N_6526);
and U7196 (N_7196,N_6648,N_6858);
xnor U7197 (N_7197,N_6571,N_6763);
and U7198 (N_7198,N_6649,N_6960);
xnor U7199 (N_7199,N_6586,N_6855);
nor U7200 (N_7200,N_6913,N_6772);
nand U7201 (N_7201,N_6860,N_6869);
xnor U7202 (N_7202,N_6761,N_6863);
and U7203 (N_7203,N_6872,N_6839);
or U7204 (N_7204,N_6518,N_6602);
nand U7205 (N_7205,N_6660,N_6615);
nor U7206 (N_7206,N_6644,N_6647);
nand U7207 (N_7207,N_6943,N_6725);
and U7208 (N_7208,N_6751,N_6737);
xor U7209 (N_7209,N_6719,N_6774);
nand U7210 (N_7210,N_6974,N_6537);
or U7211 (N_7211,N_6951,N_6687);
or U7212 (N_7212,N_6581,N_6887);
and U7213 (N_7213,N_6964,N_6611);
and U7214 (N_7214,N_6898,N_6962);
nand U7215 (N_7215,N_6876,N_6572);
and U7216 (N_7216,N_6682,N_6634);
nor U7217 (N_7217,N_6530,N_6938);
and U7218 (N_7218,N_6902,N_6770);
nand U7219 (N_7219,N_6582,N_6934);
nand U7220 (N_7220,N_6600,N_6890);
and U7221 (N_7221,N_6852,N_6503);
nand U7222 (N_7222,N_6508,N_6588);
and U7223 (N_7223,N_6650,N_6685);
xnor U7224 (N_7224,N_6548,N_6533);
nor U7225 (N_7225,N_6814,N_6784);
xnor U7226 (N_7226,N_6859,N_6793);
or U7227 (N_7227,N_6694,N_6893);
or U7228 (N_7228,N_6501,N_6897);
nor U7229 (N_7229,N_6567,N_6928);
or U7230 (N_7230,N_6757,N_6891);
and U7231 (N_7231,N_6849,N_6861);
xnor U7232 (N_7232,N_6925,N_6901);
nand U7233 (N_7233,N_6946,N_6927);
and U7234 (N_7234,N_6726,N_6957);
nor U7235 (N_7235,N_6892,N_6771);
xor U7236 (N_7236,N_6506,N_6638);
or U7237 (N_7237,N_6527,N_6744);
nand U7238 (N_7238,N_6722,N_6833);
xnor U7239 (N_7239,N_6577,N_6512);
xor U7240 (N_7240,N_6842,N_6911);
nor U7241 (N_7241,N_6967,N_6550);
nand U7242 (N_7242,N_6791,N_6741);
or U7243 (N_7243,N_6515,N_6740);
nand U7244 (N_7244,N_6949,N_6798);
or U7245 (N_7245,N_6854,N_6808);
nor U7246 (N_7246,N_6846,N_6752);
xor U7247 (N_7247,N_6782,N_6723);
nand U7248 (N_7248,N_6666,N_6867);
or U7249 (N_7249,N_6552,N_6777);
xor U7250 (N_7250,N_6853,N_6940);
or U7251 (N_7251,N_6894,N_6950);
and U7252 (N_7252,N_6514,N_6791);
nor U7253 (N_7253,N_6906,N_6882);
and U7254 (N_7254,N_6627,N_6591);
nand U7255 (N_7255,N_6741,N_6889);
or U7256 (N_7256,N_6711,N_6894);
xor U7257 (N_7257,N_6944,N_6653);
xor U7258 (N_7258,N_6794,N_6787);
nand U7259 (N_7259,N_6896,N_6996);
or U7260 (N_7260,N_6808,N_6572);
nand U7261 (N_7261,N_6783,N_6802);
xnor U7262 (N_7262,N_6673,N_6809);
nor U7263 (N_7263,N_6899,N_6775);
xnor U7264 (N_7264,N_6582,N_6592);
nand U7265 (N_7265,N_6628,N_6992);
xnor U7266 (N_7266,N_6876,N_6616);
or U7267 (N_7267,N_6805,N_6511);
nor U7268 (N_7268,N_6644,N_6957);
xor U7269 (N_7269,N_6773,N_6697);
and U7270 (N_7270,N_6782,N_6625);
nor U7271 (N_7271,N_6514,N_6854);
and U7272 (N_7272,N_6600,N_6834);
xnor U7273 (N_7273,N_6631,N_6899);
xnor U7274 (N_7274,N_6774,N_6867);
xor U7275 (N_7275,N_6929,N_6736);
and U7276 (N_7276,N_6804,N_6958);
or U7277 (N_7277,N_6718,N_6855);
and U7278 (N_7278,N_6908,N_6828);
and U7279 (N_7279,N_6581,N_6526);
xor U7280 (N_7280,N_6740,N_6630);
and U7281 (N_7281,N_6962,N_6601);
and U7282 (N_7282,N_6517,N_6771);
nand U7283 (N_7283,N_6674,N_6872);
nor U7284 (N_7284,N_6622,N_6789);
or U7285 (N_7285,N_6845,N_6640);
nand U7286 (N_7286,N_6558,N_6725);
nor U7287 (N_7287,N_6943,N_6575);
or U7288 (N_7288,N_6503,N_6557);
nand U7289 (N_7289,N_6667,N_6931);
nor U7290 (N_7290,N_6516,N_6530);
or U7291 (N_7291,N_6696,N_6925);
and U7292 (N_7292,N_6690,N_6584);
and U7293 (N_7293,N_6799,N_6841);
or U7294 (N_7294,N_6974,N_6901);
nor U7295 (N_7295,N_6640,N_6973);
nor U7296 (N_7296,N_6579,N_6801);
nor U7297 (N_7297,N_6714,N_6596);
or U7298 (N_7298,N_6755,N_6656);
xnor U7299 (N_7299,N_6627,N_6595);
nand U7300 (N_7300,N_6991,N_6856);
nand U7301 (N_7301,N_6942,N_6861);
and U7302 (N_7302,N_6651,N_6654);
xor U7303 (N_7303,N_6638,N_6784);
nand U7304 (N_7304,N_6862,N_6851);
nand U7305 (N_7305,N_6601,N_6767);
nand U7306 (N_7306,N_6644,N_6804);
nand U7307 (N_7307,N_6876,N_6991);
and U7308 (N_7308,N_6838,N_6942);
and U7309 (N_7309,N_6792,N_6764);
nor U7310 (N_7310,N_6734,N_6619);
xnor U7311 (N_7311,N_6628,N_6655);
and U7312 (N_7312,N_6685,N_6696);
nor U7313 (N_7313,N_6597,N_6672);
and U7314 (N_7314,N_6739,N_6958);
nand U7315 (N_7315,N_6631,N_6961);
nor U7316 (N_7316,N_6704,N_6988);
nor U7317 (N_7317,N_6992,N_6756);
and U7318 (N_7318,N_6761,N_6838);
nor U7319 (N_7319,N_6802,N_6509);
and U7320 (N_7320,N_6722,N_6860);
and U7321 (N_7321,N_6806,N_6778);
nor U7322 (N_7322,N_6949,N_6957);
xnor U7323 (N_7323,N_6517,N_6752);
nand U7324 (N_7324,N_6742,N_6626);
nor U7325 (N_7325,N_6870,N_6771);
or U7326 (N_7326,N_6710,N_6613);
nor U7327 (N_7327,N_6568,N_6693);
nor U7328 (N_7328,N_6848,N_6900);
or U7329 (N_7329,N_6573,N_6875);
or U7330 (N_7330,N_6862,N_6624);
xnor U7331 (N_7331,N_6865,N_6902);
and U7332 (N_7332,N_6632,N_6937);
or U7333 (N_7333,N_6971,N_6571);
xor U7334 (N_7334,N_6913,N_6709);
nor U7335 (N_7335,N_6761,N_6643);
xor U7336 (N_7336,N_6780,N_6792);
or U7337 (N_7337,N_6814,N_6654);
nor U7338 (N_7338,N_6998,N_6851);
nand U7339 (N_7339,N_6877,N_6594);
nand U7340 (N_7340,N_6730,N_6983);
xor U7341 (N_7341,N_6929,N_6762);
xnor U7342 (N_7342,N_6575,N_6897);
and U7343 (N_7343,N_6956,N_6616);
nand U7344 (N_7344,N_6652,N_6891);
or U7345 (N_7345,N_6513,N_6994);
nand U7346 (N_7346,N_6745,N_6791);
and U7347 (N_7347,N_6504,N_6634);
and U7348 (N_7348,N_6994,N_6709);
xor U7349 (N_7349,N_6760,N_6976);
and U7350 (N_7350,N_6983,N_6524);
or U7351 (N_7351,N_6566,N_6853);
nand U7352 (N_7352,N_6617,N_6708);
or U7353 (N_7353,N_6722,N_6793);
nor U7354 (N_7354,N_6705,N_6633);
nand U7355 (N_7355,N_6861,N_6581);
xor U7356 (N_7356,N_6843,N_6630);
xor U7357 (N_7357,N_6585,N_6888);
nand U7358 (N_7358,N_6688,N_6828);
nand U7359 (N_7359,N_6688,N_6738);
xor U7360 (N_7360,N_6967,N_6803);
nor U7361 (N_7361,N_6838,N_6839);
nand U7362 (N_7362,N_6919,N_6885);
nand U7363 (N_7363,N_6753,N_6735);
or U7364 (N_7364,N_6779,N_6756);
and U7365 (N_7365,N_6515,N_6974);
nor U7366 (N_7366,N_6835,N_6634);
and U7367 (N_7367,N_6878,N_6974);
nor U7368 (N_7368,N_6523,N_6770);
or U7369 (N_7369,N_6995,N_6510);
or U7370 (N_7370,N_6505,N_6828);
or U7371 (N_7371,N_6945,N_6516);
xor U7372 (N_7372,N_6882,N_6839);
nand U7373 (N_7373,N_6963,N_6669);
and U7374 (N_7374,N_6504,N_6891);
and U7375 (N_7375,N_6970,N_6643);
and U7376 (N_7376,N_6572,N_6721);
xor U7377 (N_7377,N_6706,N_6561);
or U7378 (N_7378,N_6937,N_6529);
nor U7379 (N_7379,N_6604,N_6729);
xnor U7380 (N_7380,N_6778,N_6898);
nand U7381 (N_7381,N_6793,N_6814);
nand U7382 (N_7382,N_6629,N_6797);
or U7383 (N_7383,N_6739,N_6578);
nand U7384 (N_7384,N_6912,N_6622);
nor U7385 (N_7385,N_6827,N_6957);
nor U7386 (N_7386,N_6707,N_6560);
nor U7387 (N_7387,N_6980,N_6777);
nor U7388 (N_7388,N_6530,N_6756);
nor U7389 (N_7389,N_6900,N_6920);
and U7390 (N_7390,N_6836,N_6958);
nor U7391 (N_7391,N_6766,N_6581);
and U7392 (N_7392,N_6561,N_6583);
xnor U7393 (N_7393,N_6568,N_6517);
xor U7394 (N_7394,N_6978,N_6822);
or U7395 (N_7395,N_6667,N_6801);
or U7396 (N_7396,N_6689,N_6667);
nor U7397 (N_7397,N_6953,N_6915);
xnor U7398 (N_7398,N_6872,N_6978);
nand U7399 (N_7399,N_6566,N_6793);
nor U7400 (N_7400,N_6579,N_6838);
or U7401 (N_7401,N_6540,N_6840);
xor U7402 (N_7402,N_6676,N_6647);
or U7403 (N_7403,N_6644,N_6623);
xor U7404 (N_7404,N_6866,N_6677);
or U7405 (N_7405,N_6911,N_6938);
and U7406 (N_7406,N_6879,N_6891);
nand U7407 (N_7407,N_6767,N_6650);
nand U7408 (N_7408,N_6888,N_6986);
or U7409 (N_7409,N_6801,N_6543);
or U7410 (N_7410,N_6654,N_6516);
or U7411 (N_7411,N_6620,N_6879);
nand U7412 (N_7412,N_6585,N_6843);
nor U7413 (N_7413,N_6671,N_6697);
nand U7414 (N_7414,N_6597,N_6945);
and U7415 (N_7415,N_6978,N_6930);
and U7416 (N_7416,N_6703,N_6866);
xor U7417 (N_7417,N_6946,N_6766);
xor U7418 (N_7418,N_6728,N_6772);
nand U7419 (N_7419,N_6571,N_6980);
or U7420 (N_7420,N_6807,N_6814);
nand U7421 (N_7421,N_6552,N_6676);
nor U7422 (N_7422,N_6929,N_6636);
and U7423 (N_7423,N_6512,N_6515);
nand U7424 (N_7424,N_6770,N_6841);
or U7425 (N_7425,N_6919,N_6746);
nand U7426 (N_7426,N_6711,N_6579);
nor U7427 (N_7427,N_6740,N_6550);
and U7428 (N_7428,N_6787,N_6696);
or U7429 (N_7429,N_6660,N_6682);
nor U7430 (N_7430,N_6777,N_6565);
and U7431 (N_7431,N_6876,N_6878);
and U7432 (N_7432,N_6942,N_6652);
nor U7433 (N_7433,N_6714,N_6842);
and U7434 (N_7434,N_6870,N_6506);
xor U7435 (N_7435,N_6850,N_6800);
or U7436 (N_7436,N_6589,N_6971);
and U7437 (N_7437,N_6694,N_6728);
xnor U7438 (N_7438,N_6829,N_6867);
and U7439 (N_7439,N_6937,N_6528);
and U7440 (N_7440,N_6737,N_6565);
xnor U7441 (N_7441,N_6535,N_6752);
nor U7442 (N_7442,N_6697,N_6547);
nand U7443 (N_7443,N_6909,N_6990);
and U7444 (N_7444,N_6831,N_6893);
and U7445 (N_7445,N_6815,N_6625);
or U7446 (N_7446,N_6730,N_6700);
xor U7447 (N_7447,N_6933,N_6763);
or U7448 (N_7448,N_6991,N_6828);
or U7449 (N_7449,N_6719,N_6781);
and U7450 (N_7450,N_6975,N_6520);
and U7451 (N_7451,N_6907,N_6606);
or U7452 (N_7452,N_6942,N_6633);
and U7453 (N_7453,N_6610,N_6656);
or U7454 (N_7454,N_6574,N_6630);
and U7455 (N_7455,N_6650,N_6754);
and U7456 (N_7456,N_6841,N_6854);
nor U7457 (N_7457,N_6644,N_6616);
and U7458 (N_7458,N_6954,N_6843);
nor U7459 (N_7459,N_6557,N_6945);
xor U7460 (N_7460,N_6739,N_6670);
or U7461 (N_7461,N_6661,N_6635);
xor U7462 (N_7462,N_6687,N_6800);
or U7463 (N_7463,N_6870,N_6660);
and U7464 (N_7464,N_6976,N_6663);
or U7465 (N_7465,N_6506,N_6953);
nor U7466 (N_7466,N_6606,N_6925);
and U7467 (N_7467,N_6714,N_6649);
and U7468 (N_7468,N_6976,N_6500);
or U7469 (N_7469,N_6996,N_6821);
nor U7470 (N_7470,N_6529,N_6931);
nor U7471 (N_7471,N_6896,N_6738);
nand U7472 (N_7472,N_6902,N_6718);
or U7473 (N_7473,N_6976,N_6594);
nor U7474 (N_7474,N_6831,N_6881);
nand U7475 (N_7475,N_6903,N_6682);
nor U7476 (N_7476,N_6990,N_6627);
nor U7477 (N_7477,N_6955,N_6755);
and U7478 (N_7478,N_6905,N_6627);
or U7479 (N_7479,N_6754,N_6848);
and U7480 (N_7480,N_6553,N_6625);
or U7481 (N_7481,N_6750,N_6931);
or U7482 (N_7482,N_6553,N_6802);
and U7483 (N_7483,N_6618,N_6507);
xor U7484 (N_7484,N_6830,N_6655);
nand U7485 (N_7485,N_6782,N_6758);
xnor U7486 (N_7486,N_6885,N_6915);
or U7487 (N_7487,N_6974,N_6875);
or U7488 (N_7488,N_6502,N_6525);
nand U7489 (N_7489,N_6790,N_6789);
nor U7490 (N_7490,N_6744,N_6542);
nor U7491 (N_7491,N_6927,N_6907);
and U7492 (N_7492,N_6625,N_6803);
and U7493 (N_7493,N_6697,N_6543);
or U7494 (N_7494,N_6963,N_6789);
xnor U7495 (N_7495,N_6812,N_6893);
xnor U7496 (N_7496,N_6777,N_6896);
and U7497 (N_7497,N_6680,N_6866);
and U7498 (N_7498,N_6543,N_6753);
or U7499 (N_7499,N_6997,N_6823);
and U7500 (N_7500,N_7417,N_7367);
nand U7501 (N_7501,N_7499,N_7168);
nor U7502 (N_7502,N_7223,N_7271);
xor U7503 (N_7503,N_7146,N_7306);
nand U7504 (N_7504,N_7218,N_7401);
nand U7505 (N_7505,N_7495,N_7066);
nand U7506 (N_7506,N_7015,N_7154);
nor U7507 (N_7507,N_7174,N_7031);
xnor U7508 (N_7508,N_7055,N_7228);
nor U7509 (N_7509,N_7370,N_7105);
nor U7510 (N_7510,N_7485,N_7314);
nor U7511 (N_7511,N_7175,N_7237);
and U7512 (N_7512,N_7402,N_7321);
or U7513 (N_7513,N_7336,N_7125);
nor U7514 (N_7514,N_7246,N_7091);
xnor U7515 (N_7515,N_7042,N_7085);
or U7516 (N_7516,N_7061,N_7384);
nand U7517 (N_7517,N_7007,N_7373);
nand U7518 (N_7518,N_7347,N_7473);
nor U7519 (N_7519,N_7358,N_7132);
and U7520 (N_7520,N_7150,N_7455);
and U7521 (N_7521,N_7123,N_7117);
nand U7522 (N_7522,N_7204,N_7101);
and U7523 (N_7523,N_7012,N_7129);
or U7524 (N_7524,N_7393,N_7440);
xor U7525 (N_7525,N_7106,N_7379);
nor U7526 (N_7526,N_7395,N_7279);
and U7527 (N_7527,N_7059,N_7380);
and U7528 (N_7528,N_7263,N_7090);
nor U7529 (N_7529,N_7067,N_7002);
nor U7530 (N_7530,N_7303,N_7397);
and U7531 (N_7531,N_7369,N_7310);
xor U7532 (N_7532,N_7199,N_7104);
nand U7533 (N_7533,N_7164,N_7259);
and U7534 (N_7534,N_7392,N_7311);
nand U7535 (N_7535,N_7028,N_7122);
or U7536 (N_7536,N_7309,N_7365);
xnor U7537 (N_7537,N_7188,N_7006);
or U7538 (N_7538,N_7346,N_7148);
and U7539 (N_7539,N_7343,N_7337);
or U7540 (N_7540,N_7060,N_7348);
nor U7541 (N_7541,N_7222,N_7029);
nand U7542 (N_7542,N_7131,N_7464);
nor U7543 (N_7543,N_7269,N_7069);
or U7544 (N_7544,N_7338,N_7377);
or U7545 (N_7545,N_7144,N_7004);
xnor U7546 (N_7546,N_7082,N_7041);
nor U7547 (N_7547,N_7458,N_7272);
and U7548 (N_7548,N_7229,N_7138);
or U7549 (N_7549,N_7344,N_7315);
nor U7550 (N_7550,N_7200,N_7330);
or U7551 (N_7551,N_7077,N_7439);
xnor U7552 (N_7552,N_7316,N_7239);
nor U7553 (N_7553,N_7176,N_7366);
xor U7554 (N_7554,N_7327,N_7189);
xor U7555 (N_7555,N_7307,N_7065);
nand U7556 (N_7556,N_7203,N_7036);
xnor U7557 (N_7557,N_7385,N_7430);
and U7558 (N_7558,N_7312,N_7224);
xor U7559 (N_7559,N_7488,N_7213);
nor U7560 (N_7560,N_7420,N_7083);
or U7561 (N_7561,N_7103,N_7320);
and U7562 (N_7562,N_7045,N_7340);
nor U7563 (N_7563,N_7319,N_7406);
and U7564 (N_7564,N_7288,N_7086);
nand U7565 (N_7565,N_7474,N_7447);
and U7566 (N_7566,N_7167,N_7301);
nor U7567 (N_7567,N_7257,N_7054);
xnor U7568 (N_7568,N_7182,N_7496);
xor U7569 (N_7569,N_7266,N_7451);
or U7570 (N_7570,N_7362,N_7022);
nor U7571 (N_7571,N_7360,N_7375);
xor U7572 (N_7572,N_7357,N_7179);
nand U7573 (N_7573,N_7049,N_7116);
nand U7574 (N_7574,N_7145,N_7481);
or U7575 (N_7575,N_7489,N_7412);
xor U7576 (N_7576,N_7039,N_7151);
and U7577 (N_7577,N_7172,N_7419);
nand U7578 (N_7578,N_7326,N_7147);
nand U7579 (N_7579,N_7113,N_7165);
nand U7580 (N_7580,N_7097,N_7410);
nand U7581 (N_7581,N_7442,N_7256);
or U7582 (N_7582,N_7003,N_7159);
and U7583 (N_7583,N_7134,N_7483);
or U7584 (N_7584,N_7026,N_7497);
nand U7585 (N_7585,N_7196,N_7099);
or U7586 (N_7586,N_7100,N_7011);
or U7587 (N_7587,N_7403,N_7355);
nand U7588 (N_7588,N_7274,N_7124);
and U7589 (N_7589,N_7471,N_7453);
nor U7590 (N_7590,N_7056,N_7209);
xnor U7591 (N_7591,N_7277,N_7480);
or U7592 (N_7592,N_7490,N_7191);
xnor U7593 (N_7593,N_7034,N_7032);
nand U7594 (N_7594,N_7305,N_7241);
or U7595 (N_7595,N_7023,N_7308);
xnor U7596 (N_7596,N_7024,N_7426);
nor U7597 (N_7597,N_7160,N_7155);
or U7598 (N_7598,N_7247,N_7329);
xnor U7599 (N_7599,N_7267,N_7292);
xnor U7600 (N_7600,N_7166,N_7244);
xor U7601 (N_7601,N_7432,N_7405);
nand U7602 (N_7602,N_7341,N_7467);
nand U7603 (N_7603,N_7363,N_7391);
xor U7604 (N_7604,N_7071,N_7300);
nand U7605 (N_7605,N_7240,N_7163);
or U7606 (N_7606,N_7018,N_7364);
xor U7607 (N_7607,N_7141,N_7293);
or U7608 (N_7608,N_7486,N_7394);
or U7609 (N_7609,N_7411,N_7291);
nor U7610 (N_7610,N_7462,N_7177);
nand U7611 (N_7611,N_7051,N_7111);
or U7612 (N_7612,N_7334,N_7457);
xor U7613 (N_7613,N_7479,N_7073);
xor U7614 (N_7614,N_7020,N_7170);
xor U7615 (N_7615,N_7361,N_7252);
xnor U7616 (N_7616,N_7043,N_7242);
or U7617 (N_7617,N_7408,N_7470);
and U7618 (N_7618,N_7156,N_7050);
xor U7619 (N_7619,N_7038,N_7378);
xnor U7620 (N_7620,N_7452,N_7202);
and U7621 (N_7621,N_7494,N_7121);
and U7622 (N_7622,N_7478,N_7416);
nor U7623 (N_7623,N_7492,N_7227);
and U7624 (N_7624,N_7047,N_7450);
or U7625 (N_7625,N_7352,N_7044);
and U7626 (N_7626,N_7468,N_7389);
or U7627 (N_7627,N_7404,N_7013);
or U7628 (N_7628,N_7008,N_7372);
or U7629 (N_7629,N_7214,N_7424);
nor U7630 (N_7630,N_7217,N_7413);
or U7631 (N_7631,N_7040,N_7078);
and U7632 (N_7632,N_7057,N_7110);
nand U7633 (N_7633,N_7205,N_7254);
nor U7634 (N_7634,N_7445,N_7118);
xor U7635 (N_7635,N_7048,N_7127);
and U7636 (N_7636,N_7409,N_7251);
nand U7637 (N_7637,N_7287,N_7114);
and U7638 (N_7638,N_7025,N_7181);
nor U7639 (N_7639,N_7475,N_7349);
xor U7640 (N_7640,N_7456,N_7030);
and U7641 (N_7641,N_7192,N_7318);
nand U7642 (N_7642,N_7286,N_7368);
nor U7643 (N_7643,N_7425,N_7046);
nand U7644 (N_7644,N_7328,N_7339);
and U7645 (N_7645,N_7037,N_7422);
or U7646 (N_7646,N_7284,N_7211);
nor U7647 (N_7647,N_7295,N_7035);
nand U7648 (N_7648,N_7215,N_7236);
xor U7649 (N_7649,N_7137,N_7415);
xor U7650 (N_7650,N_7275,N_7102);
nand U7651 (N_7651,N_7076,N_7108);
and U7652 (N_7652,N_7437,N_7444);
xnor U7653 (N_7653,N_7281,N_7493);
and U7654 (N_7654,N_7245,N_7075);
nor U7655 (N_7655,N_7201,N_7084);
nor U7656 (N_7656,N_7414,N_7356);
and U7657 (N_7657,N_7472,N_7407);
or U7658 (N_7658,N_7443,N_7289);
and U7659 (N_7659,N_7427,N_7072);
nand U7660 (N_7660,N_7477,N_7353);
and U7661 (N_7661,N_7198,N_7001);
and U7662 (N_7662,N_7280,N_7098);
nand U7663 (N_7663,N_7441,N_7207);
and U7664 (N_7664,N_7232,N_7431);
xnor U7665 (N_7665,N_7359,N_7482);
or U7666 (N_7666,N_7139,N_7476);
nor U7667 (N_7667,N_7152,N_7469);
or U7668 (N_7668,N_7178,N_7382);
nor U7669 (N_7669,N_7171,N_7087);
nor U7670 (N_7670,N_7064,N_7019);
nor U7671 (N_7671,N_7354,N_7323);
and U7672 (N_7672,N_7221,N_7079);
xnor U7673 (N_7673,N_7313,N_7350);
nor U7674 (N_7674,N_7225,N_7268);
and U7675 (N_7675,N_7063,N_7283);
and U7676 (N_7676,N_7017,N_7193);
nor U7677 (N_7677,N_7088,N_7262);
nand U7678 (N_7678,N_7235,N_7345);
and U7679 (N_7679,N_7081,N_7317);
nand U7680 (N_7680,N_7460,N_7115);
xnor U7681 (N_7681,N_7226,N_7058);
nand U7682 (N_7682,N_7302,N_7094);
nor U7683 (N_7683,N_7095,N_7351);
nor U7684 (N_7684,N_7398,N_7248);
xnor U7685 (N_7685,N_7261,N_7264);
nand U7686 (N_7686,N_7187,N_7454);
or U7687 (N_7687,N_7169,N_7142);
xnor U7688 (N_7688,N_7273,N_7461);
nand U7689 (N_7689,N_7183,N_7296);
nor U7690 (N_7690,N_7068,N_7119);
nand U7691 (N_7691,N_7333,N_7190);
nand U7692 (N_7692,N_7230,N_7208);
nand U7693 (N_7693,N_7325,N_7487);
xor U7694 (N_7694,N_7297,N_7184);
and U7695 (N_7695,N_7285,N_7276);
and U7696 (N_7696,N_7396,N_7161);
nand U7697 (N_7697,N_7436,N_7429);
nand U7698 (N_7698,N_7173,N_7428);
nand U7699 (N_7699,N_7096,N_7206);
or U7700 (N_7700,N_7324,N_7386);
nand U7701 (N_7701,N_7219,N_7290);
or U7702 (N_7702,N_7158,N_7112);
nand U7703 (N_7703,N_7162,N_7120);
xor U7704 (N_7704,N_7298,N_7136);
and U7705 (N_7705,N_7400,N_7143);
xor U7706 (N_7706,N_7130,N_7089);
and U7707 (N_7707,N_7265,N_7423);
or U7708 (N_7708,N_7238,N_7135);
nor U7709 (N_7709,N_7128,N_7016);
nand U7710 (N_7710,N_7234,N_7080);
or U7711 (N_7711,N_7126,N_7216);
nand U7712 (N_7712,N_7140,N_7459);
nand U7713 (N_7713,N_7438,N_7399);
nand U7714 (N_7714,N_7435,N_7033);
nor U7715 (N_7715,N_7231,N_7342);
or U7716 (N_7716,N_7374,N_7304);
xor U7717 (N_7717,N_7092,N_7133);
nor U7718 (N_7718,N_7249,N_7433);
nand U7719 (N_7719,N_7331,N_7010);
and U7720 (N_7720,N_7498,N_7255);
nand U7721 (N_7721,N_7278,N_7027);
xnor U7722 (N_7722,N_7322,N_7212);
and U7723 (N_7723,N_7463,N_7009);
and U7724 (N_7724,N_7093,N_7000);
nor U7725 (N_7725,N_7109,N_7258);
and U7726 (N_7726,N_7074,N_7107);
xnor U7727 (N_7727,N_7388,N_7465);
xnor U7728 (N_7728,N_7185,N_7186);
nor U7729 (N_7729,N_7197,N_7053);
or U7730 (N_7730,N_7421,N_7390);
or U7731 (N_7731,N_7335,N_7195);
or U7732 (N_7732,N_7233,N_7194);
xnor U7733 (N_7733,N_7270,N_7243);
and U7734 (N_7734,N_7014,N_7449);
xor U7735 (N_7735,N_7376,N_7332);
nand U7736 (N_7736,N_7149,N_7070);
nand U7737 (N_7737,N_7299,N_7253);
and U7738 (N_7738,N_7021,N_7383);
and U7739 (N_7739,N_7371,N_7157);
nor U7740 (N_7740,N_7250,N_7220);
nand U7741 (N_7741,N_7294,N_7484);
and U7742 (N_7742,N_7260,N_7153);
and U7743 (N_7743,N_7446,N_7052);
xor U7744 (N_7744,N_7062,N_7387);
or U7745 (N_7745,N_7381,N_7491);
and U7746 (N_7746,N_7005,N_7210);
and U7747 (N_7747,N_7180,N_7434);
xor U7748 (N_7748,N_7418,N_7282);
or U7749 (N_7749,N_7448,N_7466);
xor U7750 (N_7750,N_7153,N_7048);
nand U7751 (N_7751,N_7350,N_7090);
and U7752 (N_7752,N_7387,N_7002);
nor U7753 (N_7753,N_7304,N_7473);
nand U7754 (N_7754,N_7127,N_7111);
nor U7755 (N_7755,N_7042,N_7391);
nand U7756 (N_7756,N_7352,N_7405);
and U7757 (N_7757,N_7417,N_7318);
xnor U7758 (N_7758,N_7467,N_7364);
nand U7759 (N_7759,N_7189,N_7289);
or U7760 (N_7760,N_7044,N_7371);
xor U7761 (N_7761,N_7248,N_7080);
and U7762 (N_7762,N_7330,N_7244);
nor U7763 (N_7763,N_7371,N_7251);
and U7764 (N_7764,N_7050,N_7425);
nor U7765 (N_7765,N_7478,N_7127);
nand U7766 (N_7766,N_7135,N_7170);
nor U7767 (N_7767,N_7370,N_7234);
and U7768 (N_7768,N_7005,N_7089);
or U7769 (N_7769,N_7372,N_7336);
and U7770 (N_7770,N_7206,N_7440);
nor U7771 (N_7771,N_7308,N_7328);
nand U7772 (N_7772,N_7334,N_7016);
or U7773 (N_7773,N_7384,N_7360);
nor U7774 (N_7774,N_7132,N_7265);
nor U7775 (N_7775,N_7271,N_7292);
or U7776 (N_7776,N_7278,N_7133);
or U7777 (N_7777,N_7338,N_7182);
xnor U7778 (N_7778,N_7309,N_7092);
xor U7779 (N_7779,N_7018,N_7059);
nor U7780 (N_7780,N_7238,N_7436);
nor U7781 (N_7781,N_7052,N_7346);
nor U7782 (N_7782,N_7489,N_7245);
or U7783 (N_7783,N_7156,N_7161);
nand U7784 (N_7784,N_7368,N_7042);
or U7785 (N_7785,N_7310,N_7300);
xnor U7786 (N_7786,N_7418,N_7132);
or U7787 (N_7787,N_7275,N_7094);
nand U7788 (N_7788,N_7091,N_7457);
and U7789 (N_7789,N_7377,N_7374);
xor U7790 (N_7790,N_7135,N_7071);
xor U7791 (N_7791,N_7136,N_7434);
and U7792 (N_7792,N_7032,N_7339);
nor U7793 (N_7793,N_7419,N_7491);
and U7794 (N_7794,N_7156,N_7357);
nor U7795 (N_7795,N_7484,N_7192);
and U7796 (N_7796,N_7061,N_7211);
nor U7797 (N_7797,N_7031,N_7317);
xor U7798 (N_7798,N_7170,N_7205);
and U7799 (N_7799,N_7426,N_7329);
xnor U7800 (N_7800,N_7376,N_7381);
xor U7801 (N_7801,N_7167,N_7492);
and U7802 (N_7802,N_7403,N_7085);
nor U7803 (N_7803,N_7140,N_7069);
nor U7804 (N_7804,N_7214,N_7148);
or U7805 (N_7805,N_7157,N_7131);
and U7806 (N_7806,N_7470,N_7253);
nor U7807 (N_7807,N_7127,N_7370);
or U7808 (N_7808,N_7234,N_7359);
nor U7809 (N_7809,N_7456,N_7261);
nor U7810 (N_7810,N_7478,N_7293);
nor U7811 (N_7811,N_7477,N_7251);
or U7812 (N_7812,N_7460,N_7282);
nand U7813 (N_7813,N_7223,N_7478);
nand U7814 (N_7814,N_7064,N_7456);
xor U7815 (N_7815,N_7247,N_7347);
nor U7816 (N_7816,N_7489,N_7295);
xor U7817 (N_7817,N_7011,N_7380);
nor U7818 (N_7818,N_7336,N_7090);
nor U7819 (N_7819,N_7403,N_7385);
or U7820 (N_7820,N_7064,N_7281);
nor U7821 (N_7821,N_7191,N_7185);
or U7822 (N_7822,N_7440,N_7369);
nand U7823 (N_7823,N_7189,N_7404);
nand U7824 (N_7824,N_7024,N_7481);
and U7825 (N_7825,N_7150,N_7385);
and U7826 (N_7826,N_7278,N_7404);
nand U7827 (N_7827,N_7198,N_7086);
or U7828 (N_7828,N_7136,N_7132);
or U7829 (N_7829,N_7310,N_7246);
and U7830 (N_7830,N_7188,N_7061);
nand U7831 (N_7831,N_7274,N_7452);
and U7832 (N_7832,N_7207,N_7123);
or U7833 (N_7833,N_7453,N_7062);
and U7834 (N_7834,N_7482,N_7216);
xnor U7835 (N_7835,N_7324,N_7140);
nand U7836 (N_7836,N_7300,N_7374);
or U7837 (N_7837,N_7068,N_7396);
xor U7838 (N_7838,N_7237,N_7025);
and U7839 (N_7839,N_7220,N_7054);
nor U7840 (N_7840,N_7455,N_7047);
nand U7841 (N_7841,N_7057,N_7174);
nand U7842 (N_7842,N_7185,N_7131);
xor U7843 (N_7843,N_7445,N_7468);
xnor U7844 (N_7844,N_7332,N_7028);
nor U7845 (N_7845,N_7361,N_7475);
and U7846 (N_7846,N_7078,N_7202);
xor U7847 (N_7847,N_7426,N_7302);
nor U7848 (N_7848,N_7120,N_7410);
nor U7849 (N_7849,N_7242,N_7333);
nor U7850 (N_7850,N_7498,N_7034);
and U7851 (N_7851,N_7029,N_7053);
nand U7852 (N_7852,N_7231,N_7034);
nor U7853 (N_7853,N_7043,N_7181);
nand U7854 (N_7854,N_7231,N_7463);
nand U7855 (N_7855,N_7245,N_7242);
xnor U7856 (N_7856,N_7252,N_7071);
xor U7857 (N_7857,N_7085,N_7051);
nor U7858 (N_7858,N_7028,N_7069);
and U7859 (N_7859,N_7276,N_7144);
xor U7860 (N_7860,N_7499,N_7171);
nor U7861 (N_7861,N_7212,N_7431);
or U7862 (N_7862,N_7024,N_7325);
nor U7863 (N_7863,N_7371,N_7263);
nand U7864 (N_7864,N_7017,N_7437);
or U7865 (N_7865,N_7147,N_7103);
nand U7866 (N_7866,N_7167,N_7024);
or U7867 (N_7867,N_7124,N_7097);
and U7868 (N_7868,N_7302,N_7448);
nor U7869 (N_7869,N_7315,N_7380);
or U7870 (N_7870,N_7346,N_7281);
nor U7871 (N_7871,N_7316,N_7066);
nor U7872 (N_7872,N_7324,N_7183);
nand U7873 (N_7873,N_7358,N_7392);
and U7874 (N_7874,N_7288,N_7461);
nand U7875 (N_7875,N_7104,N_7055);
xnor U7876 (N_7876,N_7290,N_7176);
and U7877 (N_7877,N_7140,N_7427);
nand U7878 (N_7878,N_7445,N_7295);
nor U7879 (N_7879,N_7363,N_7360);
nor U7880 (N_7880,N_7242,N_7236);
or U7881 (N_7881,N_7345,N_7479);
or U7882 (N_7882,N_7233,N_7036);
nand U7883 (N_7883,N_7203,N_7426);
and U7884 (N_7884,N_7046,N_7453);
nand U7885 (N_7885,N_7224,N_7483);
nand U7886 (N_7886,N_7168,N_7295);
or U7887 (N_7887,N_7278,N_7142);
nor U7888 (N_7888,N_7443,N_7466);
nor U7889 (N_7889,N_7323,N_7083);
and U7890 (N_7890,N_7166,N_7374);
nor U7891 (N_7891,N_7059,N_7251);
xnor U7892 (N_7892,N_7006,N_7028);
or U7893 (N_7893,N_7067,N_7474);
or U7894 (N_7894,N_7129,N_7103);
nor U7895 (N_7895,N_7428,N_7185);
and U7896 (N_7896,N_7317,N_7197);
and U7897 (N_7897,N_7197,N_7163);
nand U7898 (N_7898,N_7140,N_7251);
or U7899 (N_7899,N_7241,N_7490);
and U7900 (N_7900,N_7189,N_7117);
and U7901 (N_7901,N_7290,N_7223);
and U7902 (N_7902,N_7200,N_7122);
nand U7903 (N_7903,N_7077,N_7363);
nor U7904 (N_7904,N_7446,N_7347);
nor U7905 (N_7905,N_7231,N_7209);
xnor U7906 (N_7906,N_7461,N_7095);
nand U7907 (N_7907,N_7064,N_7373);
xnor U7908 (N_7908,N_7227,N_7447);
or U7909 (N_7909,N_7138,N_7052);
or U7910 (N_7910,N_7308,N_7276);
or U7911 (N_7911,N_7252,N_7374);
xnor U7912 (N_7912,N_7304,N_7168);
and U7913 (N_7913,N_7058,N_7248);
nor U7914 (N_7914,N_7290,N_7433);
nand U7915 (N_7915,N_7371,N_7328);
or U7916 (N_7916,N_7443,N_7100);
nand U7917 (N_7917,N_7170,N_7452);
nor U7918 (N_7918,N_7215,N_7199);
or U7919 (N_7919,N_7171,N_7465);
nor U7920 (N_7920,N_7161,N_7114);
and U7921 (N_7921,N_7218,N_7134);
and U7922 (N_7922,N_7213,N_7010);
and U7923 (N_7923,N_7457,N_7392);
or U7924 (N_7924,N_7448,N_7250);
or U7925 (N_7925,N_7295,N_7072);
nor U7926 (N_7926,N_7099,N_7407);
and U7927 (N_7927,N_7035,N_7189);
nor U7928 (N_7928,N_7353,N_7499);
and U7929 (N_7929,N_7490,N_7359);
nor U7930 (N_7930,N_7326,N_7127);
nor U7931 (N_7931,N_7028,N_7337);
and U7932 (N_7932,N_7140,N_7469);
or U7933 (N_7933,N_7274,N_7276);
and U7934 (N_7934,N_7135,N_7464);
nor U7935 (N_7935,N_7183,N_7138);
and U7936 (N_7936,N_7341,N_7090);
and U7937 (N_7937,N_7481,N_7000);
and U7938 (N_7938,N_7207,N_7474);
or U7939 (N_7939,N_7044,N_7244);
and U7940 (N_7940,N_7203,N_7018);
and U7941 (N_7941,N_7326,N_7496);
and U7942 (N_7942,N_7318,N_7041);
xor U7943 (N_7943,N_7112,N_7006);
nand U7944 (N_7944,N_7352,N_7211);
xnor U7945 (N_7945,N_7344,N_7356);
and U7946 (N_7946,N_7423,N_7052);
and U7947 (N_7947,N_7192,N_7479);
nand U7948 (N_7948,N_7184,N_7300);
nor U7949 (N_7949,N_7447,N_7036);
nor U7950 (N_7950,N_7423,N_7454);
nand U7951 (N_7951,N_7382,N_7268);
and U7952 (N_7952,N_7051,N_7028);
xnor U7953 (N_7953,N_7354,N_7357);
xnor U7954 (N_7954,N_7275,N_7254);
or U7955 (N_7955,N_7249,N_7451);
nand U7956 (N_7956,N_7398,N_7343);
and U7957 (N_7957,N_7202,N_7499);
or U7958 (N_7958,N_7484,N_7073);
xor U7959 (N_7959,N_7236,N_7087);
nand U7960 (N_7960,N_7156,N_7141);
xnor U7961 (N_7961,N_7168,N_7037);
nor U7962 (N_7962,N_7354,N_7099);
xor U7963 (N_7963,N_7081,N_7025);
and U7964 (N_7964,N_7286,N_7140);
nor U7965 (N_7965,N_7109,N_7041);
nand U7966 (N_7966,N_7215,N_7443);
nand U7967 (N_7967,N_7101,N_7307);
and U7968 (N_7968,N_7423,N_7453);
or U7969 (N_7969,N_7452,N_7034);
xor U7970 (N_7970,N_7169,N_7161);
xnor U7971 (N_7971,N_7032,N_7273);
and U7972 (N_7972,N_7432,N_7426);
xor U7973 (N_7973,N_7278,N_7410);
nor U7974 (N_7974,N_7080,N_7496);
nor U7975 (N_7975,N_7386,N_7082);
or U7976 (N_7976,N_7467,N_7047);
or U7977 (N_7977,N_7473,N_7010);
nand U7978 (N_7978,N_7411,N_7043);
and U7979 (N_7979,N_7391,N_7347);
xor U7980 (N_7980,N_7228,N_7417);
nor U7981 (N_7981,N_7058,N_7016);
nor U7982 (N_7982,N_7150,N_7099);
nand U7983 (N_7983,N_7035,N_7044);
and U7984 (N_7984,N_7339,N_7340);
nand U7985 (N_7985,N_7455,N_7435);
nand U7986 (N_7986,N_7130,N_7402);
xnor U7987 (N_7987,N_7367,N_7326);
xor U7988 (N_7988,N_7340,N_7352);
nor U7989 (N_7989,N_7236,N_7300);
and U7990 (N_7990,N_7280,N_7302);
and U7991 (N_7991,N_7315,N_7166);
or U7992 (N_7992,N_7033,N_7101);
xnor U7993 (N_7993,N_7227,N_7498);
nand U7994 (N_7994,N_7253,N_7021);
or U7995 (N_7995,N_7428,N_7424);
xnor U7996 (N_7996,N_7120,N_7239);
or U7997 (N_7997,N_7343,N_7182);
and U7998 (N_7998,N_7432,N_7253);
nor U7999 (N_7999,N_7108,N_7398);
nor U8000 (N_8000,N_7871,N_7914);
nor U8001 (N_8001,N_7899,N_7893);
and U8002 (N_8002,N_7793,N_7586);
and U8003 (N_8003,N_7666,N_7556);
nand U8004 (N_8004,N_7768,N_7579);
nand U8005 (N_8005,N_7534,N_7938);
and U8006 (N_8006,N_7807,N_7997);
and U8007 (N_8007,N_7826,N_7640);
or U8008 (N_8008,N_7731,N_7702);
nor U8009 (N_8009,N_7798,N_7719);
xor U8010 (N_8010,N_7708,N_7848);
nand U8011 (N_8011,N_7890,N_7921);
nand U8012 (N_8012,N_7979,N_7663);
or U8013 (N_8013,N_7673,N_7897);
and U8014 (N_8014,N_7757,N_7846);
nand U8015 (N_8015,N_7932,N_7632);
nor U8016 (N_8016,N_7576,N_7670);
nand U8017 (N_8017,N_7995,N_7954);
or U8018 (N_8018,N_7736,N_7989);
nor U8019 (N_8019,N_7644,N_7805);
or U8020 (N_8020,N_7516,N_7974);
and U8021 (N_8021,N_7955,N_7896);
nor U8022 (N_8022,N_7623,N_7967);
xor U8023 (N_8023,N_7841,N_7711);
or U8024 (N_8024,N_7922,N_7513);
and U8025 (N_8025,N_7924,N_7966);
xnor U8026 (N_8026,N_7879,N_7747);
xnor U8027 (N_8027,N_7937,N_7642);
xor U8028 (N_8028,N_7951,N_7873);
or U8029 (N_8029,N_7574,N_7754);
xnor U8030 (N_8030,N_7880,N_7520);
or U8031 (N_8031,N_7615,N_7972);
or U8032 (N_8032,N_7588,N_7506);
nand U8033 (N_8033,N_7943,N_7699);
nand U8034 (N_8034,N_7996,N_7763);
or U8035 (N_8035,N_7847,N_7878);
xor U8036 (N_8036,N_7650,N_7696);
and U8037 (N_8037,N_7869,N_7787);
xnor U8038 (N_8038,N_7664,N_7915);
nor U8039 (N_8039,N_7529,N_7705);
nor U8040 (N_8040,N_7601,N_7949);
and U8041 (N_8041,N_7849,N_7602);
nor U8042 (N_8042,N_7964,N_7544);
or U8043 (N_8043,N_7882,N_7976);
nand U8044 (N_8044,N_7629,N_7676);
nand U8045 (N_8045,N_7850,N_7773);
nand U8046 (N_8046,N_7660,N_7678);
nor U8047 (N_8047,N_7761,N_7988);
nand U8048 (N_8048,N_7825,N_7746);
and U8049 (N_8049,N_7780,N_7679);
nor U8050 (N_8050,N_7628,N_7695);
and U8051 (N_8051,N_7947,N_7818);
nor U8052 (N_8052,N_7504,N_7712);
and U8053 (N_8053,N_7889,N_7740);
or U8054 (N_8054,N_7521,N_7620);
xor U8055 (N_8055,N_7503,N_7875);
and U8056 (N_8056,N_7950,N_7684);
nor U8057 (N_8057,N_7830,N_7583);
or U8058 (N_8058,N_7892,N_7565);
and U8059 (N_8059,N_7727,N_7852);
or U8060 (N_8060,N_7570,N_7549);
and U8061 (N_8061,N_7874,N_7527);
or U8062 (N_8062,N_7796,N_7739);
or U8063 (N_8063,N_7828,N_7721);
nor U8064 (N_8064,N_7764,N_7683);
or U8065 (N_8065,N_7567,N_7649);
and U8066 (N_8066,N_7609,N_7838);
or U8067 (N_8067,N_7605,N_7621);
or U8068 (N_8068,N_7571,N_7547);
xnor U8069 (N_8069,N_7677,N_7606);
or U8070 (N_8070,N_7982,N_7541);
nor U8071 (N_8071,N_7991,N_7919);
xor U8072 (N_8072,N_7612,N_7963);
nor U8073 (N_8073,N_7548,N_7797);
nand U8074 (N_8074,N_7782,N_7858);
nand U8075 (N_8075,N_7905,N_7618);
and U8076 (N_8076,N_7868,N_7774);
and U8077 (N_8077,N_7697,N_7627);
and U8078 (N_8078,N_7888,N_7595);
nand U8079 (N_8079,N_7812,N_7901);
xor U8080 (N_8080,N_7610,N_7753);
or U8081 (N_8081,N_7877,N_7758);
or U8082 (N_8082,N_7759,N_7604);
nor U8083 (N_8083,N_7713,N_7543);
xor U8084 (N_8084,N_7953,N_7528);
xor U8085 (N_8085,N_7575,N_7509);
xor U8086 (N_8086,N_7795,N_7693);
xor U8087 (N_8087,N_7940,N_7735);
nor U8088 (N_8088,N_7732,N_7994);
and U8089 (N_8089,N_7800,N_7540);
or U8090 (N_8090,N_7904,N_7857);
xor U8091 (N_8091,N_7985,N_7524);
or U8092 (N_8092,N_7522,N_7933);
or U8093 (N_8093,N_7661,N_7745);
xor U8094 (N_8094,N_7537,N_7827);
xor U8095 (N_8095,N_7760,N_7655);
nand U8096 (N_8096,N_7853,N_7809);
nand U8097 (N_8097,N_7834,N_7998);
nor U8098 (N_8098,N_7785,N_7784);
and U8099 (N_8099,N_7854,N_7801);
and U8100 (N_8100,N_7856,N_7952);
xor U8101 (N_8101,N_7505,N_7842);
nand U8102 (N_8102,N_7687,N_7883);
xnor U8103 (N_8103,N_7934,N_7755);
xor U8104 (N_8104,N_7639,N_7941);
and U8105 (N_8105,N_7778,N_7862);
xor U8106 (N_8106,N_7659,N_7859);
nand U8107 (N_8107,N_7930,N_7597);
nand U8108 (N_8108,N_7598,N_7726);
nand U8109 (N_8109,N_7552,N_7700);
nand U8110 (N_8110,N_7555,N_7822);
xnor U8111 (N_8111,N_7566,N_7756);
or U8112 (N_8112,N_7686,N_7500);
nor U8113 (N_8113,N_7971,N_7900);
xor U8114 (N_8114,N_7851,N_7990);
nand U8115 (N_8115,N_7630,N_7762);
and U8116 (N_8116,N_7562,N_7886);
nor U8117 (N_8117,N_7923,N_7561);
nor U8118 (N_8118,N_7614,N_7531);
xor U8119 (N_8119,N_7682,N_7738);
and U8120 (N_8120,N_7652,N_7594);
nor U8121 (N_8121,N_7777,N_7843);
xor U8122 (N_8122,N_7987,N_7631);
nand U8123 (N_8123,N_7589,N_7600);
nand U8124 (N_8124,N_7675,N_7510);
nand U8125 (N_8125,N_7730,N_7634);
nor U8126 (N_8126,N_7884,N_7918);
and U8127 (N_8127,N_7837,N_7910);
or U8128 (N_8128,N_7672,N_7765);
or U8129 (N_8129,N_7819,N_7958);
xor U8130 (N_8130,N_7962,N_7554);
xor U8131 (N_8131,N_7944,N_7743);
or U8132 (N_8132,N_7936,N_7821);
nor U8133 (N_8133,N_7641,N_7722);
or U8134 (N_8134,N_7526,N_7569);
nor U8135 (N_8135,N_7833,N_7820);
or U8136 (N_8136,N_7978,N_7863);
xnor U8137 (N_8137,N_7720,N_7654);
nor U8138 (N_8138,N_7692,N_7816);
and U8139 (N_8139,N_7839,N_7592);
nor U8140 (N_8140,N_7578,N_7885);
xor U8141 (N_8141,N_7624,N_7802);
and U8142 (N_8142,N_7993,N_7551);
xor U8143 (N_8143,N_7902,N_7909);
xor U8144 (N_8144,N_7917,N_7959);
or U8145 (N_8145,N_7724,N_7519);
nor U8146 (N_8146,N_7653,N_7891);
or U8147 (N_8147,N_7704,N_7744);
nand U8148 (N_8148,N_7626,N_7643);
nand U8149 (N_8149,N_7908,N_7969);
nor U8150 (N_8150,N_7694,N_7749);
xor U8151 (N_8151,N_7748,N_7590);
nand U8152 (N_8152,N_7518,N_7961);
nand U8153 (N_8153,N_7895,N_7742);
or U8154 (N_8154,N_7535,N_7790);
and U8155 (N_8155,N_7898,N_7515);
nor U8156 (N_8156,N_7771,N_7690);
nand U8157 (N_8157,N_7808,N_7667);
nor U8158 (N_8158,N_7983,N_7789);
nor U8159 (N_8159,N_7968,N_7783);
nand U8160 (N_8160,N_7925,N_7617);
nor U8161 (N_8161,N_7876,N_7999);
nor U8162 (N_8162,N_7907,N_7714);
xor U8163 (N_8163,N_7866,N_7814);
nor U8164 (N_8164,N_7647,N_7530);
and U8165 (N_8165,N_7633,N_7836);
nor U8166 (N_8166,N_7920,N_7867);
xnor U8167 (N_8167,N_7638,N_7558);
and U8168 (N_8168,N_7733,N_7636);
nor U8169 (N_8169,N_7542,N_7582);
nand U8170 (N_8170,N_7502,N_7546);
nand U8171 (N_8171,N_7929,N_7946);
nor U8172 (N_8172,N_7706,N_7703);
nand U8173 (N_8173,N_7957,N_7593);
and U8174 (N_8174,N_7545,N_7646);
xnor U8175 (N_8175,N_7855,N_7913);
xor U8176 (N_8176,N_7750,N_7935);
and U8177 (N_8177,N_7781,N_7973);
or U8178 (N_8178,N_7525,N_7734);
and U8179 (N_8179,N_7861,N_7927);
and U8180 (N_8180,N_7810,N_7779);
or U8181 (N_8181,N_7645,N_7553);
and U8182 (N_8182,N_7906,N_7970);
nand U8183 (N_8183,N_7517,N_7911);
and U8184 (N_8184,N_7662,N_7532);
nand U8185 (N_8185,N_7536,N_7523);
or U8186 (N_8186,N_7926,N_7607);
or U8187 (N_8187,N_7685,N_7680);
nand U8188 (N_8188,N_7715,N_7539);
nand U8189 (N_8189,N_7572,N_7668);
nor U8190 (N_8190,N_7619,N_7823);
xor U8191 (N_8191,N_7651,N_7587);
or U8192 (N_8192,N_7689,N_7507);
and U8193 (N_8193,N_7603,N_7865);
nor U8194 (N_8194,N_7728,N_7718);
xnor U8195 (N_8195,N_7608,N_7709);
nand U8196 (N_8196,N_7635,N_7584);
nand U8197 (N_8197,N_7948,N_7701);
or U8198 (N_8198,N_7698,N_7591);
nor U8199 (N_8199,N_7975,N_7956);
and U8200 (N_8200,N_7717,N_7960);
xor U8201 (N_8201,N_7665,N_7835);
xnor U8202 (N_8202,N_7573,N_7580);
and U8203 (N_8203,N_7710,N_7860);
or U8204 (N_8204,N_7533,N_7840);
nand U8205 (N_8205,N_7725,N_7766);
nor U8206 (N_8206,N_7776,N_7894);
nand U8207 (N_8207,N_7563,N_7829);
or U8208 (N_8208,N_7585,N_7656);
xnor U8209 (N_8209,N_7928,N_7775);
nand U8210 (N_8210,N_7648,N_7658);
and U8211 (N_8211,N_7577,N_7737);
nand U8212 (N_8212,N_7799,N_7550);
nor U8213 (N_8213,N_7945,N_7688);
nor U8214 (N_8214,N_7804,N_7872);
nand U8215 (N_8215,N_7716,N_7832);
or U8216 (N_8216,N_7707,N_7512);
xnor U8217 (N_8217,N_7881,N_7931);
nand U8218 (N_8218,N_7752,N_7511);
and U8219 (N_8219,N_7811,N_7751);
nor U8220 (N_8220,N_7965,N_7559);
and U8221 (N_8221,N_7916,N_7870);
nor U8222 (N_8222,N_7613,N_7813);
or U8223 (N_8223,N_7912,N_7581);
nand U8224 (N_8224,N_7669,N_7611);
or U8225 (N_8225,N_7981,N_7501);
xnor U8226 (N_8226,N_7599,N_7942);
and U8227 (N_8227,N_7514,N_7806);
and U8228 (N_8228,N_7625,N_7674);
and U8229 (N_8229,N_7729,N_7723);
nand U8230 (N_8230,N_7791,N_7788);
xor U8231 (N_8231,N_7817,N_7980);
and U8232 (N_8232,N_7616,N_7864);
and U8233 (N_8233,N_7741,N_7769);
nor U8234 (N_8234,N_7538,N_7831);
nor U8235 (N_8235,N_7767,N_7824);
nand U8236 (N_8236,N_7786,N_7622);
and U8237 (N_8237,N_7596,N_7792);
xnor U8238 (N_8238,N_7986,N_7815);
xnor U8239 (N_8239,N_7657,N_7691);
xor U8240 (N_8240,N_7977,N_7564);
or U8241 (N_8241,N_7803,N_7794);
nand U8242 (N_8242,N_7984,N_7770);
nor U8243 (N_8243,N_7671,N_7508);
nand U8244 (N_8244,N_7844,N_7887);
xnor U8245 (N_8245,N_7845,N_7939);
xor U8246 (N_8246,N_7637,N_7557);
xor U8247 (N_8247,N_7681,N_7568);
nand U8248 (N_8248,N_7903,N_7992);
xor U8249 (N_8249,N_7560,N_7772);
and U8250 (N_8250,N_7597,N_7809);
or U8251 (N_8251,N_7802,N_7760);
nand U8252 (N_8252,N_7680,N_7712);
xnor U8253 (N_8253,N_7963,N_7800);
nor U8254 (N_8254,N_7665,N_7574);
or U8255 (N_8255,N_7803,N_7564);
nor U8256 (N_8256,N_7892,N_7800);
xor U8257 (N_8257,N_7911,N_7936);
xor U8258 (N_8258,N_7839,N_7652);
or U8259 (N_8259,N_7685,N_7997);
or U8260 (N_8260,N_7686,N_7657);
nand U8261 (N_8261,N_7865,N_7791);
nor U8262 (N_8262,N_7978,N_7922);
or U8263 (N_8263,N_7737,N_7755);
and U8264 (N_8264,N_7531,N_7880);
nor U8265 (N_8265,N_7623,N_7626);
xor U8266 (N_8266,N_7850,N_7920);
xnor U8267 (N_8267,N_7506,N_7958);
nor U8268 (N_8268,N_7538,N_7669);
xor U8269 (N_8269,N_7836,N_7877);
and U8270 (N_8270,N_7701,N_7589);
xnor U8271 (N_8271,N_7705,N_7709);
xor U8272 (N_8272,N_7746,N_7936);
and U8273 (N_8273,N_7605,N_7618);
nor U8274 (N_8274,N_7868,N_7557);
nand U8275 (N_8275,N_7969,N_7911);
nand U8276 (N_8276,N_7691,N_7830);
or U8277 (N_8277,N_7588,N_7644);
xnor U8278 (N_8278,N_7907,N_7629);
or U8279 (N_8279,N_7597,N_7945);
or U8280 (N_8280,N_7502,N_7737);
nor U8281 (N_8281,N_7848,N_7951);
nor U8282 (N_8282,N_7837,N_7556);
and U8283 (N_8283,N_7528,N_7695);
nand U8284 (N_8284,N_7958,N_7969);
or U8285 (N_8285,N_7962,N_7819);
nand U8286 (N_8286,N_7957,N_7888);
or U8287 (N_8287,N_7610,N_7510);
or U8288 (N_8288,N_7941,N_7594);
nor U8289 (N_8289,N_7679,N_7843);
or U8290 (N_8290,N_7615,N_7616);
nand U8291 (N_8291,N_7691,N_7555);
nor U8292 (N_8292,N_7661,N_7570);
nor U8293 (N_8293,N_7925,N_7638);
nand U8294 (N_8294,N_7675,N_7890);
nor U8295 (N_8295,N_7531,N_7567);
and U8296 (N_8296,N_7700,N_7832);
and U8297 (N_8297,N_7784,N_7883);
xnor U8298 (N_8298,N_7919,N_7657);
nor U8299 (N_8299,N_7625,N_7952);
nor U8300 (N_8300,N_7619,N_7825);
xor U8301 (N_8301,N_7954,N_7955);
xor U8302 (N_8302,N_7723,N_7921);
nand U8303 (N_8303,N_7875,N_7880);
and U8304 (N_8304,N_7807,N_7944);
xnor U8305 (N_8305,N_7704,N_7664);
nand U8306 (N_8306,N_7717,N_7583);
nor U8307 (N_8307,N_7809,N_7608);
and U8308 (N_8308,N_7502,N_7878);
nor U8309 (N_8309,N_7936,N_7727);
or U8310 (N_8310,N_7938,N_7963);
or U8311 (N_8311,N_7795,N_7688);
xnor U8312 (N_8312,N_7687,N_7772);
nor U8313 (N_8313,N_7957,N_7554);
or U8314 (N_8314,N_7880,N_7762);
nor U8315 (N_8315,N_7669,N_7542);
nor U8316 (N_8316,N_7630,N_7857);
or U8317 (N_8317,N_7589,N_7758);
and U8318 (N_8318,N_7640,N_7642);
xnor U8319 (N_8319,N_7597,N_7590);
nor U8320 (N_8320,N_7727,N_7725);
and U8321 (N_8321,N_7822,N_7877);
and U8322 (N_8322,N_7728,N_7542);
and U8323 (N_8323,N_7943,N_7883);
nor U8324 (N_8324,N_7666,N_7825);
nor U8325 (N_8325,N_7543,N_7659);
xor U8326 (N_8326,N_7943,N_7718);
nor U8327 (N_8327,N_7513,N_7517);
nand U8328 (N_8328,N_7989,N_7906);
xnor U8329 (N_8329,N_7977,N_7554);
xor U8330 (N_8330,N_7880,N_7943);
or U8331 (N_8331,N_7946,N_7900);
xnor U8332 (N_8332,N_7987,N_7713);
or U8333 (N_8333,N_7520,N_7712);
nor U8334 (N_8334,N_7675,N_7871);
and U8335 (N_8335,N_7814,N_7984);
nor U8336 (N_8336,N_7716,N_7609);
xnor U8337 (N_8337,N_7729,N_7853);
xor U8338 (N_8338,N_7899,N_7834);
xnor U8339 (N_8339,N_7534,N_7862);
and U8340 (N_8340,N_7805,N_7872);
or U8341 (N_8341,N_7643,N_7869);
or U8342 (N_8342,N_7698,N_7587);
and U8343 (N_8343,N_7676,N_7607);
nor U8344 (N_8344,N_7651,N_7778);
nor U8345 (N_8345,N_7594,N_7623);
nor U8346 (N_8346,N_7742,N_7702);
nand U8347 (N_8347,N_7549,N_7877);
and U8348 (N_8348,N_7721,N_7659);
nor U8349 (N_8349,N_7508,N_7816);
nand U8350 (N_8350,N_7676,N_7829);
or U8351 (N_8351,N_7965,N_7595);
xnor U8352 (N_8352,N_7720,N_7501);
nand U8353 (N_8353,N_7947,N_7567);
nor U8354 (N_8354,N_7558,N_7547);
xnor U8355 (N_8355,N_7947,N_7677);
or U8356 (N_8356,N_7553,N_7682);
and U8357 (N_8357,N_7839,N_7963);
nor U8358 (N_8358,N_7996,N_7578);
xor U8359 (N_8359,N_7576,N_7988);
nand U8360 (N_8360,N_7868,N_7571);
nand U8361 (N_8361,N_7516,N_7657);
nand U8362 (N_8362,N_7686,N_7631);
xor U8363 (N_8363,N_7672,N_7666);
and U8364 (N_8364,N_7611,N_7952);
nand U8365 (N_8365,N_7868,N_7550);
nand U8366 (N_8366,N_7707,N_7964);
or U8367 (N_8367,N_7877,N_7735);
xor U8368 (N_8368,N_7955,N_7525);
xnor U8369 (N_8369,N_7955,N_7707);
and U8370 (N_8370,N_7545,N_7560);
or U8371 (N_8371,N_7672,N_7583);
xor U8372 (N_8372,N_7671,N_7515);
xnor U8373 (N_8373,N_7569,N_7761);
xnor U8374 (N_8374,N_7869,N_7845);
nand U8375 (N_8375,N_7649,N_7924);
or U8376 (N_8376,N_7971,N_7910);
or U8377 (N_8377,N_7963,N_7921);
and U8378 (N_8378,N_7793,N_7883);
nand U8379 (N_8379,N_7824,N_7778);
nor U8380 (N_8380,N_7673,N_7893);
nor U8381 (N_8381,N_7708,N_7671);
or U8382 (N_8382,N_7761,N_7701);
xnor U8383 (N_8383,N_7788,N_7783);
and U8384 (N_8384,N_7712,N_7579);
xor U8385 (N_8385,N_7671,N_7913);
and U8386 (N_8386,N_7610,N_7664);
nor U8387 (N_8387,N_7657,N_7891);
nand U8388 (N_8388,N_7908,N_7721);
or U8389 (N_8389,N_7536,N_7549);
and U8390 (N_8390,N_7591,N_7635);
and U8391 (N_8391,N_7630,N_7622);
xor U8392 (N_8392,N_7857,N_7861);
nand U8393 (N_8393,N_7636,N_7926);
and U8394 (N_8394,N_7840,N_7929);
and U8395 (N_8395,N_7684,N_7691);
nand U8396 (N_8396,N_7790,N_7916);
nand U8397 (N_8397,N_7563,N_7776);
nor U8398 (N_8398,N_7906,N_7690);
nor U8399 (N_8399,N_7645,N_7879);
or U8400 (N_8400,N_7961,N_7721);
or U8401 (N_8401,N_7660,N_7684);
nor U8402 (N_8402,N_7727,N_7600);
and U8403 (N_8403,N_7665,N_7996);
and U8404 (N_8404,N_7539,N_7880);
xnor U8405 (N_8405,N_7631,N_7681);
and U8406 (N_8406,N_7808,N_7962);
nor U8407 (N_8407,N_7711,N_7912);
xnor U8408 (N_8408,N_7868,N_7618);
xor U8409 (N_8409,N_7555,N_7890);
xor U8410 (N_8410,N_7670,N_7951);
or U8411 (N_8411,N_7568,N_7534);
or U8412 (N_8412,N_7510,N_7698);
nor U8413 (N_8413,N_7609,N_7789);
nand U8414 (N_8414,N_7894,N_7962);
and U8415 (N_8415,N_7960,N_7753);
xor U8416 (N_8416,N_7721,N_7820);
and U8417 (N_8417,N_7760,N_7536);
or U8418 (N_8418,N_7930,N_7660);
nor U8419 (N_8419,N_7981,N_7721);
nor U8420 (N_8420,N_7854,N_7743);
and U8421 (N_8421,N_7784,N_7869);
nand U8422 (N_8422,N_7972,N_7911);
nor U8423 (N_8423,N_7771,N_7672);
nand U8424 (N_8424,N_7706,N_7657);
or U8425 (N_8425,N_7927,N_7992);
and U8426 (N_8426,N_7559,N_7929);
xnor U8427 (N_8427,N_7623,N_7853);
or U8428 (N_8428,N_7867,N_7559);
or U8429 (N_8429,N_7754,N_7601);
nor U8430 (N_8430,N_7673,N_7979);
or U8431 (N_8431,N_7874,N_7764);
or U8432 (N_8432,N_7997,N_7779);
nand U8433 (N_8433,N_7664,N_7707);
xnor U8434 (N_8434,N_7901,N_7916);
and U8435 (N_8435,N_7706,N_7638);
and U8436 (N_8436,N_7638,N_7728);
xor U8437 (N_8437,N_7890,N_7556);
or U8438 (N_8438,N_7686,N_7725);
xnor U8439 (N_8439,N_7932,N_7879);
or U8440 (N_8440,N_7721,N_7992);
nand U8441 (N_8441,N_7700,N_7574);
xor U8442 (N_8442,N_7666,N_7567);
nand U8443 (N_8443,N_7876,N_7753);
nor U8444 (N_8444,N_7827,N_7800);
nor U8445 (N_8445,N_7908,N_7785);
or U8446 (N_8446,N_7547,N_7814);
or U8447 (N_8447,N_7981,N_7951);
and U8448 (N_8448,N_7543,N_7662);
xor U8449 (N_8449,N_7554,N_7569);
and U8450 (N_8450,N_7760,N_7931);
or U8451 (N_8451,N_7610,N_7952);
xnor U8452 (N_8452,N_7843,N_7604);
xor U8453 (N_8453,N_7826,N_7593);
nand U8454 (N_8454,N_7638,N_7537);
nor U8455 (N_8455,N_7717,N_7936);
nand U8456 (N_8456,N_7907,N_7841);
and U8457 (N_8457,N_7679,N_7829);
and U8458 (N_8458,N_7856,N_7502);
xnor U8459 (N_8459,N_7578,N_7835);
nor U8460 (N_8460,N_7522,N_7710);
nand U8461 (N_8461,N_7787,N_7545);
nor U8462 (N_8462,N_7870,N_7763);
xnor U8463 (N_8463,N_7672,N_7504);
and U8464 (N_8464,N_7555,N_7664);
nor U8465 (N_8465,N_7755,N_7701);
or U8466 (N_8466,N_7666,N_7725);
nand U8467 (N_8467,N_7952,N_7656);
and U8468 (N_8468,N_7508,N_7704);
nor U8469 (N_8469,N_7507,N_7741);
nand U8470 (N_8470,N_7734,N_7683);
or U8471 (N_8471,N_7743,N_7679);
xnor U8472 (N_8472,N_7898,N_7745);
nand U8473 (N_8473,N_7630,N_7759);
nor U8474 (N_8474,N_7586,N_7879);
and U8475 (N_8475,N_7745,N_7954);
nor U8476 (N_8476,N_7803,N_7553);
nor U8477 (N_8477,N_7676,N_7904);
or U8478 (N_8478,N_7802,N_7677);
and U8479 (N_8479,N_7561,N_7545);
or U8480 (N_8480,N_7657,N_7716);
xor U8481 (N_8481,N_7875,N_7538);
nand U8482 (N_8482,N_7602,N_7554);
xor U8483 (N_8483,N_7968,N_7733);
xor U8484 (N_8484,N_7778,N_7773);
nor U8485 (N_8485,N_7998,N_7699);
nor U8486 (N_8486,N_7988,N_7722);
xnor U8487 (N_8487,N_7675,N_7509);
nand U8488 (N_8488,N_7917,N_7839);
and U8489 (N_8489,N_7753,N_7809);
nor U8490 (N_8490,N_7870,N_7758);
or U8491 (N_8491,N_7638,N_7667);
nor U8492 (N_8492,N_7839,N_7567);
nand U8493 (N_8493,N_7945,N_7643);
nor U8494 (N_8494,N_7626,N_7656);
nand U8495 (N_8495,N_7691,N_7692);
nor U8496 (N_8496,N_7728,N_7688);
or U8497 (N_8497,N_7901,N_7926);
or U8498 (N_8498,N_7971,N_7509);
nor U8499 (N_8499,N_7906,N_7880);
xor U8500 (N_8500,N_8141,N_8021);
nor U8501 (N_8501,N_8387,N_8150);
nor U8502 (N_8502,N_8067,N_8123);
nand U8503 (N_8503,N_8298,N_8216);
xnor U8504 (N_8504,N_8202,N_8461);
or U8505 (N_8505,N_8147,N_8170);
nand U8506 (N_8506,N_8175,N_8048);
and U8507 (N_8507,N_8481,N_8005);
and U8508 (N_8508,N_8222,N_8498);
or U8509 (N_8509,N_8133,N_8327);
nand U8510 (N_8510,N_8331,N_8218);
and U8511 (N_8511,N_8277,N_8169);
or U8512 (N_8512,N_8024,N_8151);
xor U8513 (N_8513,N_8430,N_8051);
nor U8514 (N_8514,N_8310,N_8267);
nor U8515 (N_8515,N_8392,N_8064);
xor U8516 (N_8516,N_8456,N_8107);
xor U8517 (N_8517,N_8217,N_8220);
and U8518 (N_8518,N_8370,N_8432);
xor U8519 (N_8519,N_8292,N_8382);
or U8520 (N_8520,N_8032,N_8452);
xor U8521 (N_8521,N_8045,N_8022);
nor U8522 (N_8522,N_8187,N_8201);
nand U8523 (N_8523,N_8479,N_8489);
xnor U8524 (N_8524,N_8078,N_8384);
nor U8525 (N_8525,N_8403,N_8282);
and U8526 (N_8526,N_8443,N_8468);
nor U8527 (N_8527,N_8495,N_8070);
xor U8528 (N_8528,N_8463,N_8129);
nor U8529 (N_8529,N_8484,N_8247);
and U8530 (N_8530,N_8029,N_8288);
nor U8531 (N_8531,N_8320,N_8254);
and U8532 (N_8532,N_8341,N_8271);
or U8533 (N_8533,N_8446,N_8246);
nand U8534 (N_8534,N_8156,N_8033);
nand U8535 (N_8535,N_8016,N_8465);
or U8536 (N_8536,N_8460,N_8130);
nand U8537 (N_8537,N_8091,N_8287);
nand U8538 (N_8538,N_8454,N_8080);
nor U8539 (N_8539,N_8050,N_8372);
and U8540 (N_8540,N_8226,N_8198);
and U8541 (N_8541,N_8058,N_8181);
nand U8542 (N_8542,N_8017,N_8233);
nor U8543 (N_8543,N_8306,N_8371);
nand U8544 (N_8544,N_8332,N_8411);
xnor U8545 (N_8545,N_8240,N_8335);
nand U8546 (N_8546,N_8180,N_8093);
or U8547 (N_8547,N_8265,N_8023);
nor U8548 (N_8548,N_8345,N_8027);
or U8549 (N_8549,N_8099,N_8472);
and U8550 (N_8550,N_8183,N_8348);
nor U8551 (N_8551,N_8380,N_8199);
and U8552 (N_8552,N_8098,N_8128);
nand U8553 (N_8553,N_8235,N_8423);
nor U8554 (N_8554,N_8073,N_8194);
or U8555 (N_8555,N_8088,N_8476);
or U8556 (N_8556,N_8179,N_8054);
xor U8557 (N_8557,N_8367,N_8121);
or U8558 (N_8558,N_8111,N_8471);
and U8559 (N_8559,N_8487,N_8044);
nor U8560 (N_8560,N_8291,N_8100);
and U8561 (N_8561,N_8440,N_8285);
xnor U8562 (N_8562,N_8263,N_8264);
nand U8563 (N_8563,N_8072,N_8492);
xor U8564 (N_8564,N_8449,N_8231);
nand U8565 (N_8565,N_8075,N_8459);
nand U8566 (N_8566,N_8256,N_8318);
nor U8567 (N_8567,N_8322,N_8122);
xnor U8568 (N_8568,N_8182,N_8002);
nor U8569 (N_8569,N_8165,N_8205);
nor U8570 (N_8570,N_8178,N_8259);
xnor U8571 (N_8571,N_8297,N_8353);
or U8572 (N_8572,N_8293,N_8125);
nand U8573 (N_8573,N_8092,N_8059);
nand U8574 (N_8574,N_8251,N_8046);
xor U8575 (N_8575,N_8011,N_8262);
nand U8576 (N_8576,N_8162,N_8168);
nor U8577 (N_8577,N_8209,N_8397);
xor U8578 (N_8578,N_8171,N_8117);
xnor U8579 (N_8579,N_8356,N_8010);
and U8580 (N_8580,N_8349,N_8069);
xor U8581 (N_8581,N_8142,N_8284);
nor U8582 (N_8582,N_8238,N_8085);
nand U8583 (N_8583,N_8483,N_8193);
xor U8584 (N_8584,N_8307,N_8490);
and U8585 (N_8585,N_8061,N_8152);
and U8586 (N_8586,N_8211,N_8290);
and U8587 (N_8587,N_8486,N_8427);
or U8588 (N_8588,N_8361,N_8300);
nand U8589 (N_8589,N_8145,N_8467);
nand U8590 (N_8590,N_8242,N_8225);
nor U8591 (N_8591,N_8040,N_8477);
nand U8592 (N_8592,N_8418,N_8478);
and U8593 (N_8593,N_8079,N_8034);
xor U8594 (N_8594,N_8227,N_8338);
or U8595 (N_8595,N_8491,N_8358);
or U8596 (N_8596,N_8261,N_8049);
and U8597 (N_8597,N_8223,N_8144);
xor U8598 (N_8598,N_8224,N_8499);
xor U8599 (N_8599,N_8406,N_8312);
nand U8600 (N_8600,N_8112,N_8028);
xnor U8601 (N_8601,N_8043,N_8239);
nand U8602 (N_8602,N_8082,N_8410);
nand U8603 (N_8603,N_8425,N_8055);
xnor U8604 (N_8604,N_8401,N_8375);
nor U8605 (N_8605,N_8294,N_8433);
xor U8606 (N_8606,N_8270,N_8068);
nand U8607 (N_8607,N_8031,N_8053);
and U8608 (N_8608,N_8097,N_8429);
xnor U8609 (N_8609,N_8347,N_8116);
nor U8610 (N_8610,N_8391,N_8083);
nor U8611 (N_8611,N_8455,N_8090);
nand U8612 (N_8612,N_8396,N_8381);
or U8613 (N_8613,N_8374,N_8369);
nor U8614 (N_8614,N_8114,N_8385);
or U8615 (N_8615,N_8436,N_8280);
nor U8616 (N_8616,N_8435,N_8431);
xnor U8617 (N_8617,N_8008,N_8106);
or U8618 (N_8618,N_8388,N_8036);
nor U8619 (N_8619,N_8038,N_8377);
nand U8620 (N_8620,N_8464,N_8422);
xor U8621 (N_8621,N_8351,N_8173);
or U8622 (N_8622,N_8447,N_8241);
nor U8623 (N_8623,N_8081,N_8434);
nand U8624 (N_8624,N_8163,N_8143);
and U8625 (N_8625,N_8444,N_8442);
and U8626 (N_8626,N_8333,N_8445);
and U8627 (N_8627,N_8230,N_8376);
xnor U8628 (N_8628,N_8373,N_8286);
nand U8629 (N_8629,N_8278,N_8204);
xnor U8630 (N_8630,N_8042,N_8243);
and U8631 (N_8631,N_8109,N_8462);
nand U8632 (N_8632,N_8065,N_8323);
and U8633 (N_8633,N_8189,N_8400);
xnor U8634 (N_8634,N_8482,N_8200);
and U8635 (N_8635,N_8428,N_8488);
nand U8636 (N_8636,N_8138,N_8249);
nand U8637 (N_8637,N_8139,N_8328);
nand U8638 (N_8638,N_8126,N_8309);
nand U8639 (N_8639,N_8157,N_8184);
xor U8640 (N_8640,N_8301,N_8340);
nand U8641 (N_8641,N_8304,N_8299);
nand U8642 (N_8642,N_8413,N_8172);
and U8643 (N_8643,N_8132,N_8269);
nor U8644 (N_8644,N_8394,N_8103);
nand U8645 (N_8645,N_8296,N_8237);
and U8646 (N_8646,N_8450,N_8366);
nand U8647 (N_8647,N_8245,N_8190);
or U8648 (N_8648,N_8494,N_8314);
xor U8649 (N_8649,N_8208,N_8496);
or U8650 (N_8650,N_8383,N_8120);
nor U8651 (N_8651,N_8363,N_8316);
or U8652 (N_8652,N_8086,N_8137);
and U8653 (N_8653,N_8339,N_8066);
or U8654 (N_8654,N_8398,N_8195);
nand U8655 (N_8655,N_8234,N_8077);
nor U8656 (N_8656,N_8134,N_8215);
or U8657 (N_8657,N_8283,N_8355);
or U8658 (N_8658,N_8272,N_8037);
and U8659 (N_8659,N_8281,N_8244);
nand U8660 (N_8660,N_8337,N_8015);
nand U8661 (N_8661,N_8003,N_8101);
xnor U8662 (N_8662,N_8453,N_8009);
nor U8663 (N_8663,N_8343,N_8104);
and U8664 (N_8664,N_8035,N_8052);
nand U8665 (N_8665,N_8305,N_8319);
nand U8666 (N_8666,N_8229,N_8480);
and U8667 (N_8667,N_8212,N_8047);
nand U8668 (N_8668,N_8188,N_8260);
nor U8669 (N_8669,N_8219,N_8395);
nor U8670 (N_8670,N_8315,N_8119);
nand U8671 (N_8671,N_8095,N_8415);
and U8672 (N_8672,N_8336,N_8466);
and U8673 (N_8673,N_8252,N_8160);
nor U8674 (N_8674,N_8146,N_8041);
and U8675 (N_8675,N_8108,N_8007);
and U8676 (N_8676,N_8360,N_8390);
or U8677 (N_8677,N_8324,N_8148);
or U8678 (N_8678,N_8342,N_8470);
and U8679 (N_8679,N_8062,N_8105);
nor U8680 (N_8680,N_8438,N_8001);
nor U8681 (N_8681,N_8404,N_8325);
nand U8682 (N_8682,N_8115,N_8253);
and U8683 (N_8683,N_8174,N_8127);
or U8684 (N_8684,N_8354,N_8196);
xor U8685 (N_8685,N_8057,N_8191);
xor U8686 (N_8686,N_8063,N_8378);
and U8687 (N_8687,N_8096,N_8417);
and U8688 (N_8688,N_8154,N_8056);
nor U8689 (N_8689,N_8039,N_8451);
nand U8690 (N_8690,N_8250,N_8419);
or U8691 (N_8691,N_8135,N_8493);
or U8692 (N_8692,N_8030,N_8273);
and U8693 (N_8693,N_8131,N_8248);
or U8694 (N_8694,N_8421,N_8074);
xnor U8695 (N_8695,N_8457,N_8311);
or U8696 (N_8696,N_8350,N_8159);
nand U8697 (N_8697,N_8026,N_8266);
xor U8698 (N_8698,N_8275,N_8303);
and U8699 (N_8699,N_8025,N_8386);
and U8700 (N_8700,N_8221,N_8414);
nor U8701 (N_8701,N_8020,N_8110);
nand U8702 (N_8702,N_8214,N_8321);
nor U8703 (N_8703,N_8402,N_8153);
xnor U8704 (N_8704,N_8176,N_8274);
xor U8705 (N_8705,N_8076,N_8364);
and U8706 (N_8706,N_8424,N_8213);
nor U8707 (N_8707,N_8308,N_8161);
and U8708 (N_8708,N_8158,N_8149);
nor U8709 (N_8709,N_8087,N_8448);
or U8710 (N_8710,N_8426,N_8060);
nor U8711 (N_8711,N_8207,N_8018);
xor U8712 (N_8712,N_8408,N_8210);
nor U8713 (N_8713,N_8441,N_8469);
or U8714 (N_8714,N_8228,N_8439);
xnor U8715 (N_8715,N_8236,N_8167);
xnor U8716 (N_8716,N_8203,N_8405);
xor U8717 (N_8717,N_8407,N_8416);
nor U8718 (N_8718,N_8255,N_8268);
nand U8719 (N_8719,N_8185,N_8412);
xor U8720 (N_8720,N_8399,N_8497);
and U8721 (N_8721,N_8013,N_8136);
or U8722 (N_8722,N_8155,N_8313);
xnor U8723 (N_8723,N_8118,N_8326);
or U8724 (N_8724,N_8258,N_8232);
nor U8725 (N_8725,N_8357,N_8389);
and U8726 (N_8726,N_8485,N_8102);
nand U8727 (N_8727,N_8006,N_8302);
nor U8728 (N_8728,N_8071,N_8000);
or U8729 (N_8729,N_8166,N_8359);
nand U8730 (N_8730,N_8379,N_8004);
nand U8731 (N_8731,N_8276,N_8334);
xor U8732 (N_8732,N_8140,N_8362);
nor U8733 (N_8733,N_8197,N_8368);
xnor U8734 (N_8734,N_8089,N_8164);
and U8735 (N_8735,N_8346,N_8473);
nor U8736 (N_8736,N_8186,N_8420);
and U8737 (N_8737,N_8019,N_8409);
nand U8738 (N_8738,N_8317,N_8289);
nand U8739 (N_8739,N_8393,N_8084);
and U8740 (N_8740,N_8458,N_8012);
and U8741 (N_8741,N_8094,N_8352);
nand U8742 (N_8742,N_8475,N_8295);
nand U8743 (N_8743,N_8279,N_8474);
nor U8744 (N_8744,N_8344,N_8124);
xor U8745 (N_8745,N_8365,N_8014);
nand U8746 (N_8746,N_8177,N_8437);
nor U8747 (N_8747,N_8113,N_8329);
nand U8748 (N_8748,N_8257,N_8330);
nand U8749 (N_8749,N_8192,N_8206);
nor U8750 (N_8750,N_8156,N_8398);
nor U8751 (N_8751,N_8020,N_8041);
and U8752 (N_8752,N_8198,N_8372);
xor U8753 (N_8753,N_8222,N_8264);
or U8754 (N_8754,N_8304,N_8263);
or U8755 (N_8755,N_8233,N_8456);
nor U8756 (N_8756,N_8316,N_8126);
xnor U8757 (N_8757,N_8108,N_8009);
nor U8758 (N_8758,N_8410,N_8347);
and U8759 (N_8759,N_8102,N_8401);
nand U8760 (N_8760,N_8220,N_8057);
nand U8761 (N_8761,N_8327,N_8058);
xnor U8762 (N_8762,N_8380,N_8023);
or U8763 (N_8763,N_8147,N_8348);
nand U8764 (N_8764,N_8440,N_8027);
nand U8765 (N_8765,N_8034,N_8283);
nand U8766 (N_8766,N_8054,N_8193);
xnor U8767 (N_8767,N_8220,N_8327);
nand U8768 (N_8768,N_8282,N_8304);
nand U8769 (N_8769,N_8345,N_8031);
xor U8770 (N_8770,N_8414,N_8095);
or U8771 (N_8771,N_8423,N_8344);
nand U8772 (N_8772,N_8440,N_8356);
nand U8773 (N_8773,N_8344,N_8318);
nor U8774 (N_8774,N_8164,N_8462);
nand U8775 (N_8775,N_8155,N_8145);
and U8776 (N_8776,N_8345,N_8016);
nand U8777 (N_8777,N_8109,N_8350);
nand U8778 (N_8778,N_8027,N_8031);
nor U8779 (N_8779,N_8390,N_8343);
xor U8780 (N_8780,N_8276,N_8454);
and U8781 (N_8781,N_8333,N_8421);
nor U8782 (N_8782,N_8352,N_8015);
xnor U8783 (N_8783,N_8442,N_8078);
and U8784 (N_8784,N_8314,N_8324);
xnor U8785 (N_8785,N_8201,N_8182);
xor U8786 (N_8786,N_8324,N_8491);
xnor U8787 (N_8787,N_8392,N_8007);
or U8788 (N_8788,N_8177,N_8217);
or U8789 (N_8789,N_8295,N_8029);
or U8790 (N_8790,N_8126,N_8485);
xor U8791 (N_8791,N_8018,N_8445);
and U8792 (N_8792,N_8220,N_8241);
nor U8793 (N_8793,N_8241,N_8197);
xor U8794 (N_8794,N_8448,N_8404);
or U8795 (N_8795,N_8174,N_8077);
nor U8796 (N_8796,N_8245,N_8354);
nand U8797 (N_8797,N_8047,N_8311);
or U8798 (N_8798,N_8277,N_8244);
nor U8799 (N_8799,N_8159,N_8026);
nand U8800 (N_8800,N_8091,N_8092);
and U8801 (N_8801,N_8411,N_8082);
xnor U8802 (N_8802,N_8267,N_8232);
xor U8803 (N_8803,N_8205,N_8399);
nand U8804 (N_8804,N_8208,N_8058);
xor U8805 (N_8805,N_8383,N_8249);
xor U8806 (N_8806,N_8034,N_8041);
nand U8807 (N_8807,N_8454,N_8048);
and U8808 (N_8808,N_8235,N_8189);
or U8809 (N_8809,N_8321,N_8406);
and U8810 (N_8810,N_8129,N_8452);
and U8811 (N_8811,N_8405,N_8010);
or U8812 (N_8812,N_8345,N_8357);
or U8813 (N_8813,N_8480,N_8228);
nand U8814 (N_8814,N_8290,N_8009);
nand U8815 (N_8815,N_8252,N_8417);
xnor U8816 (N_8816,N_8453,N_8445);
nor U8817 (N_8817,N_8314,N_8176);
and U8818 (N_8818,N_8032,N_8076);
or U8819 (N_8819,N_8050,N_8216);
and U8820 (N_8820,N_8376,N_8309);
and U8821 (N_8821,N_8154,N_8312);
and U8822 (N_8822,N_8467,N_8185);
or U8823 (N_8823,N_8039,N_8217);
xnor U8824 (N_8824,N_8237,N_8187);
nor U8825 (N_8825,N_8250,N_8329);
or U8826 (N_8826,N_8305,N_8101);
or U8827 (N_8827,N_8348,N_8377);
and U8828 (N_8828,N_8022,N_8134);
and U8829 (N_8829,N_8221,N_8428);
xnor U8830 (N_8830,N_8267,N_8468);
or U8831 (N_8831,N_8297,N_8444);
nor U8832 (N_8832,N_8323,N_8259);
nand U8833 (N_8833,N_8140,N_8448);
and U8834 (N_8834,N_8429,N_8292);
or U8835 (N_8835,N_8275,N_8174);
nor U8836 (N_8836,N_8329,N_8303);
nor U8837 (N_8837,N_8388,N_8376);
or U8838 (N_8838,N_8022,N_8123);
xor U8839 (N_8839,N_8305,N_8004);
and U8840 (N_8840,N_8285,N_8434);
or U8841 (N_8841,N_8436,N_8153);
nand U8842 (N_8842,N_8436,N_8367);
xor U8843 (N_8843,N_8453,N_8027);
nor U8844 (N_8844,N_8259,N_8409);
xnor U8845 (N_8845,N_8281,N_8345);
nand U8846 (N_8846,N_8306,N_8218);
or U8847 (N_8847,N_8157,N_8413);
and U8848 (N_8848,N_8118,N_8376);
or U8849 (N_8849,N_8364,N_8284);
nor U8850 (N_8850,N_8178,N_8461);
and U8851 (N_8851,N_8456,N_8136);
xor U8852 (N_8852,N_8304,N_8382);
nand U8853 (N_8853,N_8170,N_8234);
xnor U8854 (N_8854,N_8254,N_8391);
xor U8855 (N_8855,N_8226,N_8329);
nand U8856 (N_8856,N_8425,N_8443);
and U8857 (N_8857,N_8498,N_8051);
nand U8858 (N_8858,N_8049,N_8436);
nand U8859 (N_8859,N_8342,N_8317);
xor U8860 (N_8860,N_8044,N_8357);
and U8861 (N_8861,N_8257,N_8414);
nor U8862 (N_8862,N_8350,N_8364);
nor U8863 (N_8863,N_8071,N_8085);
nand U8864 (N_8864,N_8418,N_8289);
nor U8865 (N_8865,N_8474,N_8057);
nor U8866 (N_8866,N_8356,N_8126);
and U8867 (N_8867,N_8356,N_8192);
xor U8868 (N_8868,N_8301,N_8488);
and U8869 (N_8869,N_8144,N_8312);
nor U8870 (N_8870,N_8432,N_8406);
nor U8871 (N_8871,N_8030,N_8349);
nor U8872 (N_8872,N_8059,N_8206);
nor U8873 (N_8873,N_8286,N_8170);
xor U8874 (N_8874,N_8235,N_8242);
or U8875 (N_8875,N_8067,N_8223);
or U8876 (N_8876,N_8225,N_8100);
nor U8877 (N_8877,N_8022,N_8082);
and U8878 (N_8878,N_8172,N_8111);
and U8879 (N_8879,N_8252,N_8432);
and U8880 (N_8880,N_8111,N_8170);
nand U8881 (N_8881,N_8392,N_8190);
and U8882 (N_8882,N_8129,N_8045);
nor U8883 (N_8883,N_8349,N_8316);
nand U8884 (N_8884,N_8433,N_8181);
xor U8885 (N_8885,N_8344,N_8207);
nand U8886 (N_8886,N_8317,N_8483);
and U8887 (N_8887,N_8079,N_8354);
xor U8888 (N_8888,N_8451,N_8037);
and U8889 (N_8889,N_8424,N_8160);
and U8890 (N_8890,N_8174,N_8457);
or U8891 (N_8891,N_8381,N_8067);
nand U8892 (N_8892,N_8447,N_8138);
xor U8893 (N_8893,N_8080,N_8260);
nand U8894 (N_8894,N_8408,N_8330);
nand U8895 (N_8895,N_8268,N_8362);
nand U8896 (N_8896,N_8028,N_8490);
nor U8897 (N_8897,N_8398,N_8187);
xnor U8898 (N_8898,N_8328,N_8204);
and U8899 (N_8899,N_8254,N_8317);
or U8900 (N_8900,N_8384,N_8231);
nand U8901 (N_8901,N_8080,N_8235);
and U8902 (N_8902,N_8294,N_8199);
xor U8903 (N_8903,N_8074,N_8326);
nor U8904 (N_8904,N_8334,N_8161);
nor U8905 (N_8905,N_8069,N_8134);
nand U8906 (N_8906,N_8170,N_8442);
xnor U8907 (N_8907,N_8000,N_8327);
nor U8908 (N_8908,N_8105,N_8280);
xnor U8909 (N_8909,N_8467,N_8033);
xor U8910 (N_8910,N_8236,N_8350);
and U8911 (N_8911,N_8330,N_8082);
xnor U8912 (N_8912,N_8335,N_8201);
xnor U8913 (N_8913,N_8229,N_8362);
xnor U8914 (N_8914,N_8235,N_8378);
or U8915 (N_8915,N_8416,N_8174);
and U8916 (N_8916,N_8466,N_8307);
nand U8917 (N_8917,N_8159,N_8387);
nor U8918 (N_8918,N_8371,N_8156);
nor U8919 (N_8919,N_8047,N_8334);
xor U8920 (N_8920,N_8190,N_8396);
nor U8921 (N_8921,N_8313,N_8166);
nand U8922 (N_8922,N_8200,N_8244);
and U8923 (N_8923,N_8138,N_8342);
nor U8924 (N_8924,N_8148,N_8078);
and U8925 (N_8925,N_8307,N_8168);
nand U8926 (N_8926,N_8071,N_8126);
nor U8927 (N_8927,N_8387,N_8426);
and U8928 (N_8928,N_8364,N_8108);
xor U8929 (N_8929,N_8290,N_8032);
and U8930 (N_8930,N_8341,N_8055);
and U8931 (N_8931,N_8494,N_8325);
nand U8932 (N_8932,N_8337,N_8309);
nand U8933 (N_8933,N_8199,N_8459);
nand U8934 (N_8934,N_8480,N_8233);
nand U8935 (N_8935,N_8090,N_8464);
xor U8936 (N_8936,N_8033,N_8206);
xnor U8937 (N_8937,N_8431,N_8351);
nor U8938 (N_8938,N_8481,N_8082);
and U8939 (N_8939,N_8256,N_8272);
and U8940 (N_8940,N_8206,N_8168);
nand U8941 (N_8941,N_8229,N_8288);
xor U8942 (N_8942,N_8323,N_8199);
nand U8943 (N_8943,N_8332,N_8496);
nand U8944 (N_8944,N_8133,N_8176);
nor U8945 (N_8945,N_8290,N_8416);
or U8946 (N_8946,N_8229,N_8465);
xor U8947 (N_8947,N_8147,N_8128);
nand U8948 (N_8948,N_8305,N_8080);
nand U8949 (N_8949,N_8325,N_8420);
or U8950 (N_8950,N_8083,N_8270);
and U8951 (N_8951,N_8409,N_8034);
and U8952 (N_8952,N_8384,N_8388);
nor U8953 (N_8953,N_8122,N_8203);
nand U8954 (N_8954,N_8364,N_8227);
xnor U8955 (N_8955,N_8392,N_8309);
and U8956 (N_8956,N_8033,N_8163);
nor U8957 (N_8957,N_8387,N_8481);
nand U8958 (N_8958,N_8482,N_8487);
and U8959 (N_8959,N_8498,N_8431);
xnor U8960 (N_8960,N_8388,N_8161);
nand U8961 (N_8961,N_8124,N_8001);
or U8962 (N_8962,N_8384,N_8058);
and U8963 (N_8963,N_8218,N_8087);
xor U8964 (N_8964,N_8218,N_8073);
and U8965 (N_8965,N_8068,N_8174);
and U8966 (N_8966,N_8244,N_8254);
xnor U8967 (N_8967,N_8019,N_8331);
nor U8968 (N_8968,N_8379,N_8224);
nand U8969 (N_8969,N_8453,N_8476);
nor U8970 (N_8970,N_8262,N_8159);
xor U8971 (N_8971,N_8143,N_8149);
xor U8972 (N_8972,N_8169,N_8006);
nand U8973 (N_8973,N_8100,N_8242);
nor U8974 (N_8974,N_8200,N_8045);
nand U8975 (N_8975,N_8049,N_8104);
and U8976 (N_8976,N_8278,N_8345);
xnor U8977 (N_8977,N_8355,N_8207);
nand U8978 (N_8978,N_8075,N_8165);
and U8979 (N_8979,N_8146,N_8236);
or U8980 (N_8980,N_8373,N_8085);
nor U8981 (N_8981,N_8001,N_8199);
or U8982 (N_8982,N_8293,N_8128);
or U8983 (N_8983,N_8367,N_8192);
xnor U8984 (N_8984,N_8490,N_8353);
xor U8985 (N_8985,N_8302,N_8121);
and U8986 (N_8986,N_8060,N_8469);
or U8987 (N_8987,N_8246,N_8282);
or U8988 (N_8988,N_8179,N_8133);
and U8989 (N_8989,N_8288,N_8403);
or U8990 (N_8990,N_8172,N_8346);
xnor U8991 (N_8991,N_8371,N_8043);
nor U8992 (N_8992,N_8019,N_8376);
nand U8993 (N_8993,N_8363,N_8418);
nor U8994 (N_8994,N_8352,N_8214);
or U8995 (N_8995,N_8257,N_8415);
nor U8996 (N_8996,N_8474,N_8223);
or U8997 (N_8997,N_8382,N_8442);
xor U8998 (N_8998,N_8188,N_8349);
nand U8999 (N_8999,N_8283,N_8258);
nor U9000 (N_9000,N_8969,N_8564);
nand U9001 (N_9001,N_8750,N_8796);
or U9002 (N_9002,N_8849,N_8847);
or U9003 (N_9003,N_8701,N_8804);
nand U9004 (N_9004,N_8655,N_8767);
nand U9005 (N_9005,N_8613,N_8630);
nor U9006 (N_9006,N_8947,N_8580);
nor U9007 (N_9007,N_8853,N_8720);
or U9008 (N_9008,N_8915,N_8734);
and U9009 (N_9009,N_8911,N_8755);
nor U9010 (N_9010,N_8574,N_8709);
nand U9011 (N_9011,N_8653,N_8743);
or U9012 (N_9012,N_8700,N_8550);
nand U9013 (N_9013,N_8839,N_8760);
nand U9014 (N_9014,N_8593,N_8799);
nand U9015 (N_9015,N_8888,N_8906);
xnor U9016 (N_9016,N_8551,N_8667);
nor U9017 (N_9017,N_8506,N_8628);
xor U9018 (N_9018,N_8617,N_8811);
nand U9019 (N_9019,N_8985,N_8671);
and U9020 (N_9020,N_8723,N_8900);
xor U9021 (N_9021,N_8511,N_8705);
or U9022 (N_9022,N_8817,N_8589);
nand U9023 (N_9023,N_8855,N_8591);
nor U9024 (N_9024,N_8757,N_8739);
or U9025 (N_9025,N_8941,N_8946);
nor U9026 (N_9026,N_8963,N_8980);
nand U9027 (N_9027,N_8658,N_8531);
nor U9028 (N_9028,N_8710,N_8590);
and U9029 (N_9029,N_8548,N_8534);
or U9030 (N_9030,N_8992,N_8523);
xnor U9031 (N_9031,N_8942,N_8549);
and U9032 (N_9032,N_8851,N_8738);
and U9033 (N_9033,N_8508,N_8538);
and U9034 (N_9034,N_8611,N_8844);
nor U9035 (N_9035,N_8514,N_8596);
or U9036 (N_9036,N_8692,N_8708);
and U9037 (N_9037,N_8547,N_8892);
and U9038 (N_9038,N_8570,N_8520);
xnor U9039 (N_9039,N_8938,N_8983);
nand U9040 (N_9040,N_8780,N_8869);
nor U9041 (N_9041,N_8977,N_8573);
nand U9042 (N_9042,N_8790,N_8503);
or U9043 (N_9043,N_8663,N_8877);
nand U9044 (N_9044,N_8659,N_8553);
nand U9045 (N_9045,N_8937,N_8896);
xnor U9046 (N_9046,N_8861,N_8837);
nand U9047 (N_9047,N_8815,N_8766);
or U9048 (N_9048,N_8558,N_8955);
xor U9049 (N_9049,N_8859,N_8545);
nand U9050 (N_9050,N_8620,N_8812);
nor U9051 (N_9051,N_8836,N_8651);
nand U9052 (N_9052,N_8940,N_8879);
xor U9053 (N_9053,N_8609,N_8685);
and U9054 (N_9054,N_8563,N_8552);
xor U9055 (N_9055,N_8825,N_8819);
nor U9056 (N_9056,N_8582,N_8728);
or U9057 (N_9057,N_8826,N_8525);
nand U9058 (N_9058,N_8987,N_8914);
nor U9059 (N_9059,N_8677,N_8908);
and U9060 (N_9060,N_8857,N_8647);
and U9061 (N_9061,N_8731,N_8950);
or U9062 (N_9062,N_8643,N_8560);
and U9063 (N_9063,N_8943,N_8664);
nor U9064 (N_9064,N_8704,N_8962);
nand U9065 (N_9065,N_8972,N_8541);
or U9066 (N_9066,N_8827,N_8850);
xnor U9067 (N_9067,N_8936,N_8800);
or U9068 (N_9068,N_8607,N_8583);
xnor U9069 (N_9069,N_8681,N_8572);
or U9070 (N_9070,N_8781,N_8510);
nor U9071 (N_9071,N_8882,N_8626);
nand U9072 (N_9072,N_8559,N_8627);
nand U9073 (N_9073,N_8810,N_8842);
or U9074 (N_9074,N_8921,N_8518);
xnor U9075 (N_9075,N_8522,N_8587);
xor U9076 (N_9076,N_8832,N_8668);
nand U9077 (N_9077,N_8689,N_8999);
and U9078 (N_9078,N_8762,N_8695);
and U9079 (N_9079,N_8752,N_8984);
or U9080 (N_9080,N_8814,N_8678);
and U9081 (N_9081,N_8960,N_8579);
and U9082 (N_9082,N_8935,N_8660);
xnor U9083 (N_9083,N_8504,N_8828);
xnor U9084 (N_9084,N_8698,N_8649);
or U9085 (N_9085,N_8872,N_8612);
or U9086 (N_9086,N_8576,N_8666);
nor U9087 (N_9087,N_8761,N_8745);
nand U9088 (N_9088,N_8951,N_8638);
nor U9089 (N_9089,N_8665,N_8656);
nor U9090 (N_9090,N_8772,N_8569);
or U9091 (N_9091,N_8715,N_8833);
and U9092 (N_9092,N_8897,N_8532);
nand U9093 (N_9093,N_8845,N_8903);
and U9094 (N_9094,N_8932,N_8934);
nor U9095 (N_9095,N_8952,N_8764);
xnor U9096 (N_9096,N_8916,N_8675);
nand U9097 (N_9097,N_8929,N_8634);
xor U9098 (N_9098,N_8961,N_8517);
and U9099 (N_9099,N_8867,N_8501);
and U9100 (N_9100,N_8994,N_8834);
xnor U9101 (N_9101,N_8797,N_8824);
and U9102 (N_9102,N_8979,N_8838);
nand U9103 (N_9103,N_8618,N_8778);
nor U9104 (N_9104,N_8688,N_8744);
and U9105 (N_9105,N_8543,N_8907);
nand U9106 (N_9106,N_8735,N_8615);
nand U9107 (N_9107,N_8724,N_8751);
or U9108 (N_9108,N_8650,N_8565);
nand U9109 (N_9109,N_8595,N_8995);
xnor U9110 (N_9110,N_8904,N_8939);
and U9111 (N_9111,N_8561,N_8753);
xor U9112 (N_9112,N_8927,N_8530);
and U9113 (N_9113,N_8736,N_8502);
or U9114 (N_9114,N_8680,N_8703);
xor U9115 (N_9115,N_8672,N_8599);
xor U9116 (N_9116,N_8697,N_8923);
xor U9117 (N_9117,N_8604,N_8562);
xnor U9118 (N_9118,N_8805,N_8798);
or U9119 (N_9119,N_8614,N_8537);
nand U9120 (N_9120,N_8557,N_8910);
xnor U9121 (N_9121,N_8873,N_8765);
or U9122 (N_9122,N_8990,N_8718);
or U9123 (N_9123,N_8644,N_8567);
xor U9124 (N_9124,N_8661,N_8600);
nor U9125 (N_9125,N_8917,N_8632);
or U9126 (N_9126,N_8544,N_8528);
and U9127 (N_9127,N_8775,N_8740);
and U9128 (N_9128,N_8893,N_8535);
nor U9129 (N_9129,N_8747,N_8807);
nor U9130 (N_9130,N_8894,N_8821);
or U9131 (N_9131,N_8625,N_8875);
nor U9132 (N_9132,N_8577,N_8905);
nand U9133 (N_9133,N_8782,N_8633);
or U9134 (N_9134,N_8787,N_8997);
xor U9135 (N_9135,N_8973,N_8868);
or U9136 (N_9136,N_8788,N_8746);
and U9137 (N_9137,N_8806,N_8533);
nand U9138 (N_9138,N_8512,N_8694);
xnor U9139 (N_9139,N_8652,N_8670);
nand U9140 (N_9140,N_8726,N_8902);
nor U9141 (N_9141,N_8895,N_8919);
nor U9142 (N_9142,N_8930,N_8621);
and U9143 (N_9143,N_8616,N_8500);
or U9144 (N_9144,N_8793,N_8759);
or U9145 (N_9145,N_8707,N_8640);
nand U9146 (N_9146,N_8729,N_8948);
or U9147 (N_9147,N_8684,N_8974);
nand U9148 (N_9148,N_8770,N_8792);
xnor U9149 (N_9149,N_8699,N_8989);
xnor U9150 (N_9150,N_8870,N_8555);
or U9151 (N_9151,N_8737,N_8721);
nand U9152 (N_9152,N_8673,N_8880);
and U9153 (N_9153,N_8635,N_8642);
nand U9154 (N_9154,N_8529,N_8803);
nor U9155 (N_9155,N_8794,N_8509);
nor U9156 (N_9156,N_8711,N_8889);
xor U9157 (N_9157,N_8901,N_8820);
or U9158 (N_9158,N_8871,N_8823);
and U9159 (N_9159,N_8791,N_8993);
nor U9160 (N_9160,N_8818,N_8748);
nand U9161 (N_9161,N_8777,N_8513);
nand U9162 (N_9162,N_8779,N_8505);
nor U9163 (N_9163,N_8978,N_8968);
nand U9164 (N_9164,N_8648,N_8885);
and U9165 (N_9165,N_8769,N_8816);
xnor U9166 (N_9166,N_8702,N_8860);
or U9167 (N_9167,N_8749,N_8540);
and U9168 (N_9168,N_8575,N_8959);
xor U9169 (N_9169,N_8776,N_8571);
xnor U9170 (N_9170,N_8608,N_8840);
nor U9171 (N_9171,N_8696,N_8713);
and U9172 (N_9172,N_8848,N_8965);
nand U9173 (N_9173,N_8975,N_8601);
or U9174 (N_9174,N_8730,N_8536);
nor U9175 (N_9175,N_8878,N_8988);
nor U9176 (N_9176,N_8866,N_8515);
xor U9177 (N_9177,N_8890,N_8725);
nor U9178 (N_9178,N_8958,N_8898);
nor U9179 (N_9179,N_8841,N_8773);
nand U9180 (N_9180,N_8886,N_8542);
xor U9181 (N_9181,N_8578,N_8913);
xor U9182 (N_9182,N_8588,N_8843);
nor U9183 (N_9183,N_8598,N_8683);
or U9184 (N_9184,N_8996,N_8981);
or U9185 (N_9185,N_8756,N_8956);
nor U9186 (N_9186,N_8581,N_8741);
xnor U9187 (N_9187,N_8526,N_8594);
or U9188 (N_9188,N_8846,N_8891);
and U9189 (N_9189,N_8830,N_8516);
xor U9190 (N_9190,N_8603,N_8933);
and U9191 (N_9191,N_8771,N_8622);
and U9192 (N_9192,N_8610,N_8592);
xnor U9193 (N_9193,N_8964,N_8733);
nor U9194 (N_9194,N_8554,N_8645);
and U9195 (N_9195,N_8662,N_8768);
and U9196 (N_9196,N_8602,N_8864);
nand U9197 (N_9197,N_8970,N_8691);
xor U9198 (N_9198,N_8931,N_8527);
or U9199 (N_9199,N_8763,N_8953);
and U9200 (N_9200,N_8966,N_8909);
or U9201 (N_9201,N_8546,N_8912);
and U9202 (N_9202,N_8856,N_8971);
nor U9203 (N_9203,N_8887,N_8802);
and U9204 (N_9204,N_8784,N_8920);
and U9205 (N_9205,N_8874,N_8881);
and U9206 (N_9206,N_8858,N_8682);
or U9207 (N_9207,N_8883,N_8945);
nor U9208 (N_9208,N_8597,N_8637);
or U9209 (N_9209,N_8801,N_8646);
nor U9210 (N_9210,N_8566,N_8783);
nor U9211 (N_9211,N_8654,N_8605);
or U9212 (N_9212,N_8986,N_8899);
and U9213 (N_9213,N_8928,N_8991);
nand U9214 (N_9214,N_8586,N_8884);
or U9215 (N_9215,N_8606,N_8924);
nand U9216 (N_9216,N_8519,N_8922);
xor U9217 (N_9217,N_8629,N_8507);
or U9218 (N_9218,N_8829,N_8727);
or U9219 (N_9219,N_8865,N_8717);
nand U9220 (N_9220,N_8669,N_8852);
nand U9221 (N_9221,N_8789,N_8679);
and U9222 (N_9222,N_8876,N_8631);
and U9223 (N_9223,N_8786,N_8624);
xnor U9224 (N_9224,N_8641,N_8774);
nor U9225 (N_9225,N_8785,N_8918);
xor U9226 (N_9226,N_8693,N_8926);
or U9227 (N_9227,N_8687,N_8809);
xnor U9228 (N_9228,N_8957,N_8944);
nand U9229 (N_9229,N_8639,N_8716);
or U9230 (N_9230,N_8862,N_8822);
nand U9231 (N_9231,N_8854,N_8585);
or U9232 (N_9232,N_8998,N_8863);
xor U9233 (N_9233,N_8674,N_8706);
and U9234 (N_9234,N_8714,N_8719);
xor U9235 (N_9235,N_8556,N_8690);
nand U9236 (N_9236,N_8949,N_8619);
xnor U9237 (N_9237,N_8831,N_8732);
nand U9238 (N_9238,N_8758,N_8657);
xnor U9239 (N_9239,N_8524,N_8976);
xnor U9240 (N_9240,N_8742,N_8584);
and U9241 (N_9241,N_8686,N_8808);
nor U9242 (N_9242,N_8925,N_8539);
and U9243 (N_9243,N_8636,N_8722);
nor U9244 (N_9244,N_8835,N_8568);
nor U9245 (N_9245,N_8712,N_8795);
xnor U9246 (N_9246,N_8521,N_8967);
nor U9247 (N_9247,N_8954,N_8754);
or U9248 (N_9248,N_8813,N_8676);
xnor U9249 (N_9249,N_8623,N_8982);
nor U9250 (N_9250,N_8595,N_8909);
xnor U9251 (N_9251,N_8589,N_8689);
or U9252 (N_9252,N_8687,N_8798);
xnor U9253 (N_9253,N_8697,N_8982);
nor U9254 (N_9254,N_8746,N_8564);
xor U9255 (N_9255,N_8822,N_8787);
or U9256 (N_9256,N_8697,N_8964);
nor U9257 (N_9257,N_8842,N_8557);
or U9258 (N_9258,N_8727,N_8907);
xnor U9259 (N_9259,N_8580,N_8923);
and U9260 (N_9260,N_8758,N_8861);
and U9261 (N_9261,N_8912,N_8948);
or U9262 (N_9262,N_8733,N_8760);
or U9263 (N_9263,N_8642,N_8648);
xor U9264 (N_9264,N_8711,N_8559);
nor U9265 (N_9265,N_8981,N_8591);
xor U9266 (N_9266,N_8690,N_8720);
and U9267 (N_9267,N_8585,N_8896);
xnor U9268 (N_9268,N_8861,N_8710);
nor U9269 (N_9269,N_8526,N_8786);
or U9270 (N_9270,N_8709,N_8844);
xor U9271 (N_9271,N_8589,N_8705);
or U9272 (N_9272,N_8762,N_8541);
or U9273 (N_9273,N_8901,N_8957);
or U9274 (N_9274,N_8809,N_8993);
or U9275 (N_9275,N_8987,N_8831);
nor U9276 (N_9276,N_8706,N_8654);
or U9277 (N_9277,N_8622,N_8583);
xor U9278 (N_9278,N_8976,N_8710);
xnor U9279 (N_9279,N_8883,N_8595);
nand U9280 (N_9280,N_8563,N_8715);
nor U9281 (N_9281,N_8738,N_8807);
nor U9282 (N_9282,N_8756,N_8975);
and U9283 (N_9283,N_8752,N_8779);
nor U9284 (N_9284,N_8868,N_8835);
xor U9285 (N_9285,N_8503,N_8991);
xnor U9286 (N_9286,N_8591,N_8727);
nor U9287 (N_9287,N_8920,N_8614);
and U9288 (N_9288,N_8643,N_8718);
nand U9289 (N_9289,N_8910,N_8786);
nor U9290 (N_9290,N_8650,N_8741);
xnor U9291 (N_9291,N_8694,N_8888);
xor U9292 (N_9292,N_8719,N_8500);
or U9293 (N_9293,N_8707,N_8830);
nand U9294 (N_9294,N_8928,N_8924);
or U9295 (N_9295,N_8732,N_8525);
xnor U9296 (N_9296,N_8568,N_8719);
xnor U9297 (N_9297,N_8564,N_8667);
nor U9298 (N_9298,N_8560,N_8887);
and U9299 (N_9299,N_8866,N_8671);
xor U9300 (N_9300,N_8910,N_8621);
and U9301 (N_9301,N_8760,N_8629);
and U9302 (N_9302,N_8886,N_8754);
nor U9303 (N_9303,N_8593,N_8977);
nand U9304 (N_9304,N_8531,N_8500);
or U9305 (N_9305,N_8635,N_8766);
nor U9306 (N_9306,N_8873,N_8827);
and U9307 (N_9307,N_8782,N_8720);
xor U9308 (N_9308,N_8520,N_8649);
nand U9309 (N_9309,N_8903,N_8823);
and U9310 (N_9310,N_8754,N_8527);
nor U9311 (N_9311,N_8523,N_8561);
or U9312 (N_9312,N_8811,N_8595);
and U9313 (N_9313,N_8534,N_8567);
or U9314 (N_9314,N_8759,N_8541);
and U9315 (N_9315,N_8970,N_8876);
nor U9316 (N_9316,N_8818,N_8990);
nand U9317 (N_9317,N_8903,N_8584);
nor U9318 (N_9318,N_8766,N_8995);
nor U9319 (N_9319,N_8535,N_8991);
or U9320 (N_9320,N_8874,N_8811);
nand U9321 (N_9321,N_8595,N_8621);
and U9322 (N_9322,N_8831,N_8752);
nor U9323 (N_9323,N_8929,N_8949);
xor U9324 (N_9324,N_8783,N_8641);
nand U9325 (N_9325,N_8740,N_8501);
nand U9326 (N_9326,N_8569,N_8624);
and U9327 (N_9327,N_8995,N_8809);
nor U9328 (N_9328,N_8819,N_8741);
or U9329 (N_9329,N_8827,N_8592);
or U9330 (N_9330,N_8869,N_8768);
or U9331 (N_9331,N_8777,N_8940);
nand U9332 (N_9332,N_8581,N_8752);
or U9333 (N_9333,N_8671,N_8708);
nand U9334 (N_9334,N_8936,N_8634);
nand U9335 (N_9335,N_8571,N_8639);
or U9336 (N_9336,N_8697,N_8546);
nor U9337 (N_9337,N_8814,N_8960);
or U9338 (N_9338,N_8529,N_8924);
xor U9339 (N_9339,N_8934,N_8852);
nor U9340 (N_9340,N_8768,N_8634);
nor U9341 (N_9341,N_8578,N_8809);
xnor U9342 (N_9342,N_8979,N_8530);
nor U9343 (N_9343,N_8514,N_8545);
nand U9344 (N_9344,N_8692,N_8722);
or U9345 (N_9345,N_8746,N_8888);
xor U9346 (N_9346,N_8920,N_8765);
or U9347 (N_9347,N_8575,N_8920);
nor U9348 (N_9348,N_8511,N_8791);
nand U9349 (N_9349,N_8771,N_8975);
or U9350 (N_9350,N_8782,N_8863);
xor U9351 (N_9351,N_8838,N_8642);
or U9352 (N_9352,N_8623,N_8793);
and U9353 (N_9353,N_8976,N_8711);
nor U9354 (N_9354,N_8632,N_8775);
xor U9355 (N_9355,N_8675,N_8896);
xnor U9356 (N_9356,N_8929,N_8681);
or U9357 (N_9357,N_8728,N_8522);
xnor U9358 (N_9358,N_8507,N_8895);
nand U9359 (N_9359,N_8576,N_8635);
nor U9360 (N_9360,N_8524,N_8679);
or U9361 (N_9361,N_8625,N_8881);
or U9362 (N_9362,N_8570,N_8687);
or U9363 (N_9363,N_8886,N_8794);
or U9364 (N_9364,N_8771,N_8641);
nor U9365 (N_9365,N_8671,N_8811);
nor U9366 (N_9366,N_8553,N_8929);
nand U9367 (N_9367,N_8577,N_8679);
and U9368 (N_9368,N_8879,N_8531);
or U9369 (N_9369,N_8788,N_8968);
xnor U9370 (N_9370,N_8829,N_8556);
nor U9371 (N_9371,N_8943,N_8897);
xor U9372 (N_9372,N_8534,N_8813);
nand U9373 (N_9373,N_8656,N_8673);
xnor U9374 (N_9374,N_8863,N_8675);
nor U9375 (N_9375,N_8508,N_8545);
nor U9376 (N_9376,N_8575,N_8594);
nand U9377 (N_9377,N_8607,N_8734);
nand U9378 (N_9378,N_8792,N_8532);
xor U9379 (N_9379,N_8865,N_8750);
nor U9380 (N_9380,N_8971,N_8799);
nand U9381 (N_9381,N_8835,N_8620);
nand U9382 (N_9382,N_8736,N_8912);
nor U9383 (N_9383,N_8539,N_8576);
and U9384 (N_9384,N_8911,N_8556);
or U9385 (N_9385,N_8978,N_8676);
and U9386 (N_9386,N_8744,N_8668);
nand U9387 (N_9387,N_8921,N_8875);
xnor U9388 (N_9388,N_8948,N_8561);
nor U9389 (N_9389,N_8889,N_8541);
and U9390 (N_9390,N_8638,N_8785);
nor U9391 (N_9391,N_8957,N_8891);
nand U9392 (N_9392,N_8883,N_8669);
nor U9393 (N_9393,N_8934,N_8747);
and U9394 (N_9394,N_8646,N_8825);
nand U9395 (N_9395,N_8639,N_8836);
or U9396 (N_9396,N_8651,N_8505);
and U9397 (N_9397,N_8703,N_8783);
xor U9398 (N_9398,N_8844,N_8898);
and U9399 (N_9399,N_8899,N_8529);
or U9400 (N_9400,N_8819,N_8972);
xnor U9401 (N_9401,N_8725,N_8807);
xnor U9402 (N_9402,N_8983,N_8774);
and U9403 (N_9403,N_8645,N_8564);
and U9404 (N_9404,N_8778,N_8712);
and U9405 (N_9405,N_8815,N_8826);
or U9406 (N_9406,N_8529,N_8585);
and U9407 (N_9407,N_8625,N_8690);
xnor U9408 (N_9408,N_8915,N_8652);
xor U9409 (N_9409,N_8543,N_8932);
xnor U9410 (N_9410,N_8717,N_8898);
and U9411 (N_9411,N_8596,N_8952);
xor U9412 (N_9412,N_8604,N_8869);
nand U9413 (N_9413,N_8536,N_8975);
xor U9414 (N_9414,N_8665,N_8950);
nand U9415 (N_9415,N_8639,N_8736);
nor U9416 (N_9416,N_8994,N_8538);
nand U9417 (N_9417,N_8970,N_8524);
and U9418 (N_9418,N_8650,N_8634);
nand U9419 (N_9419,N_8594,N_8793);
and U9420 (N_9420,N_8897,N_8827);
nor U9421 (N_9421,N_8663,N_8533);
nor U9422 (N_9422,N_8678,N_8534);
nand U9423 (N_9423,N_8881,N_8991);
and U9424 (N_9424,N_8645,N_8966);
or U9425 (N_9425,N_8813,N_8761);
and U9426 (N_9426,N_8877,N_8979);
nor U9427 (N_9427,N_8704,N_8668);
nand U9428 (N_9428,N_8936,N_8897);
nand U9429 (N_9429,N_8905,N_8847);
nor U9430 (N_9430,N_8637,N_8651);
xor U9431 (N_9431,N_8863,N_8700);
nand U9432 (N_9432,N_8760,N_8786);
or U9433 (N_9433,N_8746,N_8775);
nand U9434 (N_9434,N_8508,N_8725);
nand U9435 (N_9435,N_8678,N_8593);
and U9436 (N_9436,N_8775,N_8925);
or U9437 (N_9437,N_8975,N_8634);
nand U9438 (N_9438,N_8952,N_8671);
nand U9439 (N_9439,N_8952,N_8553);
and U9440 (N_9440,N_8984,N_8533);
nor U9441 (N_9441,N_8845,N_8765);
nor U9442 (N_9442,N_8923,N_8834);
and U9443 (N_9443,N_8877,N_8983);
nand U9444 (N_9444,N_8567,N_8584);
nor U9445 (N_9445,N_8672,N_8540);
or U9446 (N_9446,N_8704,N_8676);
nand U9447 (N_9447,N_8738,N_8626);
or U9448 (N_9448,N_8811,N_8869);
nand U9449 (N_9449,N_8967,N_8653);
or U9450 (N_9450,N_8994,N_8848);
nand U9451 (N_9451,N_8778,N_8857);
nand U9452 (N_9452,N_8806,N_8631);
nand U9453 (N_9453,N_8613,N_8546);
xnor U9454 (N_9454,N_8549,N_8530);
or U9455 (N_9455,N_8660,N_8782);
nor U9456 (N_9456,N_8515,N_8725);
nor U9457 (N_9457,N_8640,N_8754);
xor U9458 (N_9458,N_8667,N_8555);
xnor U9459 (N_9459,N_8816,N_8871);
and U9460 (N_9460,N_8768,N_8826);
and U9461 (N_9461,N_8620,N_8604);
nand U9462 (N_9462,N_8661,N_8941);
and U9463 (N_9463,N_8587,N_8501);
nor U9464 (N_9464,N_8642,N_8510);
or U9465 (N_9465,N_8880,N_8934);
and U9466 (N_9466,N_8877,N_8875);
or U9467 (N_9467,N_8860,N_8639);
nor U9468 (N_9468,N_8596,N_8963);
nand U9469 (N_9469,N_8586,N_8523);
nor U9470 (N_9470,N_8911,N_8871);
or U9471 (N_9471,N_8535,N_8574);
and U9472 (N_9472,N_8597,N_8616);
or U9473 (N_9473,N_8866,N_8707);
or U9474 (N_9474,N_8617,N_8538);
and U9475 (N_9475,N_8665,N_8585);
or U9476 (N_9476,N_8888,N_8870);
or U9477 (N_9477,N_8886,N_8796);
and U9478 (N_9478,N_8899,N_8705);
nor U9479 (N_9479,N_8560,N_8595);
and U9480 (N_9480,N_8638,N_8747);
or U9481 (N_9481,N_8649,N_8699);
xnor U9482 (N_9482,N_8702,N_8508);
nand U9483 (N_9483,N_8695,N_8956);
xnor U9484 (N_9484,N_8856,N_8781);
nand U9485 (N_9485,N_8511,N_8798);
xnor U9486 (N_9486,N_8825,N_8995);
or U9487 (N_9487,N_8596,N_8811);
xor U9488 (N_9488,N_8857,N_8937);
xnor U9489 (N_9489,N_8501,N_8858);
nor U9490 (N_9490,N_8834,N_8635);
and U9491 (N_9491,N_8523,N_8569);
or U9492 (N_9492,N_8833,N_8794);
xor U9493 (N_9493,N_8712,N_8857);
and U9494 (N_9494,N_8687,N_8510);
nor U9495 (N_9495,N_8570,N_8824);
nor U9496 (N_9496,N_8732,N_8519);
nand U9497 (N_9497,N_8942,N_8678);
and U9498 (N_9498,N_8752,N_8552);
or U9499 (N_9499,N_8678,N_8621);
nor U9500 (N_9500,N_9144,N_9108);
and U9501 (N_9501,N_9048,N_9275);
and U9502 (N_9502,N_9153,N_9191);
nand U9503 (N_9503,N_9478,N_9098);
or U9504 (N_9504,N_9129,N_9374);
or U9505 (N_9505,N_9002,N_9387);
nand U9506 (N_9506,N_9282,N_9423);
or U9507 (N_9507,N_9458,N_9262);
or U9508 (N_9508,N_9040,N_9461);
nor U9509 (N_9509,N_9091,N_9428);
nor U9510 (N_9510,N_9354,N_9308);
xnor U9511 (N_9511,N_9126,N_9210);
and U9512 (N_9512,N_9231,N_9135);
nand U9513 (N_9513,N_9044,N_9024);
and U9514 (N_9514,N_9399,N_9127);
or U9515 (N_9515,N_9172,N_9036);
nor U9516 (N_9516,N_9485,N_9476);
xor U9517 (N_9517,N_9031,N_9186);
and U9518 (N_9518,N_9089,N_9358);
or U9519 (N_9519,N_9487,N_9051);
xnor U9520 (N_9520,N_9407,N_9234);
and U9521 (N_9521,N_9214,N_9004);
or U9522 (N_9522,N_9371,N_9199);
or U9523 (N_9523,N_9090,N_9192);
or U9524 (N_9524,N_9263,N_9321);
nand U9525 (N_9525,N_9253,N_9203);
nand U9526 (N_9526,N_9352,N_9027);
and U9527 (N_9527,N_9236,N_9136);
or U9528 (N_9528,N_9306,N_9402);
and U9529 (N_9529,N_9336,N_9220);
xnor U9530 (N_9530,N_9472,N_9109);
nor U9531 (N_9531,N_9166,N_9412);
nor U9532 (N_9532,N_9015,N_9491);
or U9533 (N_9533,N_9367,N_9303);
nand U9534 (N_9534,N_9490,N_9056);
nand U9535 (N_9535,N_9190,N_9185);
nand U9536 (N_9536,N_9330,N_9137);
nand U9537 (N_9537,N_9099,N_9328);
nand U9538 (N_9538,N_9322,N_9212);
and U9539 (N_9539,N_9179,N_9434);
or U9540 (N_9540,N_9157,N_9416);
xnor U9541 (N_9541,N_9104,N_9200);
nor U9542 (N_9542,N_9421,N_9224);
nor U9543 (N_9543,N_9218,N_9161);
xnor U9544 (N_9544,N_9267,N_9429);
xor U9545 (N_9545,N_9147,N_9064);
or U9546 (N_9546,N_9038,N_9011);
and U9547 (N_9547,N_9023,N_9414);
nand U9548 (N_9548,N_9084,N_9233);
and U9549 (N_9549,N_9128,N_9422);
and U9550 (N_9550,N_9007,N_9279);
xor U9551 (N_9551,N_9103,N_9286);
and U9552 (N_9552,N_9426,N_9356);
or U9553 (N_9553,N_9293,N_9162);
nor U9554 (N_9554,N_9409,N_9152);
xnor U9555 (N_9555,N_9255,N_9287);
and U9556 (N_9556,N_9397,N_9146);
nor U9557 (N_9557,N_9140,N_9093);
or U9558 (N_9558,N_9442,N_9375);
xnor U9559 (N_9559,N_9009,N_9380);
nor U9560 (N_9560,N_9341,N_9379);
xnor U9561 (N_9561,N_9346,N_9068);
or U9562 (N_9562,N_9437,N_9047);
or U9563 (N_9563,N_9060,N_9022);
and U9564 (N_9564,N_9453,N_9457);
or U9565 (N_9565,N_9494,N_9368);
or U9566 (N_9566,N_9350,N_9477);
or U9567 (N_9567,N_9062,N_9150);
nor U9568 (N_9568,N_9325,N_9235);
nor U9569 (N_9569,N_9378,N_9469);
and U9570 (N_9570,N_9497,N_9259);
nand U9571 (N_9571,N_9138,N_9017);
and U9572 (N_9572,N_9055,N_9329);
or U9573 (N_9573,N_9493,N_9467);
xor U9574 (N_9574,N_9296,N_9304);
nand U9575 (N_9575,N_9386,N_9438);
or U9576 (N_9576,N_9213,N_9250);
nand U9577 (N_9577,N_9447,N_9254);
and U9578 (N_9578,N_9065,N_9488);
nand U9579 (N_9579,N_9499,N_9141);
xnor U9580 (N_9580,N_9156,N_9433);
xnor U9581 (N_9581,N_9432,N_9041);
or U9582 (N_9582,N_9001,N_9405);
or U9583 (N_9583,N_9169,N_9343);
or U9584 (N_9584,N_9435,N_9174);
and U9585 (N_9585,N_9280,N_9077);
and U9586 (N_9586,N_9183,N_9462);
nor U9587 (N_9587,N_9202,N_9324);
nand U9588 (N_9588,N_9078,N_9201);
nand U9589 (N_9589,N_9456,N_9290);
xor U9590 (N_9590,N_9193,N_9082);
or U9591 (N_9591,N_9197,N_9427);
nor U9592 (N_9592,N_9468,N_9385);
xnor U9593 (N_9593,N_9283,N_9219);
or U9594 (N_9594,N_9326,N_9408);
xor U9595 (N_9595,N_9340,N_9317);
xnor U9596 (N_9596,N_9301,N_9067);
xor U9597 (N_9597,N_9208,N_9252);
or U9598 (N_9598,N_9349,N_9071);
or U9599 (N_9599,N_9059,N_9281);
xor U9600 (N_9600,N_9095,N_9413);
and U9601 (N_9601,N_9195,N_9332);
xor U9602 (N_9602,N_9466,N_9285);
xnor U9603 (N_9603,N_9394,N_9196);
nand U9604 (N_9604,N_9066,N_9403);
nand U9605 (N_9605,N_9297,N_9276);
xor U9606 (N_9606,N_9215,N_9204);
and U9607 (N_9607,N_9498,N_9081);
nand U9608 (N_9608,N_9242,N_9481);
or U9609 (N_9609,N_9061,N_9076);
xor U9610 (N_9610,N_9222,N_9168);
or U9611 (N_9611,N_9258,N_9362);
or U9612 (N_9612,N_9240,N_9339);
or U9613 (N_9613,N_9319,N_9058);
nor U9614 (N_9614,N_9268,N_9016);
and U9615 (N_9615,N_9406,N_9392);
xor U9616 (N_9616,N_9446,N_9028);
nand U9617 (N_9617,N_9357,N_9014);
or U9618 (N_9618,N_9449,N_9360);
and U9619 (N_9619,N_9483,N_9170);
nand U9620 (N_9620,N_9010,N_9298);
xnor U9621 (N_9621,N_9480,N_9101);
nor U9622 (N_9622,N_9134,N_9230);
or U9623 (N_9623,N_9092,N_9313);
nor U9624 (N_9624,N_9307,N_9132);
nand U9625 (N_9625,N_9418,N_9455);
nor U9626 (N_9626,N_9316,N_9050);
and U9627 (N_9627,N_9188,N_9112);
and U9628 (N_9628,N_9390,N_9160);
xnor U9629 (N_9629,N_9159,N_9443);
and U9630 (N_9630,N_9072,N_9334);
xor U9631 (N_9631,N_9400,N_9115);
xor U9632 (N_9632,N_9436,N_9155);
nor U9633 (N_9633,N_9391,N_9118);
and U9634 (N_9634,N_9335,N_9232);
nand U9635 (N_9635,N_9020,N_9289);
or U9636 (N_9636,N_9452,N_9331);
or U9637 (N_9637,N_9277,N_9454);
nand U9638 (N_9638,N_9270,N_9474);
nor U9639 (N_9639,N_9294,N_9292);
nor U9640 (N_9640,N_9100,N_9083);
nand U9641 (N_9641,N_9345,N_9122);
or U9642 (N_9642,N_9419,N_9227);
and U9643 (N_9643,N_9229,N_9046);
nand U9644 (N_9644,N_9080,N_9105);
or U9645 (N_9645,N_9029,N_9180);
xor U9646 (N_9646,N_9035,N_9139);
nand U9647 (N_9647,N_9221,N_9353);
xnor U9648 (N_9648,N_9266,N_9057);
or U9649 (N_9649,N_9151,N_9376);
or U9650 (N_9650,N_9181,N_9264);
nand U9651 (N_9651,N_9019,N_9440);
and U9652 (N_9652,N_9359,N_9310);
nor U9653 (N_9653,N_9417,N_9125);
xor U9654 (N_9654,N_9021,N_9177);
nor U9655 (N_9655,N_9025,N_9216);
nor U9656 (N_9656,N_9464,N_9288);
nor U9657 (N_9657,N_9384,N_9261);
xor U9658 (N_9658,N_9030,N_9300);
and U9659 (N_9659,N_9256,N_9148);
or U9660 (N_9660,N_9154,N_9420);
and U9661 (N_9661,N_9363,N_9410);
or U9662 (N_9662,N_9039,N_9311);
xnor U9663 (N_9663,N_9053,N_9257);
nand U9664 (N_9664,N_9470,N_9096);
and U9665 (N_9665,N_9333,N_9026);
xnor U9666 (N_9666,N_9238,N_9320);
and U9667 (N_9667,N_9088,N_9079);
and U9668 (N_9668,N_9106,N_9463);
nor U9669 (N_9669,N_9198,N_9355);
xor U9670 (N_9670,N_9113,N_9111);
and U9671 (N_9671,N_9373,N_9465);
nor U9672 (N_9672,N_9338,N_9348);
nor U9673 (N_9673,N_9475,N_9393);
nor U9674 (N_9674,N_9178,N_9396);
or U9675 (N_9675,N_9094,N_9209);
nor U9676 (N_9676,N_9175,N_9271);
and U9677 (N_9677,N_9187,N_9381);
xnor U9678 (N_9678,N_9239,N_9295);
or U9679 (N_9679,N_9251,N_9123);
nand U9680 (N_9680,N_9116,N_9247);
or U9681 (N_9681,N_9228,N_9377);
nor U9682 (N_9682,N_9073,N_9342);
and U9683 (N_9683,N_9365,N_9244);
and U9684 (N_9684,N_9459,N_9473);
and U9685 (N_9685,N_9347,N_9448);
nand U9686 (N_9686,N_9370,N_9163);
or U9687 (N_9687,N_9114,N_9173);
or U9688 (N_9688,N_9102,N_9149);
and U9689 (N_9689,N_9085,N_9070);
nand U9690 (N_9690,N_9107,N_9404);
nand U9691 (N_9691,N_9217,N_9291);
and U9692 (N_9692,N_9164,N_9124);
or U9693 (N_9693,N_9006,N_9309);
or U9694 (N_9694,N_9351,N_9237);
or U9695 (N_9695,N_9415,N_9344);
and U9696 (N_9696,N_9005,N_9411);
or U9697 (N_9697,N_9119,N_9142);
nand U9698 (N_9698,N_9158,N_9189);
nand U9699 (N_9699,N_9063,N_9226);
nand U9700 (N_9700,N_9207,N_9312);
nand U9701 (N_9701,N_9364,N_9492);
and U9702 (N_9702,N_9120,N_9034);
nand U9703 (N_9703,N_9241,N_9305);
nor U9704 (N_9704,N_9143,N_9398);
and U9705 (N_9705,N_9012,N_9382);
nand U9706 (N_9706,N_9097,N_9495);
nor U9707 (N_9707,N_9260,N_9145);
and U9708 (N_9708,N_9315,N_9327);
or U9709 (N_9709,N_9431,N_9171);
and U9710 (N_9710,N_9117,N_9032);
or U9711 (N_9711,N_9206,N_9450);
or U9712 (N_9712,N_9372,N_9049);
nand U9713 (N_9713,N_9430,N_9245);
nor U9714 (N_9714,N_9424,N_9318);
and U9715 (N_9715,N_9008,N_9075);
and U9716 (N_9716,N_9389,N_9013);
xor U9717 (N_9717,N_9074,N_9274);
and U9718 (N_9718,N_9033,N_9087);
and U9719 (N_9719,N_9043,N_9278);
nor U9720 (N_9720,N_9369,N_9489);
and U9721 (N_9721,N_9225,N_9337);
xnor U9722 (N_9722,N_9484,N_9110);
and U9723 (N_9723,N_9479,N_9052);
xnor U9724 (N_9724,N_9086,N_9176);
xor U9725 (N_9725,N_9482,N_9302);
xnor U9726 (N_9726,N_9441,N_9323);
nand U9727 (N_9727,N_9211,N_9401);
nor U9728 (N_9728,N_9243,N_9000);
nor U9729 (N_9729,N_9246,N_9042);
nor U9730 (N_9730,N_9194,N_9269);
or U9731 (N_9731,N_9018,N_9439);
or U9732 (N_9732,N_9445,N_9265);
xnor U9733 (N_9733,N_9496,N_9223);
or U9734 (N_9734,N_9471,N_9366);
nand U9735 (N_9735,N_9037,N_9069);
nor U9736 (N_9736,N_9249,N_9272);
or U9737 (N_9737,N_9121,N_9383);
xnor U9738 (N_9738,N_9314,N_9133);
and U9739 (N_9739,N_9273,N_9299);
or U9740 (N_9740,N_9451,N_9131);
nor U9741 (N_9741,N_9444,N_9284);
xor U9742 (N_9742,N_9361,N_9388);
xnor U9743 (N_9743,N_9003,N_9460);
or U9744 (N_9744,N_9425,N_9182);
and U9745 (N_9745,N_9167,N_9205);
nor U9746 (N_9746,N_9184,N_9045);
nand U9747 (N_9747,N_9486,N_9130);
and U9748 (N_9748,N_9395,N_9248);
or U9749 (N_9749,N_9165,N_9054);
xor U9750 (N_9750,N_9160,N_9348);
xnor U9751 (N_9751,N_9311,N_9146);
nand U9752 (N_9752,N_9296,N_9235);
nor U9753 (N_9753,N_9027,N_9441);
and U9754 (N_9754,N_9079,N_9371);
or U9755 (N_9755,N_9484,N_9233);
nand U9756 (N_9756,N_9340,N_9256);
nand U9757 (N_9757,N_9411,N_9456);
or U9758 (N_9758,N_9493,N_9084);
and U9759 (N_9759,N_9030,N_9113);
nor U9760 (N_9760,N_9325,N_9101);
nand U9761 (N_9761,N_9145,N_9314);
or U9762 (N_9762,N_9242,N_9152);
nor U9763 (N_9763,N_9153,N_9380);
xor U9764 (N_9764,N_9254,N_9313);
xnor U9765 (N_9765,N_9366,N_9127);
nand U9766 (N_9766,N_9405,N_9392);
and U9767 (N_9767,N_9366,N_9000);
and U9768 (N_9768,N_9291,N_9170);
nor U9769 (N_9769,N_9258,N_9010);
nand U9770 (N_9770,N_9408,N_9086);
or U9771 (N_9771,N_9348,N_9125);
xor U9772 (N_9772,N_9326,N_9461);
or U9773 (N_9773,N_9454,N_9208);
xnor U9774 (N_9774,N_9026,N_9467);
and U9775 (N_9775,N_9211,N_9222);
nor U9776 (N_9776,N_9007,N_9065);
or U9777 (N_9777,N_9072,N_9441);
xor U9778 (N_9778,N_9379,N_9459);
and U9779 (N_9779,N_9065,N_9344);
nand U9780 (N_9780,N_9008,N_9190);
nand U9781 (N_9781,N_9051,N_9145);
nor U9782 (N_9782,N_9126,N_9146);
and U9783 (N_9783,N_9410,N_9414);
nand U9784 (N_9784,N_9138,N_9227);
nor U9785 (N_9785,N_9384,N_9036);
or U9786 (N_9786,N_9139,N_9249);
xor U9787 (N_9787,N_9296,N_9009);
nor U9788 (N_9788,N_9429,N_9030);
or U9789 (N_9789,N_9371,N_9108);
or U9790 (N_9790,N_9260,N_9139);
nand U9791 (N_9791,N_9116,N_9478);
xor U9792 (N_9792,N_9218,N_9100);
nand U9793 (N_9793,N_9217,N_9466);
nor U9794 (N_9794,N_9231,N_9080);
xnor U9795 (N_9795,N_9006,N_9387);
nand U9796 (N_9796,N_9143,N_9235);
nor U9797 (N_9797,N_9341,N_9405);
or U9798 (N_9798,N_9383,N_9428);
nand U9799 (N_9799,N_9339,N_9471);
nand U9800 (N_9800,N_9042,N_9001);
and U9801 (N_9801,N_9142,N_9287);
and U9802 (N_9802,N_9067,N_9189);
xnor U9803 (N_9803,N_9390,N_9001);
nand U9804 (N_9804,N_9290,N_9075);
nor U9805 (N_9805,N_9180,N_9244);
nand U9806 (N_9806,N_9080,N_9098);
and U9807 (N_9807,N_9152,N_9443);
nor U9808 (N_9808,N_9370,N_9005);
nor U9809 (N_9809,N_9241,N_9009);
xnor U9810 (N_9810,N_9437,N_9416);
xnor U9811 (N_9811,N_9013,N_9173);
nand U9812 (N_9812,N_9404,N_9220);
and U9813 (N_9813,N_9261,N_9436);
xor U9814 (N_9814,N_9113,N_9462);
or U9815 (N_9815,N_9334,N_9098);
nand U9816 (N_9816,N_9449,N_9247);
xor U9817 (N_9817,N_9148,N_9478);
xnor U9818 (N_9818,N_9028,N_9312);
nand U9819 (N_9819,N_9109,N_9172);
and U9820 (N_9820,N_9443,N_9030);
nor U9821 (N_9821,N_9361,N_9280);
xor U9822 (N_9822,N_9173,N_9315);
nand U9823 (N_9823,N_9212,N_9224);
and U9824 (N_9824,N_9329,N_9155);
or U9825 (N_9825,N_9001,N_9276);
and U9826 (N_9826,N_9416,N_9093);
xor U9827 (N_9827,N_9391,N_9034);
and U9828 (N_9828,N_9368,N_9055);
xnor U9829 (N_9829,N_9044,N_9190);
or U9830 (N_9830,N_9417,N_9281);
nand U9831 (N_9831,N_9400,N_9273);
nand U9832 (N_9832,N_9310,N_9429);
xnor U9833 (N_9833,N_9145,N_9348);
nor U9834 (N_9834,N_9073,N_9158);
nor U9835 (N_9835,N_9392,N_9051);
and U9836 (N_9836,N_9333,N_9264);
xor U9837 (N_9837,N_9484,N_9199);
and U9838 (N_9838,N_9397,N_9438);
nor U9839 (N_9839,N_9085,N_9398);
nand U9840 (N_9840,N_9259,N_9278);
nor U9841 (N_9841,N_9059,N_9336);
nor U9842 (N_9842,N_9333,N_9351);
nor U9843 (N_9843,N_9125,N_9030);
xor U9844 (N_9844,N_9454,N_9098);
nor U9845 (N_9845,N_9138,N_9040);
xnor U9846 (N_9846,N_9124,N_9271);
nand U9847 (N_9847,N_9210,N_9160);
and U9848 (N_9848,N_9127,N_9242);
xnor U9849 (N_9849,N_9460,N_9127);
nor U9850 (N_9850,N_9441,N_9016);
or U9851 (N_9851,N_9353,N_9171);
nand U9852 (N_9852,N_9330,N_9209);
nor U9853 (N_9853,N_9269,N_9267);
nand U9854 (N_9854,N_9128,N_9186);
nor U9855 (N_9855,N_9201,N_9338);
and U9856 (N_9856,N_9081,N_9206);
and U9857 (N_9857,N_9439,N_9463);
nor U9858 (N_9858,N_9150,N_9159);
or U9859 (N_9859,N_9073,N_9152);
xnor U9860 (N_9860,N_9239,N_9134);
xor U9861 (N_9861,N_9175,N_9202);
nor U9862 (N_9862,N_9394,N_9374);
xor U9863 (N_9863,N_9251,N_9141);
and U9864 (N_9864,N_9123,N_9166);
xor U9865 (N_9865,N_9279,N_9016);
or U9866 (N_9866,N_9095,N_9067);
nor U9867 (N_9867,N_9478,N_9014);
xor U9868 (N_9868,N_9360,N_9153);
or U9869 (N_9869,N_9122,N_9415);
nand U9870 (N_9870,N_9206,N_9167);
nand U9871 (N_9871,N_9313,N_9064);
nand U9872 (N_9872,N_9287,N_9097);
and U9873 (N_9873,N_9342,N_9447);
nor U9874 (N_9874,N_9466,N_9156);
or U9875 (N_9875,N_9289,N_9282);
and U9876 (N_9876,N_9031,N_9019);
nor U9877 (N_9877,N_9327,N_9062);
nand U9878 (N_9878,N_9281,N_9085);
nor U9879 (N_9879,N_9296,N_9343);
xor U9880 (N_9880,N_9025,N_9098);
xor U9881 (N_9881,N_9144,N_9485);
nand U9882 (N_9882,N_9089,N_9234);
nand U9883 (N_9883,N_9074,N_9449);
and U9884 (N_9884,N_9024,N_9015);
nand U9885 (N_9885,N_9013,N_9194);
nor U9886 (N_9886,N_9209,N_9248);
and U9887 (N_9887,N_9061,N_9267);
nor U9888 (N_9888,N_9018,N_9019);
nor U9889 (N_9889,N_9377,N_9051);
nand U9890 (N_9890,N_9205,N_9187);
or U9891 (N_9891,N_9272,N_9415);
xnor U9892 (N_9892,N_9423,N_9448);
nor U9893 (N_9893,N_9482,N_9410);
nor U9894 (N_9894,N_9390,N_9125);
nor U9895 (N_9895,N_9408,N_9046);
or U9896 (N_9896,N_9086,N_9143);
nor U9897 (N_9897,N_9037,N_9443);
xor U9898 (N_9898,N_9117,N_9229);
nand U9899 (N_9899,N_9041,N_9439);
and U9900 (N_9900,N_9355,N_9438);
xor U9901 (N_9901,N_9099,N_9281);
and U9902 (N_9902,N_9282,N_9067);
nand U9903 (N_9903,N_9006,N_9166);
xor U9904 (N_9904,N_9358,N_9333);
nand U9905 (N_9905,N_9164,N_9347);
and U9906 (N_9906,N_9395,N_9101);
and U9907 (N_9907,N_9403,N_9495);
nand U9908 (N_9908,N_9374,N_9402);
xor U9909 (N_9909,N_9404,N_9179);
nand U9910 (N_9910,N_9011,N_9237);
and U9911 (N_9911,N_9159,N_9399);
and U9912 (N_9912,N_9478,N_9479);
nand U9913 (N_9913,N_9103,N_9378);
xor U9914 (N_9914,N_9022,N_9252);
nand U9915 (N_9915,N_9019,N_9456);
nand U9916 (N_9916,N_9252,N_9214);
nand U9917 (N_9917,N_9136,N_9264);
nand U9918 (N_9918,N_9026,N_9087);
nand U9919 (N_9919,N_9114,N_9256);
xor U9920 (N_9920,N_9290,N_9187);
and U9921 (N_9921,N_9348,N_9191);
xnor U9922 (N_9922,N_9406,N_9484);
or U9923 (N_9923,N_9158,N_9130);
xnor U9924 (N_9924,N_9235,N_9449);
or U9925 (N_9925,N_9262,N_9399);
or U9926 (N_9926,N_9020,N_9363);
and U9927 (N_9927,N_9154,N_9281);
nor U9928 (N_9928,N_9097,N_9020);
or U9929 (N_9929,N_9007,N_9010);
nor U9930 (N_9930,N_9141,N_9124);
nand U9931 (N_9931,N_9138,N_9298);
nand U9932 (N_9932,N_9053,N_9481);
nor U9933 (N_9933,N_9447,N_9247);
or U9934 (N_9934,N_9131,N_9152);
and U9935 (N_9935,N_9494,N_9008);
nand U9936 (N_9936,N_9081,N_9188);
xnor U9937 (N_9937,N_9103,N_9074);
and U9938 (N_9938,N_9024,N_9327);
and U9939 (N_9939,N_9274,N_9082);
nor U9940 (N_9940,N_9145,N_9326);
and U9941 (N_9941,N_9130,N_9250);
nor U9942 (N_9942,N_9119,N_9410);
nand U9943 (N_9943,N_9180,N_9433);
xor U9944 (N_9944,N_9071,N_9478);
nor U9945 (N_9945,N_9091,N_9020);
nor U9946 (N_9946,N_9365,N_9098);
nand U9947 (N_9947,N_9000,N_9297);
xnor U9948 (N_9948,N_9166,N_9116);
and U9949 (N_9949,N_9459,N_9298);
and U9950 (N_9950,N_9159,N_9388);
and U9951 (N_9951,N_9216,N_9472);
and U9952 (N_9952,N_9441,N_9056);
and U9953 (N_9953,N_9305,N_9044);
nand U9954 (N_9954,N_9291,N_9452);
nand U9955 (N_9955,N_9200,N_9409);
nor U9956 (N_9956,N_9468,N_9247);
xnor U9957 (N_9957,N_9405,N_9382);
xnor U9958 (N_9958,N_9285,N_9128);
and U9959 (N_9959,N_9059,N_9261);
or U9960 (N_9960,N_9388,N_9015);
or U9961 (N_9961,N_9393,N_9141);
or U9962 (N_9962,N_9108,N_9406);
nor U9963 (N_9963,N_9200,N_9471);
and U9964 (N_9964,N_9361,N_9495);
nand U9965 (N_9965,N_9387,N_9102);
xnor U9966 (N_9966,N_9409,N_9261);
nand U9967 (N_9967,N_9243,N_9384);
or U9968 (N_9968,N_9314,N_9139);
nor U9969 (N_9969,N_9017,N_9165);
nor U9970 (N_9970,N_9385,N_9428);
nor U9971 (N_9971,N_9477,N_9334);
xor U9972 (N_9972,N_9103,N_9178);
and U9973 (N_9973,N_9235,N_9471);
nand U9974 (N_9974,N_9476,N_9047);
nand U9975 (N_9975,N_9347,N_9040);
nor U9976 (N_9976,N_9212,N_9111);
nor U9977 (N_9977,N_9181,N_9359);
nor U9978 (N_9978,N_9255,N_9423);
nor U9979 (N_9979,N_9117,N_9163);
or U9980 (N_9980,N_9004,N_9000);
nand U9981 (N_9981,N_9453,N_9109);
and U9982 (N_9982,N_9343,N_9249);
xnor U9983 (N_9983,N_9220,N_9288);
or U9984 (N_9984,N_9388,N_9211);
nor U9985 (N_9985,N_9258,N_9231);
nand U9986 (N_9986,N_9390,N_9055);
nor U9987 (N_9987,N_9105,N_9466);
or U9988 (N_9988,N_9065,N_9297);
and U9989 (N_9989,N_9356,N_9327);
nor U9990 (N_9990,N_9469,N_9366);
nor U9991 (N_9991,N_9107,N_9066);
nand U9992 (N_9992,N_9061,N_9403);
nor U9993 (N_9993,N_9202,N_9461);
and U9994 (N_9994,N_9002,N_9299);
or U9995 (N_9995,N_9203,N_9214);
xor U9996 (N_9996,N_9445,N_9272);
nand U9997 (N_9997,N_9255,N_9092);
xnor U9998 (N_9998,N_9031,N_9207);
nor U9999 (N_9999,N_9018,N_9237);
nor U10000 (N_10000,N_9726,N_9871);
xor U10001 (N_10001,N_9949,N_9741);
nand U10002 (N_10002,N_9884,N_9752);
nand U10003 (N_10003,N_9642,N_9984);
nor U10004 (N_10004,N_9763,N_9745);
nand U10005 (N_10005,N_9848,N_9817);
or U10006 (N_10006,N_9699,N_9679);
nor U10007 (N_10007,N_9598,N_9669);
and U10008 (N_10008,N_9887,N_9862);
xnor U10009 (N_10009,N_9988,N_9544);
nor U10010 (N_10010,N_9830,N_9567);
and U10011 (N_10011,N_9849,N_9935);
and U10012 (N_10012,N_9555,N_9764);
or U10013 (N_10013,N_9729,N_9748);
or U10014 (N_10014,N_9537,N_9633);
nand U10015 (N_10015,N_9969,N_9883);
xor U10016 (N_10016,N_9979,N_9782);
xor U10017 (N_10017,N_9973,N_9966);
and U10018 (N_10018,N_9825,N_9823);
nand U10019 (N_10019,N_9593,N_9793);
or U10020 (N_10020,N_9612,N_9886);
nand U10021 (N_10021,N_9677,N_9521);
nor U10022 (N_10022,N_9785,N_9653);
nor U10023 (N_10023,N_9970,N_9736);
nor U10024 (N_10024,N_9889,N_9892);
or U10025 (N_10025,N_9963,N_9919);
xnor U10026 (N_10026,N_9820,N_9561);
and U10027 (N_10027,N_9655,N_9890);
or U10028 (N_10028,N_9874,N_9922);
xnor U10029 (N_10029,N_9602,N_9542);
nor U10030 (N_10030,N_9802,N_9814);
or U10031 (N_10031,N_9512,N_9599);
or U10032 (N_10032,N_9604,N_9821);
xnor U10033 (N_10033,N_9616,N_9519);
and U10034 (N_10034,N_9836,N_9549);
and U10035 (N_10035,N_9943,N_9906);
nor U10036 (N_10036,N_9701,N_9639);
nor U10037 (N_10037,N_9546,N_9797);
nor U10038 (N_10038,N_9765,N_9995);
or U10039 (N_10039,N_9875,N_9826);
nand U10040 (N_10040,N_9667,N_9925);
and U10041 (N_10041,N_9861,N_9559);
or U10042 (N_10042,N_9796,N_9761);
and U10043 (N_10043,N_9510,N_9557);
or U10044 (N_10044,N_9914,N_9800);
nand U10045 (N_10045,N_9754,N_9937);
nor U10046 (N_10046,N_9756,N_9877);
nor U10047 (N_10047,N_9851,N_9762);
or U10048 (N_10048,N_9854,N_9516);
and U10049 (N_10049,N_9834,N_9835);
nand U10050 (N_10050,N_9606,N_9938);
and U10051 (N_10051,N_9531,N_9879);
nor U10052 (N_10052,N_9977,N_9818);
nand U10053 (N_10053,N_9511,N_9520);
xnor U10054 (N_10054,N_9528,N_9571);
and U10055 (N_10055,N_9737,N_9658);
nand U10056 (N_10056,N_9790,N_9775);
or U10057 (N_10057,N_9880,N_9731);
xnor U10058 (N_10058,N_9572,N_9698);
nor U10059 (N_10059,N_9855,N_9619);
nor U10060 (N_10060,N_9523,N_9624);
nor U10061 (N_10061,N_9507,N_9703);
and U10062 (N_10062,N_9589,N_9878);
xor U10063 (N_10063,N_9586,N_9770);
or U10064 (N_10064,N_9740,N_9873);
nor U10065 (N_10065,N_9530,N_9755);
and U10066 (N_10066,N_9615,N_9921);
xor U10067 (N_10067,N_9535,N_9576);
and U10068 (N_10068,N_9863,N_9634);
and U10069 (N_10069,N_9774,N_9915);
nand U10070 (N_10070,N_9804,N_9700);
or U10071 (N_10071,N_9758,N_9665);
nand U10072 (N_10072,N_9888,N_9690);
nor U10073 (N_10073,N_9730,N_9974);
or U10074 (N_10074,N_9526,N_9905);
xnor U10075 (N_10075,N_9986,N_9859);
or U10076 (N_10076,N_9837,N_9601);
nor U10077 (N_10077,N_9828,N_9850);
nor U10078 (N_10078,N_9842,N_9527);
or U10079 (N_10079,N_9684,N_9923);
nand U10080 (N_10080,N_9882,N_9865);
or U10081 (N_10081,N_9926,N_9524);
xnor U10082 (N_10082,N_9723,N_9934);
xnor U10083 (N_10083,N_9907,N_9975);
nand U10084 (N_10084,N_9678,N_9607);
xnor U10085 (N_10085,N_9832,N_9783);
and U10086 (N_10086,N_9733,N_9917);
and U10087 (N_10087,N_9674,N_9773);
or U10088 (N_10088,N_9972,N_9580);
xnor U10089 (N_10089,N_9771,N_9694);
and U10090 (N_10090,N_9960,N_9794);
xor U10091 (N_10091,N_9806,N_9784);
or U10092 (N_10092,N_9786,N_9628);
or U10093 (N_10093,N_9803,N_9812);
xnor U10094 (N_10094,N_9727,N_9680);
or U10095 (N_10095,N_9807,N_9713);
nand U10096 (N_10096,N_9902,N_9953);
nor U10097 (N_10097,N_9931,N_9920);
and U10098 (N_10098,N_9985,N_9757);
or U10099 (N_10099,N_9776,N_9725);
or U10100 (N_10100,N_9716,N_9739);
nor U10101 (N_10101,N_9857,N_9569);
or U10102 (N_10102,N_9671,N_9629);
nor U10103 (N_10103,N_9659,N_9707);
nor U10104 (N_10104,N_9839,N_9676);
or U10105 (N_10105,N_9635,N_9864);
nand U10106 (N_10106,N_9867,N_9662);
and U10107 (N_10107,N_9735,N_9556);
nand U10108 (N_10108,N_9632,N_9971);
nor U10109 (N_10109,N_9651,N_9640);
nor U10110 (N_10110,N_9637,N_9533);
nand U10111 (N_10111,N_9989,N_9687);
xor U10112 (N_10112,N_9792,N_9691);
nand U10113 (N_10113,N_9605,N_9688);
xnor U10114 (N_10114,N_9706,N_9777);
and U10115 (N_10115,N_9978,N_9541);
nor U10116 (N_10116,N_9976,N_9927);
nor U10117 (N_10117,N_9718,N_9646);
and U10118 (N_10118,N_9568,N_9621);
nand U10119 (N_10119,N_9538,N_9996);
nor U10120 (N_10120,N_9901,N_9709);
xnor U10121 (N_10121,N_9566,N_9750);
xor U10122 (N_10122,N_9734,N_9636);
xnor U10123 (N_10123,N_9910,N_9697);
or U10124 (N_10124,N_9983,N_9643);
xnor U10125 (N_10125,N_9553,N_9992);
xor U10126 (N_10126,N_9565,N_9772);
xnor U10127 (N_10127,N_9964,N_9824);
xnor U10128 (N_10128,N_9591,N_9522);
nor U10129 (N_10129,N_9578,N_9916);
or U10130 (N_10130,N_9501,N_9894);
or U10131 (N_10131,N_9540,N_9574);
nor U10132 (N_10132,N_9603,N_9592);
and U10133 (N_10133,N_9810,N_9841);
xnor U10134 (N_10134,N_9705,N_9847);
or U10135 (N_10135,N_9717,N_9503);
xnor U10136 (N_10136,N_9958,N_9728);
nand U10137 (N_10137,N_9618,N_9860);
or U10138 (N_10138,N_9672,N_9525);
nor U10139 (N_10139,N_9505,N_9575);
nor U10140 (N_10140,N_9627,N_9959);
nor U10141 (N_10141,N_9647,N_9950);
nand U10142 (N_10142,N_9630,N_9715);
or U10143 (N_10143,N_9809,N_9551);
and U10144 (N_10144,N_9760,N_9869);
and U10145 (N_10145,N_9896,N_9767);
xor U10146 (N_10146,N_9661,N_9948);
or U10147 (N_10147,N_9930,N_9500);
or U10148 (N_10148,N_9840,N_9582);
or U10149 (N_10149,N_9766,N_9881);
xor U10150 (N_10150,N_9614,N_9673);
nand U10151 (N_10151,N_9811,N_9868);
and U10152 (N_10152,N_9514,N_9808);
xor U10153 (N_10153,N_9594,N_9696);
nor U10154 (N_10154,N_9722,N_9670);
nor U10155 (N_10155,N_9648,N_9581);
nand U10156 (N_10156,N_9998,N_9831);
xor U10157 (N_10157,N_9652,N_9845);
xor U10158 (N_10158,N_9595,N_9852);
nor U10159 (N_10159,N_9918,N_9704);
or U10160 (N_10160,N_9720,N_9719);
xnor U10161 (N_10161,N_9798,N_9560);
and U10162 (N_10162,N_9795,N_9675);
nor U10163 (N_10163,N_9980,N_9749);
nor U10164 (N_10164,N_9638,N_9954);
nand U10165 (N_10165,N_9819,N_9957);
nand U10166 (N_10166,N_9912,N_9732);
or U10167 (N_10167,N_9945,N_9746);
and U10168 (N_10168,N_9649,N_9965);
or U10169 (N_10169,N_9872,N_9866);
or U10170 (N_10170,N_9843,N_9801);
xor U10171 (N_10171,N_9885,N_9534);
and U10172 (N_10172,N_9844,N_9816);
xnor U10173 (N_10173,N_9562,N_9623);
xor U10174 (N_10174,N_9631,N_9579);
and U10175 (N_10175,N_9666,N_9588);
or U10176 (N_10176,N_9558,N_9508);
and U10177 (N_10177,N_9714,N_9870);
or U10178 (N_10178,N_9547,N_9759);
nand U10179 (N_10179,N_9781,N_9693);
nor U10180 (N_10180,N_9611,N_9554);
nor U10181 (N_10181,N_9686,N_9682);
nand U10182 (N_10182,N_9813,N_9504);
xor U10183 (N_10183,N_9600,N_9897);
nand U10184 (N_10184,N_9552,N_9550);
or U10185 (N_10185,N_9517,N_9903);
nand U10186 (N_10186,N_9518,N_9545);
or U10187 (N_10187,N_9822,N_9981);
nand U10188 (N_10188,N_9827,N_9940);
nor U10189 (N_10189,N_9532,N_9590);
nand U10190 (N_10190,N_9644,N_9904);
or U10191 (N_10191,N_9788,N_9791);
and U10192 (N_10192,N_9645,N_9641);
or U10193 (N_10193,N_9967,N_9702);
xnor U10194 (N_10194,N_9656,N_9622);
xnor U10195 (N_10195,N_9721,N_9805);
and U10196 (N_10196,N_9924,N_9584);
xnor U10197 (N_10197,N_9929,N_9539);
nor U10198 (N_10198,N_9753,N_9608);
nor U10199 (N_10199,N_9617,N_9650);
xnor U10200 (N_10200,N_9587,N_9942);
xnor U10201 (N_10201,N_9577,N_9899);
and U10202 (N_10202,N_9529,N_9654);
nor U10203 (N_10203,N_9898,N_9932);
and U10204 (N_10204,N_9900,N_9893);
nor U10205 (N_10205,N_9913,N_9597);
or U10206 (N_10206,N_9968,N_9911);
or U10207 (N_10207,N_9928,N_9583);
nand U10208 (N_10208,N_9955,N_9509);
and U10209 (N_10209,N_9543,N_9909);
nor U10210 (N_10210,N_9742,N_9952);
and U10211 (N_10211,N_9668,N_9993);
or U10212 (N_10212,N_9609,N_9939);
nand U10213 (N_10213,N_9692,N_9683);
nand U10214 (N_10214,N_9596,N_9738);
xnor U10215 (N_10215,N_9962,N_9712);
or U10216 (N_10216,N_9513,N_9563);
or U10217 (N_10217,N_9570,N_9858);
nor U10218 (N_10218,N_9711,N_9990);
nand U10219 (N_10219,N_9573,N_9710);
nand U10220 (N_10220,N_9799,N_9502);
or U10221 (N_10221,N_9779,N_9724);
or U10222 (N_10222,N_9564,N_9789);
xnor U10223 (N_10223,N_9876,N_9944);
and U10224 (N_10224,N_9620,N_9780);
and U10225 (N_10225,N_9895,N_9689);
xor U10226 (N_10226,N_9613,N_9838);
and U10227 (N_10227,N_9956,N_9506);
and U10228 (N_10228,N_9994,N_9685);
xnor U10229 (N_10229,N_9947,N_9536);
nor U10230 (N_10230,N_9936,N_9626);
and U10231 (N_10231,N_9768,N_9951);
nand U10232 (N_10232,N_9846,N_9787);
nor U10233 (N_10233,N_9663,N_9856);
and U10234 (N_10234,N_9853,N_9908);
nor U10235 (N_10235,N_9941,N_9744);
nand U10236 (N_10236,N_9778,N_9891);
nor U10237 (N_10237,N_9997,N_9829);
xor U10238 (N_10238,N_9751,N_9664);
or U10239 (N_10239,N_9999,N_9747);
nor U10240 (N_10240,N_9681,N_9548);
xor U10241 (N_10241,N_9695,N_9515);
and U10242 (N_10242,N_9585,N_9933);
nor U10243 (N_10243,N_9833,N_9991);
nor U10244 (N_10244,N_9610,N_9961);
nor U10245 (N_10245,N_9982,N_9946);
nor U10246 (N_10246,N_9743,N_9769);
or U10247 (N_10247,N_9987,N_9625);
xnor U10248 (N_10248,N_9657,N_9708);
nand U10249 (N_10249,N_9815,N_9660);
nand U10250 (N_10250,N_9706,N_9502);
or U10251 (N_10251,N_9959,N_9697);
or U10252 (N_10252,N_9957,N_9954);
nor U10253 (N_10253,N_9807,N_9520);
and U10254 (N_10254,N_9903,N_9885);
nor U10255 (N_10255,N_9552,N_9883);
xor U10256 (N_10256,N_9806,N_9890);
or U10257 (N_10257,N_9676,N_9556);
and U10258 (N_10258,N_9939,N_9561);
and U10259 (N_10259,N_9805,N_9586);
and U10260 (N_10260,N_9986,N_9609);
nand U10261 (N_10261,N_9633,N_9788);
and U10262 (N_10262,N_9504,N_9873);
nand U10263 (N_10263,N_9852,N_9654);
or U10264 (N_10264,N_9596,N_9782);
nor U10265 (N_10265,N_9607,N_9871);
nand U10266 (N_10266,N_9745,N_9774);
nand U10267 (N_10267,N_9676,N_9783);
nor U10268 (N_10268,N_9810,N_9975);
nand U10269 (N_10269,N_9665,N_9820);
and U10270 (N_10270,N_9597,N_9856);
nand U10271 (N_10271,N_9823,N_9616);
or U10272 (N_10272,N_9555,N_9747);
and U10273 (N_10273,N_9819,N_9583);
or U10274 (N_10274,N_9662,N_9720);
nor U10275 (N_10275,N_9601,N_9627);
or U10276 (N_10276,N_9927,N_9968);
nor U10277 (N_10277,N_9597,N_9948);
nand U10278 (N_10278,N_9664,N_9640);
xnor U10279 (N_10279,N_9896,N_9620);
or U10280 (N_10280,N_9754,N_9772);
and U10281 (N_10281,N_9926,N_9705);
and U10282 (N_10282,N_9586,N_9948);
nand U10283 (N_10283,N_9636,N_9813);
or U10284 (N_10284,N_9763,N_9704);
or U10285 (N_10285,N_9507,N_9589);
and U10286 (N_10286,N_9558,N_9866);
nor U10287 (N_10287,N_9864,N_9657);
nand U10288 (N_10288,N_9956,N_9707);
nand U10289 (N_10289,N_9869,N_9957);
nand U10290 (N_10290,N_9870,N_9997);
and U10291 (N_10291,N_9822,N_9971);
nand U10292 (N_10292,N_9800,N_9610);
nor U10293 (N_10293,N_9909,N_9868);
or U10294 (N_10294,N_9524,N_9559);
nand U10295 (N_10295,N_9995,N_9662);
nand U10296 (N_10296,N_9508,N_9891);
nand U10297 (N_10297,N_9883,N_9729);
and U10298 (N_10298,N_9761,N_9577);
nand U10299 (N_10299,N_9753,N_9782);
or U10300 (N_10300,N_9788,N_9566);
nand U10301 (N_10301,N_9612,N_9789);
or U10302 (N_10302,N_9966,N_9945);
or U10303 (N_10303,N_9953,N_9957);
or U10304 (N_10304,N_9520,N_9801);
nor U10305 (N_10305,N_9603,N_9716);
nand U10306 (N_10306,N_9606,N_9890);
nor U10307 (N_10307,N_9891,N_9522);
or U10308 (N_10308,N_9608,N_9555);
nand U10309 (N_10309,N_9838,N_9570);
or U10310 (N_10310,N_9913,N_9574);
nor U10311 (N_10311,N_9534,N_9863);
xnor U10312 (N_10312,N_9826,N_9838);
nand U10313 (N_10313,N_9630,N_9848);
nand U10314 (N_10314,N_9611,N_9645);
xnor U10315 (N_10315,N_9869,N_9925);
nand U10316 (N_10316,N_9597,N_9807);
or U10317 (N_10317,N_9501,N_9963);
and U10318 (N_10318,N_9539,N_9831);
nor U10319 (N_10319,N_9698,N_9790);
nand U10320 (N_10320,N_9528,N_9910);
and U10321 (N_10321,N_9727,N_9574);
xnor U10322 (N_10322,N_9644,N_9677);
and U10323 (N_10323,N_9889,N_9902);
nand U10324 (N_10324,N_9501,N_9654);
xor U10325 (N_10325,N_9621,N_9906);
nor U10326 (N_10326,N_9811,N_9762);
or U10327 (N_10327,N_9758,N_9606);
nor U10328 (N_10328,N_9721,N_9529);
nor U10329 (N_10329,N_9618,N_9982);
and U10330 (N_10330,N_9752,N_9650);
nor U10331 (N_10331,N_9991,N_9845);
or U10332 (N_10332,N_9768,N_9579);
and U10333 (N_10333,N_9755,N_9861);
nand U10334 (N_10334,N_9897,N_9875);
and U10335 (N_10335,N_9775,N_9992);
nor U10336 (N_10336,N_9782,N_9542);
nor U10337 (N_10337,N_9715,N_9856);
and U10338 (N_10338,N_9503,N_9522);
xnor U10339 (N_10339,N_9945,N_9597);
nor U10340 (N_10340,N_9647,N_9784);
xnor U10341 (N_10341,N_9909,N_9634);
and U10342 (N_10342,N_9933,N_9521);
nor U10343 (N_10343,N_9526,N_9925);
and U10344 (N_10344,N_9693,N_9713);
and U10345 (N_10345,N_9587,N_9917);
and U10346 (N_10346,N_9716,N_9546);
and U10347 (N_10347,N_9827,N_9543);
xnor U10348 (N_10348,N_9819,N_9641);
nor U10349 (N_10349,N_9576,N_9604);
or U10350 (N_10350,N_9785,N_9859);
or U10351 (N_10351,N_9957,N_9598);
nor U10352 (N_10352,N_9562,N_9978);
nand U10353 (N_10353,N_9953,N_9730);
and U10354 (N_10354,N_9732,N_9955);
nand U10355 (N_10355,N_9623,N_9712);
nand U10356 (N_10356,N_9916,N_9940);
nand U10357 (N_10357,N_9989,N_9854);
xnor U10358 (N_10358,N_9813,N_9521);
or U10359 (N_10359,N_9788,N_9728);
nor U10360 (N_10360,N_9522,N_9730);
nor U10361 (N_10361,N_9696,N_9704);
and U10362 (N_10362,N_9764,N_9647);
nand U10363 (N_10363,N_9764,N_9708);
or U10364 (N_10364,N_9961,N_9592);
or U10365 (N_10365,N_9557,N_9753);
nand U10366 (N_10366,N_9739,N_9602);
nand U10367 (N_10367,N_9513,N_9530);
xor U10368 (N_10368,N_9701,N_9764);
xor U10369 (N_10369,N_9808,N_9999);
and U10370 (N_10370,N_9519,N_9582);
or U10371 (N_10371,N_9894,N_9697);
nor U10372 (N_10372,N_9915,N_9891);
xnor U10373 (N_10373,N_9700,N_9901);
nand U10374 (N_10374,N_9529,N_9514);
or U10375 (N_10375,N_9985,N_9769);
or U10376 (N_10376,N_9951,N_9884);
and U10377 (N_10377,N_9758,N_9938);
xnor U10378 (N_10378,N_9786,N_9579);
xnor U10379 (N_10379,N_9988,N_9936);
xor U10380 (N_10380,N_9603,N_9807);
nor U10381 (N_10381,N_9826,N_9723);
and U10382 (N_10382,N_9569,N_9558);
nor U10383 (N_10383,N_9665,N_9872);
nand U10384 (N_10384,N_9849,N_9861);
nor U10385 (N_10385,N_9996,N_9619);
nand U10386 (N_10386,N_9545,N_9777);
xor U10387 (N_10387,N_9500,N_9582);
xnor U10388 (N_10388,N_9615,N_9708);
nor U10389 (N_10389,N_9779,N_9716);
nor U10390 (N_10390,N_9899,N_9694);
xor U10391 (N_10391,N_9550,N_9596);
nand U10392 (N_10392,N_9992,N_9977);
nand U10393 (N_10393,N_9685,N_9862);
nor U10394 (N_10394,N_9627,N_9842);
xnor U10395 (N_10395,N_9572,N_9836);
xor U10396 (N_10396,N_9681,N_9765);
or U10397 (N_10397,N_9534,N_9935);
nor U10398 (N_10398,N_9750,N_9721);
and U10399 (N_10399,N_9654,N_9908);
xnor U10400 (N_10400,N_9680,N_9670);
nand U10401 (N_10401,N_9745,N_9909);
nor U10402 (N_10402,N_9948,N_9930);
xor U10403 (N_10403,N_9975,N_9843);
nand U10404 (N_10404,N_9596,N_9797);
and U10405 (N_10405,N_9511,N_9781);
xor U10406 (N_10406,N_9985,N_9715);
nor U10407 (N_10407,N_9733,N_9552);
and U10408 (N_10408,N_9609,N_9711);
xnor U10409 (N_10409,N_9635,N_9792);
nor U10410 (N_10410,N_9795,N_9596);
xnor U10411 (N_10411,N_9639,N_9842);
xnor U10412 (N_10412,N_9658,N_9579);
nor U10413 (N_10413,N_9830,N_9854);
nand U10414 (N_10414,N_9814,N_9909);
or U10415 (N_10415,N_9710,N_9738);
and U10416 (N_10416,N_9876,N_9714);
or U10417 (N_10417,N_9930,N_9802);
xnor U10418 (N_10418,N_9584,N_9819);
nand U10419 (N_10419,N_9762,N_9910);
and U10420 (N_10420,N_9614,N_9802);
or U10421 (N_10421,N_9608,N_9913);
xnor U10422 (N_10422,N_9819,N_9973);
nor U10423 (N_10423,N_9509,N_9902);
or U10424 (N_10424,N_9502,N_9751);
xnor U10425 (N_10425,N_9559,N_9550);
nand U10426 (N_10426,N_9792,N_9694);
and U10427 (N_10427,N_9936,N_9995);
or U10428 (N_10428,N_9549,N_9936);
and U10429 (N_10429,N_9998,N_9533);
or U10430 (N_10430,N_9995,N_9838);
and U10431 (N_10431,N_9520,N_9979);
nor U10432 (N_10432,N_9722,N_9550);
nor U10433 (N_10433,N_9810,N_9979);
or U10434 (N_10434,N_9787,N_9913);
and U10435 (N_10435,N_9638,N_9517);
nand U10436 (N_10436,N_9694,N_9838);
or U10437 (N_10437,N_9778,N_9755);
xor U10438 (N_10438,N_9870,N_9549);
xnor U10439 (N_10439,N_9512,N_9544);
and U10440 (N_10440,N_9993,N_9742);
nand U10441 (N_10441,N_9680,N_9785);
xor U10442 (N_10442,N_9642,N_9826);
xnor U10443 (N_10443,N_9924,N_9783);
and U10444 (N_10444,N_9933,N_9820);
nand U10445 (N_10445,N_9826,N_9714);
nand U10446 (N_10446,N_9919,N_9617);
xor U10447 (N_10447,N_9831,N_9529);
and U10448 (N_10448,N_9551,N_9631);
and U10449 (N_10449,N_9677,N_9908);
nand U10450 (N_10450,N_9825,N_9752);
xnor U10451 (N_10451,N_9816,N_9940);
xor U10452 (N_10452,N_9778,N_9507);
nand U10453 (N_10453,N_9587,N_9729);
and U10454 (N_10454,N_9640,N_9694);
and U10455 (N_10455,N_9651,N_9643);
xor U10456 (N_10456,N_9650,N_9698);
xor U10457 (N_10457,N_9927,N_9678);
xor U10458 (N_10458,N_9693,N_9938);
nand U10459 (N_10459,N_9919,N_9573);
nand U10460 (N_10460,N_9979,N_9564);
or U10461 (N_10461,N_9613,N_9774);
and U10462 (N_10462,N_9521,N_9841);
nor U10463 (N_10463,N_9996,N_9807);
and U10464 (N_10464,N_9867,N_9877);
nand U10465 (N_10465,N_9722,N_9578);
nand U10466 (N_10466,N_9951,N_9717);
and U10467 (N_10467,N_9723,N_9685);
or U10468 (N_10468,N_9614,N_9801);
xor U10469 (N_10469,N_9500,N_9955);
and U10470 (N_10470,N_9588,N_9822);
and U10471 (N_10471,N_9968,N_9942);
xor U10472 (N_10472,N_9662,N_9562);
nand U10473 (N_10473,N_9877,N_9802);
and U10474 (N_10474,N_9631,N_9899);
and U10475 (N_10475,N_9800,N_9624);
xnor U10476 (N_10476,N_9630,N_9956);
and U10477 (N_10477,N_9627,N_9666);
nor U10478 (N_10478,N_9869,N_9658);
nand U10479 (N_10479,N_9664,N_9592);
nor U10480 (N_10480,N_9860,N_9980);
and U10481 (N_10481,N_9628,N_9805);
and U10482 (N_10482,N_9791,N_9596);
or U10483 (N_10483,N_9682,N_9890);
and U10484 (N_10484,N_9537,N_9961);
nor U10485 (N_10485,N_9728,N_9547);
nand U10486 (N_10486,N_9877,N_9796);
xnor U10487 (N_10487,N_9890,N_9619);
or U10488 (N_10488,N_9856,N_9757);
nand U10489 (N_10489,N_9890,N_9973);
xor U10490 (N_10490,N_9583,N_9899);
or U10491 (N_10491,N_9990,N_9932);
xnor U10492 (N_10492,N_9809,N_9927);
xor U10493 (N_10493,N_9757,N_9841);
nand U10494 (N_10494,N_9537,N_9892);
nor U10495 (N_10495,N_9929,N_9564);
nor U10496 (N_10496,N_9837,N_9543);
nand U10497 (N_10497,N_9679,N_9660);
nor U10498 (N_10498,N_9508,N_9923);
xnor U10499 (N_10499,N_9744,N_9808);
or U10500 (N_10500,N_10117,N_10041);
nand U10501 (N_10501,N_10161,N_10307);
xor U10502 (N_10502,N_10459,N_10098);
and U10503 (N_10503,N_10067,N_10440);
xnor U10504 (N_10504,N_10004,N_10039);
nor U10505 (N_10505,N_10411,N_10034);
nand U10506 (N_10506,N_10460,N_10447);
nor U10507 (N_10507,N_10236,N_10484);
xor U10508 (N_10508,N_10010,N_10432);
or U10509 (N_10509,N_10172,N_10265);
or U10510 (N_10510,N_10143,N_10452);
and U10511 (N_10511,N_10349,N_10178);
xnor U10512 (N_10512,N_10188,N_10366);
and U10513 (N_10513,N_10457,N_10306);
or U10514 (N_10514,N_10225,N_10289);
and U10515 (N_10515,N_10191,N_10492);
xor U10516 (N_10516,N_10419,N_10444);
and U10517 (N_10517,N_10019,N_10243);
and U10518 (N_10518,N_10248,N_10240);
and U10519 (N_10519,N_10399,N_10121);
and U10520 (N_10520,N_10094,N_10272);
or U10521 (N_10521,N_10130,N_10007);
xor U10522 (N_10522,N_10071,N_10477);
xnor U10523 (N_10523,N_10220,N_10209);
xor U10524 (N_10524,N_10138,N_10278);
or U10525 (N_10525,N_10346,N_10403);
nor U10526 (N_10526,N_10396,N_10320);
or U10527 (N_10527,N_10028,N_10398);
or U10528 (N_10528,N_10113,N_10033);
or U10529 (N_10529,N_10479,N_10343);
and U10530 (N_10530,N_10057,N_10302);
nand U10531 (N_10531,N_10131,N_10363);
and U10532 (N_10532,N_10458,N_10401);
xor U10533 (N_10533,N_10304,N_10173);
nor U10534 (N_10534,N_10352,N_10029);
nor U10535 (N_10535,N_10405,N_10323);
nand U10536 (N_10536,N_10005,N_10160);
and U10537 (N_10537,N_10342,N_10139);
and U10538 (N_10538,N_10371,N_10031);
and U10539 (N_10539,N_10074,N_10192);
and U10540 (N_10540,N_10449,N_10042);
nand U10541 (N_10541,N_10495,N_10344);
or U10542 (N_10542,N_10051,N_10456);
xor U10543 (N_10543,N_10322,N_10169);
nor U10544 (N_10544,N_10496,N_10165);
xor U10545 (N_10545,N_10470,N_10391);
or U10546 (N_10546,N_10497,N_10217);
nand U10547 (N_10547,N_10055,N_10214);
and U10548 (N_10548,N_10354,N_10068);
or U10549 (N_10549,N_10049,N_10083);
xor U10550 (N_10550,N_10390,N_10355);
xor U10551 (N_10551,N_10327,N_10455);
and U10552 (N_10552,N_10294,N_10095);
or U10553 (N_10553,N_10413,N_10158);
nand U10554 (N_10554,N_10485,N_10284);
or U10555 (N_10555,N_10246,N_10385);
and U10556 (N_10556,N_10312,N_10003);
nor U10557 (N_10557,N_10205,N_10065);
and U10558 (N_10558,N_10383,N_10233);
nand U10559 (N_10559,N_10333,N_10252);
nor U10560 (N_10560,N_10461,N_10254);
or U10561 (N_10561,N_10287,N_10100);
nand U10562 (N_10562,N_10199,N_10176);
nor U10563 (N_10563,N_10469,N_10271);
or U10564 (N_10564,N_10298,N_10081);
nand U10565 (N_10565,N_10086,N_10367);
or U10566 (N_10566,N_10101,N_10221);
or U10567 (N_10567,N_10238,N_10446);
nor U10568 (N_10568,N_10465,N_10219);
xor U10569 (N_10569,N_10097,N_10054);
nand U10570 (N_10570,N_10499,N_10247);
nand U10571 (N_10571,N_10187,N_10303);
nand U10572 (N_10572,N_10464,N_10080);
and U10573 (N_10573,N_10291,N_10185);
or U10574 (N_10574,N_10112,N_10009);
and U10575 (N_10575,N_10197,N_10227);
nor U10576 (N_10576,N_10076,N_10114);
nor U10577 (N_10577,N_10285,N_10082);
xor U10578 (N_10578,N_10276,N_10239);
nor U10579 (N_10579,N_10436,N_10293);
nand U10580 (N_10580,N_10070,N_10423);
nand U10581 (N_10581,N_10348,N_10351);
nand U10582 (N_10582,N_10230,N_10339);
nor U10583 (N_10583,N_10017,N_10373);
nand U10584 (N_10584,N_10262,N_10153);
xor U10585 (N_10585,N_10453,N_10353);
and U10586 (N_10586,N_10483,N_10222);
nor U10587 (N_10587,N_10384,N_10229);
xor U10588 (N_10588,N_10395,N_10059);
and U10589 (N_10589,N_10183,N_10430);
nand U10590 (N_10590,N_10151,N_10001);
nand U10591 (N_10591,N_10467,N_10155);
nor U10592 (N_10592,N_10345,N_10089);
and U10593 (N_10593,N_10073,N_10388);
nand U10594 (N_10594,N_10266,N_10387);
or U10595 (N_10595,N_10494,N_10426);
xor U10596 (N_10596,N_10107,N_10370);
or U10597 (N_10597,N_10179,N_10206);
nand U10598 (N_10598,N_10011,N_10027);
and U10599 (N_10599,N_10000,N_10428);
nand U10600 (N_10600,N_10475,N_10064);
xnor U10601 (N_10601,N_10324,N_10148);
nor U10602 (N_10602,N_10021,N_10232);
nor U10603 (N_10603,N_10048,N_10462);
and U10604 (N_10604,N_10487,N_10002);
xnor U10605 (N_10605,N_10256,N_10255);
nor U10606 (N_10606,N_10066,N_10317);
and U10607 (N_10607,N_10441,N_10063);
nand U10608 (N_10608,N_10123,N_10099);
and U10609 (N_10609,N_10044,N_10120);
nand U10610 (N_10610,N_10418,N_10136);
or U10611 (N_10611,N_10115,N_10326);
and U10612 (N_10612,N_10321,N_10024);
nand U10613 (N_10613,N_10415,N_10164);
or U10614 (N_10614,N_10159,N_10092);
nand U10615 (N_10615,N_10290,N_10362);
or U10616 (N_10616,N_10407,N_10110);
and U10617 (N_10617,N_10231,N_10282);
nor U10618 (N_10618,N_10375,N_10102);
xor U10619 (N_10619,N_10319,N_10075);
or U10620 (N_10620,N_10315,N_10380);
and U10621 (N_10621,N_10417,N_10147);
and U10622 (N_10622,N_10168,N_10128);
nor U10623 (N_10623,N_10141,N_10486);
and U10624 (N_10624,N_10313,N_10196);
nor U10625 (N_10625,N_10267,N_10329);
or U10626 (N_10626,N_10061,N_10087);
and U10627 (N_10627,N_10166,N_10184);
nor U10628 (N_10628,N_10406,N_10400);
or U10629 (N_10629,N_10275,N_10498);
nor U10630 (N_10630,N_10242,N_10263);
nand U10631 (N_10631,N_10394,N_10218);
and U10632 (N_10632,N_10376,N_10295);
nor U10633 (N_10633,N_10198,N_10338);
xor U10634 (N_10634,N_10364,N_10281);
or U10635 (N_10635,N_10170,N_10045);
and U10636 (N_10636,N_10157,N_10473);
nor U10637 (N_10637,N_10186,N_10274);
or U10638 (N_10638,N_10062,N_10251);
and U10639 (N_10639,N_10250,N_10125);
or U10640 (N_10640,N_10253,N_10325);
nand U10641 (N_10641,N_10018,N_10382);
and U10642 (N_10642,N_10189,N_10269);
xnor U10643 (N_10643,N_10069,N_10493);
nor U10644 (N_10644,N_10084,N_10297);
nor U10645 (N_10645,N_10361,N_10026);
nor U10646 (N_10646,N_10305,N_10127);
nand U10647 (N_10647,N_10369,N_10480);
and U10648 (N_10648,N_10410,N_10133);
nand U10649 (N_10649,N_10234,N_10414);
nor U10650 (N_10650,N_10038,N_10207);
and U10651 (N_10651,N_10438,N_10341);
nor U10652 (N_10652,N_10052,N_10202);
and U10653 (N_10653,N_10135,N_10137);
and U10654 (N_10654,N_10091,N_10105);
nor U10655 (N_10655,N_10194,N_10235);
or U10656 (N_10656,N_10213,N_10118);
nand U10657 (N_10657,N_10175,N_10163);
or U10658 (N_10658,N_10488,N_10204);
nor U10659 (N_10659,N_10442,N_10037);
xor U10660 (N_10660,N_10443,N_10434);
or U10661 (N_10661,N_10360,N_10020);
or U10662 (N_10662,N_10425,N_10122);
and U10663 (N_10663,N_10016,N_10310);
xnor U10664 (N_10664,N_10119,N_10350);
xor U10665 (N_10665,N_10124,N_10299);
xnor U10666 (N_10666,N_10145,N_10181);
or U10667 (N_10667,N_10015,N_10149);
xnor U10668 (N_10668,N_10211,N_10273);
or U10669 (N_10669,N_10331,N_10193);
or U10670 (N_10670,N_10481,N_10212);
nor U10671 (N_10671,N_10190,N_10357);
xnor U10672 (N_10672,N_10022,N_10103);
nor U10673 (N_10673,N_10144,N_10337);
or U10674 (N_10674,N_10402,N_10241);
or U10675 (N_10675,N_10270,N_10142);
xor U10676 (N_10676,N_10301,N_10226);
or U10677 (N_10677,N_10359,N_10090);
nor U10678 (N_10678,N_10358,N_10283);
nor U10679 (N_10679,N_10468,N_10182);
nor U10680 (N_10680,N_10330,N_10146);
nand U10681 (N_10681,N_10008,N_10152);
nor U10682 (N_10682,N_10032,N_10108);
nand U10683 (N_10683,N_10318,N_10311);
or U10684 (N_10684,N_10264,N_10316);
or U10685 (N_10685,N_10215,N_10424);
nor U10686 (N_10686,N_10463,N_10258);
or U10687 (N_10687,N_10379,N_10368);
nor U10688 (N_10688,N_10445,N_10286);
nand U10689 (N_10689,N_10047,N_10261);
nor U10690 (N_10690,N_10386,N_10309);
xnor U10691 (N_10691,N_10056,N_10340);
xor U10692 (N_10692,N_10435,N_10377);
or U10693 (N_10693,N_10195,N_10454);
xnor U10694 (N_10694,N_10132,N_10334);
or U10695 (N_10695,N_10431,N_10035);
and U10696 (N_10696,N_10288,N_10156);
or U10697 (N_10697,N_10374,N_10397);
xor U10698 (N_10698,N_10466,N_10471);
and U10699 (N_10699,N_10308,N_10347);
and U10700 (N_10700,N_10208,N_10277);
nor U10701 (N_10701,N_10096,N_10292);
nor U10702 (N_10702,N_10356,N_10201);
or U10703 (N_10703,N_10328,N_10237);
nor U10704 (N_10704,N_10408,N_10088);
xnor U10705 (N_10705,N_10180,N_10392);
nor U10706 (N_10706,N_10420,N_10072);
and U10707 (N_10707,N_10116,N_10154);
nor U10708 (N_10708,N_10314,N_10216);
or U10709 (N_10709,N_10177,N_10476);
and U10710 (N_10710,N_10409,N_10381);
xor U10711 (N_10711,N_10060,N_10279);
or U10712 (N_10712,N_10260,N_10259);
or U10713 (N_10713,N_10421,N_10489);
nor U10714 (N_10714,N_10104,N_10058);
or U10715 (N_10715,N_10013,N_10245);
nand U10716 (N_10716,N_10474,N_10404);
and U10717 (N_10717,N_10257,N_10300);
and U10718 (N_10718,N_10043,N_10249);
nand U10719 (N_10719,N_10450,N_10053);
and U10720 (N_10720,N_10224,N_10296);
nand U10721 (N_10721,N_10244,N_10046);
nor U10722 (N_10722,N_10437,N_10014);
nand U10723 (N_10723,N_10111,N_10150);
nor U10724 (N_10724,N_10280,N_10490);
nor U10725 (N_10725,N_10167,N_10223);
xnor U10726 (N_10726,N_10389,N_10422);
and U10727 (N_10727,N_10040,N_10030);
and U10728 (N_10728,N_10429,N_10482);
nand U10729 (N_10729,N_10079,N_10085);
or U10730 (N_10730,N_10203,N_10025);
nor U10731 (N_10731,N_10472,N_10134);
xnor U10732 (N_10732,N_10210,N_10393);
and U10733 (N_10733,N_10416,N_10378);
nand U10734 (N_10734,N_10200,N_10174);
or U10735 (N_10735,N_10336,N_10106);
and U10736 (N_10736,N_10171,N_10126);
or U10737 (N_10737,N_10335,N_10491);
or U10738 (N_10738,N_10078,N_10412);
xnor U10739 (N_10739,N_10372,N_10332);
nor U10740 (N_10740,N_10427,N_10228);
xor U10741 (N_10741,N_10433,N_10140);
nand U10742 (N_10742,N_10023,N_10162);
and U10743 (N_10743,N_10006,N_10448);
and U10744 (N_10744,N_10268,N_10451);
or U10745 (N_10745,N_10036,N_10077);
xor U10746 (N_10746,N_10093,N_10109);
or U10747 (N_10747,N_10050,N_10478);
and U10748 (N_10748,N_10012,N_10439);
or U10749 (N_10749,N_10129,N_10365);
nor U10750 (N_10750,N_10335,N_10029);
or U10751 (N_10751,N_10105,N_10488);
xor U10752 (N_10752,N_10263,N_10426);
xor U10753 (N_10753,N_10063,N_10215);
xnor U10754 (N_10754,N_10164,N_10248);
and U10755 (N_10755,N_10049,N_10134);
and U10756 (N_10756,N_10290,N_10377);
or U10757 (N_10757,N_10043,N_10227);
and U10758 (N_10758,N_10142,N_10239);
nand U10759 (N_10759,N_10436,N_10310);
or U10760 (N_10760,N_10442,N_10084);
nand U10761 (N_10761,N_10326,N_10109);
nor U10762 (N_10762,N_10030,N_10075);
and U10763 (N_10763,N_10244,N_10472);
nand U10764 (N_10764,N_10119,N_10101);
nand U10765 (N_10765,N_10241,N_10360);
nor U10766 (N_10766,N_10448,N_10022);
nor U10767 (N_10767,N_10480,N_10396);
or U10768 (N_10768,N_10264,N_10296);
nor U10769 (N_10769,N_10165,N_10133);
nand U10770 (N_10770,N_10090,N_10297);
or U10771 (N_10771,N_10196,N_10197);
and U10772 (N_10772,N_10162,N_10383);
xnor U10773 (N_10773,N_10258,N_10115);
nand U10774 (N_10774,N_10173,N_10406);
nand U10775 (N_10775,N_10191,N_10197);
nor U10776 (N_10776,N_10281,N_10465);
or U10777 (N_10777,N_10149,N_10490);
and U10778 (N_10778,N_10225,N_10099);
nor U10779 (N_10779,N_10163,N_10394);
nor U10780 (N_10780,N_10386,N_10271);
nand U10781 (N_10781,N_10162,N_10064);
nor U10782 (N_10782,N_10119,N_10479);
or U10783 (N_10783,N_10481,N_10157);
or U10784 (N_10784,N_10035,N_10096);
xnor U10785 (N_10785,N_10076,N_10371);
nor U10786 (N_10786,N_10260,N_10340);
xnor U10787 (N_10787,N_10281,N_10059);
and U10788 (N_10788,N_10145,N_10110);
nand U10789 (N_10789,N_10318,N_10499);
or U10790 (N_10790,N_10202,N_10097);
or U10791 (N_10791,N_10052,N_10170);
nand U10792 (N_10792,N_10055,N_10379);
or U10793 (N_10793,N_10121,N_10168);
nand U10794 (N_10794,N_10147,N_10154);
nor U10795 (N_10795,N_10168,N_10172);
or U10796 (N_10796,N_10228,N_10110);
nand U10797 (N_10797,N_10273,N_10405);
nand U10798 (N_10798,N_10436,N_10308);
and U10799 (N_10799,N_10016,N_10136);
xor U10800 (N_10800,N_10326,N_10014);
xnor U10801 (N_10801,N_10105,N_10108);
and U10802 (N_10802,N_10293,N_10301);
nor U10803 (N_10803,N_10322,N_10083);
or U10804 (N_10804,N_10185,N_10377);
and U10805 (N_10805,N_10303,N_10292);
nor U10806 (N_10806,N_10183,N_10349);
and U10807 (N_10807,N_10184,N_10402);
nor U10808 (N_10808,N_10420,N_10176);
and U10809 (N_10809,N_10147,N_10081);
nor U10810 (N_10810,N_10386,N_10007);
nand U10811 (N_10811,N_10197,N_10147);
nor U10812 (N_10812,N_10342,N_10425);
nand U10813 (N_10813,N_10187,N_10398);
nand U10814 (N_10814,N_10095,N_10126);
and U10815 (N_10815,N_10121,N_10410);
xnor U10816 (N_10816,N_10227,N_10259);
xnor U10817 (N_10817,N_10172,N_10432);
or U10818 (N_10818,N_10253,N_10340);
nor U10819 (N_10819,N_10010,N_10026);
nor U10820 (N_10820,N_10461,N_10399);
xor U10821 (N_10821,N_10252,N_10018);
nand U10822 (N_10822,N_10453,N_10364);
or U10823 (N_10823,N_10176,N_10023);
nand U10824 (N_10824,N_10152,N_10412);
nand U10825 (N_10825,N_10025,N_10424);
and U10826 (N_10826,N_10214,N_10425);
nor U10827 (N_10827,N_10201,N_10192);
and U10828 (N_10828,N_10379,N_10012);
or U10829 (N_10829,N_10207,N_10243);
nor U10830 (N_10830,N_10046,N_10497);
and U10831 (N_10831,N_10205,N_10206);
xor U10832 (N_10832,N_10134,N_10275);
nand U10833 (N_10833,N_10422,N_10470);
and U10834 (N_10834,N_10418,N_10226);
or U10835 (N_10835,N_10157,N_10485);
and U10836 (N_10836,N_10161,N_10159);
and U10837 (N_10837,N_10324,N_10021);
nor U10838 (N_10838,N_10499,N_10363);
nand U10839 (N_10839,N_10128,N_10211);
and U10840 (N_10840,N_10264,N_10456);
nand U10841 (N_10841,N_10023,N_10486);
nand U10842 (N_10842,N_10445,N_10452);
xnor U10843 (N_10843,N_10318,N_10045);
or U10844 (N_10844,N_10036,N_10324);
xnor U10845 (N_10845,N_10464,N_10416);
or U10846 (N_10846,N_10327,N_10108);
xnor U10847 (N_10847,N_10264,N_10124);
nor U10848 (N_10848,N_10493,N_10445);
and U10849 (N_10849,N_10080,N_10484);
or U10850 (N_10850,N_10061,N_10236);
xnor U10851 (N_10851,N_10320,N_10012);
nor U10852 (N_10852,N_10479,N_10104);
nand U10853 (N_10853,N_10069,N_10005);
xor U10854 (N_10854,N_10181,N_10053);
xor U10855 (N_10855,N_10343,N_10024);
xor U10856 (N_10856,N_10401,N_10103);
and U10857 (N_10857,N_10426,N_10393);
nand U10858 (N_10858,N_10061,N_10210);
xor U10859 (N_10859,N_10193,N_10170);
and U10860 (N_10860,N_10098,N_10380);
nand U10861 (N_10861,N_10288,N_10032);
or U10862 (N_10862,N_10229,N_10029);
nor U10863 (N_10863,N_10483,N_10281);
and U10864 (N_10864,N_10460,N_10265);
xnor U10865 (N_10865,N_10488,N_10171);
nor U10866 (N_10866,N_10429,N_10457);
and U10867 (N_10867,N_10066,N_10106);
nor U10868 (N_10868,N_10348,N_10317);
nand U10869 (N_10869,N_10081,N_10231);
nor U10870 (N_10870,N_10143,N_10167);
or U10871 (N_10871,N_10054,N_10174);
nor U10872 (N_10872,N_10281,N_10264);
nand U10873 (N_10873,N_10250,N_10060);
nand U10874 (N_10874,N_10352,N_10092);
nand U10875 (N_10875,N_10165,N_10334);
or U10876 (N_10876,N_10365,N_10362);
and U10877 (N_10877,N_10083,N_10289);
or U10878 (N_10878,N_10276,N_10011);
nand U10879 (N_10879,N_10241,N_10126);
or U10880 (N_10880,N_10366,N_10485);
or U10881 (N_10881,N_10389,N_10143);
nand U10882 (N_10882,N_10338,N_10036);
or U10883 (N_10883,N_10461,N_10096);
xor U10884 (N_10884,N_10473,N_10387);
and U10885 (N_10885,N_10069,N_10001);
nand U10886 (N_10886,N_10371,N_10379);
nand U10887 (N_10887,N_10044,N_10440);
and U10888 (N_10888,N_10314,N_10000);
nand U10889 (N_10889,N_10340,N_10003);
xor U10890 (N_10890,N_10428,N_10279);
xnor U10891 (N_10891,N_10027,N_10427);
xor U10892 (N_10892,N_10171,N_10096);
xor U10893 (N_10893,N_10116,N_10234);
or U10894 (N_10894,N_10443,N_10023);
and U10895 (N_10895,N_10379,N_10351);
nor U10896 (N_10896,N_10451,N_10393);
nand U10897 (N_10897,N_10450,N_10426);
nand U10898 (N_10898,N_10342,N_10178);
xor U10899 (N_10899,N_10415,N_10453);
nor U10900 (N_10900,N_10228,N_10321);
nor U10901 (N_10901,N_10058,N_10068);
nand U10902 (N_10902,N_10406,N_10401);
or U10903 (N_10903,N_10123,N_10261);
and U10904 (N_10904,N_10399,N_10330);
xnor U10905 (N_10905,N_10176,N_10041);
nor U10906 (N_10906,N_10124,N_10472);
or U10907 (N_10907,N_10177,N_10443);
and U10908 (N_10908,N_10307,N_10106);
xnor U10909 (N_10909,N_10185,N_10289);
nor U10910 (N_10910,N_10418,N_10296);
nand U10911 (N_10911,N_10119,N_10197);
nand U10912 (N_10912,N_10388,N_10457);
or U10913 (N_10913,N_10215,N_10050);
nor U10914 (N_10914,N_10470,N_10010);
or U10915 (N_10915,N_10080,N_10424);
and U10916 (N_10916,N_10046,N_10257);
nand U10917 (N_10917,N_10302,N_10009);
and U10918 (N_10918,N_10121,N_10344);
nor U10919 (N_10919,N_10166,N_10416);
nor U10920 (N_10920,N_10350,N_10004);
nor U10921 (N_10921,N_10285,N_10066);
or U10922 (N_10922,N_10300,N_10163);
nor U10923 (N_10923,N_10453,N_10246);
nand U10924 (N_10924,N_10069,N_10017);
and U10925 (N_10925,N_10323,N_10057);
nor U10926 (N_10926,N_10493,N_10162);
nand U10927 (N_10927,N_10204,N_10011);
nand U10928 (N_10928,N_10445,N_10128);
and U10929 (N_10929,N_10325,N_10287);
and U10930 (N_10930,N_10046,N_10369);
nand U10931 (N_10931,N_10420,N_10412);
xor U10932 (N_10932,N_10416,N_10447);
xor U10933 (N_10933,N_10442,N_10433);
and U10934 (N_10934,N_10294,N_10289);
and U10935 (N_10935,N_10419,N_10253);
or U10936 (N_10936,N_10383,N_10207);
xor U10937 (N_10937,N_10264,N_10390);
xnor U10938 (N_10938,N_10310,N_10179);
or U10939 (N_10939,N_10286,N_10160);
or U10940 (N_10940,N_10043,N_10484);
and U10941 (N_10941,N_10005,N_10351);
nor U10942 (N_10942,N_10359,N_10481);
or U10943 (N_10943,N_10304,N_10421);
xnor U10944 (N_10944,N_10373,N_10395);
nand U10945 (N_10945,N_10005,N_10391);
and U10946 (N_10946,N_10064,N_10426);
or U10947 (N_10947,N_10495,N_10181);
nand U10948 (N_10948,N_10117,N_10093);
xnor U10949 (N_10949,N_10107,N_10483);
and U10950 (N_10950,N_10076,N_10414);
or U10951 (N_10951,N_10285,N_10488);
nor U10952 (N_10952,N_10124,N_10486);
or U10953 (N_10953,N_10486,N_10332);
or U10954 (N_10954,N_10266,N_10308);
and U10955 (N_10955,N_10031,N_10343);
and U10956 (N_10956,N_10148,N_10177);
and U10957 (N_10957,N_10479,N_10243);
nand U10958 (N_10958,N_10202,N_10251);
xor U10959 (N_10959,N_10394,N_10499);
xor U10960 (N_10960,N_10056,N_10079);
and U10961 (N_10961,N_10245,N_10405);
or U10962 (N_10962,N_10472,N_10117);
and U10963 (N_10963,N_10448,N_10146);
nor U10964 (N_10964,N_10432,N_10194);
nand U10965 (N_10965,N_10280,N_10135);
nor U10966 (N_10966,N_10397,N_10193);
nor U10967 (N_10967,N_10372,N_10377);
and U10968 (N_10968,N_10348,N_10374);
xnor U10969 (N_10969,N_10361,N_10255);
and U10970 (N_10970,N_10294,N_10060);
xnor U10971 (N_10971,N_10192,N_10444);
xor U10972 (N_10972,N_10266,N_10366);
nor U10973 (N_10973,N_10282,N_10483);
or U10974 (N_10974,N_10002,N_10302);
and U10975 (N_10975,N_10067,N_10102);
or U10976 (N_10976,N_10389,N_10351);
xor U10977 (N_10977,N_10047,N_10072);
nand U10978 (N_10978,N_10445,N_10028);
or U10979 (N_10979,N_10294,N_10174);
nand U10980 (N_10980,N_10192,N_10177);
and U10981 (N_10981,N_10270,N_10417);
nand U10982 (N_10982,N_10333,N_10453);
and U10983 (N_10983,N_10365,N_10078);
nor U10984 (N_10984,N_10216,N_10099);
nor U10985 (N_10985,N_10462,N_10144);
nor U10986 (N_10986,N_10323,N_10483);
and U10987 (N_10987,N_10351,N_10230);
nand U10988 (N_10988,N_10049,N_10012);
xnor U10989 (N_10989,N_10353,N_10152);
nor U10990 (N_10990,N_10187,N_10478);
xor U10991 (N_10991,N_10442,N_10458);
xnor U10992 (N_10992,N_10219,N_10271);
xnor U10993 (N_10993,N_10260,N_10020);
nand U10994 (N_10994,N_10240,N_10176);
nor U10995 (N_10995,N_10020,N_10453);
xnor U10996 (N_10996,N_10014,N_10312);
nor U10997 (N_10997,N_10163,N_10008);
nand U10998 (N_10998,N_10141,N_10385);
and U10999 (N_10999,N_10330,N_10467);
xnor U11000 (N_11000,N_10820,N_10952);
nor U11001 (N_11001,N_10953,N_10742);
nand U11002 (N_11002,N_10984,N_10580);
nand U11003 (N_11003,N_10515,N_10655);
or U11004 (N_11004,N_10922,N_10665);
xor U11005 (N_11005,N_10969,N_10573);
xnor U11006 (N_11006,N_10816,N_10618);
xor U11007 (N_11007,N_10638,N_10623);
and U11008 (N_11008,N_10729,N_10710);
nor U11009 (N_11009,N_10595,N_10990);
and U11010 (N_11010,N_10712,N_10872);
xnor U11011 (N_11011,N_10502,N_10724);
xnor U11012 (N_11012,N_10869,N_10643);
and U11013 (N_11013,N_10864,N_10589);
nand U11014 (N_11014,N_10855,N_10661);
xor U11015 (N_11015,N_10780,N_10648);
or U11016 (N_11016,N_10908,N_10613);
nor U11017 (N_11017,N_10582,N_10559);
xor U11018 (N_11018,N_10528,N_10839);
nand U11019 (N_11019,N_10663,N_10609);
nor U11020 (N_11020,N_10994,N_10986);
nand U11021 (N_11021,N_10856,N_10555);
nor U11022 (N_11022,N_10616,N_10877);
or U11023 (N_11023,N_10996,N_10772);
nand U11024 (N_11024,N_10716,N_10862);
or U11025 (N_11025,N_10921,N_10823);
nand U11026 (N_11026,N_10951,N_10619);
or U11027 (N_11027,N_10646,N_10781);
nand U11028 (N_11028,N_10628,N_10548);
or U11029 (N_11029,N_10658,N_10596);
xnor U11030 (N_11030,N_10827,N_10622);
or U11031 (N_11031,N_10846,N_10909);
and U11032 (N_11032,N_10644,N_10681);
and U11033 (N_11033,N_10833,N_10972);
xnor U11034 (N_11034,N_10999,N_10983);
nand U11035 (N_11035,N_10543,N_10552);
and U11036 (N_11036,N_10894,N_10945);
nor U11037 (N_11037,N_10874,N_10568);
or U11038 (N_11038,N_10949,N_10562);
nor U11039 (N_11039,N_10586,N_10521);
nor U11040 (N_11040,N_10795,N_10517);
nand U11041 (N_11041,N_10919,N_10660);
and U11042 (N_11042,N_10906,N_10767);
nand U11043 (N_11043,N_10858,N_10747);
xnor U11044 (N_11044,N_10868,N_10762);
and U11045 (N_11045,N_10933,N_10640);
nor U11046 (N_11046,N_10849,N_10903);
or U11047 (N_11047,N_10806,N_10717);
and U11048 (N_11048,N_10898,N_10695);
nor U11049 (N_11049,N_10981,N_10722);
nor U11050 (N_11050,N_10691,N_10626);
nor U11051 (N_11051,N_10575,N_10977);
nand U11052 (N_11052,N_10798,N_10939);
nor U11053 (N_11053,N_10536,N_10549);
xor U11054 (N_11054,N_10936,N_10597);
xor U11055 (N_11055,N_10918,N_10963);
nand U11056 (N_11056,N_10965,N_10591);
xnor U11057 (N_11057,N_10859,N_10624);
and U11058 (N_11058,N_10531,N_10671);
nor U11059 (N_11059,N_10927,N_10875);
nand U11060 (N_11060,N_10571,N_10669);
nor U11061 (N_11061,N_10841,N_10789);
xor U11062 (N_11062,N_10887,N_10572);
and U11063 (N_11063,N_10873,N_10593);
and U11064 (N_11064,N_10885,N_10773);
or U11065 (N_11065,N_10602,N_10700);
and U11066 (N_11066,N_10689,N_10917);
nand U11067 (N_11067,N_10588,N_10730);
xnor U11068 (N_11068,N_10960,N_10967);
or U11069 (N_11069,N_10749,N_10824);
and U11070 (N_11070,N_10755,N_10687);
nor U11071 (N_11071,N_10692,N_10649);
nand U11072 (N_11072,N_10514,N_10895);
and U11073 (N_11073,N_10561,N_10956);
and U11074 (N_11074,N_10802,N_10932);
and U11075 (N_11075,N_10664,N_10629);
nand U11076 (N_11076,N_10534,N_10707);
or U11077 (N_11077,N_10690,N_10611);
xor U11078 (N_11078,N_10520,N_10954);
xnor U11079 (N_11079,N_10708,N_10889);
or U11080 (N_11080,N_10535,N_10667);
xor U11081 (N_11081,N_10975,N_10878);
and U11082 (N_11082,N_10844,N_10938);
nand U11083 (N_11083,N_10857,N_10713);
xnor U11084 (N_11084,N_10529,N_10679);
and U11085 (N_11085,N_10530,N_10594);
xor U11086 (N_11086,N_10533,N_10653);
xnor U11087 (N_11087,N_10746,N_10714);
or U11088 (N_11088,N_10578,N_10888);
nand U11089 (N_11089,N_10947,N_10860);
xnor U11090 (N_11090,N_10641,N_10847);
or U11091 (N_11091,N_10739,N_10754);
or U11092 (N_11092,N_10843,N_10786);
xor U11093 (N_11093,N_10705,N_10513);
xnor U11094 (N_11094,N_10735,N_10782);
and U11095 (N_11095,N_10867,N_10992);
xnor U11096 (N_11096,N_10923,N_10913);
and U11097 (N_11097,N_10720,N_10545);
nand U11098 (N_11098,N_10757,N_10674);
nor U11099 (N_11099,N_10850,N_10505);
or U11100 (N_11100,N_10801,N_10651);
nor U11101 (N_11101,N_10542,N_10673);
or U11102 (N_11102,N_10733,N_10775);
and U11103 (N_11103,N_10685,N_10501);
and U11104 (N_11104,N_10592,N_10701);
xnor U11105 (N_11105,N_10518,N_10962);
xor U11106 (N_11106,N_10740,N_10627);
xnor U11107 (N_11107,N_10605,N_10851);
or U11108 (N_11108,N_10812,N_10853);
or U11109 (N_11109,N_10794,N_10998);
nor U11110 (N_11110,N_10916,N_10924);
nor U11111 (N_11111,N_10828,N_10905);
or U11112 (N_11112,N_10564,N_10751);
or U11113 (N_11113,N_10512,N_10752);
nor U11114 (N_11114,N_10978,N_10737);
nor U11115 (N_11115,N_10866,N_10769);
nand U11116 (N_11116,N_10809,N_10944);
nor U11117 (N_11117,N_10756,N_10583);
nor U11118 (N_11118,N_10870,N_10834);
xor U11119 (N_11119,N_10968,N_10630);
nor U11120 (N_11120,N_10930,N_10576);
nand U11121 (N_11121,N_10524,N_10694);
nand U11122 (N_11122,N_10584,N_10937);
and U11123 (N_11123,N_10760,N_10987);
nor U11124 (N_11124,N_10980,N_10509);
nand U11125 (N_11125,N_10790,N_10715);
and U11126 (N_11126,N_10709,N_10519);
nor U11127 (N_11127,N_10693,N_10523);
or U11128 (N_11128,N_10800,N_10610);
nor U11129 (N_11129,N_10865,N_10632);
nor U11130 (N_11130,N_10558,N_10814);
nor U11131 (N_11131,N_10527,N_10808);
nand U11132 (N_11132,N_10907,N_10743);
nor U11133 (N_11133,N_10768,N_10662);
nor U11134 (N_11134,N_10604,N_10970);
xnor U11135 (N_11135,N_10642,N_10884);
and U11136 (N_11136,N_10810,N_10961);
xnor U11137 (N_11137,N_10506,N_10959);
and U11138 (N_11138,N_10979,N_10826);
xnor U11139 (N_11139,N_10861,N_10606);
nand U11140 (N_11140,N_10753,N_10910);
xnor U11141 (N_11141,N_10837,N_10680);
and U11142 (N_11142,N_10647,N_10522);
nand U11143 (N_11143,N_10797,N_10706);
or U11144 (N_11144,N_10946,N_10718);
and U11145 (N_11145,N_10645,N_10832);
xnor U11146 (N_11146,N_10882,N_10886);
xor U11147 (N_11147,N_10848,N_10796);
or U11148 (N_11148,N_10904,N_10654);
nor U11149 (N_11149,N_10745,N_10852);
nor U11150 (N_11150,N_10553,N_10516);
xnor U11151 (N_11151,N_10982,N_10625);
and U11152 (N_11152,N_10929,N_10891);
nand U11153 (N_11153,N_10551,N_10639);
and U11154 (N_11154,N_10510,N_10985);
or U11155 (N_11155,N_10764,N_10902);
nand U11156 (N_11156,N_10803,N_10758);
nand U11157 (N_11157,N_10703,N_10504);
nor U11158 (N_11158,N_10598,N_10668);
and U11159 (N_11159,N_10765,N_10600);
nor U11160 (N_11160,N_10620,N_10615);
and U11161 (N_11161,N_10854,N_10900);
nand U11162 (N_11162,N_10670,N_10581);
and U11163 (N_11163,N_10704,N_10770);
xor U11164 (N_11164,N_10881,N_10955);
nor U11165 (N_11165,N_10500,N_10822);
or U11166 (N_11166,N_10508,N_10896);
nor U11167 (N_11167,N_10819,N_10744);
nor U11168 (N_11168,N_10799,N_10731);
or U11169 (N_11169,N_10911,N_10935);
or U11170 (N_11170,N_10883,N_10554);
or U11171 (N_11171,N_10840,N_10567);
xnor U11172 (N_11172,N_10776,N_10541);
xnor U11173 (N_11173,N_10991,N_10652);
nor U11174 (N_11174,N_10817,N_10728);
or U11175 (N_11175,N_10880,N_10791);
and U11176 (N_11176,N_10940,N_10719);
and U11177 (N_11177,N_10777,N_10988);
or U11178 (N_11178,N_10599,N_10783);
xor U11179 (N_11179,N_10876,N_10792);
and U11180 (N_11180,N_10557,N_10948);
nor U11181 (N_11181,N_10579,N_10787);
xnor U11182 (N_11182,N_10574,N_10560);
nand U11183 (N_11183,N_10778,N_10995);
nor U11184 (N_11184,N_10964,N_10973);
and U11185 (N_11185,N_10813,N_10732);
and U11186 (N_11186,N_10723,N_10784);
and U11187 (N_11187,N_10811,N_10788);
and U11188 (N_11188,N_10612,N_10925);
xor U11189 (N_11189,N_10637,N_10537);
and U11190 (N_11190,N_10971,N_10943);
xor U11191 (N_11191,N_10766,N_10556);
nor U11192 (N_11192,N_10656,N_10761);
nor U11193 (N_11193,N_10678,N_10565);
xor U11194 (N_11194,N_10748,N_10771);
nor U11195 (N_11195,N_10818,N_10912);
xnor U11196 (N_11196,N_10577,N_10897);
nor U11197 (N_11197,N_10901,N_10711);
nand U11198 (N_11198,N_10928,N_10566);
nand U11199 (N_11199,N_10807,N_10734);
nand U11200 (N_11200,N_10763,N_10525);
xor U11201 (N_11201,N_10950,N_10688);
xnor U11202 (N_11202,N_10635,N_10942);
xnor U11203 (N_11203,N_10750,N_10958);
or U11204 (N_11204,N_10633,N_10511);
and U11205 (N_11205,N_10829,N_10830);
xnor U11206 (N_11206,N_10759,N_10831);
xnor U11207 (N_11207,N_10621,N_10585);
and U11208 (N_11208,N_10532,N_10957);
nand U11209 (N_11209,N_10997,N_10893);
and U11210 (N_11210,N_10974,N_10603);
nor U11211 (N_11211,N_10682,N_10779);
or U11212 (N_11212,N_10926,N_10871);
and U11213 (N_11213,N_10634,N_10587);
or U11214 (N_11214,N_10540,N_10569);
xnor U11215 (N_11215,N_10617,N_10920);
and U11216 (N_11216,N_10546,N_10785);
and U11217 (N_11217,N_10845,N_10697);
nand U11218 (N_11218,N_10590,N_10989);
nor U11219 (N_11219,N_10815,N_10507);
xnor U11220 (N_11220,N_10838,N_10683);
nand U11221 (N_11221,N_10699,N_10915);
and U11222 (N_11222,N_10736,N_10698);
nand U11223 (N_11223,N_10934,N_10677);
nor U11224 (N_11224,N_10890,N_10804);
xnor U11225 (N_11225,N_10741,N_10676);
xor U11226 (N_11226,N_10636,N_10821);
nor U11227 (N_11227,N_10702,N_10608);
nor U11228 (N_11228,N_10657,N_10503);
or U11229 (N_11229,N_10805,N_10550);
xnor U11230 (N_11230,N_10899,N_10563);
nand U11231 (N_11231,N_10526,N_10659);
nand U11232 (N_11232,N_10842,N_10672);
and U11233 (N_11233,N_10914,N_10725);
nor U11234 (N_11234,N_10993,N_10863);
or U11235 (N_11235,N_10650,N_10721);
nand U11236 (N_11236,N_10879,N_10631);
and U11237 (N_11237,N_10727,N_10825);
nand U11238 (N_11238,N_10696,N_10675);
nor U11239 (N_11239,N_10547,N_10941);
nor U11240 (N_11240,N_10614,N_10835);
or U11241 (N_11241,N_10544,N_10966);
or U11242 (N_11242,N_10836,N_10686);
xnor U11243 (N_11243,N_10601,N_10931);
or U11244 (N_11244,N_10684,N_10538);
xor U11245 (N_11245,N_10607,N_10726);
and U11246 (N_11246,N_10539,N_10666);
nand U11247 (N_11247,N_10892,N_10570);
or U11248 (N_11248,N_10976,N_10738);
nor U11249 (N_11249,N_10774,N_10793);
nand U11250 (N_11250,N_10643,N_10567);
xnor U11251 (N_11251,N_10569,N_10980);
nor U11252 (N_11252,N_10739,N_10883);
or U11253 (N_11253,N_10912,N_10503);
or U11254 (N_11254,N_10765,N_10927);
or U11255 (N_11255,N_10580,N_10685);
nor U11256 (N_11256,N_10566,N_10613);
xnor U11257 (N_11257,N_10966,N_10547);
nor U11258 (N_11258,N_10592,N_10904);
nand U11259 (N_11259,N_10840,N_10559);
nand U11260 (N_11260,N_10853,N_10757);
nand U11261 (N_11261,N_10695,N_10854);
xor U11262 (N_11262,N_10629,N_10939);
or U11263 (N_11263,N_10674,N_10673);
xor U11264 (N_11264,N_10507,N_10841);
nand U11265 (N_11265,N_10675,N_10764);
nor U11266 (N_11266,N_10564,N_10523);
and U11267 (N_11267,N_10767,N_10729);
or U11268 (N_11268,N_10989,N_10837);
nand U11269 (N_11269,N_10736,N_10746);
xor U11270 (N_11270,N_10944,N_10593);
xnor U11271 (N_11271,N_10719,N_10679);
or U11272 (N_11272,N_10618,N_10603);
nor U11273 (N_11273,N_10614,N_10640);
nor U11274 (N_11274,N_10799,N_10951);
xnor U11275 (N_11275,N_10550,N_10694);
nand U11276 (N_11276,N_10912,N_10569);
or U11277 (N_11277,N_10614,N_10667);
and U11278 (N_11278,N_10908,N_10948);
and U11279 (N_11279,N_10598,N_10739);
or U11280 (N_11280,N_10801,N_10645);
nand U11281 (N_11281,N_10790,N_10968);
and U11282 (N_11282,N_10591,N_10793);
nand U11283 (N_11283,N_10750,N_10569);
xnor U11284 (N_11284,N_10520,N_10554);
xor U11285 (N_11285,N_10742,N_10621);
nand U11286 (N_11286,N_10911,N_10541);
xnor U11287 (N_11287,N_10508,N_10768);
nand U11288 (N_11288,N_10511,N_10702);
nand U11289 (N_11289,N_10898,N_10574);
nand U11290 (N_11290,N_10579,N_10841);
or U11291 (N_11291,N_10824,N_10952);
xor U11292 (N_11292,N_10731,N_10779);
and U11293 (N_11293,N_10688,N_10610);
and U11294 (N_11294,N_10931,N_10720);
xor U11295 (N_11295,N_10918,N_10740);
nor U11296 (N_11296,N_10710,N_10766);
nor U11297 (N_11297,N_10529,N_10551);
and U11298 (N_11298,N_10678,N_10836);
xor U11299 (N_11299,N_10579,N_10572);
nor U11300 (N_11300,N_10707,N_10810);
xor U11301 (N_11301,N_10616,N_10664);
nor U11302 (N_11302,N_10720,N_10640);
xnor U11303 (N_11303,N_10806,N_10501);
and U11304 (N_11304,N_10575,N_10522);
or U11305 (N_11305,N_10522,N_10979);
xor U11306 (N_11306,N_10836,N_10910);
nor U11307 (N_11307,N_10980,N_10637);
xnor U11308 (N_11308,N_10524,N_10641);
nor U11309 (N_11309,N_10866,N_10549);
xnor U11310 (N_11310,N_10708,N_10831);
or U11311 (N_11311,N_10958,N_10565);
nand U11312 (N_11312,N_10678,N_10893);
nand U11313 (N_11313,N_10669,N_10769);
nor U11314 (N_11314,N_10838,N_10567);
or U11315 (N_11315,N_10515,N_10542);
and U11316 (N_11316,N_10882,N_10931);
xor U11317 (N_11317,N_10795,N_10685);
and U11318 (N_11318,N_10651,N_10572);
nand U11319 (N_11319,N_10587,N_10816);
nand U11320 (N_11320,N_10684,N_10679);
xor U11321 (N_11321,N_10791,N_10702);
and U11322 (N_11322,N_10887,N_10786);
nand U11323 (N_11323,N_10803,N_10914);
nor U11324 (N_11324,N_10934,N_10884);
and U11325 (N_11325,N_10555,N_10664);
nor U11326 (N_11326,N_10657,N_10829);
xnor U11327 (N_11327,N_10901,N_10974);
nor U11328 (N_11328,N_10775,N_10971);
xor U11329 (N_11329,N_10669,N_10817);
and U11330 (N_11330,N_10689,N_10616);
xor U11331 (N_11331,N_10648,N_10518);
xnor U11332 (N_11332,N_10781,N_10760);
or U11333 (N_11333,N_10671,N_10760);
xor U11334 (N_11334,N_10730,N_10565);
nor U11335 (N_11335,N_10796,N_10716);
nor U11336 (N_11336,N_10984,N_10548);
or U11337 (N_11337,N_10508,N_10782);
and U11338 (N_11338,N_10993,N_10641);
nor U11339 (N_11339,N_10668,N_10999);
and U11340 (N_11340,N_10768,N_10769);
nand U11341 (N_11341,N_10544,N_10954);
or U11342 (N_11342,N_10903,N_10887);
or U11343 (N_11343,N_10850,N_10507);
or U11344 (N_11344,N_10736,N_10683);
xor U11345 (N_11345,N_10603,N_10726);
nand U11346 (N_11346,N_10844,N_10617);
nor U11347 (N_11347,N_10780,N_10911);
or U11348 (N_11348,N_10639,N_10641);
nand U11349 (N_11349,N_10540,N_10684);
or U11350 (N_11350,N_10808,N_10869);
and U11351 (N_11351,N_10755,N_10564);
nor U11352 (N_11352,N_10918,N_10519);
xnor U11353 (N_11353,N_10591,N_10898);
or U11354 (N_11354,N_10786,N_10937);
and U11355 (N_11355,N_10676,N_10776);
xnor U11356 (N_11356,N_10651,N_10721);
xnor U11357 (N_11357,N_10888,N_10630);
xor U11358 (N_11358,N_10923,N_10658);
and U11359 (N_11359,N_10647,N_10857);
nor U11360 (N_11360,N_10711,N_10801);
nor U11361 (N_11361,N_10792,N_10571);
nand U11362 (N_11362,N_10684,N_10552);
and U11363 (N_11363,N_10735,N_10727);
and U11364 (N_11364,N_10547,N_10853);
and U11365 (N_11365,N_10560,N_10975);
and U11366 (N_11366,N_10966,N_10945);
nand U11367 (N_11367,N_10792,N_10951);
nand U11368 (N_11368,N_10561,N_10911);
nand U11369 (N_11369,N_10600,N_10907);
and U11370 (N_11370,N_10752,N_10925);
xnor U11371 (N_11371,N_10601,N_10851);
nor U11372 (N_11372,N_10959,N_10995);
nor U11373 (N_11373,N_10602,N_10787);
and U11374 (N_11374,N_10869,N_10814);
and U11375 (N_11375,N_10945,N_10616);
or U11376 (N_11376,N_10949,N_10517);
nand U11377 (N_11377,N_10918,N_10589);
nor U11378 (N_11378,N_10712,N_10775);
nor U11379 (N_11379,N_10800,N_10909);
nand U11380 (N_11380,N_10630,N_10523);
nor U11381 (N_11381,N_10661,N_10592);
and U11382 (N_11382,N_10517,N_10990);
xor U11383 (N_11383,N_10629,N_10631);
xnor U11384 (N_11384,N_10820,N_10859);
xor U11385 (N_11385,N_10665,N_10821);
nor U11386 (N_11386,N_10508,N_10515);
xor U11387 (N_11387,N_10707,N_10899);
xor U11388 (N_11388,N_10781,N_10792);
nor U11389 (N_11389,N_10508,N_10678);
or U11390 (N_11390,N_10885,N_10906);
xnor U11391 (N_11391,N_10613,N_10868);
or U11392 (N_11392,N_10783,N_10857);
nand U11393 (N_11393,N_10637,N_10571);
xnor U11394 (N_11394,N_10509,N_10633);
nor U11395 (N_11395,N_10714,N_10741);
xnor U11396 (N_11396,N_10513,N_10520);
and U11397 (N_11397,N_10636,N_10860);
nand U11398 (N_11398,N_10928,N_10983);
nand U11399 (N_11399,N_10594,N_10833);
nor U11400 (N_11400,N_10634,N_10859);
nor U11401 (N_11401,N_10820,N_10933);
or U11402 (N_11402,N_10869,N_10656);
xnor U11403 (N_11403,N_10719,N_10783);
and U11404 (N_11404,N_10523,N_10623);
and U11405 (N_11405,N_10748,N_10876);
and U11406 (N_11406,N_10550,N_10792);
nor U11407 (N_11407,N_10927,N_10968);
and U11408 (N_11408,N_10582,N_10766);
or U11409 (N_11409,N_10609,N_10736);
and U11410 (N_11410,N_10812,N_10979);
or U11411 (N_11411,N_10892,N_10988);
xor U11412 (N_11412,N_10569,N_10847);
and U11413 (N_11413,N_10910,N_10640);
nor U11414 (N_11414,N_10922,N_10567);
nand U11415 (N_11415,N_10676,N_10668);
and U11416 (N_11416,N_10986,N_10622);
nand U11417 (N_11417,N_10522,N_10618);
or U11418 (N_11418,N_10799,N_10909);
nor U11419 (N_11419,N_10575,N_10525);
nor U11420 (N_11420,N_10678,N_10648);
nor U11421 (N_11421,N_10766,N_10613);
xor U11422 (N_11422,N_10751,N_10754);
xor U11423 (N_11423,N_10835,N_10986);
nor U11424 (N_11424,N_10887,N_10796);
nand U11425 (N_11425,N_10958,N_10634);
and U11426 (N_11426,N_10865,N_10758);
xor U11427 (N_11427,N_10986,N_10970);
or U11428 (N_11428,N_10842,N_10657);
xnor U11429 (N_11429,N_10562,N_10838);
or U11430 (N_11430,N_10646,N_10638);
and U11431 (N_11431,N_10815,N_10736);
and U11432 (N_11432,N_10876,N_10910);
and U11433 (N_11433,N_10523,N_10998);
xnor U11434 (N_11434,N_10562,N_10818);
or U11435 (N_11435,N_10872,N_10515);
nand U11436 (N_11436,N_10714,N_10774);
xor U11437 (N_11437,N_10711,N_10927);
xor U11438 (N_11438,N_10905,N_10830);
xor U11439 (N_11439,N_10936,N_10893);
or U11440 (N_11440,N_10796,N_10665);
nand U11441 (N_11441,N_10585,N_10767);
nor U11442 (N_11442,N_10810,N_10978);
nand U11443 (N_11443,N_10555,N_10848);
xor U11444 (N_11444,N_10600,N_10781);
or U11445 (N_11445,N_10532,N_10992);
nand U11446 (N_11446,N_10814,N_10564);
nand U11447 (N_11447,N_10577,N_10860);
xor U11448 (N_11448,N_10593,N_10871);
nand U11449 (N_11449,N_10730,N_10547);
nand U11450 (N_11450,N_10894,N_10794);
nand U11451 (N_11451,N_10536,N_10567);
xor U11452 (N_11452,N_10815,N_10959);
xnor U11453 (N_11453,N_10504,N_10939);
nor U11454 (N_11454,N_10729,N_10664);
and U11455 (N_11455,N_10928,N_10597);
nor U11456 (N_11456,N_10972,N_10599);
xor U11457 (N_11457,N_10533,N_10785);
xnor U11458 (N_11458,N_10528,N_10905);
nor U11459 (N_11459,N_10587,N_10726);
or U11460 (N_11460,N_10965,N_10888);
and U11461 (N_11461,N_10685,N_10694);
nand U11462 (N_11462,N_10529,N_10790);
and U11463 (N_11463,N_10732,N_10581);
nor U11464 (N_11464,N_10740,N_10548);
or U11465 (N_11465,N_10684,N_10960);
nand U11466 (N_11466,N_10952,N_10629);
nor U11467 (N_11467,N_10725,N_10699);
and U11468 (N_11468,N_10678,N_10711);
nand U11469 (N_11469,N_10535,N_10800);
nand U11470 (N_11470,N_10880,N_10737);
nor U11471 (N_11471,N_10806,N_10695);
xnor U11472 (N_11472,N_10596,N_10734);
nand U11473 (N_11473,N_10858,N_10573);
or U11474 (N_11474,N_10829,N_10795);
nor U11475 (N_11475,N_10629,N_10524);
xor U11476 (N_11476,N_10594,N_10976);
xnor U11477 (N_11477,N_10898,N_10747);
and U11478 (N_11478,N_10825,N_10704);
nand U11479 (N_11479,N_10568,N_10824);
nand U11480 (N_11480,N_10884,N_10643);
or U11481 (N_11481,N_10876,N_10563);
nor U11482 (N_11482,N_10707,N_10996);
or U11483 (N_11483,N_10680,N_10683);
and U11484 (N_11484,N_10747,N_10845);
nand U11485 (N_11485,N_10861,N_10771);
or U11486 (N_11486,N_10868,N_10688);
nor U11487 (N_11487,N_10960,N_10959);
or U11488 (N_11488,N_10508,N_10524);
xor U11489 (N_11489,N_10931,N_10838);
and U11490 (N_11490,N_10940,N_10926);
or U11491 (N_11491,N_10988,N_10797);
nor U11492 (N_11492,N_10869,N_10966);
nand U11493 (N_11493,N_10839,N_10891);
nand U11494 (N_11494,N_10913,N_10725);
and U11495 (N_11495,N_10814,N_10997);
or U11496 (N_11496,N_10877,N_10683);
nand U11497 (N_11497,N_10751,N_10774);
nor U11498 (N_11498,N_10616,N_10623);
nor U11499 (N_11499,N_10582,N_10926);
nand U11500 (N_11500,N_11239,N_11131);
or U11501 (N_11501,N_11110,N_11419);
and U11502 (N_11502,N_11322,N_11281);
and U11503 (N_11503,N_11207,N_11233);
nand U11504 (N_11504,N_11438,N_11160);
and U11505 (N_11505,N_11264,N_11128);
and U11506 (N_11506,N_11367,N_11388);
xor U11507 (N_11507,N_11404,N_11448);
nor U11508 (N_11508,N_11187,N_11302);
and U11509 (N_11509,N_11284,N_11338);
and U11510 (N_11510,N_11313,N_11396);
and U11511 (N_11511,N_11356,N_11097);
nor U11512 (N_11512,N_11330,N_11359);
and U11513 (N_11513,N_11236,N_11149);
or U11514 (N_11514,N_11267,N_11420);
nand U11515 (N_11515,N_11455,N_11259);
xnor U11516 (N_11516,N_11253,N_11415);
nor U11517 (N_11517,N_11288,N_11465);
nand U11518 (N_11518,N_11057,N_11375);
nand U11519 (N_11519,N_11241,N_11273);
xor U11520 (N_11520,N_11445,N_11218);
nor U11521 (N_11521,N_11073,N_11077);
or U11522 (N_11522,N_11026,N_11215);
xor U11523 (N_11523,N_11368,N_11378);
and U11524 (N_11524,N_11055,N_11462);
and U11525 (N_11525,N_11498,N_11031);
or U11526 (N_11526,N_11488,N_11047);
or U11527 (N_11527,N_11230,N_11252);
nor U11528 (N_11528,N_11016,N_11470);
xor U11529 (N_11529,N_11039,N_11352);
nand U11530 (N_11530,N_11483,N_11166);
or U11531 (N_11531,N_11350,N_11494);
and U11532 (N_11532,N_11070,N_11435);
or U11533 (N_11533,N_11290,N_11472);
nor U11534 (N_11534,N_11229,N_11030);
and U11535 (N_11535,N_11254,N_11314);
or U11536 (N_11536,N_11004,N_11021);
xor U11537 (N_11537,N_11122,N_11422);
nand U11538 (N_11538,N_11399,N_11117);
xnor U11539 (N_11539,N_11118,N_11286);
xnor U11540 (N_11540,N_11373,N_11268);
nand U11541 (N_11541,N_11289,N_11456);
and U11542 (N_11542,N_11072,N_11403);
and U11543 (N_11543,N_11180,N_11499);
xnor U11544 (N_11544,N_11402,N_11217);
or U11545 (N_11545,N_11023,N_11351);
nor U11546 (N_11546,N_11140,N_11418);
nor U11547 (N_11547,N_11221,N_11119);
nor U11548 (N_11548,N_11009,N_11410);
xor U11549 (N_11549,N_11431,N_11088);
nand U11550 (N_11550,N_11293,N_11349);
nand U11551 (N_11551,N_11015,N_11183);
nand U11552 (N_11552,N_11371,N_11346);
nor U11553 (N_11553,N_11365,N_11269);
or U11554 (N_11554,N_11204,N_11277);
or U11555 (N_11555,N_11051,N_11075);
nand U11556 (N_11556,N_11082,N_11222);
or U11557 (N_11557,N_11407,N_11176);
nor U11558 (N_11558,N_11411,N_11335);
nor U11559 (N_11559,N_11428,N_11491);
or U11560 (N_11560,N_11405,N_11423);
and U11561 (N_11561,N_11340,N_11094);
nand U11562 (N_11562,N_11372,N_11048);
nor U11563 (N_11563,N_11478,N_11050);
or U11564 (N_11564,N_11102,N_11341);
xnor U11565 (N_11565,N_11374,N_11476);
and U11566 (N_11566,N_11090,N_11200);
nor U11567 (N_11567,N_11487,N_11164);
nor U11568 (N_11568,N_11464,N_11091);
nor U11569 (N_11569,N_11364,N_11300);
and U11570 (N_11570,N_11135,N_11171);
xor U11571 (N_11571,N_11362,N_11467);
or U11572 (N_11572,N_11353,N_11227);
nand U11573 (N_11573,N_11209,N_11142);
and U11574 (N_11574,N_11439,N_11401);
xnor U11575 (N_11575,N_11201,N_11390);
nand U11576 (N_11576,N_11005,N_11260);
and U11577 (N_11577,N_11473,N_11296);
nand U11578 (N_11578,N_11248,N_11025);
or U11579 (N_11579,N_11336,N_11497);
and U11580 (N_11580,N_11033,N_11147);
xnor U11581 (N_11581,N_11111,N_11173);
nor U11582 (N_11582,N_11242,N_11427);
nor U11583 (N_11583,N_11042,N_11451);
or U11584 (N_11584,N_11079,N_11076);
and U11585 (N_11585,N_11249,N_11141);
xor U11586 (N_11586,N_11484,N_11060);
or U11587 (N_11587,N_11255,N_11417);
or U11588 (N_11588,N_11468,N_11295);
nand U11589 (N_11589,N_11316,N_11308);
and U11590 (N_11590,N_11449,N_11436);
or U11591 (N_11591,N_11337,N_11447);
nand U11592 (N_11592,N_11089,N_11324);
nand U11593 (N_11593,N_11460,N_11188);
nand U11594 (N_11594,N_11257,N_11041);
xnor U11595 (N_11595,N_11101,N_11019);
xnor U11596 (N_11596,N_11315,N_11413);
nor U11597 (N_11597,N_11245,N_11064);
or U11598 (N_11598,N_11272,N_11162);
nand U11599 (N_11599,N_11360,N_11262);
nand U11600 (N_11600,N_11294,N_11344);
and U11601 (N_11601,N_11120,N_11062);
or U11602 (N_11602,N_11022,N_11095);
nand U11603 (N_11603,N_11471,N_11145);
and U11604 (N_11604,N_11112,N_11458);
nand U11605 (N_11605,N_11168,N_11186);
and U11606 (N_11606,N_11163,N_11225);
or U11607 (N_11607,N_11292,N_11012);
or U11608 (N_11608,N_11475,N_11244);
or U11609 (N_11609,N_11114,N_11212);
and U11610 (N_11610,N_11202,N_11325);
nor U11611 (N_11611,N_11053,N_11197);
nor U11612 (N_11612,N_11307,N_11136);
or U11613 (N_11613,N_11138,N_11379);
or U11614 (N_11614,N_11087,N_11394);
or U11615 (N_11615,N_11006,N_11078);
nand U11616 (N_11616,N_11063,N_11074);
nand U11617 (N_11617,N_11066,N_11126);
or U11618 (N_11618,N_11010,N_11243);
nand U11619 (N_11619,N_11309,N_11266);
nand U11620 (N_11620,N_11305,N_11208);
or U11621 (N_11621,N_11256,N_11446);
xor U11622 (N_11622,N_11450,N_11152);
nand U11623 (N_11623,N_11065,N_11412);
or U11624 (N_11624,N_11098,N_11382);
xnor U11625 (N_11625,N_11107,N_11151);
xor U11626 (N_11626,N_11220,N_11115);
xor U11627 (N_11627,N_11291,N_11270);
nand U11628 (N_11628,N_11032,N_11157);
nor U11629 (N_11629,N_11106,N_11170);
and U11630 (N_11630,N_11370,N_11306);
and U11631 (N_11631,N_11093,N_11490);
nor U11632 (N_11632,N_11381,N_11061);
nand U11633 (N_11633,N_11392,N_11461);
xnor U11634 (N_11634,N_11194,N_11361);
or U11635 (N_11635,N_11219,N_11214);
or U11636 (N_11636,N_11132,N_11304);
nor U11637 (N_11637,N_11329,N_11024);
xor U11638 (N_11638,N_11043,N_11232);
xnor U11639 (N_11639,N_11092,N_11384);
nor U11640 (N_11640,N_11210,N_11040);
and U11641 (N_11641,N_11251,N_11081);
or U11642 (N_11642,N_11285,N_11333);
nor U11643 (N_11643,N_11196,N_11358);
xor U11644 (N_11644,N_11020,N_11137);
xnor U11645 (N_11645,N_11059,N_11319);
nand U11646 (N_11646,N_11044,N_11086);
nor U11647 (N_11647,N_11071,N_11426);
xor U11648 (N_11648,N_11363,N_11165);
nor U11649 (N_11649,N_11246,N_11454);
xor U11650 (N_11650,N_11134,N_11148);
nor U11651 (N_11651,N_11393,N_11357);
or U11652 (N_11652,N_11211,N_11496);
xnor U11653 (N_11653,N_11100,N_11181);
and U11654 (N_11654,N_11398,N_11424);
nor U11655 (N_11655,N_11027,N_11345);
and U11656 (N_11656,N_11018,N_11013);
and U11657 (N_11657,N_11317,N_11011);
nand U11658 (N_11658,N_11105,N_11058);
or U11659 (N_11659,N_11299,N_11195);
nand U11660 (N_11660,N_11193,N_11429);
xnor U11661 (N_11661,N_11334,N_11441);
nand U11662 (N_11662,N_11355,N_11125);
or U11663 (N_11663,N_11282,N_11113);
nand U11664 (N_11664,N_11109,N_11469);
and U11665 (N_11665,N_11366,N_11437);
nor U11666 (N_11666,N_11421,N_11150);
and U11667 (N_11667,N_11096,N_11103);
xor U11668 (N_11668,N_11213,N_11321);
xnor U11669 (N_11669,N_11143,N_11271);
xor U11670 (N_11670,N_11347,N_11444);
nand U11671 (N_11671,N_11395,N_11226);
nor U11672 (N_11672,N_11133,N_11342);
and U11673 (N_11673,N_11014,N_11432);
and U11674 (N_11674,N_11199,N_11108);
nand U11675 (N_11675,N_11430,N_11198);
and U11676 (N_11676,N_11167,N_11332);
and U11677 (N_11677,N_11283,N_11493);
or U11678 (N_11678,N_11159,N_11301);
or U11679 (N_11679,N_11425,N_11084);
nor U11680 (N_11680,N_11386,N_11276);
nand U11681 (N_11681,N_11279,N_11320);
and U11682 (N_11682,N_11069,N_11278);
nand U11683 (N_11683,N_11191,N_11129);
nand U11684 (N_11684,N_11234,N_11068);
nand U11685 (N_11685,N_11104,N_11017);
nor U11686 (N_11686,N_11224,N_11377);
xnor U11687 (N_11687,N_11443,N_11231);
or U11688 (N_11688,N_11085,N_11029);
or U11689 (N_11689,N_11459,N_11369);
or U11690 (N_11690,N_11139,N_11007);
or U11691 (N_11691,N_11144,N_11121);
xor U11692 (N_11692,N_11127,N_11035);
and U11693 (N_11693,N_11156,N_11002);
xor U11694 (N_11694,N_11327,N_11153);
or U11695 (N_11695,N_11312,N_11380);
xnor U11696 (N_11696,N_11206,N_11116);
nor U11697 (N_11697,N_11326,N_11343);
nand U11698 (N_11698,N_11049,N_11480);
or U11699 (N_11699,N_11339,N_11036);
nor U11700 (N_11700,N_11034,N_11434);
nor U11701 (N_11701,N_11038,N_11080);
nand U11702 (N_11702,N_11328,N_11177);
nand U11703 (N_11703,N_11182,N_11400);
xor U11704 (N_11704,N_11099,N_11190);
nor U11705 (N_11705,N_11385,N_11169);
xor U11706 (N_11706,N_11261,N_11263);
and U11707 (N_11707,N_11247,N_11311);
xor U11708 (N_11708,N_11178,N_11205);
and U11709 (N_11709,N_11083,N_11397);
nor U11710 (N_11710,N_11442,N_11323);
nand U11711 (N_11711,N_11482,N_11406);
nor U11712 (N_11712,N_11489,N_11154);
and U11713 (N_11713,N_11237,N_11495);
nand U11714 (N_11714,N_11216,N_11008);
xnor U11715 (N_11715,N_11389,N_11240);
nor U11716 (N_11716,N_11067,N_11433);
and U11717 (N_11717,N_11172,N_11185);
and U11718 (N_11718,N_11000,N_11223);
xnor U11719 (N_11719,N_11001,N_11045);
or U11720 (N_11720,N_11056,N_11477);
nor U11721 (N_11721,N_11161,N_11481);
or U11722 (N_11722,N_11228,N_11189);
or U11723 (N_11723,N_11123,N_11440);
nor U11724 (N_11724,N_11146,N_11287);
or U11725 (N_11725,N_11130,N_11463);
xnor U11726 (N_11726,N_11158,N_11457);
nand U11727 (N_11727,N_11348,N_11124);
or U11728 (N_11728,N_11376,N_11175);
nand U11729 (N_11729,N_11354,N_11318);
and U11730 (N_11730,N_11387,N_11258);
nand U11731 (N_11731,N_11192,N_11474);
or U11732 (N_11732,N_11238,N_11408);
nand U11733 (N_11733,N_11303,N_11275);
xnor U11734 (N_11734,N_11310,N_11298);
and U11735 (N_11735,N_11280,N_11184);
nor U11736 (N_11736,N_11391,N_11486);
nor U11737 (N_11737,N_11235,N_11452);
nor U11738 (N_11738,N_11052,N_11155);
xor U11739 (N_11739,N_11174,N_11453);
nand U11740 (N_11740,N_11331,N_11492);
nand U11741 (N_11741,N_11485,N_11037);
nor U11742 (N_11742,N_11250,N_11179);
or U11743 (N_11743,N_11274,N_11265);
or U11744 (N_11744,N_11479,N_11466);
nand U11745 (N_11745,N_11046,N_11297);
xnor U11746 (N_11746,N_11003,N_11409);
or U11747 (N_11747,N_11203,N_11416);
and U11748 (N_11748,N_11028,N_11054);
and U11749 (N_11749,N_11414,N_11383);
and U11750 (N_11750,N_11106,N_11206);
xnor U11751 (N_11751,N_11057,N_11482);
nor U11752 (N_11752,N_11090,N_11452);
or U11753 (N_11753,N_11308,N_11291);
nand U11754 (N_11754,N_11482,N_11225);
nand U11755 (N_11755,N_11113,N_11268);
nor U11756 (N_11756,N_11264,N_11075);
nand U11757 (N_11757,N_11282,N_11008);
xor U11758 (N_11758,N_11319,N_11180);
nand U11759 (N_11759,N_11178,N_11094);
and U11760 (N_11760,N_11047,N_11414);
nor U11761 (N_11761,N_11133,N_11191);
and U11762 (N_11762,N_11224,N_11087);
or U11763 (N_11763,N_11098,N_11490);
xnor U11764 (N_11764,N_11365,N_11377);
and U11765 (N_11765,N_11401,N_11029);
nand U11766 (N_11766,N_11083,N_11429);
or U11767 (N_11767,N_11495,N_11222);
or U11768 (N_11768,N_11331,N_11094);
and U11769 (N_11769,N_11093,N_11461);
xnor U11770 (N_11770,N_11015,N_11405);
xor U11771 (N_11771,N_11093,N_11402);
or U11772 (N_11772,N_11256,N_11442);
and U11773 (N_11773,N_11015,N_11326);
nand U11774 (N_11774,N_11356,N_11025);
or U11775 (N_11775,N_11274,N_11176);
or U11776 (N_11776,N_11246,N_11245);
xnor U11777 (N_11777,N_11489,N_11063);
and U11778 (N_11778,N_11359,N_11344);
nor U11779 (N_11779,N_11260,N_11240);
nand U11780 (N_11780,N_11404,N_11380);
nor U11781 (N_11781,N_11461,N_11390);
nand U11782 (N_11782,N_11088,N_11021);
and U11783 (N_11783,N_11416,N_11470);
nor U11784 (N_11784,N_11001,N_11434);
or U11785 (N_11785,N_11041,N_11303);
and U11786 (N_11786,N_11318,N_11370);
nand U11787 (N_11787,N_11379,N_11460);
and U11788 (N_11788,N_11200,N_11054);
nand U11789 (N_11789,N_11048,N_11066);
nand U11790 (N_11790,N_11350,N_11139);
xnor U11791 (N_11791,N_11043,N_11442);
nand U11792 (N_11792,N_11098,N_11493);
or U11793 (N_11793,N_11445,N_11496);
xor U11794 (N_11794,N_11330,N_11203);
nand U11795 (N_11795,N_11336,N_11476);
or U11796 (N_11796,N_11444,N_11178);
and U11797 (N_11797,N_11105,N_11446);
xor U11798 (N_11798,N_11307,N_11263);
nand U11799 (N_11799,N_11325,N_11208);
nand U11800 (N_11800,N_11073,N_11118);
nor U11801 (N_11801,N_11214,N_11471);
or U11802 (N_11802,N_11183,N_11495);
nor U11803 (N_11803,N_11192,N_11242);
nor U11804 (N_11804,N_11428,N_11341);
nand U11805 (N_11805,N_11109,N_11348);
nand U11806 (N_11806,N_11166,N_11396);
nor U11807 (N_11807,N_11411,N_11292);
nand U11808 (N_11808,N_11112,N_11473);
and U11809 (N_11809,N_11170,N_11318);
xor U11810 (N_11810,N_11036,N_11302);
and U11811 (N_11811,N_11284,N_11153);
xnor U11812 (N_11812,N_11240,N_11252);
and U11813 (N_11813,N_11122,N_11431);
and U11814 (N_11814,N_11071,N_11132);
or U11815 (N_11815,N_11014,N_11229);
nand U11816 (N_11816,N_11481,N_11167);
nor U11817 (N_11817,N_11128,N_11262);
nor U11818 (N_11818,N_11432,N_11412);
and U11819 (N_11819,N_11035,N_11450);
xnor U11820 (N_11820,N_11410,N_11461);
xor U11821 (N_11821,N_11279,N_11261);
nand U11822 (N_11822,N_11304,N_11032);
xor U11823 (N_11823,N_11130,N_11063);
xor U11824 (N_11824,N_11462,N_11076);
or U11825 (N_11825,N_11368,N_11186);
nand U11826 (N_11826,N_11317,N_11321);
or U11827 (N_11827,N_11437,N_11430);
nand U11828 (N_11828,N_11286,N_11356);
or U11829 (N_11829,N_11357,N_11349);
xor U11830 (N_11830,N_11398,N_11209);
xor U11831 (N_11831,N_11137,N_11377);
xor U11832 (N_11832,N_11172,N_11067);
nand U11833 (N_11833,N_11318,N_11388);
nor U11834 (N_11834,N_11415,N_11097);
or U11835 (N_11835,N_11026,N_11189);
xor U11836 (N_11836,N_11042,N_11435);
or U11837 (N_11837,N_11051,N_11090);
nand U11838 (N_11838,N_11214,N_11107);
nor U11839 (N_11839,N_11031,N_11185);
and U11840 (N_11840,N_11402,N_11191);
nor U11841 (N_11841,N_11310,N_11414);
or U11842 (N_11842,N_11104,N_11014);
xnor U11843 (N_11843,N_11182,N_11197);
xor U11844 (N_11844,N_11455,N_11376);
nand U11845 (N_11845,N_11438,N_11237);
or U11846 (N_11846,N_11256,N_11486);
xor U11847 (N_11847,N_11476,N_11231);
and U11848 (N_11848,N_11271,N_11027);
nand U11849 (N_11849,N_11353,N_11057);
or U11850 (N_11850,N_11192,N_11285);
nand U11851 (N_11851,N_11067,N_11233);
and U11852 (N_11852,N_11446,N_11054);
xor U11853 (N_11853,N_11069,N_11131);
or U11854 (N_11854,N_11051,N_11435);
and U11855 (N_11855,N_11281,N_11341);
and U11856 (N_11856,N_11069,N_11297);
or U11857 (N_11857,N_11422,N_11116);
or U11858 (N_11858,N_11105,N_11235);
and U11859 (N_11859,N_11467,N_11373);
xor U11860 (N_11860,N_11356,N_11004);
nand U11861 (N_11861,N_11204,N_11232);
or U11862 (N_11862,N_11170,N_11302);
nor U11863 (N_11863,N_11160,N_11127);
or U11864 (N_11864,N_11037,N_11234);
nand U11865 (N_11865,N_11212,N_11225);
or U11866 (N_11866,N_11464,N_11178);
and U11867 (N_11867,N_11240,N_11143);
or U11868 (N_11868,N_11111,N_11249);
or U11869 (N_11869,N_11035,N_11070);
nor U11870 (N_11870,N_11266,N_11297);
or U11871 (N_11871,N_11057,N_11263);
nand U11872 (N_11872,N_11114,N_11098);
xor U11873 (N_11873,N_11278,N_11492);
and U11874 (N_11874,N_11204,N_11291);
and U11875 (N_11875,N_11025,N_11084);
nor U11876 (N_11876,N_11230,N_11028);
nor U11877 (N_11877,N_11476,N_11414);
or U11878 (N_11878,N_11365,N_11357);
nor U11879 (N_11879,N_11457,N_11294);
and U11880 (N_11880,N_11040,N_11296);
xor U11881 (N_11881,N_11109,N_11114);
xnor U11882 (N_11882,N_11216,N_11288);
nor U11883 (N_11883,N_11078,N_11013);
and U11884 (N_11884,N_11216,N_11267);
or U11885 (N_11885,N_11112,N_11224);
nor U11886 (N_11886,N_11463,N_11433);
or U11887 (N_11887,N_11272,N_11115);
and U11888 (N_11888,N_11212,N_11023);
nand U11889 (N_11889,N_11005,N_11086);
xor U11890 (N_11890,N_11224,N_11211);
nand U11891 (N_11891,N_11176,N_11285);
nor U11892 (N_11892,N_11241,N_11231);
or U11893 (N_11893,N_11208,N_11412);
nand U11894 (N_11894,N_11388,N_11236);
or U11895 (N_11895,N_11479,N_11273);
nor U11896 (N_11896,N_11001,N_11069);
and U11897 (N_11897,N_11488,N_11297);
nand U11898 (N_11898,N_11055,N_11196);
nand U11899 (N_11899,N_11481,N_11362);
and U11900 (N_11900,N_11367,N_11209);
nor U11901 (N_11901,N_11180,N_11089);
nor U11902 (N_11902,N_11420,N_11183);
or U11903 (N_11903,N_11471,N_11175);
nand U11904 (N_11904,N_11420,N_11292);
nand U11905 (N_11905,N_11206,N_11494);
nand U11906 (N_11906,N_11396,N_11329);
and U11907 (N_11907,N_11215,N_11474);
or U11908 (N_11908,N_11141,N_11357);
or U11909 (N_11909,N_11410,N_11102);
nand U11910 (N_11910,N_11148,N_11255);
or U11911 (N_11911,N_11429,N_11265);
xnor U11912 (N_11912,N_11249,N_11391);
or U11913 (N_11913,N_11281,N_11121);
nand U11914 (N_11914,N_11473,N_11219);
nand U11915 (N_11915,N_11108,N_11254);
nand U11916 (N_11916,N_11147,N_11424);
nor U11917 (N_11917,N_11194,N_11190);
or U11918 (N_11918,N_11285,N_11097);
xor U11919 (N_11919,N_11023,N_11497);
or U11920 (N_11920,N_11371,N_11477);
xor U11921 (N_11921,N_11293,N_11150);
xor U11922 (N_11922,N_11198,N_11226);
nand U11923 (N_11923,N_11317,N_11413);
nor U11924 (N_11924,N_11238,N_11293);
and U11925 (N_11925,N_11297,N_11067);
and U11926 (N_11926,N_11024,N_11456);
and U11927 (N_11927,N_11318,N_11101);
xor U11928 (N_11928,N_11157,N_11398);
xnor U11929 (N_11929,N_11035,N_11391);
nor U11930 (N_11930,N_11495,N_11358);
and U11931 (N_11931,N_11109,N_11455);
and U11932 (N_11932,N_11229,N_11396);
and U11933 (N_11933,N_11172,N_11462);
and U11934 (N_11934,N_11128,N_11411);
xor U11935 (N_11935,N_11430,N_11097);
nand U11936 (N_11936,N_11025,N_11068);
and U11937 (N_11937,N_11292,N_11058);
nand U11938 (N_11938,N_11245,N_11088);
or U11939 (N_11939,N_11013,N_11016);
and U11940 (N_11940,N_11313,N_11440);
and U11941 (N_11941,N_11474,N_11092);
or U11942 (N_11942,N_11159,N_11397);
xnor U11943 (N_11943,N_11033,N_11028);
or U11944 (N_11944,N_11460,N_11061);
or U11945 (N_11945,N_11160,N_11274);
and U11946 (N_11946,N_11285,N_11246);
nand U11947 (N_11947,N_11113,N_11353);
xor U11948 (N_11948,N_11190,N_11398);
nor U11949 (N_11949,N_11123,N_11173);
xor U11950 (N_11950,N_11084,N_11273);
xor U11951 (N_11951,N_11381,N_11001);
nor U11952 (N_11952,N_11353,N_11191);
and U11953 (N_11953,N_11499,N_11040);
or U11954 (N_11954,N_11448,N_11195);
or U11955 (N_11955,N_11343,N_11345);
or U11956 (N_11956,N_11317,N_11060);
and U11957 (N_11957,N_11282,N_11335);
xnor U11958 (N_11958,N_11336,N_11260);
nor U11959 (N_11959,N_11034,N_11228);
nand U11960 (N_11960,N_11076,N_11000);
xor U11961 (N_11961,N_11192,N_11108);
and U11962 (N_11962,N_11114,N_11284);
and U11963 (N_11963,N_11448,N_11252);
and U11964 (N_11964,N_11247,N_11107);
nor U11965 (N_11965,N_11047,N_11021);
or U11966 (N_11966,N_11046,N_11178);
xor U11967 (N_11967,N_11167,N_11336);
nand U11968 (N_11968,N_11003,N_11345);
nand U11969 (N_11969,N_11438,N_11487);
and U11970 (N_11970,N_11243,N_11063);
nor U11971 (N_11971,N_11009,N_11129);
or U11972 (N_11972,N_11070,N_11053);
xor U11973 (N_11973,N_11141,N_11202);
nor U11974 (N_11974,N_11044,N_11280);
and U11975 (N_11975,N_11263,N_11182);
or U11976 (N_11976,N_11116,N_11252);
nor U11977 (N_11977,N_11066,N_11381);
and U11978 (N_11978,N_11116,N_11343);
nand U11979 (N_11979,N_11113,N_11329);
xnor U11980 (N_11980,N_11002,N_11010);
nor U11981 (N_11981,N_11269,N_11113);
or U11982 (N_11982,N_11335,N_11221);
or U11983 (N_11983,N_11135,N_11276);
or U11984 (N_11984,N_11111,N_11005);
nand U11985 (N_11985,N_11474,N_11014);
xor U11986 (N_11986,N_11276,N_11437);
xnor U11987 (N_11987,N_11159,N_11256);
nor U11988 (N_11988,N_11066,N_11036);
and U11989 (N_11989,N_11345,N_11289);
xnor U11990 (N_11990,N_11150,N_11286);
xnor U11991 (N_11991,N_11133,N_11300);
nor U11992 (N_11992,N_11385,N_11480);
xor U11993 (N_11993,N_11468,N_11177);
xnor U11994 (N_11994,N_11470,N_11127);
or U11995 (N_11995,N_11292,N_11392);
xor U11996 (N_11996,N_11173,N_11082);
or U11997 (N_11997,N_11147,N_11003);
xnor U11998 (N_11998,N_11302,N_11024);
and U11999 (N_11999,N_11118,N_11319);
and U12000 (N_12000,N_11871,N_11684);
xor U12001 (N_12001,N_11618,N_11769);
and U12002 (N_12002,N_11735,N_11675);
nor U12003 (N_12003,N_11580,N_11765);
and U12004 (N_12004,N_11702,N_11514);
and U12005 (N_12005,N_11650,N_11801);
nor U12006 (N_12006,N_11756,N_11969);
or U12007 (N_12007,N_11809,N_11577);
nand U12008 (N_12008,N_11530,N_11639);
and U12009 (N_12009,N_11778,N_11668);
xor U12010 (N_12010,N_11763,N_11951);
or U12011 (N_12011,N_11926,N_11761);
and U12012 (N_12012,N_11842,N_11641);
or U12013 (N_12013,N_11958,N_11510);
nor U12014 (N_12014,N_11712,N_11538);
nand U12015 (N_12015,N_11725,N_11894);
xor U12016 (N_12016,N_11938,N_11543);
and U12017 (N_12017,N_11664,N_11706);
and U12018 (N_12018,N_11630,N_11906);
and U12019 (N_12019,N_11805,N_11784);
nand U12020 (N_12020,N_11662,N_11539);
xor U12021 (N_12021,N_11716,N_11825);
xor U12022 (N_12022,N_11655,N_11652);
nor U12023 (N_12023,N_11867,N_11983);
or U12024 (N_12024,N_11707,N_11857);
nor U12025 (N_12025,N_11837,N_11633);
nand U12026 (N_12026,N_11518,N_11748);
xnor U12027 (N_12027,N_11612,N_11690);
nand U12028 (N_12028,N_11705,N_11513);
nand U12029 (N_12029,N_11903,N_11767);
nand U12030 (N_12030,N_11579,N_11509);
or U12031 (N_12031,N_11930,N_11853);
nor U12032 (N_12032,N_11807,N_11814);
xor U12033 (N_12033,N_11944,N_11952);
and U12034 (N_12034,N_11519,N_11792);
xnor U12035 (N_12035,N_11540,N_11526);
xor U12036 (N_12036,N_11967,N_11770);
or U12037 (N_12037,N_11892,N_11987);
or U12038 (N_12038,N_11847,N_11762);
nor U12039 (N_12039,N_11573,N_11615);
nor U12040 (N_12040,N_11833,N_11681);
and U12041 (N_12041,N_11605,N_11920);
nand U12042 (N_12042,N_11891,N_11563);
or U12043 (N_12043,N_11817,N_11759);
or U12044 (N_12044,N_11985,N_11672);
xor U12045 (N_12045,N_11811,N_11787);
nand U12046 (N_12046,N_11528,N_11890);
xnor U12047 (N_12047,N_11934,N_11553);
nor U12048 (N_12048,N_11758,N_11585);
xnor U12049 (N_12049,N_11597,N_11546);
or U12050 (N_12050,N_11941,N_11711);
and U12051 (N_12051,N_11824,N_11856);
nor U12052 (N_12052,N_11960,N_11973);
xnor U12053 (N_12053,N_11704,N_11924);
xnor U12054 (N_12054,N_11834,N_11555);
nand U12055 (N_12055,N_11557,N_11986);
nand U12056 (N_12056,N_11777,N_11950);
xor U12057 (N_12057,N_11516,N_11572);
nor U12058 (N_12058,N_11932,N_11799);
or U12059 (N_12059,N_11700,N_11904);
nand U12060 (N_12060,N_11945,N_11803);
nand U12061 (N_12061,N_11689,N_11841);
nand U12062 (N_12062,N_11679,N_11603);
nor U12063 (N_12063,N_11525,N_11744);
or U12064 (N_12064,N_11593,N_11609);
nor U12065 (N_12065,N_11931,N_11974);
xor U12066 (N_12066,N_11552,N_11649);
nand U12067 (N_12067,N_11873,N_11659);
xnor U12068 (N_12068,N_11625,N_11629);
nand U12069 (N_12069,N_11502,N_11794);
or U12070 (N_12070,N_11898,N_11747);
xor U12071 (N_12071,N_11874,N_11883);
and U12072 (N_12072,N_11780,N_11547);
nand U12073 (N_12073,N_11795,N_11984);
xor U12074 (N_12074,N_11999,N_11589);
nand U12075 (N_12075,N_11644,N_11586);
nand U12076 (N_12076,N_11627,N_11512);
nand U12077 (N_12077,N_11783,N_11899);
or U12078 (N_12078,N_11750,N_11746);
or U12079 (N_12079,N_11570,N_11953);
xor U12080 (N_12080,N_11562,N_11840);
nand U12081 (N_12081,N_11743,N_11982);
nand U12082 (N_12082,N_11855,N_11910);
or U12083 (N_12083,N_11727,N_11595);
nand U12084 (N_12084,N_11879,N_11755);
and U12085 (N_12085,N_11677,N_11607);
and U12086 (N_12086,N_11949,N_11821);
xnor U12087 (N_12087,N_11617,N_11768);
or U12088 (N_12088,N_11948,N_11975);
or U12089 (N_12089,N_11893,N_11622);
nor U12090 (N_12090,N_11802,N_11541);
or U12091 (N_12091,N_11511,N_11714);
or U12092 (N_12092,N_11927,N_11507);
and U12093 (N_12093,N_11889,N_11523);
or U12094 (N_12094,N_11925,N_11631);
or U12095 (N_12095,N_11670,N_11610);
xnor U12096 (N_12096,N_11545,N_11703);
nor U12097 (N_12097,N_11506,N_11793);
xor U12098 (N_12098,N_11699,N_11872);
nand U12099 (N_12099,N_11500,N_11532);
xnor U12100 (N_12100,N_11839,N_11901);
or U12101 (N_12101,N_11749,N_11963);
nand U12102 (N_12102,N_11550,N_11708);
and U12103 (N_12103,N_11692,N_11621);
nand U12104 (N_12104,N_11537,N_11940);
nand U12105 (N_12105,N_11571,N_11544);
xor U12106 (N_12106,N_11896,N_11774);
and U12107 (N_12107,N_11905,N_11616);
nand U12108 (N_12108,N_11914,N_11567);
nand U12109 (N_12109,N_11582,N_11718);
nor U12110 (N_12110,N_11971,N_11591);
and U12111 (N_12111,N_11574,N_11776);
and U12112 (N_12112,N_11638,N_11527);
or U12113 (N_12113,N_11884,N_11788);
xor U12114 (N_12114,N_11624,N_11864);
nor U12115 (N_12115,N_11863,N_11994);
and U12116 (N_12116,N_11858,N_11740);
xnor U12117 (N_12117,N_11875,N_11671);
and U12118 (N_12118,N_11565,N_11520);
and U12119 (N_12119,N_11614,N_11870);
nand U12120 (N_12120,N_11850,N_11643);
xor U12121 (N_12121,N_11697,N_11632);
or U12122 (N_12122,N_11669,N_11815);
nor U12123 (N_12123,N_11654,N_11849);
xnor U12124 (N_12124,N_11976,N_11658);
nor U12125 (N_12125,N_11656,N_11909);
xor U12126 (N_12126,N_11843,N_11797);
and U12127 (N_12127,N_11946,N_11623);
or U12128 (N_12128,N_11937,N_11878);
or U12129 (N_12129,N_11694,N_11583);
and U12130 (N_12130,N_11868,N_11885);
nand U12131 (N_12131,N_11737,N_11647);
xnor U12132 (N_12132,N_11600,N_11628);
nor U12133 (N_12133,N_11554,N_11508);
nor U12134 (N_12134,N_11561,N_11729);
nand U12135 (N_12135,N_11559,N_11693);
or U12136 (N_12136,N_11753,N_11608);
nor U12137 (N_12137,N_11517,N_11745);
xnor U12138 (N_12138,N_11696,N_11678);
and U12139 (N_12139,N_11501,N_11653);
nand U12140 (N_12140,N_11846,N_11587);
xnor U12141 (N_12141,N_11916,N_11646);
nor U12142 (N_12142,N_11912,N_11732);
nand U12143 (N_12143,N_11535,N_11980);
or U12144 (N_12144,N_11775,N_11998);
and U12145 (N_12145,N_11876,N_11730);
and U12146 (N_12146,N_11635,N_11505);
and U12147 (N_12147,N_11859,N_11995);
nor U12148 (N_12148,N_11599,N_11789);
nand U12149 (N_12149,N_11710,N_11804);
nor U12150 (N_12150,N_11935,N_11645);
xor U12151 (N_12151,N_11606,N_11993);
nor U12152 (N_12152,N_11733,N_11503);
or U12153 (N_12153,N_11524,N_11828);
xnor U12154 (N_12154,N_11791,N_11663);
and U12155 (N_12155,N_11726,N_11685);
xor U12156 (N_12156,N_11619,N_11835);
nand U12157 (N_12157,N_11549,N_11723);
and U12158 (N_12158,N_11760,N_11590);
nor U12159 (N_12159,N_11636,N_11581);
nand U12160 (N_12160,N_11640,N_11687);
or U12161 (N_12161,N_11515,N_11683);
xor U12162 (N_12162,N_11796,N_11830);
nand U12163 (N_12163,N_11551,N_11956);
xnor U12164 (N_12164,N_11992,N_11548);
and U12165 (N_12165,N_11785,N_11522);
nor U12166 (N_12166,N_11642,N_11919);
xor U12167 (N_12167,N_11826,N_11531);
and U12168 (N_12168,N_11782,N_11578);
xnor U12169 (N_12169,N_11822,N_11997);
and U12170 (N_12170,N_11965,N_11954);
nor U12171 (N_12171,N_11720,N_11961);
xnor U12172 (N_12172,N_11991,N_11972);
nand U12173 (N_12173,N_11888,N_11584);
xor U12174 (N_12174,N_11751,N_11827);
nor U12175 (N_12175,N_11741,N_11861);
xnor U12176 (N_12176,N_11964,N_11766);
xnor U12177 (N_12177,N_11637,N_11897);
xnor U12178 (N_12178,N_11661,N_11602);
xor U12179 (N_12179,N_11979,N_11836);
or U12180 (N_12180,N_11695,N_11728);
nand U12181 (N_12181,N_11666,N_11929);
or U12182 (N_12182,N_11820,N_11988);
nor U12183 (N_12183,N_11838,N_11918);
nor U12184 (N_12184,N_11816,N_11786);
nor U12185 (N_12185,N_11757,N_11660);
nand U12186 (N_12186,N_11596,N_11854);
nor U12187 (N_12187,N_11558,N_11556);
and U12188 (N_12188,N_11739,N_11880);
xor U12189 (N_12189,N_11922,N_11911);
and U12190 (N_12190,N_11900,N_11977);
nor U12191 (N_12191,N_11813,N_11917);
or U12192 (N_12192,N_11831,N_11709);
nand U12193 (N_12193,N_11713,N_11626);
nor U12194 (N_12194,N_11754,N_11800);
xor U12195 (N_12195,N_11915,N_11611);
xnor U12196 (N_12196,N_11908,N_11594);
and U12197 (N_12197,N_11674,N_11676);
and U12198 (N_12198,N_11881,N_11772);
nand U12199 (N_12199,N_11877,N_11844);
nand U12200 (N_12200,N_11657,N_11808);
nand U12201 (N_12201,N_11968,N_11529);
xor U12202 (N_12202,N_11942,N_11569);
nor U12203 (N_12203,N_11810,N_11682);
nor U12204 (N_12204,N_11534,N_11943);
xor U12205 (N_12205,N_11978,N_11542);
xnor U12206 (N_12206,N_11701,N_11955);
or U12207 (N_12207,N_11966,N_11667);
xnor U12208 (N_12208,N_11798,N_11981);
and U12209 (N_12209,N_11691,N_11819);
xnor U12210 (N_12210,N_11939,N_11812);
and U12211 (N_12211,N_11719,N_11818);
and U12212 (N_12212,N_11568,N_11613);
nand U12213 (N_12213,N_11752,N_11990);
and U12214 (N_12214,N_11560,N_11648);
nand U12215 (N_12215,N_11575,N_11736);
nand U12216 (N_12216,N_11686,N_11970);
nor U12217 (N_12217,N_11734,N_11651);
and U12218 (N_12218,N_11742,N_11989);
or U12219 (N_12219,N_11521,N_11882);
and U12220 (N_12220,N_11923,N_11957);
and U12221 (N_12221,N_11722,N_11564);
and U12222 (N_12222,N_11869,N_11673);
nand U12223 (N_12223,N_11779,N_11790);
nand U12224 (N_12224,N_11717,N_11921);
xor U12225 (N_12225,N_11832,N_11829);
or U12226 (N_12226,N_11533,N_11866);
or U12227 (N_12227,N_11860,N_11588);
xor U12228 (N_12228,N_11886,N_11592);
and U12229 (N_12229,N_11576,N_11848);
and U12230 (N_12230,N_11738,N_11962);
nand U12231 (N_12231,N_11680,N_11634);
nor U12232 (N_12232,N_11566,N_11947);
xor U12233 (N_12233,N_11851,N_11823);
xnor U12234 (N_12234,N_11715,N_11933);
or U12235 (N_12235,N_11959,N_11852);
xnor U12236 (N_12236,N_11724,N_11698);
xor U12237 (N_12237,N_11620,N_11688);
xnor U12238 (N_12238,N_11845,N_11773);
nand U12239 (N_12239,N_11721,N_11598);
nor U12240 (N_12240,N_11601,N_11865);
and U12241 (N_12241,N_11913,N_11604);
and U12242 (N_12242,N_11902,N_11862);
nor U12243 (N_12243,N_11806,N_11887);
nand U12244 (N_12244,N_11504,N_11665);
and U12245 (N_12245,N_11781,N_11731);
or U12246 (N_12246,N_11895,N_11928);
and U12247 (N_12247,N_11771,N_11764);
xor U12248 (N_12248,N_11907,N_11996);
nor U12249 (N_12249,N_11936,N_11536);
xnor U12250 (N_12250,N_11533,N_11901);
and U12251 (N_12251,N_11709,N_11808);
and U12252 (N_12252,N_11553,N_11713);
or U12253 (N_12253,N_11707,N_11633);
xor U12254 (N_12254,N_11960,N_11806);
xnor U12255 (N_12255,N_11939,N_11860);
nand U12256 (N_12256,N_11792,N_11828);
or U12257 (N_12257,N_11585,N_11986);
xnor U12258 (N_12258,N_11585,N_11903);
or U12259 (N_12259,N_11949,N_11748);
and U12260 (N_12260,N_11942,N_11829);
nand U12261 (N_12261,N_11942,N_11798);
nor U12262 (N_12262,N_11619,N_11945);
xnor U12263 (N_12263,N_11536,N_11678);
xnor U12264 (N_12264,N_11907,N_11857);
nand U12265 (N_12265,N_11674,N_11769);
nand U12266 (N_12266,N_11512,N_11961);
xor U12267 (N_12267,N_11706,N_11739);
xnor U12268 (N_12268,N_11714,N_11723);
and U12269 (N_12269,N_11525,N_11884);
xor U12270 (N_12270,N_11978,N_11790);
nor U12271 (N_12271,N_11687,N_11866);
xnor U12272 (N_12272,N_11775,N_11563);
and U12273 (N_12273,N_11705,N_11511);
and U12274 (N_12274,N_11865,N_11580);
nor U12275 (N_12275,N_11608,N_11523);
and U12276 (N_12276,N_11637,N_11694);
xnor U12277 (N_12277,N_11633,N_11714);
nor U12278 (N_12278,N_11769,N_11933);
and U12279 (N_12279,N_11525,N_11891);
and U12280 (N_12280,N_11621,N_11721);
xor U12281 (N_12281,N_11930,N_11972);
or U12282 (N_12282,N_11585,N_11984);
nor U12283 (N_12283,N_11850,N_11890);
xnor U12284 (N_12284,N_11993,N_11774);
nand U12285 (N_12285,N_11808,N_11752);
nor U12286 (N_12286,N_11632,N_11775);
nand U12287 (N_12287,N_11523,N_11972);
xor U12288 (N_12288,N_11864,N_11507);
xnor U12289 (N_12289,N_11852,N_11992);
nor U12290 (N_12290,N_11773,N_11506);
nor U12291 (N_12291,N_11889,N_11794);
and U12292 (N_12292,N_11535,N_11902);
xor U12293 (N_12293,N_11605,N_11776);
nor U12294 (N_12294,N_11526,N_11765);
xnor U12295 (N_12295,N_11608,N_11857);
nand U12296 (N_12296,N_11673,N_11745);
and U12297 (N_12297,N_11827,N_11955);
or U12298 (N_12298,N_11813,N_11618);
xor U12299 (N_12299,N_11656,N_11605);
and U12300 (N_12300,N_11675,N_11797);
nand U12301 (N_12301,N_11791,N_11634);
xnor U12302 (N_12302,N_11566,N_11959);
and U12303 (N_12303,N_11956,N_11838);
and U12304 (N_12304,N_11573,N_11692);
or U12305 (N_12305,N_11790,N_11835);
and U12306 (N_12306,N_11752,N_11759);
xnor U12307 (N_12307,N_11840,N_11672);
or U12308 (N_12308,N_11833,N_11858);
nand U12309 (N_12309,N_11830,N_11978);
or U12310 (N_12310,N_11835,N_11818);
nor U12311 (N_12311,N_11521,N_11812);
or U12312 (N_12312,N_11942,N_11874);
nor U12313 (N_12313,N_11580,N_11648);
and U12314 (N_12314,N_11578,N_11583);
nor U12315 (N_12315,N_11757,N_11768);
and U12316 (N_12316,N_11635,N_11727);
or U12317 (N_12317,N_11729,N_11842);
nor U12318 (N_12318,N_11705,N_11691);
and U12319 (N_12319,N_11703,N_11864);
and U12320 (N_12320,N_11977,N_11866);
nand U12321 (N_12321,N_11907,N_11990);
nor U12322 (N_12322,N_11791,N_11921);
or U12323 (N_12323,N_11941,N_11924);
or U12324 (N_12324,N_11674,N_11861);
xnor U12325 (N_12325,N_11505,N_11935);
nand U12326 (N_12326,N_11526,N_11800);
xor U12327 (N_12327,N_11798,N_11644);
and U12328 (N_12328,N_11746,N_11915);
and U12329 (N_12329,N_11980,N_11990);
nor U12330 (N_12330,N_11549,N_11725);
nand U12331 (N_12331,N_11921,N_11873);
xnor U12332 (N_12332,N_11984,N_11555);
xor U12333 (N_12333,N_11868,N_11940);
nand U12334 (N_12334,N_11506,N_11591);
xor U12335 (N_12335,N_11947,N_11778);
and U12336 (N_12336,N_11904,N_11567);
nor U12337 (N_12337,N_11687,N_11920);
or U12338 (N_12338,N_11638,N_11892);
nor U12339 (N_12339,N_11760,N_11801);
xnor U12340 (N_12340,N_11751,N_11737);
or U12341 (N_12341,N_11558,N_11636);
xnor U12342 (N_12342,N_11677,N_11549);
xnor U12343 (N_12343,N_11942,N_11525);
xnor U12344 (N_12344,N_11742,N_11858);
and U12345 (N_12345,N_11879,N_11742);
xnor U12346 (N_12346,N_11733,N_11750);
nand U12347 (N_12347,N_11685,N_11917);
nor U12348 (N_12348,N_11938,N_11943);
and U12349 (N_12349,N_11823,N_11528);
nand U12350 (N_12350,N_11528,N_11748);
and U12351 (N_12351,N_11587,N_11945);
nor U12352 (N_12352,N_11867,N_11805);
and U12353 (N_12353,N_11625,N_11747);
or U12354 (N_12354,N_11994,N_11784);
or U12355 (N_12355,N_11640,N_11743);
nand U12356 (N_12356,N_11556,N_11822);
nor U12357 (N_12357,N_11843,N_11598);
nand U12358 (N_12358,N_11637,N_11794);
nor U12359 (N_12359,N_11951,N_11676);
nand U12360 (N_12360,N_11759,N_11680);
or U12361 (N_12361,N_11863,N_11587);
or U12362 (N_12362,N_11717,N_11555);
xnor U12363 (N_12363,N_11673,N_11750);
nor U12364 (N_12364,N_11743,N_11501);
nor U12365 (N_12365,N_11842,N_11816);
nand U12366 (N_12366,N_11702,N_11761);
xnor U12367 (N_12367,N_11955,N_11684);
nor U12368 (N_12368,N_11545,N_11825);
nor U12369 (N_12369,N_11734,N_11571);
or U12370 (N_12370,N_11525,N_11630);
and U12371 (N_12371,N_11528,N_11838);
and U12372 (N_12372,N_11867,N_11713);
and U12373 (N_12373,N_11605,N_11696);
nor U12374 (N_12374,N_11574,N_11829);
and U12375 (N_12375,N_11817,N_11958);
and U12376 (N_12376,N_11609,N_11537);
nand U12377 (N_12377,N_11611,N_11770);
and U12378 (N_12378,N_11845,N_11686);
nor U12379 (N_12379,N_11876,N_11949);
nor U12380 (N_12380,N_11824,N_11878);
xnor U12381 (N_12381,N_11797,N_11776);
nand U12382 (N_12382,N_11913,N_11693);
xor U12383 (N_12383,N_11828,N_11744);
nand U12384 (N_12384,N_11503,N_11623);
or U12385 (N_12385,N_11673,N_11918);
and U12386 (N_12386,N_11552,N_11857);
or U12387 (N_12387,N_11727,N_11609);
nand U12388 (N_12388,N_11513,N_11701);
xor U12389 (N_12389,N_11632,N_11597);
nand U12390 (N_12390,N_11793,N_11667);
xnor U12391 (N_12391,N_11985,N_11904);
and U12392 (N_12392,N_11781,N_11659);
and U12393 (N_12393,N_11911,N_11647);
xnor U12394 (N_12394,N_11627,N_11602);
xor U12395 (N_12395,N_11834,N_11673);
nand U12396 (N_12396,N_11874,N_11939);
and U12397 (N_12397,N_11627,N_11908);
xnor U12398 (N_12398,N_11824,N_11798);
nand U12399 (N_12399,N_11508,N_11746);
xnor U12400 (N_12400,N_11802,N_11782);
nor U12401 (N_12401,N_11578,N_11594);
nand U12402 (N_12402,N_11804,N_11518);
or U12403 (N_12403,N_11627,N_11762);
or U12404 (N_12404,N_11559,N_11665);
nand U12405 (N_12405,N_11889,N_11812);
or U12406 (N_12406,N_11575,N_11834);
or U12407 (N_12407,N_11701,N_11584);
nor U12408 (N_12408,N_11974,N_11771);
and U12409 (N_12409,N_11520,N_11926);
nand U12410 (N_12410,N_11816,N_11689);
nor U12411 (N_12411,N_11804,N_11826);
and U12412 (N_12412,N_11946,N_11709);
or U12413 (N_12413,N_11986,N_11869);
xnor U12414 (N_12414,N_11686,N_11846);
nor U12415 (N_12415,N_11654,N_11876);
and U12416 (N_12416,N_11804,N_11505);
xnor U12417 (N_12417,N_11618,N_11719);
xor U12418 (N_12418,N_11718,N_11743);
and U12419 (N_12419,N_11866,N_11696);
nand U12420 (N_12420,N_11981,N_11951);
nand U12421 (N_12421,N_11589,N_11740);
nor U12422 (N_12422,N_11622,N_11975);
or U12423 (N_12423,N_11606,N_11696);
xnor U12424 (N_12424,N_11565,N_11766);
xnor U12425 (N_12425,N_11676,N_11800);
or U12426 (N_12426,N_11882,N_11667);
and U12427 (N_12427,N_11829,N_11770);
nand U12428 (N_12428,N_11623,N_11745);
nor U12429 (N_12429,N_11636,N_11780);
xor U12430 (N_12430,N_11502,N_11862);
and U12431 (N_12431,N_11979,N_11547);
nand U12432 (N_12432,N_11969,N_11906);
xor U12433 (N_12433,N_11717,N_11632);
or U12434 (N_12434,N_11536,N_11921);
and U12435 (N_12435,N_11836,N_11783);
nor U12436 (N_12436,N_11565,N_11538);
nand U12437 (N_12437,N_11919,N_11763);
nand U12438 (N_12438,N_11770,N_11868);
or U12439 (N_12439,N_11645,N_11739);
or U12440 (N_12440,N_11696,N_11787);
nand U12441 (N_12441,N_11716,N_11672);
nor U12442 (N_12442,N_11971,N_11693);
or U12443 (N_12443,N_11796,N_11611);
nand U12444 (N_12444,N_11773,N_11649);
nand U12445 (N_12445,N_11984,N_11658);
or U12446 (N_12446,N_11683,N_11690);
xnor U12447 (N_12447,N_11877,N_11739);
nand U12448 (N_12448,N_11987,N_11571);
or U12449 (N_12449,N_11502,N_11894);
xor U12450 (N_12450,N_11583,N_11685);
nand U12451 (N_12451,N_11536,N_11643);
xnor U12452 (N_12452,N_11642,N_11988);
or U12453 (N_12453,N_11768,N_11976);
or U12454 (N_12454,N_11693,N_11967);
or U12455 (N_12455,N_11850,N_11535);
or U12456 (N_12456,N_11923,N_11985);
and U12457 (N_12457,N_11608,N_11504);
nand U12458 (N_12458,N_11993,N_11888);
or U12459 (N_12459,N_11866,N_11581);
xor U12460 (N_12460,N_11680,N_11973);
and U12461 (N_12461,N_11660,N_11719);
nand U12462 (N_12462,N_11567,N_11512);
nand U12463 (N_12463,N_11582,N_11968);
xor U12464 (N_12464,N_11970,N_11637);
and U12465 (N_12465,N_11627,N_11530);
nand U12466 (N_12466,N_11728,N_11619);
xnor U12467 (N_12467,N_11517,N_11515);
nor U12468 (N_12468,N_11985,N_11943);
or U12469 (N_12469,N_11911,N_11818);
and U12470 (N_12470,N_11974,N_11883);
nand U12471 (N_12471,N_11996,N_11706);
nand U12472 (N_12472,N_11546,N_11956);
nor U12473 (N_12473,N_11701,N_11859);
nor U12474 (N_12474,N_11742,N_11817);
nor U12475 (N_12475,N_11904,N_11752);
or U12476 (N_12476,N_11796,N_11573);
and U12477 (N_12477,N_11679,N_11795);
and U12478 (N_12478,N_11536,N_11989);
and U12479 (N_12479,N_11648,N_11825);
and U12480 (N_12480,N_11868,N_11603);
or U12481 (N_12481,N_11972,N_11894);
and U12482 (N_12482,N_11546,N_11845);
xor U12483 (N_12483,N_11891,N_11858);
and U12484 (N_12484,N_11973,N_11877);
and U12485 (N_12485,N_11673,N_11856);
or U12486 (N_12486,N_11562,N_11572);
nand U12487 (N_12487,N_11558,N_11707);
or U12488 (N_12488,N_11595,N_11552);
or U12489 (N_12489,N_11711,N_11679);
nand U12490 (N_12490,N_11833,N_11723);
nor U12491 (N_12491,N_11911,N_11802);
or U12492 (N_12492,N_11600,N_11590);
or U12493 (N_12493,N_11617,N_11962);
nand U12494 (N_12494,N_11956,N_11974);
nor U12495 (N_12495,N_11767,N_11779);
nor U12496 (N_12496,N_11628,N_11927);
xor U12497 (N_12497,N_11834,N_11860);
or U12498 (N_12498,N_11939,N_11732);
xnor U12499 (N_12499,N_11856,N_11628);
xnor U12500 (N_12500,N_12296,N_12273);
and U12501 (N_12501,N_12003,N_12269);
nand U12502 (N_12502,N_12375,N_12491);
nand U12503 (N_12503,N_12496,N_12290);
xnor U12504 (N_12504,N_12316,N_12390);
nor U12505 (N_12505,N_12358,N_12477);
nor U12506 (N_12506,N_12180,N_12445);
nand U12507 (N_12507,N_12173,N_12171);
nand U12508 (N_12508,N_12061,N_12382);
nand U12509 (N_12509,N_12054,N_12449);
nor U12510 (N_12510,N_12134,N_12387);
nand U12511 (N_12511,N_12189,N_12106);
nand U12512 (N_12512,N_12029,N_12009);
nor U12513 (N_12513,N_12367,N_12069);
or U12514 (N_12514,N_12439,N_12337);
xnor U12515 (N_12515,N_12287,N_12323);
xor U12516 (N_12516,N_12100,N_12179);
and U12517 (N_12517,N_12408,N_12192);
and U12518 (N_12518,N_12128,N_12129);
nor U12519 (N_12519,N_12056,N_12321);
nor U12520 (N_12520,N_12347,N_12348);
nand U12521 (N_12521,N_12379,N_12473);
xnor U12522 (N_12522,N_12286,N_12116);
xnor U12523 (N_12523,N_12088,N_12036);
or U12524 (N_12524,N_12410,N_12031);
nand U12525 (N_12525,N_12064,N_12083);
and U12526 (N_12526,N_12479,N_12193);
nand U12527 (N_12527,N_12455,N_12428);
xnor U12528 (N_12528,N_12080,N_12198);
and U12529 (N_12529,N_12177,N_12291);
xor U12530 (N_12530,N_12312,N_12174);
nand U12531 (N_12531,N_12463,N_12395);
or U12532 (N_12532,N_12006,N_12397);
nor U12533 (N_12533,N_12470,N_12331);
xor U12534 (N_12534,N_12049,N_12482);
xnor U12535 (N_12535,N_12362,N_12032);
and U12536 (N_12536,N_12209,N_12462);
nor U12537 (N_12537,N_12452,N_12404);
nand U12538 (N_12538,N_12188,N_12438);
xor U12539 (N_12539,N_12227,N_12097);
or U12540 (N_12540,N_12242,N_12152);
nand U12541 (N_12541,N_12051,N_12153);
or U12542 (N_12542,N_12121,N_12306);
nor U12543 (N_12543,N_12057,N_12026);
nor U12544 (N_12544,N_12386,N_12046);
nand U12545 (N_12545,N_12433,N_12266);
and U12546 (N_12546,N_12248,N_12454);
nor U12547 (N_12547,N_12494,N_12234);
and U12548 (N_12548,N_12254,N_12063);
and U12549 (N_12549,N_12341,N_12369);
nand U12550 (N_12550,N_12474,N_12424);
xnor U12551 (N_12551,N_12210,N_12246);
xnor U12552 (N_12552,N_12484,N_12401);
xor U12553 (N_12553,N_12075,N_12377);
nand U12554 (N_12554,N_12004,N_12270);
or U12555 (N_12555,N_12368,N_12344);
and U12556 (N_12556,N_12156,N_12487);
or U12557 (N_12557,N_12353,N_12374);
or U12558 (N_12558,N_12175,N_12115);
nand U12559 (N_12559,N_12238,N_12328);
xor U12560 (N_12560,N_12262,N_12154);
nand U12561 (N_12561,N_12235,N_12357);
xnor U12562 (N_12562,N_12403,N_12478);
xor U12563 (N_12563,N_12044,N_12412);
nand U12564 (N_12564,N_12010,N_12340);
nand U12565 (N_12565,N_12309,N_12371);
nand U12566 (N_12566,N_12264,N_12411);
nand U12567 (N_12567,N_12278,N_12030);
xnor U12568 (N_12568,N_12232,N_12435);
nand U12569 (N_12569,N_12355,N_12111);
and U12570 (N_12570,N_12087,N_12033);
nand U12571 (N_12571,N_12204,N_12372);
or U12572 (N_12572,N_12011,N_12140);
xnor U12573 (N_12573,N_12079,N_12440);
xor U12574 (N_12574,N_12119,N_12486);
or U12575 (N_12575,N_12142,N_12109);
and U12576 (N_12576,N_12418,N_12099);
nor U12577 (N_12577,N_12332,N_12050);
xnor U12578 (N_12578,N_12359,N_12365);
nor U12579 (N_12579,N_12441,N_12240);
or U12580 (N_12580,N_12135,N_12195);
nor U12581 (N_12581,N_12336,N_12216);
or U12582 (N_12582,N_12074,N_12320);
or U12583 (N_12583,N_12166,N_12161);
or U12584 (N_12584,N_12131,N_12190);
xnor U12585 (N_12585,N_12409,N_12400);
nor U12586 (N_12586,N_12007,N_12313);
nand U12587 (N_12587,N_12149,N_12275);
nand U12588 (N_12588,N_12257,N_12228);
xnor U12589 (N_12589,N_12416,N_12392);
xnor U12590 (N_12590,N_12151,N_12101);
and U12591 (N_12591,N_12251,N_12429);
nand U12592 (N_12592,N_12191,N_12060);
and U12593 (N_12593,N_12095,N_12324);
nor U12594 (N_12594,N_12492,N_12253);
nand U12595 (N_12595,N_12342,N_12130);
and U12596 (N_12596,N_12127,N_12094);
or U12597 (N_12597,N_12202,N_12460);
and U12598 (N_12598,N_12447,N_12233);
nor U12599 (N_12599,N_12421,N_12308);
nor U12600 (N_12600,N_12059,N_12349);
xnor U12601 (N_12601,N_12488,N_12292);
and U12602 (N_12602,N_12495,N_12393);
xor U12603 (N_12603,N_12468,N_12394);
or U12604 (N_12604,N_12098,N_12102);
or U12605 (N_12605,N_12018,N_12274);
nor U12606 (N_12606,N_12459,N_12008);
xor U12607 (N_12607,N_12081,N_12268);
nand U12608 (N_12608,N_12398,N_12304);
and U12609 (N_12609,N_12147,N_12014);
nand U12610 (N_12610,N_12295,N_12108);
nand U12611 (N_12611,N_12071,N_12105);
or U12612 (N_12612,N_12443,N_12196);
nand U12613 (N_12613,N_12072,N_12413);
and U12614 (N_12614,N_12084,N_12110);
and U12615 (N_12615,N_12381,N_12112);
and U12616 (N_12616,N_12241,N_12453);
xor U12617 (N_12617,N_12489,N_12001);
xnor U12618 (N_12618,N_12255,N_12294);
nor U12619 (N_12619,N_12226,N_12126);
nor U12620 (N_12620,N_12194,N_12045);
xnor U12621 (N_12621,N_12082,N_12422);
nand U12622 (N_12622,N_12035,N_12158);
or U12623 (N_12623,N_12258,N_12475);
nor U12624 (N_12624,N_12385,N_12338);
xnor U12625 (N_12625,N_12457,N_12466);
or U12626 (N_12626,N_12481,N_12461);
or U12627 (N_12627,N_12148,N_12176);
or U12628 (N_12628,N_12263,N_12282);
nor U12629 (N_12629,N_12444,N_12172);
and U12630 (N_12630,N_12483,N_12053);
nor U12631 (N_12631,N_12016,N_12252);
nor U12632 (N_12632,N_12005,N_12089);
and U12633 (N_12633,N_12243,N_12187);
or U12634 (N_12634,N_12334,N_12427);
or U12635 (N_12635,N_12157,N_12021);
and U12636 (N_12636,N_12327,N_12048);
nor U12637 (N_12637,N_12042,N_12467);
nand U12638 (N_12638,N_12376,N_12318);
and U12639 (N_12639,N_12213,N_12464);
nor U12640 (N_12640,N_12034,N_12025);
xnor U12641 (N_12641,N_12230,N_12093);
xnor U12642 (N_12642,N_12027,N_12448);
nand U12643 (N_12643,N_12162,N_12038);
or U12644 (N_12644,N_12039,N_12207);
nand U12645 (N_12645,N_12335,N_12271);
or U12646 (N_12646,N_12420,N_12450);
nor U12647 (N_12647,N_12378,N_12086);
xor U12648 (N_12648,N_12302,N_12247);
and U12649 (N_12649,N_12236,N_12244);
nand U12650 (N_12650,N_12123,N_12310);
or U12651 (N_12651,N_12333,N_12000);
or U12652 (N_12652,N_12345,N_12406);
nor U12653 (N_12653,N_12476,N_12017);
nand U12654 (N_12654,N_12396,N_12352);
nor U12655 (N_12655,N_12208,N_12212);
nand U12656 (N_12656,N_12297,N_12480);
nand U12657 (N_12657,N_12138,N_12360);
xor U12658 (N_12658,N_12322,N_12499);
nor U12659 (N_12659,N_12013,N_12430);
nor U12660 (N_12660,N_12419,N_12062);
nor U12661 (N_12661,N_12317,N_12144);
nor U12662 (N_12662,N_12206,N_12019);
xor U12663 (N_12663,N_12052,N_12022);
nand U12664 (N_12664,N_12145,N_12199);
and U12665 (N_12665,N_12218,N_12103);
nand U12666 (N_12666,N_12326,N_12283);
nor U12667 (N_12667,N_12136,N_12222);
or U12668 (N_12668,N_12041,N_12169);
and U12669 (N_12669,N_12389,N_12485);
nor U12670 (N_12670,N_12436,N_12301);
nand U12671 (N_12671,N_12402,N_12167);
nand U12672 (N_12672,N_12104,N_12343);
nand U12673 (N_12673,N_12002,N_12160);
and U12674 (N_12674,N_12307,N_12077);
nand U12675 (N_12675,N_12245,N_12280);
or U12676 (N_12676,N_12329,N_12465);
and U12677 (N_12677,N_12155,N_12183);
nand U12678 (N_12678,N_12137,N_12182);
and U12679 (N_12679,N_12366,N_12311);
or U12680 (N_12680,N_12350,N_12472);
nand U12681 (N_12681,N_12380,N_12250);
nand U12682 (N_12682,N_12170,N_12040);
nor U12683 (N_12683,N_12091,N_12217);
and U12684 (N_12684,N_12224,N_12107);
nor U12685 (N_12685,N_12139,N_12314);
xnor U12686 (N_12686,N_12065,N_12184);
nor U12687 (N_12687,N_12415,N_12165);
nand U12688 (N_12688,N_12164,N_12425);
or U12689 (N_12689,N_12339,N_12426);
xnor U12690 (N_12690,N_12078,N_12383);
and U12691 (N_12691,N_12351,N_12434);
nand U12692 (N_12692,N_12285,N_12361);
nand U12693 (N_12693,N_12220,N_12205);
or U12694 (N_12694,N_12047,N_12023);
and U12695 (N_12695,N_12085,N_12281);
xnor U12696 (N_12696,N_12432,N_12346);
nor U12697 (N_12697,N_12370,N_12414);
nor U12698 (N_12698,N_12260,N_12118);
and U12699 (N_12699,N_12117,N_12181);
nand U12700 (N_12700,N_12015,N_12214);
xor U12701 (N_12701,N_12237,N_12122);
or U12702 (N_12702,N_12229,N_12067);
nor U12703 (N_12703,N_12076,N_12293);
and U12704 (N_12704,N_12388,N_12090);
or U12705 (N_12705,N_12325,N_12070);
xnor U12706 (N_12706,N_12277,N_12299);
or U12707 (N_12707,N_12141,N_12120);
or U12708 (N_12708,N_12300,N_12498);
nor U12709 (N_12709,N_12456,N_12143);
and U12710 (N_12710,N_12159,N_12407);
nand U12711 (N_12711,N_12146,N_12330);
nor U12712 (N_12712,N_12219,N_12092);
and U12713 (N_12713,N_12289,N_12223);
and U12714 (N_12714,N_12305,N_12267);
nor U12715 (N_12715,N_12055,N_12451);
nor U12716 (N_12716,N_12058,N_12239);
or U12717 (N_12717,N_12020,N_12114);
nor U12718 (N_12718,N_12279,N_12132);
or U12719 (N_12719,N_12276,N_12231);
and U12720 (N_12720,N_12442,N_12469);
nand U12721 (N_12721,N_12259,N_12225);
xor U12722 (N_12722,N_12261,N_12423);
nand U12723 (N_12723,N_12288,N_12391);
nor U12724 (N_12724,N_12265,N_12356);
or U12725 (N_12725,N_12012,N_12354);
nor U12726 (N_12726,N_12471,N_12163);
or U12727 (N_12727,N_12185,N_12458);
and U12728 (N_12728,N_12073,N_12319);
xnor U12729 (N_12729,N_12197,N_12364);
nand U12730 (N_12730,N_12028,N_12203);
nor U12731 (N_12731,N_12168,N_12399);
or U12732 (N_12732,N_12215,N_12066);
or U12733 (N_12733,N_12497,N_12221);
nand U12734 (N_12734,N_12431,N_12303);
or U12735 (N_12735,N_12043,N_12113);
and U12736 (N_12736,N_12249,N_12037);
nor U12737 (N_12737,N_12490,N_12315);
and U12738 (N_12738,N_12133,N_12201);
xnor U12739 (N_12739,N_12446,N_12272);
nor U12740 (N_12740,N_12178,N_12024);
and U12741 (N_12741,N_12284,N_12363);
or U12742 (N_12742,N_12096,N_12373);
or U12743 (N_12743,N_12493,N_12200);
xor U12744 (N_12744,N_12068,N_12256);
or U12745 (N_12745,N_12125,N_12186);
xor U12746 (N_12746,N_12150,N_12124);
and U12747 (N_12747,N_12298,N_12437);
nand U12748 (N_12748,N_12384,N_12405);
nor U12749 (N_12749,N_12211,N_12417);
nand U12750 (N_12750,N_12321,N_12135);
nand U12751 (N_12751,N_12173,N_12400);
nand U12752 (N_12752,N_12195,N_12152);
xnor U12753 (N_12753,N_12245,N_12162);
and U12754 (N_12754,N_12000,N_12147);
and U12755 (N_12755,N_12120,N_12397);
xor U12756 (N_12756,N_12473,N_12324);
and U12757 (N_12757,N_12090,N_12466);
or U12758 (N_12758,N_12449,N_12101);
or U12759 (N_12759,N_12188,N_12214);
nor U12760 (N_12760,N_12065,N_12178);
nor U12761 (N_12761,N_12151,N_12304);
or U12762 (N_12762,N_12291,N_12444);
nand U12763 (N_12763,N_12124,N_12447);
nor U12764 (N_12764,N_12466,N_12023);
and U12765 (N_12765,N_12465,N_12391);
nand U12766 (N_12766,N_12158,N_12493);
xor U12767 (N_12767,N_12170,N_12342);
nand U12768 (N_12768,N_12230,N_12220);
and U12769 (N_12769,N_12461,N_12413);
nand U12770 (N_12770,N_12097,N_12185);
nand U12771 (N_12771,N_12144,N_12233);
nor U12772 (N_12772,N_12209,N_12135);
nand U12773 (N_12773,N_12118,N_12204);
nand U12774 (N_12774,N_12366,N_12492);
and U12775 (N_12775,N_12087,N_12274);
or U12776 (N_12776,N_12030,N_12272);
xor U12777 (N_12777,N_12464,N_12423);
nor U12778 (N_12778,N_12039,N_12494);
xor U12779 (N_12779,N_12316,N_12169);
nor U12780 (N_12780,N_12251,N_12304);
and U12781 (N_12781,N_12469,N_12397);
nor U12782 (N_12782,N_12485,N_12321);
and U12783 (N_12783,N_12141,N_12274);
nand U12784 (N_12784,N_12038,N_12224);
nand U12785 (N_12785,N_12151,N_12013);
xor U12786 (N_12786,N_12276,N_12101);
or U12787 (N_12787,N_12157,N_12238);
and U12788 (N_12788,N_12469,N_12050);
nor U12789 (N_12789,N_12235,N_12279);
and U12790 (N_12790,N_12429,N_12345);
nor U12791 (N_12791,N_12052,N_12074);
nor U12792 (N_12792,N_12084,N_12115);
or U12793 (N_12793,N_12082,N_12404);
or U12794 (N_12794,N_12360,N_12260);
nand U12795 (N_12795,N_12351,N_12122);
nor U12796 (N_12796,N_12108,N_12483);
xor U12797 (N_12797,N_12468,N_12170);
and U12798 (N_12798,N_12021,N_12389);
nor U12799 (N_12799,N_12207,N_12202);
nand U12800 (N_12800,N_12013,N_12225);
xnor U12801 (N_12801,N_12099,N_12341);
xnor U12802 (N_12802,N_12048,N_12285);
and U12803 (N_12803,N_12044,N_12396);
and U12804 (N_12804,N_12357,N_12416);
and U12805 (N_12805,N_12444,N_12386);
or U12806 (N_12806,N_12482,N_12083);
xnor U12807 (N_12807,N_12481,N_12168);
and U12808 (N_12808,N_12006,N_12168);
nand U12809 (N_12809,N_12446,N_12244);
xnor U12810 (N_12810,N_12346,N_12275);
xor U12811 (N_12811,N_12344,N_12332);
and U12812 (N_12812,N_12363,N_12440);
nand U12813 (N_12813,N_12009,N_12319);
nor U12814 (N_12814,N_12306,N_12383);
nand U12815 (N_12815,N_12168,N_12385);
nor U12816 (N_12816,N_12173,N_12460);
xor U12817 (N_12817,N_12062,N_12245);
nor U12818 (N_12818,N_12329,N_12227);
xnor U12819 (N_12819,N_12240,N_12161);
nor U12820 (N_12820,N_12481,N_12129);
xnor U12821 (N_12821,N_12000,N_12045);
or U12822 (N_12822,N_12238,N_12278);
nand U12823 (N_12823,N_12130,N_12171);
nand U12824 (N_12824,N_12341,N_12050);
or U12825 (N_12825,N_12090,N_12337);
and U12826 (N_12826,N_12032,N_12407);
or U12827 (N_12827,N_12341,N_12261);
and U12828 (N_12828,N_12206,N_12128);
or U12829 (N_12829,N_12383,N_12179);
or U12830 (N_12830,N_12452,N_12235);
and U12831 (N_12831,N_12388,N_12419);
or U12832 (N_12832,N_12411,N_12448);
nor U12833 (N_12833,N_12413,N_12424);
or U12834 (N_12834,N_12462,N_12384);
and U12835 (N_12835,N_12200,N_12239);
xor U12836 (N_12836,N_12102,N_12023);
xor U12837 (N_12837,N_12001,N_12003);
nor U12838 (N_12838,N_12067,N_12060);
nor U12839 (N_12839,N_12340,N_12175);
xor U12840 (N_12840,N_12470,N_12172);
nor U12841 (N_12841,N_12465,N_12240);
or U12842 (N_12842,N_12142,N_12413);
xnor U12843 (N_12843,N_12409,N_12027);
xor U12844 (N_12844,N_12332,N_12381);
xor U12845 (N_12845,N_12133,N_12109);
nand U12846 (N_12846,N_12360,N_12346);
and U12847 (N_12847,N_12294,N_12262);
or U12848 (N_12848,N_12270,N_12427);
nand U12849 (N_12849,N_12128,N_12242);
or U12850 (N_12850,N_12127,N_12027);
nor U12851 (N_12851,N_12330,N_12030);
xor U12852 (N_12852,N_12427,N_12132);
nor U12853 (N_12853,N_12004,N_12435);
and U12854 (N_12854,N_12042,N_12060);
and U12855 (N_12855,N_12412,N_12074);
xnor U12856 (N_12856,N_12043,N_12425);
nor U12857 (N_12857,N_12423,N_12206);
nor U12858 (N_12858,N_12270,N_12340);
or U12859 (N_12859,N_12035,N_12111);
nand U12860 (N_12860,N_12473,N_12079);
xor U12861 (N_12861,N_12279,N_12187);
nand U12862 (N_12862,N_12063,N_12330);
or U12863 (N_12863,N_12328,N_12243);
xnor U12864 (N_12864,N_12169,N_12335);
or U12865 (N_12865,N_12337,N_12260);
or U12866 (N_12866,N_12334,N_12128);
and U12867 (N_12867,N_12100,N_12089);
xnor U12868 (N_12868,N_12297,N_12396);
or U12869 (N_12869,N_12387,N_12194);
nand U12870 (N_12870,N_12244,N_12159);
or U12871 (N_12871,N_12374,N_12244);
and U12872 (N_12872,N_12051,N_12073);
nand U12873 (N_12873,N_12386,N_12274);
nand U12874 (N_12874,N_12157,N_12106);
xor U12875 (N_12875,N_12394,N_12464);
nand U12876 (N_12876,N_12157,N_12313);
nand U12877 (N_12877,N_12029,N_12465);
nand U12878 (N_12878,N_12084,N_12070);
xor U12879 (N_12879,N_12063,N_12055);
nor U12880 (N_12880,N_12049,N_12236);
xor U12881 (N_12881,N_12427,N_12477);
xor U12882 (N_12882,N_12082,N_12464);
or U12883 (N_12883,N_12187,N_12332);
and U12884 (N_12884,N_12404,N_12077);
nand U12885 (N_12885,N_12294,N_12455);
xnor U12886 (N_12886,N_12373,N_12151);
xnor U12887 (N_12887,N_12160,N_12347);
or U12888 (N_12888,N_12143,N_12207);
xor U12889 (N_12889,N_12407,N_12113);
nand U12890 (N_12890,N_12097,N_12266);
and U12891 (N_12891,N_12058,N_12137);
and U12892 (N_12892,N_12451,N_12327);
xnor U12893 (N_12893,N_12287,N_12166);
or U12894 (N_12894,N_12040,N_12073);
or U12895 (N_12895,N_12451,N_12036);
nand U12896 (N_12896,N_12024,N_12349);
nand U12897 (N_12897,N_12336,N_12277);
nand U12898 (N_12898,N_12364,N_12352);
nor U12899 (N_12899,N_12011,N_12242);
nor U12900 (N_12900,N_12395,N_12053);
nand U12901 (N_12901,N_12188,N_12409);
nor U12902 (N_12902,N_12320,N_12171);
or U12903 (N_12903,N_12141,N_12345);
and U12904 (N_12904,N_12394,N_12082);
nand U12905 (N_12905,N_12446,N_12119);
nor U12906 (N_12906,N_12198,N_12247);
and U12907 (N_12907,N_12141,N_12499);
or U12908 (N_12908,N_12136,N_12356);
nand U12909 (N_12909,N_12301,N_12151);
nand U12910 (N_12910,N_12055,N_12273);
and U12911 (N_12911,N_12096,N_12148);
and U12912 (N_12912,N_12280,N_12191);
nor U12913 (N_12913,N_12002,N_12236);
nand U12914 (N_12914,N_12496,N_12248);
xnor U12915 (N_12915,N_12105,N_12170);
or U12916 (N_12916,N_12044,N_12490);
and U12917 (N_12917,N_12063,N_12101);
and U12918 (N_12918,N_12106,N_12198);
xor U12919 (N_12919,N_12320,N_12484);
nand U12920 (N_12920,N_12178,N_12244);
or U12921 (N_12921,N_12150,N_12331);
nor U12922 (N_12922,N_12244,N_12052);
nor U12923 (N_12923,N_12241,N_12091);
and U12924 (N_12924,N_12254,N_12379);
and U12925 (N_12925,N_12431,N_12144);
and U12926 (N_12926,N_12081,N_12160);
or U12927 (N_12927,N_12329,N_12482);
xnor U12928 (N_12928,N_12238,N_12266);
and U12929 (N_12929,N_12498,N_12317);
xor U12930 (N_12930,N_12493,N_12201);
or U12931 (N_12931,N_12131,N_12153);
and U12932 (N_12932,N_12462,N_12029);
xnor U12933 (N_12933,N_12146,N_12271);
and U12934 (N_12934,N_12359,N_12279);
xor U12935 (N_12935,N_12002,N_12427);
xor U12936 (N_12936,N_12488,N_12149);
nor U12937 (N_12937,N_12231,N_12469);
nor U12938 (N_12938,N_12499,N_12226);
nand U12939 (N_12939,N_12041,N_12002);
or U12940 (N_12940,N_12254,N_12097);
nor U12941 (N_12941,N_12347,N_12125);
and U12942 (N_12942,N_12183,N_12445);
and U12943 (N_12943,N_12402,N_12303);
nor U12944 (N_12944,N_12284,N_12145);
nor U12945 (N_12945,N_12130,N_12380);
nor U12946 (N_12946,N_12203,N_12316);
xor U12947 (N_12947,N_12079,N_12177);
or U12948 (N_12948,N_12424,N_12000);
xor U12949 (N_12949,N_12311,N_12161);
xor U12950 (N_12950,N_12337,N_12479);
nand U12951 (N_12951,N_12352,N_12197);
xnor U12952 (N_12952,N_12196,N_12364);
nand U12953 (N_12953,N_12270,N_12013);
xnor U12954 (N_12954,N_12394,N_12035);
nand U12955 (N_12955,N_12493,N_12361);
xor U12956 (N_12956,N_12304,N_12001);
and U12957 (N_12957,N_12160,N_12053);
or U12958 (N_12958,N_12085,N_12170);
nor U12959 (N_12959,N_12122,N_12330);
and U12960 (N_12960,N_12179,N_12003);
nor U12961 (N_12961,N_12469,N_12235);
xnor U12962 (N_12962,N_12056,N_12351);
xnor U12963 (N_12963,N_12104,N_12124);
or U12964 (N_12964,N_12269,N_12225);
nor U12965 (N_12965,N_12175,N_12391);
or U12966 (N_12966,N_12274,N_12245);
or U12967 (N_12967,N_12137,N_12489);
xnor U12968 (N_12968,N_12102,N_12272);
nor U12969 (N_12969,N_12422,N_12450);
xor U12970 (N_12970,N_12251,N_12230);
and U12971 (N_12971,N_12046,N_12104);
nand U12972 (N_12972,N_12185,N_12013);
nor U12973 (N_12973,N_12039,N_12054);
nand U12974 (N_12974,N_12070,N_12346);
and U12975 (N_12975,N_12245,N_12366);
xor U12976 (N_12976,N_12261,N_12452);
nor U12977 (N_12977,N_12301,N_12270);
nand U12978 (N_12978,N_12374,N_12125);
nand U12979 (N_12979,N_12145,N_12142);
nand U12980 (N_12980,N_12317,N_12338);
nor U12981 (N_12981,N_12253,N_12015);
nand U12982 (N_12982,N_12310,N_12095);
nor U12983 (N_12983,N_12286,N_12386);
and U12984 (N_12984,N_12354,N_12003);
nand U12985 (N_12985,N_12201,N_12469);
nand U12986 (N_12986,N_12488,N_12337);
or U12987 (N_12987,N_12422,N_12418);
or U12988 (N_12988,N_12022,N_12275);
nor U12989 (N_12989,N_12481,N_12249);
nand U12990 (N_12990,N_12202,N_12375);
nand U12991 (N_12991,N_12211,N_12457);
or U12992 (N_12992,N_12310,N_12423);
xor U12993 (N_12993,N_12083,N_12203);
and U12994 (N_12994,N_12314,N_12457);
nor U12995 (N_12995,N_12273,N_12438);
nand U12996 (N_12996,N_12237,N_12371);
and U12997 (N_12997,N_12212,N_12289);
and U12998 (N_12998,N_12027,N_12144);
or U12999 (N_12999,N_12088,N_12259);
or U13000 (N_13000,N_12740,N_12757);
nor U13001 (N_13001,N_12591,N_12675);
nor U13002 (N_13002,N_12540,N_12941);
and U13003 (N_13003,N_12767,N_12866);
or U13004 (N_13004,N_12712,N_12959);
xnor U13005 (N_13005,N_12918,N_12728);
nor U13006 (N_13006,N_12636,N_12895);
and U13007 (N_13007,N_12676,N_12705);
xor U13008 (N_13008,N_12722,N_12585);
nand U13009 (N_13009,N_12642,N_12937);
nor U13010 (N_13010,N_12932,N_12853);
nand U13011 (N_13011,N_12517,N_12965);
xor U13012 (N_13012,N_12793,N_12551);
nor U13013 (N_13013,N_12758,N_12632);
xor U13014 (N_13014,N_12645,N_12592);
nor U13015 (N_13015,N_12766,N_12960);
or U13016 (N_13016,N_12610,N_12568);
or U13017 (N_13017,N_12977,N_12537);
and U13018 (N_13018,N_12673,N_12800);
nor U13019 (N_13019,N_12613,N_12761);
xnor U13020 (N_13020,N_12839,N_12683);
or U13021 (N_13021,N_12523,N_12858);
nor U13022 (N_13022,N_12648,N_12957);
xor U13023 (N_13023,N_12762,N_12899);
and U13024 (N_13024,N_12894,N_12611);
or U13025 (N_13025,N_12790,N_12527);
or U13026 (N_13026,N_12837,N_12565);
and U13027 (N_13027,N_12798,N_12542);
nand U13028 (N_13028,N_12804,N_12543);
and U13029 (N_13029,N_12562,N_12573);
or U13030 (N_13030,N_12588,N_12860);
xor U13031 (N_13031,N_12952,N_12909);
and U13032 (N_13032,N_12701,N_12943);
nor U13033 (N_13033,N_12940,N_12987);
nand U13034 (N_13034,N_12535,N_12963);
nand U13035 (N_13035,N_12521,N_12748);
and U13036 (N_13036,N_12902,N_12845);
xnor U13037 (N_13037,N_12975,N_12862);
xor U13038 (N_13038,N_12991,N_12704);
nor U13039 (N_13039,N_12802,N_12884);
nor U13040 (N_13040,N_12541,N_12631);
nor U13041 (N_13041,N_12516,N_12630);
or U13042 (N_13042,N_12928,N_12825);
nor U13043 (N_13043,N_12846,N_12984);
nor U13044 (N_13044,N_12580,N_12714);
xor U13045 (N_13045,N_12688,N_12544);
nor U13046 (N_13046,N_12737,N_12581);
nor U13047 (N_13047,N_12643,N_12951);
and U13048 (N_13048,N_12911,N_12921);
or U13049 (N_13049,N_12628,N_12560);
nand U13050 (N_13050,N_12785,N_12618);
nor U13051 (N_13051,N_12732,N_12892);
xor U13052 (N_13052,N_12603,N_12958);
or U13053 (N_13053,N_12575,N_12920);
xnor U13054 (N_13054,N_12770,N_12998);
or U13055 (N_13055,N_12811,N_12703);
nand U13056 (N_13056,N_12686,N_12882);
xor U13057 (N_13057,N_12566,N_12930);
nor U13058 (N_13058,N_12624,N_12854);
or U13059 (N_13059,N_12906,N_12679);
xnor U13060 (N_13060,N_12534,N_12731);
nor U13061 (N_13061,N_12742,N_12555);
or U13062 (N_13062,N_12794,N_12905);
nor U13063 (N_13063,N_12912,N_12914);
xor U13064 (N_13064,N_12824,N_12788);
nor U13065 (N_13065,N_12881,N_12868);
xor U13066 (N_13066,N_12848,N_12944);
and U13067 (N_13067,N_12723,N_12887);
nand U13068 (N_13068,N_12514,N_12653);
and U13069 (N_13069,N_12671,N_12572);
and U13070 (N_13070,N_12669,N_12590);
nor U13071 (N_13071,N_12769,N_12649);
and U13072 (N_13072,N_12900,N_12931);
nand U13073 (N_13073,N_12787,N_12525);
nor U13074 (N_13074,N_12996,N_12621);
and U13075 (N_13075,N_12518,N_12577);
or U13076 (N_13076,N_12847,N_12746);
and U13077 (N_13077,N_12936,N_12828);
nor U13078 (N_13078,N_12620,N_12893);
nand U13079 (N_13079,N_12609,N_12665);
xnor U13080 (N_13080,N_12536,N_12515);
or U13081 (N_13081,N_12946,N_12729);
or U13082 (N_13082,N_12771,N_12710);
nand U13083 (N_13083,N_12747,N_12834);
or U13084 (N_13084,N_12583,N_12644);
or U13085 (N_13085,N_12763,N_12961);
or U13086 (N_13086,N_12711,N_12997);
xnor U13087 (N_13087,N_12809,N_12656);
or U13088 (N_13088,N_12956,N_12744);
or U13089 (N_13089,N_12708,N_12838);
xor U13090 (N_13090,N_12614,N_12850);
nor U13091 (N_13091,N_12564,N_12657);
nor U13092 (N_13092,N_12922,N_12939);
nor U13093 (N_13093,N_12933,N_12806);
and U13094 (N_13094,N_12874,N_12780);
nor U13095 (N_13095,N_12559,N_12570);
xor U13096 (N_13096,N_12639,N_12797);
xor U13097 (N_13097,N_12813,N_12608);
nor U13098 (N_13098,N_12964,N_12992);
xor U13099 (N_13099,N_12972,N_12554);
xor U13100 (N_13100,N_12765,N_12795);
xnor U13101 (N_13101,N_12724,N_12721);
nand U13102 (N_13102,N_12883,N_12615);
and U13103 (N_13103,N_12563,N_12889);
xnor U13104 (N_13104,N_12815,N_12638);
xor U13105 (N_13105,N_12699,N_12859);
xor U13106 (N_13106,N_12971,N_12607);
or U13107 (N_13107,N_12764,N_12759);
and U13108 (N_13108,N_12947,N_12538);
nand U13109 (N_13109,N_12707,N_12955);
and U13110 (N_13110,N_12857,N_12796);
or U13111 (N_13111,N_12855,N_12807);
and U13112 (N_13112,N_12692,N_12916);
nor U13113 (N_13113,N_12550,N_12864);
nand U13114 (N_13114,N_12626,N_12879);
or U13115 (N_13115,N_12738,N_12500);
or U13116 (N_13116,N_12519,N_12617);
nand U13117 (N_13117,N_12548,N_12663);
or U13118 (N_13118,N_12924,N_12567);
or U13119 (N_13119,N_12844,N_12576);
nand U13120 (N_13120,N_12792,N_12980);
xor U13121 (N_13121,N_12784,N_12830);
and U13122 (N_13122,N_12612,N_12602);
nor U13123 (N_13123,N_12782,N_12507);
and U13124 (N_13124,N_12604,N_12768);
xor U13125 (N_13125,N_12662,N_12635);
xor U13126 (N_13126,N_12579,N_12901);
xnor U13127 (N_13127,N_12510,N_12739);
xor U13128 (N_13128,N_12741,N_12843);
or U13129 (N_13129,N_12552,N_12690);
and U13130 (N_13130,N_12973,N_12594);
nand U13131 (N_13131,N_12949,N_12664);
and U13132 (N_13132,N_12969,N_12715);
xor U13133 (N_13133,N_12826,N_12791);
and U13134 (N_13134,N_12526,N_12511);
nand U13135 (N_13135,N_12684,N_12598);
nor U13136 (N_13136,N_12896,N_12988);
nor U13137 (N_13137,N_12993,N_12942);
and U13138 (N_13138,N_12832,N_12908);
or U13139 (N_13139,N_12730,N_12650);
and U13140 (N_13140,N_12789,N_12633);
or U13141 (N_13141,N_12927,N_12781);
and U13142 (N_13142,N_12727,N_12818);
xor U13143 (N_13143,N_12655,N_12512);
and U13144 (N_13144,N_12634,N_12733);
xor U13145 (N_13145,N_12851,N_12718);
and U13146 (N_13146,N_12865,N_12524);
or U13147 (N_13147,N_12979,N_12546);
nor U13148 (N_13148,N_12503,N_12677);
or U13149 (N_13149,N_12652,N_12702);
nor U13150 (N_13150,N_12561,N_12885);
nor U13151 (N_13151,N_12532,N_12735);
or U13152 (N_13152,N_12919,N_12753);
nor U13153 (N_13153,N_12915,N_12968);
nor U13154 (N_13154,N_12775,N_12697);
and U13155 (N_13155,N_12833,N_12528);
or U13156 (N_13156,N_12817,N_12605);
and U13157 (N_13157,N_12619,N_12539);
nand U13158 (N_13158,N_12601,N_12502);
nand U13159 (N_13159,N_12827,N_12897);
nand U13160 (N_13160,N_12666,N_12982);
nor U13161 (N_13161,N_12926,N_12501);
and U13162 (N_13162,N_12668,N_12595);
and U13163 (N_13163,N_12646,N_12616);
and U13164 (N_13164,N_12903,N_12953);
and U13165 (N_13165,N_12934,N_12522);
nor U13166 (N_13166,N_12823,N_12779);
and U13167 (N_13167,N_12599,N_12876);
or U13168 (N_13168,N_12578,N_12606);
nor U13169 (N_13169,N_12681,N_12696);
nand U13170 (N_13170,N_12520,N_12651);
nand U13171 (N_13171,N_12981,N_12709);
or U13172 (N_13172,N_12553,N_12547);
nor U13173 (N_13173,N_12842,N_12533);
nor U13174 (N_13174,N_12831,N_12774);
and U13175 (N_13175,N_12877,N_12674);
and U13176 (N_13176,N_12506,N_12558);
nor U13177 (N_13177,N_12596,N_12725);
nand U13178 (N_13178,N_12716,N_12698);
nand U13179 (N_13179,N_12571,N_12967);
xor U13180 (N_13180,N_12869,N_12976);
and U13181 (N_13181,N_12871,N_12856);
and U13182 (N_13182,N_12505,N_12509);
and U13183 (N_13183,N_12962,N_12948);
or U13184 (N_13184,N_12600,N_12667);
nand U13185 (N_13185,N_12772,N_12530);
nor U13186 (N_13186,N_12863,N_12890);
or U13187 (N_13187,N_12990,N_12622);
and U13188 (N_13188,N_12945,N_12678);
nand U13189 (N_13189,N_12687,N_12529);
or U13190 (N_13190,N_12852,N_12672);
nand U13191 (N_13191,N_12907,N_12989);
xnor U13192 (N_13192,N_12808,N_12886);
nand U13193 (N_13193,N_12913,N_12584);
and U13194 (N_13194,N_12637,N_12799);
nor U13195 (N_13195,N_12810,N_12970);
nand U13196 (N_13196,N_12861,N_12891);
or U13197 (N_13197,N_12812,N_12556);
or U13198 (N_13198,N_12803,N_12814);
and U13199 (N_13199,N_12647,N_12640);
or U13200 (N_13200,N_12706,N_12875);
nand U13201 (N_13201,N_12593,N_12745);
nand U13202 (N_13202,N_12974,N_12755);
or U13203 (N_13203,N_12836,N_12660);
or U13204 (N_13204,N_12743,N_12720);
or U13205 (N_13205,N_12888,N_12878);
xor U13206 (N_13206,N_12625,N_12569);
nand U13207 (N_13207,N_12898,N_12872);
and U13208 (N_13208,N_12713,N_12999);
and U13209 (N_13209,N_12786,N_12849);
and U13210 (N_13210,N_12835,N_12950);
and U13211 (N_13211,N_12654,N_12670);
nor U13212 (N_13212,N_12819,N_12689);
xor U13213 (N_13213,N_12589,N_12917);
nor U13214 (N_13214,N_12910,N_12749);
nand U13215 (N_13215,N_12840,N_12693);
and U13216 (N_13216,N_12985,N_12751);
and U13217 (N_13217,N_12685,N_12978);
or U13218 (N_13218,N_12659,N_12661);
or U13219 (N_13219,N_12549,N_12695);
nand U13220 (N_13220,N_12776,N_12726);
nor U13221 (N_13221,N_12925,N_12904);
nand U13222 (N_13222,N_12691,N_12938);
nand U13223 (N_13223,N_12508,N_12995);
nor U13224 (N_13224,N_12641,N_12760);
nand U13225 (N_13225,N_12682,N_12719);
and U13226 (N_13226,N_12754,N_12954);
and U13227 (N_13227,N_12821,N_12777);
xnor U13228 (N_13228,N_12756,N_12829);
nor U13229 (N_13229,N_12994,N_12783);
and U13230 (N_13230,N_12822,N_12623);
nand U13231 (N_13231,N_12734,N_12700);
nor U13232 (N_13232,N_12966,N_12597);
or U13233 (N_13233,N_12929,N_12841);
or U13234 (N_13234,N_12801,N_12574);
nand U13235 (N_13235,N_12513,N_12629);
and U13236 (N_13236,N_12557,N_12880);
and U13237 (N_13237,N_12778,N_12658);
nand U13238 (N_13238,N_12805,N_12923);
or U13239 (N_13239,N_12627,N_12717);
nor U13240 (N_13240,N_12545,N_12531);
and U13241 (N_13241,N_12750,N_12736);
or U13242 (N_13242,N_12820,N_12694);
or U13243 (N_13243,N_12587,N_12816);
nand U13244 (N_13244,N_12752,N_12773);
or U13245 (N_13245,N_12983,N_12504);
xnor U13246 (N_13246,N_12586,N_12870);
and U13247 (N_13247,N_12867,N_12935);
and U13248 (N_13248,N_12680,N_12873);
nor U13249 (N_13249,N_12986,N_12582);
nand U13250 (N_13250,N_12714,N_12665);
nor U13251 (N_13251,N_12857,N_12797);
or U13252 (N_13252,N_12857,N_12663);
nand U13253 (N_13253,N_12688,N_12954);
xor U13254 (N_13254,N_12803,N_12831);
nor U13255 (N_13255,N_12955,N_12708);
xnor U13256 (N_13256,N_12891,N_12851);
nand U13257 (N_13257,N_12669,N_12583);
and U13258 (N_13258,N_12693,N_12968);
nor U13259 (N_13259,N_12558,N_12764);
nand U13260 (N_13260,N_12998,N_12704);
xor U13261 (N_13261,N_12775,N_12901);
nand U13262 (N_13262,N_12501,N_12566);
or U13263 (N_13263,N_12659,N_12834);
nor U13264 (N_13264,N_12597,N_12665);
xor U13265 (N_13265,N_12839,N_12980);
or U13266 (N_13266,N_12745,N_12684);
xnor U13267 (N_13267,N_12654,N_12767);
nor U13268 (N_13268,N_12630,N_12827);
xnor U13269 (N_13269,N_12683,N_12921);
and U13270 (N_13270,N_12804,N_12833);
nand U13271 (N_13271,N_12505,N_12769);
xnor U13272 (N_13272,N_12874,N_12697);
nand U13273 (N_13273,N_12922,N_12728);
xor U13274 (N_13274,N_12833,N_12934);
xor U13275 (N_13275,N_12857,N_12965);
nor U13276 (N_13276,N_12808,N_12813);
and U13277 (N_13277,N_12963,N_12506);
xnor U13278 (N_13278,N_12859,N_12586);
nor U13279 (N_13279,N_12737,N_12810);
xnor U13280 (N_13280,N_12603,N_12801);
and U13281 (N_13281,N_12924,N_12742);
or U13282 (N_13282,N_12748,N_12545);
nand U13283 (N_13283,N_12763,N_12670);
or U13284 (N_13284,N_12785,N_12689);
nand U13285 (N_13285,N_12842,N_12941);
nor U13286 (N_13286,N_12705,N_12557);
nor U13287 (N_13287,N_12851,N_12525);
and U13288 (N_13288,N_12704,N_12966);
and U13289 (N_13289,N_12532,N_12892);
and U13290 (N_13290,N_12722,N_12697);
xor U13291 (N_13291,N_12882,N_12532);
or U13292 (N_13292,N_12892,N_12730);
or U13293 (N_13293,N_12736,N_12868);
and U13294 (N_13294,N_12550,N_12646);
or U13295 (N_13295,N_12987,N_12890);
and U13296 (N_13296,N_12845,N_12719);
nor U13297 (N_13297,N_12884,N_12784);
nand U13298 (N_13298,N_12760,N_12897);
and U13299 (N_13299,N_12830,N_12542);
and U13300 (N_13300,N_12702,N_12538);
nor U13301 (N_13301,N_12701,N_12551);
nor U13302 (N_13302,N_12706,N_12625);
xor U13303 (N_13303,N_12693,N_12931);
nand U13304 (N_13304,N_12785,N_12692);
xor U13305 (N_13305,N_12666,N_12706);
nand U13306 (N_13306,N_12643,N_12733);
xnor U13307 (N_13307,N_12963,N_12509);
nand U13308 (N_13308,N_12510,N_12596);
or U13309 (N_13309,N_12592,N_12847);
and U13310 (N_13310,N_12820,N_12831);
or U13311 (N_13311,N_12615,N_12672);
and U13312 (N_13312,N_12607,N_12739);
nor U13313 (N_13313,N_12938,N_12886);
xor U13314 (N_13314,N_12609,N_12729);
nor U13315 (N_13315,N_12600,N_12534);
nor U13316 (N_13316,N_12720,N_12578);
xnor U13317 (N_13317,N_12539,N_12825);
and U13318 (N_13318,N_12673,N_12990);
nand U13319 (N_13319,N_12660,N_12799);
xor U13320 (N_13320,N_12732,N_12759);
nand U13321 (N_13321,N_12530,N_12705);
and U13322 (N_13322,N_12938,N_12824);
or U13323 (N_13323,N_12883,N_12634);
and U13324 (N_13324,N_12830,N_12549);
nor U13325 (N_13325,N_12514,N_12817);
nor U13326 (N_13326,N_12636,N_12974);
and U13327 (N_13327,N_12796,N_12831);
xor U13328 (N_13328,N_12688,N_12612);
xor U13329 (N_13329,N_12730,N_12809);
nand U13330 (N_13330,N_12534,N_12530);
xnor U13331 (N_13331,N_12810,N_12942);
xor U13332 (N_13332,N_12536,N_12814);
nor U13333 (N_13333,N_12519,N_12762);
nand U13334 (N_13334,N_12928,N_12817);
nor U13335 (N_13335,N_12721,N_12867);
xor U13336 (N_13336,N_12759,N_12601);
xnor U13337 (N_13337,N_12547,N_12639);
and U13338 (N_13338,N_12860,N_12572);
nand U13339 (N_13339,N_12840,N_12855);
and U13340 (N_13340,N_12659,N_12752);
nor U13341 (N_13341,N_12748,N_12527);
and U13342 (N_13342,N_12673,N_12857);
and U13343 (N_13343,N_12530,N_12891);
nor U13344 (N_13344,N_12742,N_12735);
and U13345 (N_13345,N_12993,N_12517);
and U13346 (N_13346,N_12835,N_12583);
nor U13347 (N_13347,N_12884,N_12809);
or U13348 (N_13348,N_12764,N_12819);
xnor U13349 (N_13349,N_12502,N_12870);
xnor U13350 (N_13350,N_12951,N_12589);
and U13351 (N_13351,N_12544,N_12554);
and U13352 (N_13352,N_12742,N_12529);
and U13353 (N_13353,N_12670,N_12734);
or U13354 (N_13354,N_12610,N_12546);
nand U13355 (N_13355,N_12862,N_12735);
xor U13356 (N_13356,N_12830,N_12702);
and U13357 (N_13357,N_12734,N_12577);
nor U13358 (N_13358,N_12660,N_12781);
nor U13359 (N_13359,N_12710,N_12803);
or U13360 (N_13360,N_12758,N_12910);
nand U13361 (N_13361,N_12729,N_12797);
nand U13362 (N_13362,N_12877,N_12892);
nand U13363 (N_13363,N_12968,N_12798);
and U13364 (N_13364,N_12690,N_12641);
nor U13365 (N_13365,N_12515,N_12616);
and U13366 (N_13366,N_12596,N_12899);
nand U13367 (N_13367,N_12507,N_12968);
xnor U13368 (N_13368,N_12998,N_12962);
and U13369 (N_13369,N_12657,N_12759);
nand U13370 (N_13370,N_12851,N_12886);
xor U13371 (N_13371,N_12668,N_12688);
and U13372 (N_13372,N_12787,N_12946);
and U13373 (N_13373,N_12507,N_12930);
or U13374 (N_13374,N_12656,N_12880);
and U13375 (N_13375,N_12773,N_12821);
or U13376 (N_13376,N_12759,N_12874);
xor U13377 (N_13377,N_12620,N_12723);
nor U13378 (N_13378,N_12780,N_12675);
nor U13379 (N_13379,N_12738,N_12823);
and U13380 (N_13380,N_12826,N_12738);
nand U13381 (N_13381,N_12623,N_12812);
nand U13382 (N_13382,N_12600,N_12531);
or U13383 (N_13383,N_12877,N_12799);
xnor U13384 (N_13384,N_12837,N_12757);
or U13385 (N_13385,N_12505,N_12516);
nand U13386 (N_13386,N_12834,N_12523);
nor U13387 (N_13387,N_12913,N_12981);
or U13388 (N_13388,N_12761,N_12907);
nand U13389 (N_13389,N_12621,N_12874);
and U13390 (N_13390,N_12997,N_12506);
xnor U13391 (N_13391,N_12587,N_12930);
nor U13392 (N_13392,N_12948,N_12505);
nand U13393 (N_13393,N_12840,N_12618);
nand U13394 (N_13394,N_12764,N_12538);
and U13395 (N_13395,N_12784,N_12805);
xor U13396 (N_13396,N_12899,N_12669);
xor U13397 (N_13397,N_12895,N_12973);
nand U13398 (N_13398,N_12841,N_12925);
nor U13399 (N_13399,N_12589,N_12665);
or U13400 (N_13400,N_12597,N_12611);
xnor U13401 (N_13401,N_12716,N_12558);
xor U13402 (N_13402,N_12786,N_12698);
or U13403 (N_13403,N_12544,N_12963);
or U13404 (N_13404,N_12818,N_12535);
or U13405 (N_13405,N_12817,N_12845);
nand U13406 (N_13406,N_12505,N_12641);
xor U13407 (N_13407,N_12628,N_12565);
nand U13408 (N_13408,N_12774,N_12819);
xnor U13409 (N_13409,N_12995,N_12676);
nand U13410 (N_13410,N_12735,N_12875);
nor U13411 (N_13411,N_12705,N_12583);
and U13412 (N_13412,N_12894,N_12832);
or U13413 (N_13413,N_12701,N_12757);
xnor U13414 (N_13414,N_12878,N_12543);
nor U13415 (N_13415,N_12636,N_12870);
nor U13416 (N_13416,N_12816,N_12595);
or U13417 (N_13417,N_12566,N_12954);
nor U13418 (N_13418,N_12603,N_12941);
xnor U13419 (N_13419,N_12676,N_12917);
xnor U13420 (N_13420,N_12843,N_12715);
nor U13421 (N_13421,N_12981,N_12751);
and U13422 (N_13422,N_12962,N_12684);
nor U13423 (N_13423,N_12746,N_12655);
nand U13424 (N_13424,N_12664,N_12588);
or U13425 (N_13425,N_12746,N_12896);
and U13426 (N_13426,N_12518,N_12610);
nor U13427 (N_13427,N_12823,N_12640);
nor U13428 (N_13428,N_12694,N_12552);
nor U13429 (N_13429,N_12608,N_12565);
nand U13430 (N_13430,N_12788,N_12809);
nor U13431 (N_13431,N_12558,N_12765);
nor U13432 (N_13432,N_12845,N_12635);
xor U13433 (N_13433,N_12910,N_12695);
nand U13434 (N_13434,N_12826,N_12952);
nor U13435 (N_13435,N_12737,N_12878);
xnor U13436 (N_13436,N_12766,N_12616);
or U13437 (N_13437,N_12759,N_12702);
or U13438 (N_13438,N_12889,N_12526);
or U13439 (N_13439,N_12518,N_12763);
xor U13440 (N_13440,N_12518,N_12873);
nand U13441 (N_13441,N_12732,N_12875);
and U13442 (N_13442,N_12866,N_12603);
nor U13443 (N_13443,N_12983,N_12671);
nand U13444 (N_13444,N_12928,N_12651);
and U13445 (N_13445,N_12590,N_12939);
or U13446 (N_13446,N_12648,N_12793);
and U13447 (N_13447,N_12837,N_12723);
or U13448 (N_13448,N_12883,N_12575);
xnor U13449 (N_13449,N_12659,N_12980);
nand U13450 (N_13450,N_12668,N_12697);
xor U13451 (N_13451,N_12987,N_12822);
nor U13452 (N_13452,N_12732,N_12776);
nor U13453 (N_13453,N_12849,N_12719);
nand U13454 (N_13454,N_12993,N_12624);
or U13455 (N_13455,N_12752,N_12785);
or U13456 (N_13456,N_12729,N_12997);
nand U13457 (N_13457,N_12896,N_12827);
or U13458 (N_13458,N_12552,N_12766);
and U13459 (N_13459,N_12966,N_12755);
xor U13460 (N_13460,N_12818,N_12815);
xor U13461 (N_13461,N_12502,N_12583);
nor U13462 (N_13462,N_12846,N_12601);
nor U13463 (N_13463,N_12824,N_12766);
nor U13464 (N_13464,N_12646,N_12845);
xnor U13465 (N_13465,N_12897,N_12562);
and U13466 (N_13466,N_12612,N_12797);
or U13467 (N_13467,N_12835,N_12847);
or U13468 (N_13468,N_12658,N_12545);
or U13469 (N_13469,N_12547,N_12842);
nand U13470 (N_13470,N_12735,N_12820);
xor U13471 (N_13471,N_12656,N_12943);
and U13472 (N_13472,N_12708,N_12664);
and U13473 (N_13473,N_12811,N_12835);
and U13474 (N_13474,N_12884,N_12980);
nand U13475 (N_13475,N_12661,N_12825);
xor U13476 (N_13476,N_12885,N_12534);
xnor U13477 (N_13477,N_12584,N_12780);
xor U13478 (N_13478,N_12994,N_12791);
or U13479 (N_13479,N_12523,N_12672);
nand U13480 (N_13480,N_12831,N_12861);
nand U13481 (N_13481,N_12860,N_12535);
or U13482 (N_13482,N_12947,N_12665);
xor U13483 (N_13483,N_12555,N_12889);
xnor U13484 (N_13484,N_12687,N_12599);
xnor U13485 (N_13485,N_12715,N_12834);
nand U13486 (N_13486,N_12890,N_12543);
and U13487 (N_13487,N_12881,N_12527);
xor U13488 (N_13488,N_12811,N_12944);
nor U13489 (N_13489,N_12906,N_12879);
nand U13490 (N_13490,N_12607,N_12731);
xnor U13491 (N_13491,N_12856,N_12814);
or U13492 (N_13492,N_12986,N_12797);
xnor U13493 (N_13493,N_12642,N_12553);
or U13494 (N_13494,N_12743,N_12601);
xnor U13495 (N_13495,N_12691,N_12670);
or U13496 (N_13496,N_12768,N_12817);
nand U13497 (N_13497,N_12509,N_12625);
or U13498 (N_13498,N_12544,N_12705);
or U13499 (N_13499,N_12970,N_12512);
and U13500 (N_13500,N_13163,N_13037);
nor U13501 (N_13501,N_13422,N_13354);
or U13502 (N_13502,N_13449,N_13020);
and U13503 (N_13503,N_13274,N_13092);
nand U13504 (N_13504,N_13397,N_13133);
nor U13505 (N_13505,N_13080,N_13122);
or U13506 (N_13506,N_13264,N_13138);
and U13507 (N_13507,N_13025,N_13479);
nand U13508 (N_13508,N_13343,N_13294);
nand U13509 (N_13509,N_13233,N_13091);
and U13510 (N_13510,N_13414,N_13398);
and U13511 (N_13511,N_13018,N_13200);
or U13512 (N_13512,N_13209,N_13167);
and U13513 (N_13513,N_13346,N_13110);
xnor U13514 (N_13514,N_13369,N_13436);
and U13515 (N_13515,N_13351,N_13260);
nand U13516 (N_13516,N_13427,N_13392);
or U13517 (N_13517,N_13229,N_13389);
and U13518 (N_13518,N_13453,N_13191);
or U13519 (N_13519,N_13432,N_13242);
xnor U13520 (N_13520,N_13281,N_13339);
nor U13521 (N_13521,N_13070,N_13411);
nand U13522 (N_13522,N_13442,N_13166);
xnor U13523 (N_13523,N_13055,N_13386);
xnor U13524 (N_13524,N_13207,N_13009);
xor U13525 (N_13525,N_13429,N_13017);
xor U13526 (N_13526,N_13399,N_13379);
nor U13527 (N_13527,N_13117,N_13413);
xor U13528 (N_13528,N_13099,N_13466);
xnor U13529 (N_13529,N_13243,N_13071);
xnor U13530 (N_13530,N_13363,N_13226);
nor U13531 (N_13531,N_13170,N_13309);
xnor U13532 (N_13532,N_13491,N_13296);
or U13533 (N_13533,N_13390,N_13285);
or U13534 (N_13534,N_13345,N_13056);
or U13535 (N_13535,N_13049,N_13140);
xor U13536 (N_13536,N_13341,N_13032);
and U13537 (N_13537,N_13401,N_13433);
nor U13538 (N_13538,N_13127,N_13324);
nand U13539 (N_13539,N_13195,N_13253);
xor U13540 (N_13540,N_13428,N_13284);
nor U13541 (N_13541,N_13086,N_13474);
nand U13542 (N_13542,N_13104,N_13150);
nor U13543 (N_13543,N_13035,N_13177);
or U13544 (N_13544,N_13330,N_13282);
nand U13545 (N_13545,N_13204,N_13277);
xor U13546 (N_13546,N_13265,N_13154);
xor U13547 (N_13547,N_13084,N_13459);
nand U13548 (N_13548,N_13162,N_13225);
nand U13549 (N_13549,N_13314,N_13470);
nor U13550 (N_13550,N_13161,N_13164);
nor U13551 (N_13551,N_13085,N_13289);
and U13552 (N_13552,N_13186,N_13477);
and U13553 (N_13553,N_13008,N_13248);
and U13554 (N_13554,N_13350,N_13121);
and U13555 (N_13555,N_13041,N_13423);
and U13556 (N_13556,N_13266,N_13258);
or U13557 (N_13557,N_13441,N_13238);
nor U13558 (N_13558,N_13268,N_13406);
nor U13559 (N_13559,N_13319,N_13338);
or U13560 (N_13560,N_13083,N_13439);
xnor U13561 (N_13561,N_13472,N_13081);
nor U13562 (N_13562,N_13391,N_13288);
and U13563 (N_13563,N_13444,N_13189);
nand U13564 (N_13564,N_13473,N_13030);
or U13565 (N_13565,N_13063,N_13303);
nand U13566 (N_13566,N_13403,N_13367);
or U13567 (N_13567,N_13155,N_13124);
xor U13568 (N_13568,N_13297,N_13492);
and U13569 (N_13569,N_13490,N_13058);
nand U13570 (N_13570,N_13327,N_13299);
nand U13571 (N_13571,N_13434,N_13342);
xor U13572 (N_13572,N_13286,N_13494);
xor U13573 (N_13573,N_13273,N_13072);
nor U13574 (N_13574,N_13039,N_13368);
xor U13575 (N_13575,N_13173,N_13489);
nor U13576 (N_13576,N_13196,N_13152);
and U13577 (N_13577,N_13005,N_13214);
and U13578 (N_13578,N_13144,N_13178);
nor U13579 (N_13579,N_13115,N_13456);
or U13580 (N_13580,N_13402,N_13145);
or U13581 (N_13581,N_13311,N_13486);
nand U13582 (N_13582,N_13348,N_13254);
or U13583 (N_13583,N_13159,N_13206);
xnor U13584 (N_13584,N_13371,N_13052);
nand U13585 (N_13585,N_13280,N_13272);
or U13586 (N_13586,N_13377,N_13374);
nor U13587 (N_13587,N_13292,N_13329);
nor U13588 (N_13588,N_13464,N_13216);
nand U13589 (N_13589,N_13151,N_13312);
nor U13590 (N_13590,N_13454,N_13135);
nor U13591 (N_13591,N_13300,N_13487);
nor U13592 (N_13592,N_13128,N_13340);
nand U13593 (N_13593,N_13384,N_13129);
nand U13594 (N_13594,N_13325,N_13385);
xnor U13595 (N_13595,N_13498,N_13111);
or U13596 (N_13596,N_13257,N_13307);
and U13597 (N_13597,N_13073,N_13180);
nor U13598 (N_13598,N_13499,N_13038);
xnor U13599 (N_13599,N_13010,N_13412);
nor U13600 (N_13600,N_13262,N_13451);
and U13601 (N_13601,N_13219,N_13148);
and U13602 (N_13602,N_13102,N_13076);
and U13603 (N_13603,N_13335,N_13431);
and U13604 (N_13604,N_13356,N_13157);
or U13605 (N_13605,N_13438,N_13149);
nor U13606 (N_13606,N_13134,N_13250);
nor U13607 (N_13607,N_13275,N_13347);
nand U13608 (N_13608,N_13448,N_13141);
nand U13609 (N_13609,N_13333,N_13482);
nor U13610 (N_13610,N_13131,N_13421);
and U13611 (N_13611,N_13187,N_13218);
nor U13612 (N_13612,N_13278,N_13417);
xor U13613 (N_13613,N_13308,N_13359);
or U13614 (N_13614,N_13158,N_13089);
and U13615 (N_13615,N_13425,N_13001);
nor U13616 (N_13616,N_13077,N_13251);
and U13617 (N_13617,N_13483,N_13101);
and U13618 (N_13618,N_13336,N_13269);
and U13619 (N_13619,N_13109,N_13301);
nand U13620 (N_13620,N_13156,N_13409);
nor U13621 (N_13621,N_13331,N_13042);
xor U13622 (N_13622,N_13011,N_13344);
nand U13623 (N_13623,N_13271,N_13291);
or U13624 (N_13624,N_13034,N_13227);
xor U13625 (N_13625,N_13059,N_13185);
and U13626 (N_13626,N_13194,N_13044);
nand U13627 (N_13627,N_13016,N_13255);
and U13628 (N_13628,N_13211,N_13305);
or U13629 (N_13629,N_13182,N_13310);
nor U13630 (N_13630,N_13212,N_13113);
xor U13631 (N_13631,N_13252,N_13365);
and U13632 (N_13632,N_13231,N_13051);
xor U13633 (N_13633,N_13290,N_13237);
and U13634 (N_13634,N_13328,N_13147);
and U13635 (N_13635,N_13287,N_13240);
nand U13636 (N_13636,N_13139,N_13107);
nand U13637 (N_13637,N_13267,N_13079);
xnor U13638 (N_13638,N_13452,N_13106);
and U13639 (N_13639,N_13097,N_13105);
or U13640 (N_13640,N_13137,N_13493);
xor U13641 (N_13641,N_13298,N_13192);
xnor U13642 (N_13642,N_13322,N_13024);
and U13643 (N_13643,N_13249,N_13234);
or U13644 (N_13644,N_13400,N_13090);
xor U13645 (N_13645,N_13019,N_13014);
xor U13646 (N_13646,N_13213,N_13088);
and U13647 (N_13647,N_13125,N_13096);
nor U13648 (N_13648,N_13373,N_13246);
and U13649 (N_13649,N_13376,N_13203);
or U13650 (N_13650,N_13380,N_13031);
or U13651 (N_13651,N_13228,N_13210);
and U13652 (N_13652,N_13029,N_13458);
and U13653 (N_13653,N_13215,N_13485);
nor U13654 (N_13654,N_13095,N_13455);
nor U13655 (N_13655,N_13112,N_13283);
xor U13656 (N_13656,N_13450,N_13198);
and U13657 (N_13657,N_13467,N_13496);
and U13658 (N_13658,N_13488,N_13244);
and U13659 (N_13659,N_13358,N_13108);
and U13660 (N_13660,N_13481,N_13146);
and U13661 (N_13661,N_13045,N_13181);
xnor U13662 (N_13662,N_13313,N_13028);
nand U13663 (N_13663,N_13318,N_13261);
and U13664 (N_13664,N_13387,N_13461);
and U13665 (N_13665,N_13171,N_13120);
or U13666 (N_13666,N_13160,N_13270);
and U13667 (N_13667,N_13174,N_13046);
nor U13668 (N_13668,N_13224,N_13381);
nand U13669 (N_13669,N_13446,N_13395);
xnor U13670 (N_13670,N_13142,N_13263);
xor U13671 (N_13671,N_13469,N_13202);
nor U13672 (N_13672,N_13420,N_13230);
or U13673 (N_13673,N_13362,N_13006);
or U13674 (N_13674,N_13418,N_13153);
or U13675 (N_13675,N_13419,N_13353);
xnor U13676 (N_13676,N_13114,N_13276);
and U13677 (N_13677,N_13320,N_13027);
nand U13678 (N_13678,N_13040,N_13245);
nor U13679 (N_13679,N_13256,N_13334);
nor U13680 (N_13680,N_13443,N_13116);
nand U13681 (N_13681,N_13007,N_13337);
nor U13682 (N_13682,N_13355,N_13021);
or U13683 (N_13683,N_13424,N_13103);
nor U13684 (N_13684,N_13364,N_13463);
nand U13685 (N_13685,N_13375,N_13003);
or U13686 (N_13686,N_13259,N_13415);
nor U13687 (N_13687,N_13193,N_13279);
nor U13688 (N_13688,N_13457,N_13349);
and U13689 (N_13689,N_13065,N_13220);
or U13690 (N_13690,N_13430,N_13462);
nand U13691 (N_13691,N_13062,N_13067);
nand U13692 (N_13692,N_13235,N_13304);
xnor U13693 (N_13693,N_13426,N_13082);
nand U13694 (N_13694,N_13208,N_13075);
nand U13695 (N_13695,N_13119,N_13013);
nand U13696 (N_13696,N_13495,N_13239);
nand U13697 (N_13697,N_13000,N_13370);
xnor U13698 (N_13698,N_13378,N_13136);
xnor U13699 (N_13699,N_13361,N_13471);
and U13700 (N_13700,N_13197,N_13435);
nand U13701 (N_13701,N_13100,N_13407);
nor U13702 (N_13702,N_13061,N_13047);
xor U13703 (N_13703,N_13326,N_13241);
xor U13704 (N_13704,N_13476,N_13315);
xor U13705 (N_13705,N_13168,N_13053);
xor U13706 (N_13706,N_13098,N_13004);
and U13707 (N_13707,N_13078,N_13440);
xnor U13708 (N_13708,N_13132,N_13060);
or U13709 (N_13709,N_13321,N_13205);
nor U13710 (N_13710,N_13184,N_13480);
or U13711 (N_13711,N_13468,N_13497);
xnor U13712 (N_13712,N_13360,N_13221);
and U13713 (N_13713,N_13015,N_13393);
xnor U13714 (N_13714,N_13317,N_13437);
and U13715 (N_13715,N_13460,N_13445);
xor U13716 (N_13716,N_13199,N_13465);
xnor U13717 (N_13717,N_13093,N_13183);
or U13718 (N_13718,N_13026,N_13416);
or U13719 (N_13719,N_13232,N_13316);
or U13720 (N_13720,N_13048,N_13201);
xnor U13721 (N_13721,N_13118,N_13366);
and U13722 (N_13722,N_13074,N_13169);
and U13723 (N_13723,N_13126,N_13372);
nand U13724 (N_13724,N_13302,N_13295);
or U13725 (N_13725,N_13293,N_13306);
xor U13726 (N_13726,N_13323,N_13057);
nand U13727 (N_13727,N_13188,N_13036);
nor U13728 (N_13728,N_13068,N_13002);
nor U13729 (N_13729,N_13222,N_13094);
and U13730 (N_13730,N_13130,N_13404);
or U13731 (N_13731,N_13179,N_13064);
xor U13732 (N_13732,N_13408,N_13357);
or U13733 (N_13733,N_13172,N_13066);
nor U13734 (N_13734,N_13475,N_13175);
and U13735 (N_13735,N_13352,N_13223);
xnor U13736 (N_13736,N_13087,N_13217);
nand U13737 (N_13737,N_13405,N_13388);
and U13738 (N_13738,N_13022,N_13054);
nand U13739 (N_13739,N_13332,N_13190);
nand U13740 (N_13740,N_13143,N_13484);
nor U13741 (N_13741,N_13236,N_13410);
or U13742 (N_13742,N_13247,N_13023);
nor U13743 (N_13743,N_13123,N_13050);
nand U13744 (N_13744,N_13012,N_13033);
and U13745 (N_13745,N_13165,N_13382);
xor U13746 (N_13746,N_13176,N_13396);
or U13747 (N_13747,N_13394,N_13447);
or U13748 (N_13748,N_13478,N_13043);
and U13749 (N_13749,N_13383,N_13069);
nor U13750 (N_13750,N_13099,N_13419);
xnor U13751 (N_13751,N_13242,N_13069);
or U13752 (N_13752,N_13076,N_13069);
nand U13753 (N_13753,N_13484,N_13420);
nor U13754 (N_13754,N_13188,N_13381);
and U13755 (N_13755,N_13398,N_13452);
or U13756 (N_13756,N_13385,N_13376);
nand U13757 (N_13757,N_13455,N_13468);
nor U13758 (N_13758,N_13280,N_13162);
xnor U13759 (N_13759,N_13019,N_13438);
nor U13760 (N_13760,N_13049,N_13399);
and U13761 (N_13761,N_13312,N_13053);
nand U13762 (N_13762,N_13369,N_13372);
nand U13763 (N_13763,N_13158,N_13017);
nand U13764 (N_13764,N_13430,N_13375);
nor U13765 (N_13765,N_13079,N_13158);
xnor U13766 (N_13766,N_13039,N_13366);
xor U13767 (N_13767,N_13173,N_13406);
nor U13768 (N_13768,N_13374,N_13076);
nor U13769 (N_13769,N_13075,N_13021);
nor U13770 (N_13770,N_13008,N_13375);
and U13771 (N_13771,N_13358,N_13472);
xnor U13772 (N_13772,N_13243,N_13034);
nand U13773 (N_13773,N_13188,N_13296);
or U13774 (N_13774,N_13035,N_13396);
or U13775 (N_13775,N_13270,N_13027);
xnor U13776 (N_13776,N_13304,N_13368);
xor U13777 (N_13777,N_13394,N_13063);
or U13778 (N_13778,N_13312,N_13143);
and U13779 (N_13779,N_13230,N_13011);
and U13780 (N_13780,N_13115,N_13325);
nand U13781 (N_13781,N_13310,N_13396);
nor U13782 (N_13782,N_13498,N_13339);
or U13783 (N_13783,N_13172,N_13334);
and U13784 (N_13784,N_13157,N_13067);
nor U13785 (N_13785,N_13008,N_13399);
nand U13786 (N_13786,N_13061,N_13311);
xor U13787 (N_13787,N_13473,N_13477);
nor U13788 (N_13788,N_13156,N_13163);
and U13789 (N_13789,N_13291,N_13330);
xor U13790 (N_13790,N_13053,N_13172);
nor U13791 (N_13791,N_13039,N_13127);
nand U13792 (N_13792,N_13286,N_13289);
and U13793 (N_13793,N_13208,N_13179);
or U13794 (N_13794,N_13235,N_13151);
and U13795 (N_13795,N_13071,N_13271);
nand U13796 (N_13796,N_13148,N_13315);
xnor U13797 (N_13797,N_13477,N_13454);
and U13798 (N_13798,N_13470,N_13108);
nor U13799 (N_13799,N_13421,N_13043);
nand U13800 (N_13800,N_13369,N_13286);
and U13801 (N_13801,N_13178,N_13391);
or U13802 (N_13802,N_13313,N_13090);
and U13803 (N_13803,N_13074,N_13128);
xor U13804 (N_13804,N_13470,N_13090);
and U13805 (N_13805,N_13467,N_13312);
or U13806 (N_13806,N_13385,N_13105);
and U13807 (N_13807,N_13225,N_13023);
and U13808 (N_13808,N_13004,N_13346);
nand U13809 (N_13809,N_13329,N_13039);
nand U13810 (N_13810,N_13210,N_13043);
xor U13811 (N_13811,N_13289,N_13047);
xnor U13812 (N_13812,N_13183,N_13185);
xnor U13813 (N_13813,N_13046,N_13185);
nor U13814 (N_13814,N_13182,N_13177);
or U13815 (N_13815,N_13005,N_13349);
xor U13816 (N_13816,N_13319,N_13107);
nor U13817 (N_13817,N_13178,N_13192);
xnor U13818 (N_13818,N_13210,N_13091);
or U13819 (N_13819,N_13355,N_13294);
nor U13820 (N_13820,N_13253,N_13272);
nand U13821 (N_13821,N_13161,N_13221);
nand U13822 (N_13822,N_13412,N_13308);
nand U13823 (N_13823,N_13439,N_13199);
xnor U13824 (N_13824,N_13216,N_13446);
nor U13825 (N_13825,N_13167,N_13052);
nor U13826 (N_13826,N_13394,N_13072);
nand U13827 (N_13827,N_13015,N_13358);
nor U13828 (N_13828,N_13412,N_13153);
or U13829 (N_13829,N_13316,N_13046);
nor U13830 (N_13830,N_13374,N_13322);
nor U13831 (N_13831,N_13256,N_13301);
nand U13832 (N_13832,N_13364,N_13353);
or U13833 (N_13833,N_13201,N_13197);
nor U13834 (N_13834,N_13434,N_13130);
xor U13835 (N_13835,N_13354,N_13220);
nand U13836 (N_13836,N_13196,N_13486);
xnor U13837 (N_13837,N_13106,N_13256);
nand U13838 (N_13838,N_13165,N_13483);
nor U13839 (N_13839,N_13412,N_13021);
xor U13840 (N_13840,N_13489,N_13346);
and U13841 (N_13841,N_13212,N_13174);
and U13842 (N_13842,N_13367,N_13226);
and U13843 (N_13843,N_13311,N_13437);
xor U13844 (N_13844,N_13260,N_13176);
nor U13845 (N_13845,N_13007,N_13229);
or U13846 (N_13846,N_13217,N_13037);
and U13847 (N_13847,N_13311,N_13216);
xor U13848 (N_13848,N_13399,N_13223);
or U13849 (N_13849,N_13246,N_13112);
nor U13850 (N_13850,N_13240,N_13108);
and U13851 (N_13851,N_13153,N_13057);
and U13852 (N_13852,N_13137,N_13420);
nand U13853 (N_13853,N_13456,N_13201);
xor U13854 (N_13854,N_13392,N_13447);
and U13855 (N_13855,N_13078,N_13262);
and U13856 (N_13856,N_13379,N_13273);
nor U13857 (N_13857,N_13439,N_13066);
nor U13858 (N_13858,N_13194,N_13205);
nor U13859 (N_13859,N_13365,N_13313);
xor U13860 (N_13860,N_13460,N_13326);
and U13861 (N_13861,N_13457,N_13419);
or U13862 (N_13862,N_13285,N_13116);
xor U13863 (N_13863,N_13377,N_13014);
nor U13864 (N_13864,N_13115,N_13224);
nand U13865 (N_13865,N_13231,N_13023);
nor U13866 (N_13866,N_13272,N_13357);
and U13867 (N_13867,N_13334,N_13045);
nor U13868 (N_13868,N_13093,N_13422);
or U13869 (N_13869,N_13453,N_13491);
or U13870 (N_13870,N_13108,N_13474);
or U13871 (N_13871,N_13153,N_13497);
xor U13872 (N_13872,N_13020,N_13229);
and U13873 (N_13873,N_13206,N_13285);
nor U13874 (N_13874,N_13053,N_13034);
or U13875 (N_13875,N_13146,N_13439);
nor U13876 (N_13876,N_13392,N_13487);
nand U13877 (N_13877,N_13248,N_13289);
nand U13878 (N_13878,N_13101,N_13264);
and U13879 (N_13879,N_13160,N_13394);
and U13880 (N_13880,N_13334,N_13290);
xor U13881 (N_13881,N_13256,N_13316);
nor U13882 (N_13882,N_13151,N_13307);
xor U13883 (N_13883,N_13051,N_13082);
or U13884 (N_13884,N_13230,N_13041);
or U13885 (N_13885,N_13030,N_13034);
nor U13886 (N_13886,N_13384,N_13418);
xnor U13887 (N_13887,N_13267,N_13207);
nor U13888 (N_13888,N_13399,N_13074);
or U13889 (N_13889,N_13347,N_13104);
or U13890 (N_13890,N_13402,N_13435);
xor U13891 (N_13891,N_13462,N_13144);
nor U13892 (N_13892,N_13027,N_13219);
nor U13893 (N_13893,N_13072,N_13341);
nand U13894 (N_13894,N_13042,N_13484);
or U13895 (N_13895,N_13416,N_13042);
xnor U13896 (N_13896,N_13493,N_13394);
or U13897 (N_13897,N_13325,N_13282);
nand U13898 (N_13898,N_13174,N_13445);
nor U13899 (N_13899,N_13105,N_13454);
and U13900 (N_13900,N_13150,N_13422);
nor U13901 (N_13901,N_13430,N_13030);
nor U13902 (N_13902,N_13479,N_13215);
and U13903 (N_13903,N_13140,N_13369);
xnor U13904 (N_13904,N_13311,N_13058);
or U13905 (N_13905,N_13175,N_13311);
nor U13906 (N_13906,N_13341,N_13141);
or U13907 (N_13907,N_13189,N_13332);
or U13908 (N_13908,N_13450,N_13026);
nand U13909 (N_13909,N_13431,N_13087);
and U13910 (N_13910,N_13480,N_13478);
xnor U13911 (N_13911,N_13408,N_13162);
nand U13912 (N_13912,N_13349,N_13047);
nor U13913 (N_13913,N_13056,N_13460);
xnor U13914 (N_13914,N_13256,N_13419);
and U13915 (N_13915,N_13274,N_13354);
xnor U13916 (N_13916,N_13016,N_13242);
or U13917 (N_13917,N_13396,N_13340);
xnor U13918 (N_13918,N_13194,N_13179);
nand U13919 (N_13919,N_13479,N_13254);
nor U13920 (N_13920,N_13265,N_13445);
or U13921 (N_13921,N_13360,N_13313);
nand U13922 (N_13922,N_13131,N_13309);
and U13923 (N_13923,N_13159,N_13103);
nand U13924 (N_13924,N_13273,N_13430);
and U13925 (N_13925,N_13038,N_13420);
and U13926 (N_13926,N_13385,N_13497);
xor U13927 (N_13927,N_13370,N_13183);
or U13928 (N_13928,N_13354,N_13008);
and U13929 (N_13929,N_13077,N_13192);
xnor U13930 (N_13930,N_13475,N_13213);
nor U13931 (N_13931,N_13271,N_13162);
nand U13932 (N_13932,N_13205,N_13493);
xor U13933 (N_13933,N_13129,N_13194);
and U13934 (N_13934,N_13230,N_13033);
nand U13935 (N_13935,N_13143,N_13439);
or U13936 (N_13936,N_13184,N_13157);
and U13937 (N_13937,N_13406,N_13434);
nand U13938 (N_13938,N_13450,N_13173);
or U13939 (N_13939,N_13350,N_13273);
nand U13940 (N_13940,N_13308,N_13283);
or U13941 (N_13941,N_13088,N_13419);
or U13942 (N_13942,N_13025,N_13132);
or U13943 (N_13943,N_13003,N_13179);
nor U13944 (N_13944,N_13463,N_13099);
or U13945 (N_13945,N_13128,N_13008);
and U13946 (N_13946,N_13192,N_13138);
or U13947 (N_13947,N_13477,N_13200);
and U13948 (N_13948,N_13261,N_13460);
or U13949 (N_13949,N_13152,N_13087);
nand U13950 (N_13950,N_13264,N_13031);
or U13951 (N_13951,N_13255,N_13474);
nor U13952 (N_13952,N_13319,N_13368);
nor U13953 (N_13953,N_13254,N_13225);
xor U13954 (N_13954,N_13491,N_13093);
or U13955 (N_13955,N_13377,N_13298);
or U13956 (N_13956,N_13392,N_13396);
nand U13957 (N_13957,N_13036,N_13437);
xnor U13958 (N_13958,N_13411,N_13219);
nor U13959 (N_13959,N_13459,N_13046);
nor U13960 (N_13960,N_13017,N_13376);
and U13961 (N_13961,N_13000,N_13086);
and U13962 (N_13962,N_13173,N_13281);
nand U13963 (N_13963,N_13055,N_13476);
xnor U13964 (N_13964,N_13416,N_13421);
and U13965 (N_13965,N_13228,N_13272);
xor U13966 (N_13966,N_13124,N_13255);
nor U13967 (N_13967,N_13281,N_13330);
and U13968 (N_13968,N_13047,N_13225);
nor U13969 (N_13969,N_13284,N_13367);
or U13970 (N_13970,N_13471,N_13051);
xor U13971 (N_13971,N_13374,N_13390);
xnor U13972 (N_13972,N_13340,N_13115);
or U13973 (N_13973,N_13115,N_13172);
and U13974 (N_13974,N_13146,N_13237);
or U13975 (N_13975,N_13111,N_13196);
xor U13976 (N_13976,N_13373,N_13370);
xnor U13977 (N_13977,N_13257,N_13450);
nand U13978 (N_13978,N_13166,N_13014);
xor U13979 (N_13979,N_13102,N_13449);
nand U13980 (N_13980,N_13415,N_13387);
nor U13981 (N_13981,N_13055,N_13224);
nand U13982 (N_13982,N_13364,N_13208);
xor U13983 (N_13983,N_13420,N_13029);
nor U13984 (N_13984,N_13137,N_13457);
xor U13985 (N_13985,N_13004,N_13189);
and U13986 (N_13986,N_13354,N_13342);
and U13987 (N_13987,N_13296,N_13408);
nand U13988 (N_13988,N_13056,N_13300);
nor U13989 (N_13989,N_13359,N_13234);
nor U13990 (N_13990,N_13245,N_13113);
or U13991 (N_13991,N_13024,N_13150);
nor U13992 (N_13992,N_13024,N_13253);
or U13993 (N_13993,N_13157,N_13064);
xor U13994 (N_13994,N_13405,N_13239);
and U13995 (N_13995,N_13174,N_13396);
and U13996 (N_13996,N_13442,N_13350);
or U13997 (N_13997,N_13428,N_13208);
nand U13998 (N_13998,N_13446,N_13333);
and U13999 (N_13999,N_13393,N_13014);
and U14000 (N_14000,N_13624,N_13652);
or U14001 (N_14001,N_13606,N_13585);
nor U14002 (N_14002,N_13572,N_13660);
nor U14003 (N_14003,N_13893,N_13868);
or U14004 (N_14004,N_13509,N_13937);
and U14005 (N_14005,N_13985,N_13871);
nand U14006 (N_14006,N_13850,N_13619);
xor U14007 (N_14007,N_13852,N_13865);
nor U14008 (N_14008,N_13936,N_13549);
xor U14009 (N_14009,N_13962,N_13755);
nand U14010 (N_14010,N_13862,N_13646);
xnor U14011 (N_14011,N_13861,N_13930);
nand U14012 (N_14012,N_13725,N_13820);
or U14013 (N_14013,N_13533,N_13704);
nor U14014 (N_14014,N_13955,N_13931);
or U14015 (N_14015,N_13537,N_13899);
or U14016 (N_14016,N_13544,N_13535);
nand U14017 (N_14017,N_13956,N_13680);
and U14018 (N_14018,N_13895,N_13654);
xor U14019 (N_14019,N_13612,N_13567);
and U14020 (N_14020,N_13942,N_13963);
and U14021 (N_14021,N_13501,N_13674);
or U14022 (N_14022,N_13757,N_13915);
nand U14023 (N_14023,N_13527,N_13576);
nand U14024 (N_14024,N_13629,N_13663);
or U14025 (N_14025,N_13966,N_13753);
or U14026 (N_14026,N_13591,N_13760);
and U14027 (N_14027,N_13977,N_13703);
nor U14028 (N_14028,N_13553,N_13696);
or U14029 (N_14029,N_13630,N_13858);
or U14030 (N_14030,N_13948,N_13690);
and U14031 (N_14031,N_13584,N_13994);
xnor U14032 (N_14032,N_13802,N_13919);
xnor U14033 (N_14033,N_13534,N_13961);
nand U14034 (N_14034,N_13598,N_13617);
xnor U14035 (N_14035,N_13970,N_13883);
nor U14036 (N_14036,N_13904,N_13661);
or U14037 (N_14037,N_13819,N_13752);
xnor U14038 (N_14038,N_13771,N_13679);
or U14039 (N_14039,N_13670,N_13989);
nand U14040 (N_14040,N_13859,N_13742);
nor U14041 (N_14041,N_13518,N_13816);
and U14042 (N_14042,N_13668,N_13712);
nand U14043 (N_14043,N_13664,N_13812);
nor U14044 (N_14044,N_13788,N_13596);
xor U14045 (N_14045,N_13982,N_13795);
or U14046 (N_14046,N_13647,N_13701);
nor U14047 (N_14047,N_13737,N_13929);
nor U14048 (N_14048,N_13933,N_13626);
or U14049 (N_14049,N_13876,N_13833);
nand U14050 (N_14050,N_13541,N_13902);
or U14051 (N_14051,N_13525,N_13620);
xnor U14052 (N_14052,N_13736,N_13848);
and U14053 (N_14053,N_13616,N_13558);
xnor U14054 (N_14054,N_13810,N_13784);
xor U14055 (N_14055,N_13841,N_13625);
nand U14056 (N_14056,N_13556,N_13896);
and U14057 (N_14057,N_13794,N_13838);
or U14058 (N_14058,N_13763,N_13972);
and U14059 (N_14059,N_13759,N_13706);
or U14060 (N_14060,N_13796,N_13554);
nand U14061 (N_14061,N_13638,N_13528);
xnor U14062 (N_14062,N_13540,N_13688);
or U14063 (N_14063,N_13952,N_13825);
nor U14064 (N_14064,N_13580,N_13722);
or U14065 (N_14065,N_13705,N_13949);
nand U14066 (N_14066,N_13906,N_13574);
xnor U14067 (N_14067,N_13921,N_13775);
nand U14068 (N_14068,N_13995,N_13849);
or U14069 (N_14069,N_13615,N_13939);
or U14070 (N_14070,N_13853,N_13557);
or U14071 (N_14071,N_13597,N_13740);
and U14072 (N_14072,N_13718,N_13887);
or U14073 (N_14073,N_13566,N_13683);
and U14074 (N_14074,N_13789,N_13761);
and U14075 (N_14075,N_13676,N_13953);
and U14076 (N_14076,N_13945,N_13542);
nor U14077 (N_14077,N_13691,N_13792);
xnor U14078 (N_14078,N_13925,N_13879);
and U14079 (N_14079,N_13854,N_13910);
xnor U14080 (N_14080,N_13685,N_13516);
nand U14081 (N_14081,N_13536,N_13637);
nand U14082 (N_14082,N_13918,N_13981);
and U14083 (N_14083,N_13514,N_13863);
nand U14084 (N_14084,N_13756,N_13746);
and U14085 (N_14085,N_13800,N_13716);
nand U14086 (N_14086,N_13739,N_13733);
or U14087 (N_14087,N_13748,N_13506);
nor U14088 (N_14088,N_13999,N_13967);
and U14089 (N_14089,N_13726,N_13634);
or U14090 (N_14090,N_13898,N_13824);
nand U14091 (N_14091,N_13560,N_13973);
and U14092 (N_14092,N_13988,N_13627);
xnor U14093 (N_14093,N_13545,N_13793);
nand U14094 (N_14094,N_13844,N_13837);
nor U14095 (N_14095,N_13564,N_13603);
and U14096 (N_14096,N_13957,N_13875);
or U14097 (N_14097,N_13747,N_13984);
nand U14098 (N_14098,N_13806,N_13522);
nand U14099 (N_14099,N_13734,N_13974);
nor U14100 (N_14100,N_13604,N_13743);
nand U14101 (N_14101,N_13526,N_13714);
and U14102 (N_14102,N_13878,N_13658);
nor U14103 (N_14103,N_13507,N_13531);
xnor U14104 (N_14104,N_13851,N_13735);
nor U14105 (N_14105,N_13571,N_13607);
and U14106 (N_14106,N_13959,N_13524);
nand U14107 (N_14107,N_13791,N_13642);
nor U14108 (N_14108,N_13965,N_13811);
nand U14109 (N_14109,N_13969,N_13872);
or U14110 (N_14110,N_13594,N_13723);
and U14111 (N_14111,N_13610,N_13618);
nand U14112 (N_14112,N_13890,N_13830);
xor U14113 (N_14113,N_13593,N_13997);
nand U14114 (N_14114,N_13640,N_13751);
nand U14115 (N_14115,N_13547,N_13821);
and U14116 (N_14116,N_13856,N_13870);
xor U14117 (N_14117,N_13836,N_13926);
and U14118 (N_14118,N_13903,N_13565);
and U14119 (N_14119,N_13947,N_13983);
or U14120 (N_14120,N_13608,N_13938);
and U14121 (N_14121,N_13835,N_13628);
and U14122 (N_14122,N_13840,N_13662);
xor U14123 (N_14123,N_13589,N_13729);
nand U14124 (N_14124,N_13614,N_13707);
xor U14125 (N_14125,N_13613,N_13503);
xnor U14126 (N_14126,N_13828,N_13934);
nor U14127 (N_14127,N_13991,N_13889);
nand U14128 (N_14128,N_13842,N_13866);
or U14129 (N_14129,N_13990,N_13781);
xnor U14130 (N_14130,N_13731,N_13546);
nand U14131 (N_14131,N_13592,N_13684);
and U14132 (N_14132,N_13880,N_13827);
and U14133 (N_14133,N_13745,N_13897);
nand U14134 (N_14134,N_13641,N_13960);
xnor U14135 (N_14135,N_13940,N_13801);
and U14136 (N_14136,N_13590,N_13874);
nand U14137 (N_14137,N_13699,N_13976);
nor U14138 (N_14138,N_13724,N_13667);
and U14139 (N_14139,N_13601,N_13980);
nand U14140 (N_14140,N_13754,N_13645);
xor U14141 (N_14141,N_13582,N_13877);
nand U14142 (N_14142,N_13678,N_13561);
nand U14143 (N_14143,N_13927,N_13978);
or U14144 (N_14144,N_13520,N_13888);
and U14145 (N_14145,N_13777,N_13909);
nor U14146 (N_14146,N_13932,N_13867);
and U14147 (N_14147,N_13529,N_13750);
xor U14148 (N_14148,N_13599,N_13687);
nand U14149 (N_14149,N_13798,N_13950);
xor U14150 (N_14150,N_13971,N_13884);
nor U14151 (N_14151,N_13666,N_13720);
and U14152 (N_14152,N_13728,N_13673);
or U14153 (N_14153,N_13523,N_13709);
xnor U14154 (N_14154,N_13782,N_13730);
or U14155 (N_14155,N_13935,N_13611);
nor U14156 (N_14156,N_13686,N_13986);
and U14157 (N_14157,N_13769,N_13916);
and U14158 (N_14158,N_13809,N_13573);
nor U14159 (N_14159,N_13650,N_13515);
nand U14160 (N_14160,N_13588,N_13779);
nor U14161 (N_14161,N_13539,N_13808);
xnor U14162 (N_14162,N_13787,N_13505);
nand U14163 (N_14163,N_13799,N_13968);
or U14164 (N_14164,N_13998,N_13656);
or U14165 (N_14165,N_13508,N_13568);
nor U14166 (N_14166,N_13681,N_13857);
xnor U14167 (N_14167,N_13846,N_13776);
or U14168 (N_14168,N_13822,N_13517);
nor U14169 (N_14169,N_13575,N_13738);
nand U14170 (N_14170,N_13892,N_13923);
and U14171 (N_14171,N_13710,N_13922);
xnor U14172 (N_14172,N_13804,N_13860);
nor U14173 (N_14173,N_13951,N_13913);
nand U14174 (N_14174,N_13829,N_13583);
or U14175 (N_14175,N_13511,N_13907);
nand U14176 (N_14176,N_13924,N_13803);
xor U14177 (N_14177,N_13548,N_13657);
nor U14178 (N_14178,N_13563,N_13964);
and U14179 (N_14179,N_13636,N_13832);
and U14180 (N_14180,N_13671,N_13774);
xnor U14181 (N_14181,N_13555,N_13943);
or U14182 (N_14182,N_13886,N_13677);
or U14183 (N_14183,N_13695,N_13894);
nor U14184 (N_14184,N_13831,N_13869);
or U14185 (N_14185,N_13719,N_13521);
or U14186 (N_14186,N_13783,N_13669);
and U14187 (N_14187,N_13928,N_13817);
xor U14188 (N_14188,N_13586,N_13651);
nand U14189 (N_14189,N_13911,N_13900);
or U14190 (N_14190,N_13749,N_13711);
nand U14191 (N_14191,N_13543,N_13510);
xor U14192 (N_14192,N_13605,N_13570);
nor U14193 (N_14193,N_13632,N_13655);
nand U14194 (N_14194,N_13653,N_13621);
nor U14195 (N_14195,N_13633,N_13768);
nor U14196 (N_14196,N_13659,N_13577);
or U14197 (N_14197,N_13917,N_13732);
nand U14198 (N_14198,N_13823,N_13559);
nand U14199 (N_14199,N_13532,N_13891);
xor U14200 (N_14200,N_13885,N_13905);
and U14201 (N_14201,N_13579,N_13694);
or U14202 (N_14202,N_13770,N_13500);
xor U14203 (N_14203,N_13538,N_13786);
nand U14204 (N_14204,N_13881,N_13715);
or U14205 (N_14205,N_13920,N_13958);
xnor U14206 (N_14206,N_13692,N_13530);
xnor U14207 (N_14207,N_13847,N_13697);
xnor U14208 (N_14208,N_13502,N_13993);
and U14209 (N_14209,N_13578,N_13839);
nor U14210 (N_14210,N_13675,N_13648);
nand U14211 (N_14211,N_13773,N_13805);
and U14212 (N_14212,N_13550,N_13721);
nand U14213 (N_14213,N_13941,N_13569);
nand U14214 (N_14214,N_13702,N_13882);
nor U14215 (N_14215,N_13504,N_13855);
and U14216 (N_14216,N_13797,N_13826);
or U14217 (N_14217,N_13587,N_13519);
nor U14218 (N_14218,N_13987,N_13708);
nor U14219 (N_14219,N_13562,N_13672);
nand U14220 (N_14220,N_13912,N_13551);
and U14221 (N_14221,N_13996,N_13764);
nor U14222 (N_14222,N_13766,N_13744);
nand U14223 (N_14223,N_13944,N_13992);
nand U14224 (N_14224,N_13873,N_13644);
or U14225 (N_14225,N_13649,N_13780);
nor U14226 (N_14226,N_13693,N_13689);
nand U14227 (N_14227,N_13581,N_13914);
xnor U14228 (N_14228,N_13700,N_13772);
nand U14229 (N_14229,N_13814,N_13845);
nand U14230 (N_14230,N_13595,N_13758);
nor U14231 (N_14231,N_13864,N_13682);
nor U14232 (N_14232,N_13767,N_13609);
and U14233 (N_14233,N_13979,N_13815);
or U14234 (N_14234,N_13946,N_13818);
nand U14235 (N_14235,N_13790,N_13622);
nor U14236 (N_14236,N_13954,N_13713);
nand U14237 (N_14237,N_13512,N_13623);
or U14238 (N_14238,N_13765,N_13785);
nand U14239 (N_14239,N_13727,N_13834);
and U14240 (N_14240,N_13602,N_13813);
and U14241 (N_14241,N_13635,N_13600);
and U14242 (N_14242,N_13665,N_13643);
nand U14243 (N_14243,N_13741,N_13698);
and U14244 (N_14244,N_13908,N_13762);
xor U14245 (N_14245,N_13552,N_13778);
nand U14246 (N_14246,N_13975,N_13631);
xnor U14247 (N_14247,N_13717,N_13901);
and U14248 (N_14248,N_13513,N_13843);
or U14249 (N_14249,N_13807,N_13639);
xor U14250 (N_14250,N_13989,N_13512);
or U14251 (N_14251,N_13933,N_13898);
xnor U14252 (N_14252,N_13629,N_13697);
xor U14253 (N_14253,N_13603,N_13834);
and U14254 (N_14254,N_13819,N_13672);
xnor U14255 (N_14255,N_13807,N_13883);
nand U14256 (N_14256,N_13691,N_13658);
nand U14257 (N_14257,N_13670,N_13700);
xor U14258 (N_14258,N_13874,N_13580);
or U14259 (N_14259,N_13878,N_13972);
or U14260 (N_14260,N_13995,N_13809);
and U14261 (N_14261,N_13609,N_13928);
nand U14262 (N_14262,N_13797,N_13902);
xor U14263 (N_14263,N_13906,N_13603);
nand U14264 (N_14264,N_13843,N_13968);
or U14265 (N_14265,N_13902,N_13856);
and U14266 (N_14266,N_13680,N_13787);
xor U14267 (N_14267,N_13675,N_13933);
xor U14268 (N_14268,N_13625,N_13667);
xor U14269 (N_14269,N_13690,N_13874);
or U14270 (N_14270,N_13509,N_13768);
xnor U14271 (N_14271,N_13947,N_13618);
xnor U14272 (N_14272,N_13633,N_13994);
xor U14273 (N_14273,N_13907,N_13656);
xnor U14274 (N_14274,N_13867,N_13993);
and U14275 (N_14275,N_13925,N_13802);
nor U14276 (N_14276,N_13606,N_13993);
nor U14277 (N_14277,N_13914,N_13807);
and U14278 (N_14278,N_13942,N_13665);
nor U14279 (N_14279,N_13990,N_13776);
and U14280 (N_14280,N_13889,N_13656);
and U14281 (N_14281,N_13997,N_13901);
nand U14282 (N_14282,N_13996,N_13977);
or U14283 (N_14283,N_13770,N_13542);
and U14284 (N_14284,N_13585,N_13537);
and U14285 (N_14285,N_13774,N_13750);
and U14286 (N_14286,N_13683,N_13854);
or U14287 (N_14287,N_13509,N_13844);
nor U14288 (N_14288,N_13652,N_13746);
and U14289 (N_14289,N_13858,N_13635);
and U14290 (N_14290,N_13910,N_13973);
nand U14291 (N_14291,N_13902,N_13641);
and U14292 (N_14292,N_13715,N_13601);
and U14293 (N_14293,N_13974,N_13990);
nor U14294 (N_14294,N_13937,N_13912);
xor U14295 (N_14295,N_13708,N_13732);
nor U14296 (N_14296,N_13727,N_13686);
xor U14297 (N_14297,N_13991,N_13593);
xnor U14298 (N_14298,N_13536,N_13826);
or U14299 (N_14299,N_13949,N_13526);
or U14300 (N_14300,N_13811,N_13563);
nor U14301 (N_14301,N_13872,N_13541);
xor U14302 (N_14302,N_13544,N_13928);
or U14303 (N_14303,N_13515,N_13696);
nor U14304 (N_14304,N_13553,N_13515);
and U14305 (N_14305,N_13643,N_13742);
xor U14306 (N_14306,N_13847,N_13792);
and U14307 (N_14307,N_13978,N_13767);
or U14308 (N_14308,N_13782,N_13826);
nand U14309 (N_14309,N_13530,N_13959);
xor U14310 (N_14310,N_13807,N_13577);
xnor U14311 (N_14311,N_13871,N_13792);
xnor U14312 (N_14312,N_13951,N_13798);
xnor U14313 (N_14313,N_13570,N_13662);
nor U14314 (N_14314,N_13762,N_13796);
or U14315 (N_14315,N_13557,N_13759);
nand U14316 (N_14316,N_13800,N_13836);
or U14317 (N_14317,N_13911,N_13602);
nor U14318 (N_14318,N_13881,N_13876);
and U14319 (N_14319,N_13779,N_13772);
xnor U14320 (N_14320,N_13528,N_13584);
nor U14321 (N_14321,N_13574,N_13849);
nand U14322 (N_14322,N_13531,N_13942);
nand U14323 (N_14323,N_13575,N_13803);
nor U14324 (N_14324,N_13508,N_13799);
or U14325 (N_14325,N_13890,N_13775);
xnor U14326 (N_14326,N_13767,N_13993);
xnor U14327 (N_14327,N_13840,N_13791);
nand U14328 (N_14328,N_13734,N_13807);
and U14329 (N_14329,N_13968,N_13999);
xor U14330 (N_14330,N_13580,N_13764);
and U14331 (N_14331,N_13614,N_13866);
xnor U14332 (N_14332,N_13746,N_13837);
nor U14333 (N_14333,N_13916,N_13771);
nor U14334 (N_14334,N_13887,N_13557);
nor U14335 (N_14335,N_13643,N_13755);
nand U14336 (N_14336,N_13930,N_13638);
xor U14337 (N_14337,N_13560,N_13916);
nor U14338 (N_14338,N_13531,N_13555);
or U14339 (N_14339,N_13971,N_13824);
nor U14340 (N_14340,N_13796,N_13512);
xor U14341 (N_14341,N_13793,N_13869);
and U14342 (N_14342,N_13808,N_13605);
and U14343 (N_14343,N_13725,N_13571);
xnor U14344 (N_14344,N_13894,N_13910);
and U14345 (N_14345,N_13735,N_13848);
xnor U14346 (N_14346,N_13995,N_13763);
nor U14347 (N_14347,N_13828,N_13540);
xnor U14348 (N_14348,N_13940,N_13624);
xor U14349 (N_14349,N_13783,N_13693);
nor U14350 (N_14350,N_13953,N_13874);
and U14351 (N_14351,N_13874,N_13650);
and U14352 (N_14352,N_13614,N_13512);
or U14353 (N_14353,N_13839,N_13682);
nor U14354 (N_14354,N_13681,N_13916);
nand U14355 (N_14355,N_13838,N_13619);
or U14356 (N_14356,N_13788,N_13645);
nand U14357 (N_14357,N_13882,N_13885);
and U14358 (N_14358,N_13516,N_13773);
and U14359 (N_14359,N_13628,N_13825);
and U14360 (N_14360,N_13776,N_13900);
nand U14361 (N_14361,N_13743,N_13641);
and U14362 (N_14362,N_13723,N_13794);
and U14363 (N_14363,N_13856,N_13999);
or U14364 (N_14364,N_13670,N_13520);
nor U14365 (N_14365,N_13873,N_13850);
xor U14366 (N_14366,N_13550,N_13692);
and U14367 (N_14367,N_13970,N_13995);
xor U14368 (N_14368,N_13700,N_13672);
xor U14369 (N_14369,N_13945,N_13714);
nor U14370 (N_14370,N_13893,N_13517);
and U14371 (N_14371,N_13617,N_13522);
or U14372 (N_14372,N_13909,N_13908);
nor U14373 (N_14373,N_13984,N_13563);
nor U14374 (N_14374,N_13558,N_13659);
nor U14375 (N_14375,N_13805,N_13741);
xnor U14376 (N_14376,N_13689,N_13797);
and U14377 (N_14377,N_13535,N_13866);
xnor U14378 (N_14378,N_13623,N_13855);
or U14379 (N_14379,N_13894,N_13638);
and U14380 (N_14380,N_13539,N_13949);
nand U14381 (N_14381,N_13738,N_13820);
nor U14382 (N_14382,N_13823,N_13932);
xnor U14383 (N_14383,N_13637,N_13786);
nor U14384 (N_14384,N_13866,N_13918);
xnor U14385 (N_14385,N_13875,N_13915);
xnor U14386 (N_14386,N_13693,N_13793);
nor U14387 (N_14387,N_13586,N_13994);
or U14388 (N_14388,N_13996,N_13661);
or U14389 (N_14389,N_13763,N_13795);
nor U14390 (N_14390,N_13917,N_13797);
nor U14391 (N_14391,N_13552,N_13690);
xor U14392 (N_14392,N_13954,N_13958);
nor U14393 (N_14393,N_13912,N_13842);
nand U14394 (N_14394,N_13807,N_13895);
and U14395 (N_14395,N_13612,N_13546);
and U14396 (N_14396,N_13568,N_13768);
or U14397 (N_14397,N_13636,N_13741);
and U14398 (N_14398,N_13979,N_13915);
xor U14399 (N_14399,N_13586,N_13731);
nor U14400 (N_14400,N_13693,N_13696);
or U14401 (N_14401,N_13977,N_13816);
or U14402 (N_14402,N_13752,N_13774);
nand U14403 (N_14403,N_13848,N_13859);
nor U14404 (N_14404,N_13995,N_13775);
xor U14405 (N_14405,N_13934,N_13849);
and U14406 (N_14406,N_13581,N_13784);
nor U14407 (N_14407,N_13505,N_13669);
xnor U14408 (N_14408,N_13847,N_13859);
nand U14409 (N_14409,N_13965,N_13916);
or U14410 (N_14410,N_13795,N_13605);
nand U14411 (N_14411,N_13624,N_13873);
or U14412 (N_14412,N_13941,N_13896);
and U14413 (N_14413,N_13802,N_13932);
xor U14414 (N_14414,N_13836,N_13839);
nand U14415 (N_14415,N_13545,N_13695);
nor U14416 (N_14416,N_13719,N_13861);
xor U14417 (N_14417,N_13844,N_13798);
nor U14418 (N_14418,N_13593,N_13885);
xor U14419 (N_14419,N_13941,N_13762);
nand U14420 (N_14420,N_13605,N_13726);
xor U14421 (N_14421,N_13618,N_13507);
and U14422 (N_14422,N_13662,N_13890);
nor U14423 (N_14423,N_13600,N_13542);
nand U14424 (N_14424,N_13664,N_13882);
nand U14425 (N_14425,N_13612,N_13512);
or U14426 (N_14426,N_13615,N_13898);
xnor U14427 (N_14427,N_13813,N_13675);
xor U14428 (N_14428,N_13550,N_13708);
xnor U14429 (N_14429,N_13593,N_13825);
nor U14430 (N_14430,N_13850,N_13899);
xor U14431 (N_14431,N_13698,N_13621);
and U14432 (N_14432,N_13931,N_13816);
or U14433 (N_14433,N_13924,N_13731);
and U14434 (N_14434,N_13575,N_13840);
and U14435 (N_14435,N_13655,N_13961);
xnor U14436 (N_14436,N_13529,N_13813);
nor U14437 (N_14437,N_13587,N_13854);
nor U14438 (N_14438,N_13996,N_13738);
xnor U14439 (N_14439,N_13832,N_13831);
or U14440 (N_14440,N_13555,N_13506);
nand U14441 (N_14441,N_13926,N_13567);
and U14442 (N_14442,N_13668,N_13747);
nor U14443 (N_14443,N_13537,N_13540);
nor U14444 (N_14444,N_13862,N_13769);
nand U14445 (N_14445,N_13619,N_13538);
or U14446 (N_14446,N_13641,N_13739);
nand U14447 (N_14447,N_13570,N_13839);
or U14448 (N_14448,N_13605,N_13858);
xor U14449 (N_14449,N_13833,N_13956);
or U14450 (N_14450,N_13560,N_13700);
xnor U14451 (N_14451,N_13981,N_13572);
xnor U14452 (N_14452,N_13812,N_13800);
or U14453 (N_14453,N_13551,N_13910);
or U14454 (N_14454,N_13945,N_13961);
and U14455 (N_14455,N_13817,N_13655);
nor U14456 (N_14456,N_13777,N_13689);
nand U14457 (N_14457,N_13773,N_13975);
and U14458 (N_14458,N_13551,N_13945);
nand U14459 (N_14459,N_13797,N_13895);
or U14460 (N_14460,N_13678,N_13934);
xor U14461 (N_14461,N_13928,N_13992);
xnor U14462 (N_14462,N_13570,N_13845);
nor U14463 (N_14463,N_13673,N_13595);
xor U14464 (N_14464,N_13917,N_13957);
nor U14465 (N_14465,N_13502,N_13531);
nand U14466 (N_14466,N_13783,N_13532);
or U14467 (N_14467,N_13900,N_13952);
or U14468 (N_14468,N_13747,N_13679);
nand U14469 (N_14469,N_13904,N_13790);
xnor U14470 (N_14470,N_13746,N_13754);
xor U14471 (N_14471,N_13792,N_13828);
and U14472 (N_14472,N_13854,N_13759);
and U14473 (N_14473,N_13762,N_13855);
xnor U14474 (N_14474,N_13594,N_13737);
nor U14475 (N_14475,N_13931,N_13988);
nand U14476 (N_14476,N_13878,N_13765);
nand U14477 (N_14477,N_13934,N_13923);
and U14478 (N_14478,N_13969,N_13654);
xor U14479 (N_14479,N_13933,N_13614);
xnor U14480 (N_14480,N_13585,N_13995);
nor U14481 (N_14481,N_13725,N_13819);
or U14482 (N_14482,N_13554,N_13508);
and U14483 (N_14483,N_13537,N_13992);
xor U14484 (N_14484,N_13820,N_13846);
nor U14485 (N_14485,N_13966,N_13522);
and U14486 (N_14486,N_13757,N_13618);
and U14487 (N_14487,N_13679,N_13831);
nor U14488 (N_14488,N_13796,N_13582);
xnor U14489 (N_14489,N_13801,N_13631);
nand U14490 (N_14490,N_13655,N_13612);
or U14491 (N_14491,N_13711,N_13852);
and U14492 (N_14492,N_13697,N_13870);
or U14493 (N_14493,N_13973,N_13769);
nor U14494 (N_14494,N_13971,N_13641);
nand U14495 (N_14495,N_13973,N_13556);
xnor U14496 (N_14496,N_13591,N_13702);
and U14497 (N_14497,N_13910,N_13511);
nor U14498 (N_14498,N_13721,N_13545);
nor U14499 (N_14499,N_13605,N_13575);
or U14500 (N_14500,N_14380,N_14215);
or U14501 (N_14501,N_14173,N_14175);
nor U14502 (N_14502,N_14066,N_14230);
xnor U14503 (N_14503,N_14348,N_14299);
xor U14504 (N_14504,N_14490,N_14418);
nor U14505 (N_14505,N_14459,N_14160);
nand U14506 (N_14506,N_14400,N_14322);
or U14507 (N_14507,N_14461,N_14302);
nand U14508 (N_14508,N_14038,N_14036);
xnor U14509 (N_14509,N_14248,N_14324);
nor U14510 (N_14510,N_14070,N_14243);
nor U14511 (N_14511,N_14141,N_14057);
and U14512 (N_14512,N_14359,N_14352);
or U14513 (N_14513,N_14019,N_14148);
or U14514 (N_14514,N_14481,N_14071);
nand U14515 (N_14515,N_14210,N_14336);
and U14516 (N_14516,N_14128,N_14254);
and U14517 (N_14517,N_14225,N_14365);
nor U14518 (N_14518,N_14494,N_14267);
nand U14519 (N_14519,N_14216,N_14377);
nor U14520 (N_14520,N_14350,N_14011);
xnor U14521 (N_14521,N_14339,N_14269);
and U14522 (N_14522,N_14244,N_14462);
nand U14523 (N_14523,N_14039,N_14329);
nand U14524 (N_14524,N_14064,N_14439);
nor U14525 (N_14525,N_14040,N_14079);
or U14526 (N_14526,N_14407,N_14105);
nand U14527 (N_14527,N_14233,N_14386);
nand U14528 (N_14528,N_14090,N_14209);
or U14529 (N_14529,N_14488,N_14250);
nand U14530 (N_14530,N_14154,N_14255);
and U14531 (N_14531,N_14297,N_14177);
or U14532 (N_14532,N_14021,N_14126);
nor U14533 (N_14533,N_14346,N_14344);
nand U14534 (N_14534,N_14262,N_14261);
xor U14535 (N_14535,N_14013,N_14452);
xnor U14536 (N_14536,N_14437,N_14423);
nor U14537 (N_14537,N_14296,N_14338);
nor U14538 (N_14538,N_14319,N_14016);
and U14539 (N_14539,N_14412,N_14200);
or U14540 (N_14540,N_14004,N_14231);
xor U14541 (N_14541,N_14479,N_14457);
and U14542 (N_14542,N_14181,N_14398);
xnor U14543 (N_14543,N_14211,N_14272);
and U14544 (N_14544,N_14473,N_14333);
xor U14545 (N_14545,N_14076,N_14056);
nor U14546 (N_14546,N_14208,N_14421);
nand U14547 (N_14547,N_14206,N_14080);
xor U14548 (N_14548,N_14445,N_14157);
nor U14549 (N_14549,N_14030,N_14130);
nand U14550 (N_14550,N_14472,N_14174);
xnor U14551 (N_14551,N_14107,N_14395);
nand U14552 (N_14552,N_14031,N_14098);
or U14553 (N_14553,N_14046,N_14293);
and U14554 (N_14554,N_14438,N_14342);
nor U14555 (N_14555,N_14122,N_14301);
xor U14556 (N_14556,N_14493,N_14448);
and U14557 (N_14557,N_14314,N_14073);
nand U14558 (N_14558,N_14012,N_14178);
nor U14559 (N_14559,N_14035,N_14162);
and U14560 (N_14560,N_14043,N_14218);
or U14561 (N_14561,N_14403,N_14227);
nor U14562 (N_14562,N_14343,N_14155);
nor U14563 (N_14563,N_14393,N_14025);
nand U14564 (N_14564,N_14023,N_14307);
nor U14565 (N_14565,N_14042,N_14006);
and U14566 (N_14566,N_14404,N_14228);
or U14567 (N_14567,N_14381,N_14084);
and U14568 (N_14568,N_14075,N_14153);
xor U14569 (N_14569,N_14067,N_14356);
and U14570 (N_14570,N_14102,N_14383);
and U14571 (N_14571,N_14417,N_14292);
or U14572 (N_14572,N_14465,N_14024);
nand U14573 (N_14573,N_14477,N_14353);
nand U14574 (N_14574,N_14235,N_14089);
nand U14575 (N_14575,N_14442,N_14109);
xnor U14576 (N_14576,N_14468,N_14222);
or U14577 (N_14577,N_14409,N_14320);
or U14578 (N_14578,N_14497,N_14271);
nor U14579 (N_14579,N_14123,N_14176);
xnor U14580 (N_14580,N_14480,N_14309);
xor U14581 (N_14581,N_14447,N_14366);
nor U14582 (N_14582,N_14249,N_14265);
or U14583 (N_14583,N_14145,N_14256);
and U14584 (N_14584,N_14044,N_14303);
or U14585 (N_14585,N_14323,N_14091);
nand U14586 (N_14586,N_14185,N_14048);
or U14587 (N_14587,N_14416,N_14001);
and U14588 (N_14588,N_14422,N_14028);
or U14589 (N_14589,N_14427,N_14099);
and U14590 (N_14590,N_14266,N_14186);
or U14591 (N_14591,N_14298,N_14087);
nand U14592 (N_14592,N_14092,N_14486);
nand U14593 (N_14593,N_14425,N_14283);
nand U14594 (N_14594,N_14399,N_14220);
xor U14595 (N_14595,N_14197,N_14325);
or U14596 (N_14596,N_14003,N_14041);
and U14597 (N_14597,N_14276,N_14411);
xor U14598 (N_14598,N_14124,N_14111);
nand U14599 (N_14599,N_14007,N_14410);
nand U14600 (N_14600,N_14062,N_14183);
and U14601 (N_14601,N_14096,N_14385);
and U14602 (N_14602,N_14444,N_14384);
nand U14603 (N_14603,N_14168,N_14161);
nand U14604 (N_14604,N_14115,N_14285);
nor U14605 (N_14605,N_14419,N_14002);
xnor U14606 (N_14606,N_14078,N_14396);
xor U14607 (N_14607,N_14121,N_14167);
xor U14608 (N_14608,N_14432,N_14193);
or U14609 (N_14609,N_14495,N_14300);
nor U14610 (N_14610,N_14351,N_14433);
nor U14611 (N_14611,N_14387,N_14037);
nand U14612 (N_14612,N_14072,N_14327);
or U14613 (N_14613,N_14143,N_14058);
and U14614 (N_14614,N_14182,N_14401);
and U14615 (N_14615,N_14047,N_14489);
and U14616 (N_14616,N_14196,N_14483);
or U14617 (N_14617,N_14334,N_14018);
and U14618 (N_14618,N_14372,N_14033);
nand U14619 (N_14619,N_14189,N_14147);
or U14620 (N_14620,N_14221,N_14010);
nor U14621 (N_14621,N_14190,N_14132);
or U14622 (N_14622,N_14471,N_14219);
nor U14623 (N_14623,N_14129,N_14052);
nand U14624 (N_14624,N_14156,N_14260);
and U14625 (N_14625,N_14277,N_14166);
or U14626 (N_14626,N_14382,N_14053);
nor U14627 (N_14627,N_14014,N_14345);
or U14628 (N_14628,N_14469,N_14369);
nand U14629 (N_14629,N_14083,N_14405);
nand U14630 (N_14630,N_14466,N_14360);
nor U14631 (N_14631,N_14349,N_14212);
nor U14632 (N_14632,N_14094,N_14491);
or U14633 (N_14633,N_14317,N_14009);
xnor U14634 (N_14634,N_14424,N_14364);
or U14635 (N_14635,N_14097,N_14436);
nand U14636 (N_14636,N_14355,N_14451);
xor U14637 (N_14637,N_14258,N_14275);
xnor U14638 (N_14638,N_14114,N_14051);
and U14639 (N_14639,N_14159,N_14420);
and U14640 (N_14640,N_14478,N_14117);
xor U14641 (N_14641,N_14113,N_14119);
and U14642 (N_14642,N_14453,N_14237);
and U14643 (N_14643,N_14020,N_14441);
xnor U14644 (N_14644,N_14374,N_14120);
and U14645 (N_14645,N_14476,N_14279);
or U14646 (N_14646,N_14055,N_14188);
nand U14647 (N_14647,N_14032,N_14492);
xnor U14648 (N_14648,N_14165,N_14240);
xor U14649 (N_14649,N_14000,N_14245);
nand U14650 (N_14650,N_14485,N_14487);
xnor U14651 (N_14651,N_14288,N_14458);
nand U14652 (N_14652,N_14257,N_14252);
nand U14653 (N_14653,N_14214,N_14284);
nand U14654 (N_14654,N_14063,N_14286);
nor U14655 (N_14655,N_14357,N_14194);
nor U14656 (N_14656,N_14110,N_14069);
nand U14657 (N_14657,N_14263,N_14379);
and U14658 (N_14658,N_14140,N_14311);
or U14659 (N_14659,N_14443,N_14308);
nand U14660 (N_14660,N_14354,N_14224);
and U14661 (N_14661,N_14456,N_14137);
xor U14662 (N_14662,N_14242,N_14499);
nor U14663 (N_14663,N_14118,N_14205);
nor U14664 (N_14664,N_14367,N_14074);
and U14665 (N_14665,N_14144,N_14413);
nand U14666 (N_14666,N_14455,N_14498);
nor U14667 (N_14667,N_14316,N_14049);
xnor U14668 (N_14668,N_14335,N_14232);
or U14669 (N_14669,N_14142,N_14291);
or U14670 (N_14670,N_14136,N_14373);
nand U14671 (N_14671,N_14281,N_14135);
or U14672 (N_14672,N_14065,N_14392);
and U14673 (N_14673,N_14318,N_14388);
nand U14674 (N_14674,N_14199,N_14429);
and U14675 (N_14675,N_14127,N_14305);
nand U14676 (N_14676,N_14008,N_14125);
and U14677 (N_14677,N_14446,N_14259);
nand U14678 (N_14678,N_14247,N_14376);
and U14679 (N_14679,N_14101,N_14241);
nor U14680 (N_14680,N_14394,N_14022);
nand U14681 (N_14681,N_14431,N_14146);
xnor U14682 (N_14682,N_14226,N_14192);
nand U14683 (N_14683,N_14061,N_14278);
nor U14684 (N_14684,N_14287,N_14191);
or U14685 (N_14685,N_14005,N_14229);
or U14686 (N_14686,N_14017,N_14397);
nor U14687 (N_14687,N_14034,N_14198);
nand U14688 (N_14688,N_14246,N_14310);
nor U14689 (N_14689,N_14289,N_14015);
nand U14690 (N_14690,N_14313,N_14460);
and U14691 (N_14691,N_14415,N_14390);
nand U14692 (N_14692,N_14213,N_14149);
nand U14693 (N_14693,N_14068,N_14482);
nor U14694 (N_14694,N_14450,N_14361);
or U14695 (N_14695,N_14201,N_14054);
or U14696 (N_14696,N_14434,N_14368);
nand U14697 (N_14697,N_14104,N_14470);
nand U14698 (N_14698,N_14295,N_14163);
or U14699 (N_14699,N_14108,N_14321);
and U14700 (N_14700,N_14358,N_14026);
nand U14701 (N_14701,N_14179,N_14251);
and U14702 (N_14702,N_14294,N_14408);
xnor U14703 (N_14703,N_14151,N_14059);
and U14704 (N_14704,N_14467,N_14440);
nand U14705 (N_14705,N_14152,N_14328);
xnor U14706 (N_14706,N_14081,N_14204);
xnor U14707 (N_14707,N_14391,N_14375);
xor U14708 (N_14708,N_14133,N_14164);
nor U14709 (N_14709,N_14378,N_14150);
nor U14710 (N_14710,N_14370,N_14139);
xnor U14711 (N_14711,N_14171,N_14337);
or U14712 (N_14712,N_14077,N_14389);
and U14713 (N_14713,N_14304,N_14341);
and U14714 (N_14714,N_14238,N_14426);
or U14715 (N_14715,N_14475,N_14184);
nor U14716 (N_14716,N_14274,N_14406);
and U14717 (N_14717,N_14253,N_14496);
or U14718 (N_14718,N_14428,N_14312);
nor U14719 (N_14719,N_14331,N_14463);
nand U14720 (N_14720,N_14187,N_14280);
or U14721 (N_14721,N_14449,N_14095);
or U14722 (N_14722,N_14454,N_14169);
xnor U14723 (N_14723,N_14362,N_14172);
xor U14724 (N_14724,N_14106,N_14195);
nor U14725 (N_14725,N_14085,N_14093);
nand U14726 (N_14726,N_14134,N_14340);
and U14727 (N_14727,N_14131,N_14430);
nor U14728 (N_14728,N_14207,N_14158);
nand U14729 (N_14729,N_14203,N_14402);
or U14730 (N_14730,N_14264,N_14282);
or U14731 (N_14731,N_14180,N_14273);
and U14732 (N_14732,N_14268,N_14347);
and U14733 (N_14733,N_14112,N_14330);
nand U14734 (N_14734,N_14435,N_14027);
nor U14735 (N_14735,N_14103,N_14332);
nor U14736 (N_14736,N_14315,N_14088);
nor U14737 (N_14737,N_14138,N_14050);
nor U14738 (N_14738,N_14223,N_14086);
xnor U14739 (N_14739,N_14371,N_14474);
nand U14740 (N_14740,N_14100,N_14484);
and U14741 (N_14741,N_14239,N_14234);
or U14742 (N_14742,N_14236,N_14029);
and U14743 (N_14743,N_14464,N_14060);
nor U14744 (N_14744,N_14363,N_14217);
nand U14745 (N_14745,N_14045,N_14270);
or U14746 (N_14746,N_14326,N_14414);
nand U14747 (N_14747,N_14116,N_14202);
and U14748 (N_14748,N_14082,N_14290);
nor U14749 (N_14749,N_14306,N_14170);
nor U14750 (N_14750,N_14354,N_14434);
and U14751 (N_14751,N_14029,N_14483);
xnor U14752 (N_14752,N_14465,N_14325);
and U14753 (N_14753,N_14202,N_14392);
and U14754 (N_14754,N_14285,N_14294);
nor U14755 (N_14755,N_14403,N_14394);
or U14756 (N_14756,N_14259,N_14484);
nand U14757 (N_14757,N_14450,N_14064);
or U14758 (N_14758,N_14446,N_14421);
nand U14759 (N_14759,N_14378,N_14126);
or U14760 (N_14760,N_14306,N_14054);
xor U14761 (N_14761,N_14301,N_14103);
or U14762 (N_14762,N_14012,N_14016);
xor U14763 (N_14763,N_14167,N_14412);
nor U14764 (N_14764,N_14013,N_14227);
nand U14765 (N_14765,N_14024,N_14373);
xnor U14766 (N_14766,N_14286,N_14014);
and U14767 (N_14767,N_14264,N_14449);
and U14768 (N_14768,N_14060,N_14412);
nor U14769 (N_14769,N_14076,N_14148);
or U14770 (N_14770,N_14313,N_14065);
xnor U14771 (N_14771,N_14448,N_14142);
xor U14772 (N_14772,N_14433,N_14342);
and U14773 (N_14773,N_14459,N_14475);
xnor U14774 (N_14774,N_14390,N_14498);
nor U14775 (N_14775,N_14223,N_14374);
or U14776 (N_14776,N_14187,N_14201);
xor U14777 (N_14777,N_14344,N_14154);
xor U14778 (N_14778,N_14084,N_14235);
nand U14779 (N_14779,N_14224,N_14444);
or U14780 (N_14780,N_14433,N_14410);
xnor U14781 (N_14781,N_14214,N_14414);
nand U14782 (N_14782,N_14304,N_14027);
and U14783 (N_14783,N_14267,N_14235);
xor U14784 (N_14784,N_14128,N_14226);
nand U14785 (N_14785,N_14123,N_14244);
xnor U14786 (N_14786,N_14425,N_14250);
or U14787 (N_14787,N_14076,N_14354);
or U14788 (N_14788,N_14263,N_14371);
nand U14789 (N_14789,N_14081,N_14118);
and U14790 (N_14790,N_14456,N_14295);
nand U14791 (N_14791,N_14024,N_14495);
xor U14792 (N_14792,N_14082,N_14004);
and U14793 (N_14793,N_14300,N_14240);
or U14794 (N_14794,N_14427,N_14358);
or U14795 (N_14795,N_14093,N_14181);
and U14796 (N_14796,N_14283,N_14170);
nand U14797 (N_14797,N_14309,N_14292);
nand U14798 (N_14798,N_14288,N_14143);
nor U14799 (N_14799,N_14236,N_14456);
nor U14800 (N_14800,N_14439,N_14474);
nor U14801 (N_14801,N_14137,N_14242);
xnor U14802 (N_14802,N_14008,N_14061);
nand U14803 (N_14803,N_14404,N_14499);
nand U14804 (N_14804,N_14374,N_14391);
nand U14805 (N_14805,N_14231,N_14455);
nand U14806 (N_14806,N_14171,N_14258);
nand U14807 (N_14807,N_14186,N_14040);
or U14808 (N_14808,N_14386,N_14009);
nor U14809 (N_14809,N_14071,N_14078);
nand U14810 (N_14810,N_14388,N_14125);
or U14811 (N_14811,N_14133,N_14415);
or U14812 (N_14812,N_14124,N_14010);
and U14813 (N_14813,N_14440,N_14244);
nand U14814 (N_14814,N_14178,N_14030);
nor U14815 (N_14815,N_14324,N_14224);
xor U14816 (N_14816,N_14091,N_14489);
and U14817 (N_14817,N_14052,N_14094);
nand U14818 (N_14818,N_14174,N_14260);
xor U14819 (N_14819,N_14025,N_14340);
and U14820 (N_14820,N_14370,N_14068);
xor U14821 (N_14821,N_14124,N_14355);
or U14822 (N_14822,N_14469,N_14410);
nand U14823 (N_14823,N_14388,N_14099);
or U14824 (N_14824,N_14372,N_14464);
xnor U14825 (N_14825,N_14480,N_14030);
xor U14826 (N_14826,N_14403,N_14170);
or U14827 (N_14827,N_14294,N_14030);
xnor U14828 (N_14828,N_14273,N_14141);
xnor U14829 (N_14829,N_14466,N_14035);
nand U14830 (N_14830,N_14230,N_14086);
nand U14831 (N_14831,N_14195,N_14460);
and U14832 (N_14832,N_14386,N_14054);
nor U14833 (N_14833,N_14492,N_14215);
xor U14834 (N_14834,N_14479,N_14095);
nor U14835 (N_14835,N_14382,N_14492);
nand U14836 (N_14836,N_14254,N_14257);
or U14837 (N_14837,N_14393,N_14396);
xor U14838 (N_14838,N_14427,N_14320);
and U14839 (N_14839,N_14046,N_14106);
and U14840 (N_14840,N_14136,N_14320);
nand U14841 (N_14841,N_14057,N_14329);
and U14842 (N_14842,N_14168,N_14196);
or U14843 (N_14843,N_14076,N_14314);
nand U14844 (N_14844,N_14147,N_14045);
xor U14845 (N_14845,N_14149,N_14196);
and U14846 (N_14846,N_14293,N_14131);
nor U14847 (N_14847,N_14006,N_14365);
or U14848 (N_14848,N_14324,N_14067);
nor U14849 (N_14849,N_14170,N_14265);
and U14850 (N_14850,N_14042,N_14322);
nor U14851 (N_14851,N_14309,N_14422);
and U14852 (N_14852,N_14036,N_14474);
or U14853 (N_14853,N_14063,N_14270);
nor U14854 (N_14854,N_14343,N_14221);
or U14855 (N_14855,N_14172,N_14141);
nand U14856 (N_14856,N_14202,N_14180);
or U14857 (N_14857,N_14368,N_14218);
or U14858 (N_14858,N_14180,N_14135);
xor U14859 (N_14859,N_14396,N_14110);
nand U14860 (N_14860,N_14364,N_14199);
xnor U14861 (N_14861,N_14436,N_14001);
nor U14862 (N_14862,N_14468,N_14112);
nor U14863 (N_14863,N_14070,N_14220);
or U14864 (N_14864,N_14433,N_14354);
xor U14865 (N_14865,N_14282,N_14080);
nand U14866 (N_14866,N_14096,N_14072);
and U14867 (N_14867,N_14426,N_14359);
nor U14868 (N_14868,N_14403,N_14198);
nor U14869 (N_14869,N_14393,N_14294);
or U14870 (N_14870,N_14496,N_14301);
or U14871 (N_14871,N_14006,N_14086);
and U14872 (N_14872,N_14235,N_14049);
nand U14873 (N_14873,N_14367,N_14487);
nor U14874 (N_14874,N_14286,N_14061);
nand U14875 (N_14875,N_14446,N_14295);
or U14876 (N_14876,N_14157,N_14384);
nand U14877 (N_14877,N_14210,N_14264);
or U14878 (N_14878,N_14284,N_14167);
and U14879 (N_14879,N_14173,N_14069);
nand U14880 (N_14880,N_14184,N_14285);
xnor U14881 (N_14881,N_14413,N_14054);
nor U14882 (N_14882,N_14219,N_14491);
xor U14883 (N_14883,N_14071,N_14161);
nand U14884 (N_14884,N_14478,N_14267);
nand U14885 (N_14885,N_14174,N_14359);
and U14886 (N_14886,N_14325,N_14255);
nand U14887 (N_14887,N_14278,N_14035);
or U14888 (N_14888,N_14268,N_14246);
or U14889 (N_14889,N_14297,N_14250);
nand U14890 (N_14890,N_14043,N_14301);
nor U14891 (N_14891,N_14410,N_14328);
and U14892 (N_14892,N_14472,N_14059);
or U14893 (N_14893,N_14277,N_14276);
xor U14894 (N_14894,N_14113,N_14314);
nor U14895 (N_14895,N_14136,N_14195);
and U14896 (N_14896,N_14431,N_14129);
xor U14897 (N_14897,N_14137,N_14437);
nor U14898 (N_14898,N_14276,N_14347);
nor U14899 (N_14899,N_14011,N_14043);
and U14900 (N_14900,N_14164,N_14467);
nor U14901 (N_14901,N_14161,N_14460);
xor U14902 (N_14902,N_14211,N_14171);
and U14903 (N_14903,N_14316,N_14319);
or U14904 (N_14904,N_14089,N_14083);
or U14905 (N_14905,N_14454,N_14138);
xnor U14906 (N_14906,N_14389,N_14360);
nor U14907 (N_14907,N_14027,N_14162);
or U14908 (N_14908,N_14467,N_14348);
or U14909 (N_14909,N_14033,N_14237);
or U14910 (N_14910,N_14428,N_14485);
nand U14911 (N_14911,N_14247,N_14454);
xor U14912 (N_14912,N_14108,N_14284);
xnor U14913 (N_14913,N_14169,N_14070);
nor U14914 (N_14914,N_14186,N_14417);
or U14915 (N_14915,N_14295,N_14313);
nor U14916 (N_14916,N_14467,N_14400);
xnor U14917 (N_14917,N_14283,N_14345);
nor U14918 (N_14918,N_14005,N_14398);
nor U14919 (N_14919,N_14025,N_14082);
or U14920 (N_14920,N_14460,N_14399);
or U14921 (N_14921,N_14221,N_14044);
or U14922 (N_14922,N_14342,N_14309);
nand U14923 (N_14923,N_14001,N_14134);
xnor U14924 (N_14924,N_14378,N_14028);
and U14925 (N_14925,N_14001,N_14322);
nor U14926 (N_14926,N_14060,N_14313);
xor U14927 (N_14927,N_14310,N_14011);
nand U14928 (N_14928,N_14448,N_14365);
xnor U14929 (N_14929,N_14409,N_14315);
or U14930 (N_14930,N_14381,N_14377);
or U14931 (N_14931,N_14088,N_14247);
and U14932 (N_14932,N_14403,N_14477);
xor U14933 (N_14933,N_14467,N_14460);
nor U14934 (N_14934,N_14372,N_14121);
or U14935 (N_14935,N_14424,N_14459);
or U14936 (N_14936,N_14498,N_14185);
xnor U14937 (N_14937,N_14417,N_14195);
or U14938 (N_14938,N_14189,N_14308);
nor U14939 (N_14939,N_14081,N_14107);
and U14940 (N_14940,N_14023,N_14095);
nor U14941 (N_14941,N_14104,N_14431);
xor U14942 (N_14942,N_14349,N_14248);
nor U14943 (N_14943,N_14101,N_14486);
or U14944 (N_14944,N_14054,N_14495);
nor U14945 (N_14945,N_14341,N_14473);
nor U14946 (N_14946,N_14447,N_14040);
nor U14947 (N_14947,N_14400,N_14024);
and U14948 (N_14948,N_14006,N_14080);
and U14949 (N_14949,N_14178,N_14009);
nor U14950 (N_14950,N_14051,N_14095);
or U14951 (N_14951,N_14469,N_14196);
and U14952 (N_14952,N_14387,N_14420);
nand U14953 (N_14953,N_14240,N_14155);
nor U14954 (N_14954,N_14151,N_14459);
nand U14955 (N_14955,N_14417,N_14133);
or U14956 (N_14956,N_14302,N_14345);
nor U14957 (N_14957,N_14434,N_14090);
and U14958 (N_14958,N_14139,N_14241);
or U14959 (N_14959,N_14151,N_14231);
and U14960 (N_14960,N_14014,N_14185);
and U14961 (N_14961,N_14177,N_14424);
xor U14962 (N_14962,N_14458,N_14317);
or U14963 (N_14963,N_14442,N_14388);
nor U14964 (N_14964,N_14432,N_14135);
xnor U14965 (N_14965,N_14439,N_14138);
nand U14966 (N_14966,N_14098,N_14046);
and U14967 (N_14967,N_14213,N_14286);
nor U14968 (N_14968,N_14107,N_14054);
and U14969 (N_14969,N_14205,N_14366);
nand U14970 (N_14970,N_14290,N_14481);
or U14971 (N_14971,N_14398,N_14091);
or U14972 (N_14972,N_14108,N_14218);
nand U14973 (N_14973,N_14282,N_14442);
xor U14974 (N_14974,N_14109,N_14195);
and U14975 (N_14975,N_14475,N_14192);
nand U14976 (N_14976,N_14207,N_14150);
nand U14977 (N_14977,N_14416,N_14042);
and U14978 (N_14978,N_14334,N_14432);
and U14979 (N_14979,N_14279,N_14384);
and U14980 (N_14980,N_14041,N_14434);
nor U14981 (N_14981,N_14271,N_14010);
nand U14982 (N_14982,N_14470,N_14157);
and U14983 (N_14983,N_14408,N_14164);
and U14984 (N_14984,N_14063,N_14439);
nand U14985 (N_14985,N_14344,N_14231);
and U14986 (N_14986,N_14448,N_14246);
nand U14987 (N_14987,N_14030,N_14293);
xor U14988 (N_14988,N_14321,N_14164);
and U14989 (N_14989,N_14176,N_14478);
and U14990 (N_14990,N_14061,N_14313);
or U14991 (N_14991,N_14259,N_14377);
or U14992 (N_14992,N_14112,N_14378);
or U14993 (N_14993,N_14418,N_14268);
and U14994 (N_14994,N_14173,N_14337);
xor U14995 (N_14995,N_14327,N_14117);
or U14996 (N_14996,N_14289,N_14407);
and U14997 (N_14997,N_14238,N_14495);
xor U14998 (N_14998,N_14496,N_14361);
and U14999 (N_14999,N_14424,N_14169);
or U15000 (N_15000,N_14835,N_14833);
and U15001 (N_15001,N_14872,N_14944);
and U15002 (N_15002,N_14900,N_14714);
nor U15003 (N_15003,N_14999,N_14724);
xor U15004 (N_15004,N_14920,N_14549);
and U15005 (N_15005,N_14695,N_14687);
nor U15006 (N_15006,N_14726,N_14806);
or U15007 (N_15007,N_14918,N_14517);
or U15008 (N_15008,N_14827,N_14813);
xnor U15009 (N_15009,N_14527,N_14996);
xor U15010 (N_15010,N_14853,N_14817);
nand U15011 (N_15011,N_14621,N_14728);
nor U15012 (N_15012,N_14914,N_14722);
and U15013 (N_15013,N_14622,N_14600);
or U15014 (N_15014,N_14965,N_14635);
or U15015 (N_15015,N_14694,N_14896);
nor U15016 (N_15016,N_14620,N_14788);
xnor U15017 (N_15017,N_14673,N_14768);
or U15018 (N_15018,N_14608,N_14542);
nor U15019 (N_15019,N_14789,N_14780);
or U15020 (N_15020,N_14974,N_14670);
and U15021 (N_15021,N_14590,N_14886);
xor U15022 (N_15022,N_14528,N_14681);
and U15023 (N_15023,N_14822,N_14762);
xnor U15024 (N_15024,N_14760,N_14824);
nand U15025 (N_15025,N_14649,N_14689);
xnor U15026 (N_15026,N_14516,N_14972);
xnor U15027 (N_15027,N_14633,N_14943);
xnor U15028 (N_15028,N_14950,N_14981);
nor U15029 (N_15029,N_14998,N_14556);
or U15030 (N_15030,N_14660,N_14523);
nand U15031 (N_15031,N_14561,N_14630);
xor U15032 (N_15032,N_14849,N_14603);
or U15033 (N_15033,N_14522,N_14832);
xor U15034 (N_15034,N_14671,N_14910);
or U15035 (N_15035,N_14716,N_14645);
or U15036 (N_15036,N_14513,N_14637);
xnor U15037 (N_15037,N_14717,N_14536);
xnor U15038 (N_15038,N_14905,N_14646);
nor U15039 (N_15039,N_14616,N_14672);
and U15040 (N_15040,N_14607,N_14564);
nand U15041 (N_15041,N_14837,N_14774);
or U15042 (N_15042,N_14627,N_14570);
and U15043 (N_15043,N_14738,N_14957);
and U15044 (N_15044,N_14624,N_14569);
or U15045 (N_15045,N_14558,N_14766);
and U15046 (N_15046,N_14924,N_14895);
nor U15047 (N_15047,N_14879,N_14826);
nand U15048 (N_15048,N_14869,N_14692);
or U15049 (N_15049,N_14554,N_14892);
nand U15050 (N_15050,N_14840,N_14852);
xnor U15051 (N_15051,N_14656,N_14650);
nor U15052 (N_15052,N_14787,N_14880);
nand U15053 (N_15053,N_14655,N_14956);
nand U15054 (N_15054,N_14632,N_14858);
or U15055 (N_15055,N_14613,N_14563);
nor U15056 (N_15056,N_14700,N_14825);
xnor U15057 (N_15057,N_14805,N_14983);
and U15058 (N_15058,N_14654,N_14544);
and U15059 (N_15059,N_14578,N_14702);
and U15060 (N_15060,N_14891,N_14751);
xor U15061 (N_15061,N_14752,N_14504);
or U15062 (N_15062,N_14730,N_14529);
and U15063 (N_15063,N_14969,N_14609);
and U15064 (N_15064,N_14749,N_14555);
xor U15065 (N_15065,N_14588,N_14512);
or U15066 (N_15066,N_14741,N_14810);
and U15067 (N_15067,N_14693,N_14775);
and U15068 (N_15068,N_14506,N_14740);
nand U15069 (N_15069,N_14743,N_14507);
nor U15070 (N_15070,N_14934,N_14602);
nand U15071 (N_15071,N_14785,N_14798);
nor U15072 (N_15072,N_14873,N_14992);
nor U15073 (N_15073,N_14883,N_14975);
xor U15074 (N_15074,N_14511,N_14989);
nand U15075 (N_15075,N_14970,N_14574);
nand U15076 (N_15076,N_14868,N_14525);
xor U15077 (N_15077,N_14666,N_14505);
nand U15078 (N_15078,N_14669,N_14955);
or U15079 (N_15079,N_14939,N_14809);
xnor U15080 (N_15080,N_14850,N_14978);
xnor U15081 (N_15081,N_14538,N_14927);
or U15082 (N_15082,N_14721,N_14966);
nor U15083 (N_15083,N_14857,N_14946);
and U15084 (N_15084,N_14587,N_14941);
or U15085 (N_15085,N_14893,N_14778);
nor U15086 (N_15086,N_14958,N_14770);
xnor U15087 (N_15087,N_14677,N_14793);
nand U15088 (N_15088,N_14963,N_14744);
xnor U15089 (N_15089,N_14763,N_14848);
nand U15090 (N_15090,N_14931,N_14642);
xor U15091 (N_15091,N_14546,N_14930);
xor U15092 (N_15092,N_14500,N_14962);
or U15093 (N_15093,N_14980,N_14926);
or U15094 (N_15094,N_14901,N_14796);
or U15095 (N_15095,N_14617,N_14945);
xnor U15096 (N_15096,N_14729,N_14815);
or U15097 (N_15097,N_14836,N_14884);
or U15098 (N_15098,N_14921,N_14593);
or U15099 (N_15099,N_14594,N_14948);
or U15100 (N_15100,N_14923,N_14786);
nand U15101 (N_15101,N_14909,N_14604);
or U15102 (N_15102,N_14735,N_14577);
xor U15103 (N_15103,N_14863,N_14625);
or U15104 (N_15104,N_14605,N_14547);
nand U15105 (N_15105,N_14859,N_14818);
nand U15106 (N_15106,N_14843,N_14887);
nand U15107 (N_15107,N_14720,N_14995);
or U15108 (N_15108,N_14878,N_14732);
nor U15109 (N_15109,N_14531,N_14890);
and U15110 (N_15110,N_14885,N_14585);
xnor U15111 (N_15111,N_14932,N_14701);
or U15112 (N_15112,N_14964,N_14739);
nand U15113 (N_15113,N_14711,N_14782);
xor U15114 (N_15114,N_14682,N_14658);
and U15115 (N_15115,N_14678,N_14541);
and U15116 (N_15116,N_14845,N_14875);
and U15117 (N_15117,N_14844,N_14917);
nor U15118 (N_15118,N_14942,N_14715);
nor U15119 (N_15119,N_14560,N_14937);
xor U15120 (N_15120,N_14582,N_14537);
and U15121 (N_15121,N_14540,N_14949);
nor U15122 (N_15122,N_14792,N_14897);
and U15123 (N_15123,N_14773,N_14619);
or U15124 (N_15124,N_14710,N_14733);
and U15125 (N_15125,N_14987,N_14783);
xnor U15126 (N_15126,N_14794,N_14565);
and U15127 (N_15127,N_14982,N_14601);
nor U15128 (N_15128,N_14589,N_14902);
nor U15129 (N_15129,N_14644,N_14696);
and U15130 (N_15130,N_14799,N_14518);
nand U15131 (N_15131,N_14706,N_14748);
and U15132 (N_15132,N_14545,N_14971);
or U15133 (N_15133,N_14867,N_14906);
and U15134 (N_15134,N_14712,N_14647);
and U15135 (N_15135,N_14913,N_14960);
or U15136 (N_15136,N_14509,N_14882);
and U15137 (N_15137,N_14723,N_14680);
xnor U15138 (N_15138,N_14746,N_14626);
nand U15139 (N_15139,N_14911,N_14802);
nand U15140 (N_15140,N_14583,N_14769);
nand U15141 (N_15141,N_14688,N_14756);
or U15142 (N_15142,N_14708,N_14703);
nand U15143 (N_15143,N_14719,N_14781);
xor U15144 (N_15144,N_14907,N_14567);
or U15145 (N_15145,N_14874,N_14690);
or U15146 (N_15146,N_14862,N_14997);
xnor U15147 (N_15147,N_14916,N_14830);
or U15148 (N_15148,N_14562,N_14709);
or U15149 (N_15149,N_14606,N_14663);
nand U15150 (N_15150,N_14812,N_14572);
or U15151 (N_15151,N_14979,N_14953);
xnor U15152 (N_15152,N_14842,N_14936);
nand U15153 (N_15153,N_14676,N_14508);
or U15154 (N_15154,N_14591,N_14807);
nor U15155 (N_15155,N_14940,N_14668);
xor U15156 (N_15156,N_14838,N_14990);
nor U15157 (N_15157,N_14596,N_14977);
nand U15158 (N_15158,N_14653,N_14639);
and U15159 (N_15159,N_14571,N_14651);
nand U15160 (N_15160,N_14870,N_14860);
xor U15161 (N_15161,N_14871,N_14592);
nor U15162 (N_15162,N_14904,N_14614);
nand U15163 (N_15163,N_14664,N_14535);
or U15164 (N_15164,N_14820,N_14821);
xor U15165 (N_15165,N_14846,N_14823);
nor U15166 (N_15166,N_14779,N_14800);
nand U15167 (N_15167,N_14854,N_14698);
and U15168 (N_15168,N_14801,N_14772);
and U15169 (N_15169,N_14831,N_14611);
nand U15170 (N_15170,N_14803,N_14514);
and U15171 (N_15171,N_14991,N_14580);
or U15172 (N_15172,N_14864,N_14510);
nor U15173 (N_15173,N_14573,N_14954);
and U15174 (N_15174,N_14598,N_14643);
nor U15175 (N_15175,N_14713,N_14502);
and U15176 (N_15176,N_14759,N_14521);
and U15177 (N_15177,N_14684,N_14922);
and U15178 (N_15178,N_14898,N_14777);
xnor U15179 (N_15179,N_14731,N_14612);
nand U15180 (N_15180,N_14631,N_14697);
nor U15181 (N_15181,N_14959,N_14765);
and U15182 (N_15182,N_14819,N_14986);
nor U15183 (N_15183,N_14951,N_14734);
xnor U15184 (N_15184,N_14534,N_14586);
xnor U15185 (N_15185,N_14947,N_14599);
and U15186 (N_15186,N_14581,N_14938);
xnor U15187 (N_15187,N_14550,N_14553);
nor U15188 (N_15188,N_14638,N_14704);
and U15189 (N_15189,N_14595,N_14912);
xor U15190 (N_15190,N_14961,N_14705);
and U15191 (N_15191,N_14804,N_14686);
nand U15192 (N_15192,N_14736,N_14566);
xor U15193 (N_15193,N_14662,N_14984);
nor U15194 (N_15194,N_14520,N_14866);
or U15195 (N_15195,N_14640,N_14501);
and U15196 (N_15196,N_14829,N_14707);
xnor U15197 (N_15197,N_14699,N_14532);
xnor U15198 (N_15198,N_14648,N_14559);
nor U15199 (N_15199,N_14791,N_14808);
and U15200 (N_15200,N_14967,N_14742);
or U15201 (N_15201,N_14889,N_14679);
and U15202 (N_15202,N_14899,N_14816);
and U15203 (N_15203,N_14834,N_14641);
nand U15204 (N_15204,N_14908,N_14915);
nand U15205 (N_15205,N_14552,N_14524);
or U15206 (N_15206,N_14515,N_14888);
nand U15207 (N_15207,N_14925,N_14771);
and U15208 (N_15208,N_14755,N_14795);
nor U15209 (N_15209,N_14758,N_14615);
nand U15210 (N_15210,N_14952,N_14576);
nor U15211 (N_15211,N_14675,N_14753);
or U15212 (N_15212,N_14985,N_14894);
nor U15213 (N_15213,N_14661,N_14933);
xor U15214 (N_15214,N_14935,N_14551);
and U15215 (N_15215,N_14841,N_14628);
xnor U15216 (N_15216,N_14988,N_14727);
and U15217 (N_15217,N_14636,N_14623);
and U15218 (N_15218,N_14667,N_14747);
and U15219 (N_15219,N_14618,N_14764);
xnor U15220 (N_15220,N_14851,N_14584);
or U15221 (N_15221,N_14797,N_14776);
and U15222 (N_15222,N_14579,N_14847);
nand U15223 (N_15223,N_14790,N_14750);
nor U15224 (N_15224,N_14855,N_14993);
nor U15225 (N_15225,N_14754,N_14767);
nor U15226 (N_15226,N_14610,N_14530);
nand U15227 (N_15227,N_14533,N_14657);
xor U15228 (N_15228,N_14761,N_14548);
xnor U15229 (N_15229,N_14725,N_14568);
or U15230 (N_15230,N_14526,N_14674);
xnor U15231 (N_15231,N_14659,N_14503);
nor U15232 (N_15232,N_14814,N_14691);
and U15233 (N_15233,N_14877,N_14652);
or U15234 (N_15234,N_14811,N_14861);
xnor U15235 (N_15235,N_14539,N_14881);
xor U15236 (N_15236,N_14557,N_14784);
nor U15237 (N_15237,N_14634,N_14745);
and U15238 (N_15238,N_14839,N_14856);
nand U15239 (N_15239,N_14519,N_14543);
nor U15240 (N_15240,N_14629,N_14575);
nand U15241 (N_15241,N_14685,N_14976);
or U15242 (N_15242,N_14973,N_14718);
and U15243 (N_15243,N_14968,N_14828);
or U15244 (N_15244,N_14597,N_14903);
xnor U15245 (N_15245,N_14994,N_14665);
and U15246 (N_15246,N_14929,N_14919);
nor U15247 (N_15247,N_14683,N_14928);
xor U15248 (N_15248,N_14737,N_14757);
nand U15249 (N_15249,N_14865,N_14876);
nor U15250 (N_15250,N_14537,N_14801);
nor U15251 (N_15251,N_14944,N_14930);
or U15252 (N_15252,N_14744,N_14791);
nor U15253 (N_15253,N_14840,N_14804);
or U15254 (N_15254,N_14773,N_14607);
nand U15255 (N_15255,N_14881,N_14950);
nor U15256 (N_15256,N_14966,N_14913);
xnor U15257 (N_15257,N_14955,N_14597);
nand U15258 (N_15258,N_14886,N_14660);
xor U15259 (N_15259,N_14893,N_14971);
or U15260 (N_15260,N_14799,N_14501);
and U15261 (N_15261,N_14681,N_14605);
nand U15262 (N_15262,N_14796,N_14760);
nor U15263 (N_15263,N_14721,N_14946);
nor U15264 (N_15264,N_14977,N_14558);
or U15265 (N_15265,N_14652,N_14637);
nand U15266 (N_15266,N_14859,N_14973);
nand U15267 (N_15267,N_14742,N_14903);
or U15268 (N_15268,N_14590,N_14648);
nor U15269 (N_15269,N_14539,N_14818);
or U15270 (N_15270,N_14730,N_14777);
and U15271 (N_15271,N_14669,N_14883);
and U15272 (N_15272,N_14629,N_14985);
nand U15273 (N_15273,N_14737,N_14618);
and U15274 (N_15274,N_14522,N_14892);
or U15275 (N_15275,N_14885,N_14532);
and U15276 (N_15276,N_14792,N_14747);
nor U15277 (N_15277,N_14589,N_14988);
xor U15278 (N_15278,N_14741,N_14797);
or U15279 (N_15279,N_14637,N_14659);
nand U15280 (N_15280,N_14775,N_14860);
xnor U15281 (N_15281,N_14528,N_14970);
or U15282 (N_15282,N_14979,N_14616);
nor U15283 (N_15283,N_14511,N_14881);
nand U15284 (N_15284,N_14688,N_14964);
xnor U15285 (N_15285,N_14713,N_14575);
nand U15286 (N_15286,N_14771,N_14719);
xor U15287 (N_15287,N_14852,N_14681);
or U15288 (N_15288,N_14832,N_14797);
or U15289 (N_15289,N_14528,N_14851);
and U15290 (N_15290,N_14776,N_14846);
or U15291 (N_15291,N_14627,N_14972);
and U15292 (N_15292,N_14675,N_14870);
nor U15293 (N_15293,N_14509,N_14527);
xor U15294 (N_15294,N_14780,N_14801);
xnor U15295 (N_15295,N_14579,N_14777);
and U15296 (N_15296,N_14657,N_14945);
nand U15297 (N_15297,N_14770,N_14835);
xnor U15298 (N_15298,N_14964,N_14836);
or U15299 (N_15299,N_14614,N_14897);
and U15300 (N_15300,N_14638,N_14736);
or U15301 (N_15301,N_14571,N_14960);
nand U15302 (N_15302,N_14978,N_14502);
nand U15303 (N_15303,N_14523,N_14885);
or U15304 (N_15304,N_14536,N_14654);
and U15305 (N_15305,N_14923,N_14512);
xor U15306 (N_15306,N_14535,N_14611);
or U15307 (N_15307,N_14914,N_14897);
or U15308 (N_15308,N_14984,N_14837);
nor U15309 (N_15309,N_14963,N_14578);
and U15310 (N_15310,N_14655,N_14916);
xor U15311 (N_15311,N_14748,N_14989);
nor U15312 (N_15312,N_14971,N_14592);
or U15313 (N_15313,N_14902,N_14709);
nor U15314 (N_15314,N_14528,N_14558);
nor U15315 (N_15315,N_14915,N_14906);
xor U15316 (N_15316,N_14587,N_14740);
or U15317 (N_15317,N_14947,N_14785);
nor U15318 (N_15318,N_14866,N_14530);
nand U15319 (N_15319,N_14559,N_14700);
xor U15320 (N_15320,N_14515,N_14832);
or U15321 (N_15321,N_14800,N_14774);
and U15322 (N_15322,N_14832,N_14583);
nor U15323 (N_15323,N_14698,N_14869);
xnor U15324 (N_15324,N_14628,N_14591);
xnor U15325 (N_15325,N_14777,N_14836);
or U15326 (N_15326,N_14877,N_14794);
or U15327 (N_15327,N_14588,N_14850);
xnor U15328 (N_15328,N_14962,N_14804);
nor U15329 (N_15329,N_14669,N_14968);
nor U15330 (N_15330,N_14692,N_14693);
or U15331 (N_15331,N_14853,N_14504);
xnor U15332 (N_15332,N_14694,N_14577);
xnor U15333 (N_15333,N_14718,N_14993);
nand U15334 (N_15334,N_14879,N_14809);
and U15335 (N_15335,N_14909,N_14759);
xor U15336 (N_15336,N_14742,N_14815);
and U15337 (N_15337,N_14517,N_14728);
and U15338 (N_15338,N_14908,N_14964);
nor U15339 (N_15339,N_14545,N_14931);
and U15340 (N_15340,N_14943,N_14537);
nand U15341 (N_15341,N_14649,N_14997);
or U15342 (N_15342,N_14610,N_14902);
and U15343 (N_15343,N_14674,N_14819);
nand U15344 (N_15344,N_14800,N_14821);
and U15345 (N_15345,N_14974,N_14530);
nand U15346 (N_15346,N_14527,N_14736);
or U15347 (N_15347,N_14750,N_14896);
or U15348 (N_15348,N_14741,N_14565);
and U15349 (N_15349,N_14711,N_14847);
xnor U15350 (N_15350,N_14897,N_14965);
or U15351 (N_15351,N_14513,N_14569);
nor U15352 (N_15352,N_14894,N_14582);
xnor U15353 (N_15353,N_14506,N_14635);
and U15354 (N_15354,N_14714,N_14758);
nand U15355 (N_15355,N_14663,N_14950);
nor U15356 (N_15356,N_14881,N_14991);
and U15357 (N_15357,N_14790,N_14868);
nor U15358 (N_15358,N_14973,N_14985);
xnor U15359 (N_15359,N_14815,N_14655);
nor U15360 (N_15360,N_14995,N_14673);
nor U15361 (N_15361,N_14577,N_14948);
nor U15362 (N_15362,N_14935,N_14500);
nor U15363 (N_15363,N_14574,N_14993);
xnor U15364 (N_15364,N_14843,N_14782);
nand U15365 (N_15365,N_14783,N_14569);
and U15366 (N_15366,N_14577,N_14763);
nand U15367 (N_15367,N_14746,N_14500);
nor U15368 (N_15368,N_14544,N_14997);
or U15369 (N_15369,N_14683,N_14780);
xor U15370 (N_15370,N_14573,N_14967);
and U15371 (N_15371,N_14987,N_14820);
and U15372 (N_15372,N_14760,N_14603);
nand U15373 (N_15373,N_14611,N_14949);
nor U15374 (N_15374,N_14596,N_14907);
nand U15375 (N_15375,N_14683,N_14745);
nand U15376 (N_15376,N_14641,N_14843);
nor U15377 (N_15377,N_14851,N_14576);
or U15378 (N_15378,N_14959,N_14578);
and U15379 (N_15379,N_14566,N_14624);
xor U15380 (N_15380,N_14711,N_14720);
or U15381 (N_15381,N_14950,N_14861);
or U15382 (N_15382,N_14728,N_14760);
xor U15383 (N_15383,N_14953,N_14908);
or U15384 (N_15384,N_14929,N_14672);
nand U15385 (N_15385,N_14710,N_14866);
nor U15386 (N_15386,N_14780,N_14967);
and U15387 (N_15387,N_14833,N_14672);
nor U15388 (N_15388,N_14820,N_14960);
or U15389 (N_15389,N_14875,N_14670);
and U15390 (N_15390,N_14624,N_14957);
nor U15391 (N_15391,N_14504,N_14583);
or U15392 (N_15392,N_14844,N_14936);
or U15393 (N_15393,N_14554,N_14977);
and U15394 (N_15394,N_14706,N_14637);
nand U15395 (N_15395,N_14568,N_14955);
or U15396 (N_15396,N_14984,N_14759);
nand U15397 (N_15397,N_14937,N_14623);
and U15398 (N_15398,N_14530,N_14736);
or U15399 (N_15399,N_14707,N_14555);
or U15400 (N_15400,N_14967,N_14835);
and U15401 (N_15401,N_14683,N_14907);
xnor U15402 (N_15402,N_14771,N_14659);
nor U15403 (N_15403,N_14590,N_14793);
xnor U15404 (N_15404,N_14887,N_14856);
nor U15405 (N_15405,N_14770,N_14685);
nand U15406 (N_15406,N_14708,N_14564);
or U15407 (N_15407,N_14700,N_14569);
or U15408 (N_15408,N_14522,N_14776);
nor U15409 (N_15409,N_14917,N_14811);
nand U15410 (N_15410,N_14578,N_14597);
nand U15411 (N_15411,N_14546,N_14590);
nor U15412 (N_15412,N_14513,N_14737);
and U15413 (N_15413,N_14737,N_14828);
and U15414 (N_15414,N_14821,N_14827);
nor U15415 (N_15415,N_14699,N_14542);
and U15416 (N_15416,N_14909,N_14997);
nand U15417 (N_15417,N_14695,N_14661);
or U15418 (N_15418,N_14897,N_14907);
nand U15419 (N_15419,N_14613,N_14768);
nand U15420 (N_15420,N_14792,N_14802);
or U15421 (N_15421,N_14871,N_14745);
and U15422 (N_15422,N_14649,N_14706);
and U15423 (N_15423,N_14844,N_14505);
or U15424 (N_15424,N_14600,N_14874);
or U15425 (N_15425,N_14563,N_14656);
nand U15426 (N_15426,N_14961,N_14947);
nor U15427 (N_15427,N_14810,N_14730);
xnor U15428 (N_15428,N_14653,N_14672);
nor U15429 (N_15429,N_14688,N_14968);
or U15430 (N_15430,N_14508,N_14836);
nand U15431 (N_15431,N_14714,N_14854);
or U15432 (N_15432,N_14536,N_14546);
nor U15433 (N_15433,N_14728,N_14910);
xnor U15434 (N_15434,N_14689,N_14942);
or U15435 (N_15435,N_14872,N_14652);
xor U15436 (N_15436,N_14904,N_14824);
and U15437 (N_15437,N_14601,N_14564);
xor U15438 (N_15438,N_14594,N_14858);
nand U15439 (N_15439,N_14733,N_14576);
xor U15440 (N_15440,N_14999,N_14563);
nand U15441 (N_15441,N_14830,N_14880);
and U15442 (N_15442,N_14960,N_14754);
xor U15443 (N_15443,N_14740,N_14523);
nand U15444 (N_15444,N_14787,N_14588);
nand U15445 (N_15445,N_14606,N_14828);
and U15446 (N_15446,N_14555,N_14945);
nand U15447 (N_15447,N_14980,N_14543);
nor U15448 (N_15448,N_14773,N_14560);
nand U15449 (N_15449,N_14702,N_14948);
xnor U15450 (N_15450,N_14624,N_14734);
and U15451 (N_15451,N_14886,N_14967);
xor U15452 (N_15452,N_14952,N_14668);
xor U15453 (N_15453,N_14501,N_14892);
nor U15454 (N_15454,N_14594,N_14563);
and U15455 (N_15455,N_14558,N_14912);
or U15456 (N_15456,N_14797,N_14981);
xnor U15457 (N_15457,N_14510,N_14679);
nand U15458 (N_15458,N_14714,N_14765);
nor U15459 (N_15459,N_14826,N_14715);
nand U15460 (N_15460,N_14635,N_14986);
or U15461 (N_15461,N_14754,N_14959);
nand U15462 (N_15462,N_14653,N_14598);
or U15463 (N_15463,N_14514,N_14872);
or U15464 (N_15464,N_14586,N_14626);
or U15465 (N_15465,N_14614,N_14509);
or U15466 (N_15466,N_14787,N_14607);
xor U15467 (N_15467,N_14799,N_14915);
nor U15468 (N_15468,N_14773,N_14518);
nor U15469 (N_15469,N_14772,N_14547);
nand U15470 (N_15470,N_14532,N_14768);
and U15471 (N_15471,N_14765,N_14939);
nor U15472 (N_15472,N_14910,N_14694);
and U15473 (N_15473,N_14534,N_14809);
xor U15474 (N_15474,N_14532,N_14512);
nand U15475 (N_15475,N_14616,N_14834);
nor U15476 (N_15476,N_14785,N_14672);
or U15477 (N_15477,N_14957,N_14583);
or U15478 (N_15478,N_14930,N_14863);
xnor U15479 (N_15479,N_14557,N_14595);
or U15480 (N_15480,N_14617,N_14830);
xnor U15481 (N_15481,N_14591,N_14529);
and U15482 (N_15482,N_14578,N_14699);
xnor U15483 (N_15483,N_14724,N_14923);
or U15484 (N_15484,N_14871,N_14707);
nor U15485 (N_15485,N_14609,N_14668);
nor U15486 (N_15486,N_14772,N_14694);
nor U15487 (N_15487,N_14989,N_14950);
and U15488 (N_15488,N_14622,N_14685);
or U15489 (N_15489,N_14684,N_14735);
or U15490 (N_15490,N_14646,N_14535);
or U15491 (N_15491,N_14690,N_14993);
nor U15492 (N_15492,N_14976,N_14741);
and U15493 (N_15493,N_14881,N_14772);
xor U15494 (N_15494,N_14572,N_14810);
xor U15495 (N_15495,N_14995,N_14870);
and U15496 (N_15496,N_14786,N_14527);
nor U15497 (N_15497,N_14779,N_14927);
nand U15498 (N_15498,N_14563,N_14875);
nand U15499 (N_15499,N_14668,N_14737);
nand U15500 (N_15500,N_15358,N_15030);
xnor U15501 (N_15501,N_15147,N_15036);
xnor U15502 (N_15502,N_15087,N_15433);
xor U15503 (N_15503,N_15007,N_15263);
or U15504 (N_15504,N_15101,N_15409);
nand U15505 (N_15505,N_15340,N_15023);
nand U15506 (N_15506,N_15441,N_15499);
nand U15507 (N_15507,N_15278,N_15426);
and U15508 (N_15508,N_15205,N_15172);
or U15509 (N_15509,N_15240,N_15299);
nor U15510 (N_15510,N_15292,N_15321);
nand U15511 (N_15511,N_15350,N_15148);
or U15512 (N_15512,N_15170,N_15290);
or U15513 (N_15513,N_15028,N_15199);
nand U15514 (N_15514,N_15266,N_15370);
nor U15515 (N_15515,N_15181,N_15349);
or U15516 (N_15516,N_15466,N_15438);
nand U15517 (N_15517,N_15395,N_15270);
nor U15518 (N_15518,N_15308,N_15413);
nand U15519 (N_15519,N_15243,N_15472);
nand U15520 (N_15520,N_15168,N_15360);
xor U15521 (N_15521,N_15019,N_15444);
or U15522 (N_15522,N_15232,N_15204);
nand U15523 (N_15523,N_15218,N_15480);
nor U15524 (N_15524,N_15476,N_15376);
and U15525 (N_15525,N_15038,N_15234);
and U15526 (N_15526,N_15237,N_15437);
and U15527 (N_15527,N_15104,N_15047);
nor U15528 (N_15528,N_15415,N_15462);
xor U15529 (N_15529,N_15430,N_15295);
xnor U15530 (N_15530,N_15488,N_15265);
nor U15531 (N_15531,N_15277,N_15077);
xor U15532 (N_15532,N_15364,N_15363);
or U15533 (N_15533,N_15215,N_15152);
nor U15534 (N_15534,N_15084,N_15136);
and U15535 (N_15535,N_15453,N_15303);
nor U15536 (N_15536,N_15100,N_15421);
xor U15537 (N_15537,N_15478,N_15034);
nor U15538 (N_15538,N_15387,N_15221);
xnor U15539 (N_15539,N_15056,N_15378);
and U15540 (N_15540,N_15105,N_15385);
nand U15541 (N_15541,N_15469,N_15254);
nor U15542 (N_15542,N_15442,N_15198);
or U15543 (N_15543,N_15186,N_15337);
and U15544 (N_15544,N_15106,N_15003);
or U15545 (N_15545,N_15241,N_15079);
or U15546 (N_15546,N_15236,N_15361);
nand U15547 (N_15547,N_15163,N_15146);
xnor U15548 (N_15548,N_15216,N_15396);
and U15549 (N_15549,N_15090,N_15115);
or U15550 (N_15550,N_15344,N_15195);
xor U15551 (N_15551,N_15213,N_15103);
xor U15552 (N_15552,N_15293,N_15397);
or U15553 (N_15553,N_15238,N_15155);
nor U15554 (N_15554,N_15184,N_15315);
nor U15555 (N_15555,N_15139,N_15455);
and U15556 (N_15556,N_15200,N_15123);
xnor U15557 (N_15557,N_15403,N_15039);
or U15558 (N_15558,N_15117,N_15009);
nand U15559 (N_15559,N_15020,N_15080);
or U15560 (N_15560,N_15268,N_15405);
nor U15561 (N_15561,N_15060,N_15280);
or U15562 (N_15562,N_15246,N_15468);
nand U15563 (N_15563,N_15427,N_15006);
and U15564 (N_15564,N_15000,N_15072);
nor U15565 (N_15565,N_15282,N_15096);
and U15566 (N_15566,N_15327,N_15276);
and U15567 (N_15567,N_15259,N_15332);
xnor U15568 (N_15568,N_15356,N_15484);
nor U15569 (N_15569,N_15133,N_15026);
nand U15570 (N_15570,N_15202,N_15474);
and U15571 (N_15571,N_15473,N_15368);
nand U15572 (N_15572,N_15062,N_15074);
nand U15573 (N_15573,N_15486,N_15015);
nand U15574 (N_15574,N_15330,N_15365);
or U15575 (N_15575,N_15423,N_15402);
and U15576 (N_15576,N_15301,N_15046);
and U15577 (N_15577,N_15165,N_15322);
and U15578 (N_15578,N_15461,N_15412);
or U15579 (N_15579,N_15428,N_15223);
nand U15580 (N_15580,N_15339,N_15093);
and U15581 (N_15581,N_15109,N_15312);
or U15582 (N_15582,N_15255,N_15377);
nand U15583 (N_15583,N_15177,N_15227);
and U15584 (N_15584,N_15024,N_15372);
nor U15585 (N_15585,N_15193,N_15094);
nor U15586 (N_15586,N_15121,N_15081);
or U15587 (N_15587,N_15279,N_15171);
xor U15588 (N_15588,N_15311,N_15125);
nand U15589 (N_15589,N_15424,N_15206);
xnor U15590 (N_15590,N_15188,N_15226);
and U15591 (N_15591,N_15068,N_15008);
nand U15592 (N_15592,N_15178,N_15224);
or U15593 (N_15593,N_15491,N_15353);
nand U15594 (N_15594,N_15066,N_15318);
xnor U15595 (N_15595,N_15440,N_15061);
nand U15596 (N_15596,N_15137,N_15010);
nand U15597 (N_15597,N_15314,N_15244);
nand U15598 (N_15598,N_15251,N_15054);
and U15599 (N_15599,N_15031,N_15258);
and U15600 (N_15600,N_15045,N_15425);
xor U15601 (N_15601,N_15274,N_15214);
nand U15602 (N_15602,N_15436,N_15220);
nor U15603 (N_15603,N_15497,N_15174);
nor U15604 (N_15604,N_15228,N_15013);
nor U15605 (N_15605,N_15180,N_15035);
or U15606 (N_15606,N_15448,N_15479);
or U15607 (N_15607,N_15097,N_15065);
and U15608 (N_15608,N_15154,N_15288);
xnor U15609 (N_15609,N_15328,N_15375);
and U15610 (N_15610,N_15201,N_15119);
nand U15611 (N_15611,N_15134,N_15264);
nor U15612 (N_15612,N_15306,N_15449);
and U15613 (N_15613,N_15130,N_15207);
nand U15614 (N_15614,N_15160,N_15242);
nor U15615 (N_15615,N_15173,N_15212);
nand U15616 (N_15616,N_15092,N_15294);
nor U15617 (N_15617,N_15143,N_15260);
nor U15618 (N_15618,N_15102,N_15142);
nor U15619 (N_15619,N_15298,N_15420);
and U15620 (N_15620,N_15460,N_15281);
and U15621 (N_15621,N_15132,N_15252);
nand U15622 (N_15622,N_15287,N_15037);
nor U15623 (N_15623,N_15419,N_15158);
nor U15624 (N_15624,N_15445,N_15230);
nor U15625 (N_15625,N_15225,N_15267);
nor U15626 (N_15626,N_15383,N_15369);
or U15627 (N_15627,N_15492,N_15310);
nor U15628 (N_15628,N_15192,N_15326);
or U15629 (N_15629,N_15371,N_15304);
xnor U15630 (N_15630,N_15043,N_15408);
nand U15631 (N_15631,N_15050,N_15335);
xnor U15632 (N_15632,N_15042,N_15022);
nand U15633 (N_15633,N_15189,N_15300);
or U15634 (N_15634,N_15011,N_15343);
nand U15635 (N_15635,N_15317,N_15347);
xor U15636 (N_15636,N_15359,N_15140);
nand U15637 (N_15637,N_15398,N_15012);
and U15638 (N_15638,N_15439,N_15166);
xnor U15639 (N_15639,N_15374,N_15355);
nor U15640 (N_15640,N_15495,N_15297);
xnor U15641 (N_15641,N_15078,N_15348);
nand U15642 (N_15642,N_15016,N_15307);
nand U15643 (N_15643,N_15063,N_15052);
nand U15644 (N_15644,N_15185,N_15135);
nor U15645 (N_15645,N_15144,N_15141);
nand U15646 (N_15646,N_15346,N_15336);
or U15647 (N_15647,N_15482,N_15086);
and U15648 (N_15648,N_15187,N_15058);
nand U15649 (N_15649,N_15190,N_15457);
xor U15650 (N_15650,N_15285,N_15051);
and U15651 (N_15651,N_15248,N_15329);
xor U15652 (N_15652,N_15323,N_15451);
nor U15653 (N_15653,N_15487,N_15150);
nor U15654 (N_15654,N_15429,N_15382);
or U15655 (N_15655,N_15055,N_15489);
nor U15656 (N_15656,N_15443,N_15253);
nand U15657 (N_15657,N_15032,N_15099);
nand U15658 (N_15658,N_15247,N_15291);
xnor U15659 (N_15659,N_15362,N_15319);
or U15660 (N_15660,N_15197,N_15219);
nor U15661 (N_15661,N_15183,N_15110);
nor U15662 (N_15662,N_15176,N_15229);
or U15663 (N_15663,N_15388,N_15149);
xnor U15664 (N_15664,N_15459,N_15467);
and U15665 (N_15665,N_15222,N_15194);
or U15666 (N_15666,N_15273,N_15048);
nand U15667 (N_15667,N_15416,N_15272);
nor U15668 (N_15668,N_15483,N_15076);
or U15669 (N_15669,N_15302,N_15498);
and U15670 (N_15670,N_15410,N_15334);
nor U15671 (N_15671,N_15452,N_15250);
or U15672 (N_15672,N_15394,N_15095);
and U15673 (N_15673,N_15210,N_15431);
nor U15674 (N_15674,N_15269,N_15014);
and U15675 (N_15675,N_15027,N_15153);
nor U15676 (N_15676,N_15367,N_15208);
and U15677 (N_15677,N_15033,N_15122);
nor U15678 (N_15678,N_15470,N_15475);
nor U15679 (N_15679,N_15203,N_15040);
or U15680 (N_15680,N_15384,N_15175);
nor U15681 (N_15681,N_15157,N_15390);
or U15682 (N_15682,N_15351,N_15366);
xor U15683 (N_15683,N_15284,N_15127);
nor U15684 (N_15684,N_15354,N_15156);
and U15685 (N_15685,N_15209,N_15129);
or U15686 (N_15686,N_15379,N_15116);
nor U15687 (N_15687,N_15352,N_15041);
and U15688 (N_15688,N_15271,N_15257);
nand U15689 (N_15689,N_15496,N_15456);
nand U15690 (N_15690,N_15161,N_15091);
nand U15691 (N_15691,N_15162,N_15049);
or U15692 (N_15692,N_15447,N_15381);
nand U15693 (N_15693,N_15256,N_15124);
xor U15694 (N_15694,N_15088,N_15414);
nor U15695 (N_15695,N_15465,N_15196);
or U15696 (N_15696,N_15145,N_15261);
nand U15697 (N_15697,N_15481,N_15138);
nand U15698 (N_15698,N_15417,N_15004);
and U15699 (N_15699,N_15235,N_15400);
and U15700 (N_15700,N_15411,N_15341);
and U15701 (N_15701,N_15283,N_15477);
and U15702 (N_15702,N_15182,N_15233);
nand U15703 (N_15703,N_15380,N_15073);
or U15704 (N_15704,N_15082,N_15316);
nor U15705 (N_15705,N_15446,N_15112);
nor U15706 (N_15706,N_15471,N_15111);
xor U15707 (N_15707,N_15211,N_15128);
nor U15708 (N_15708,N_15320,N_15191);
xor U15709 (N_15709,N_15159,N_15108);
nor U15710 (N_15710,N_15025,N_15164);
or U15711 (N_15711,N_15432,N_15324);
nor U15712 (N_15712,N_15107,N_15406);
xor U15713 (N_15713,N_15059,N_15085);
or U15714 (N_15714,N_15118,N_15392);
or U15715 (N_15715,N_15044,N_15490);
xnor U15716 (N_15716,N_15067,N_15002);
xnor U15717 (N_15717,N_15120,N_15069);
nand U15718 (N_15718,N_15053,N_15179);
nand U15719 (N_15719,N_15494,N_15450);
nand U15720 (N_15720,N_15309,N_15131);
or U15721 (N_15721,N_15458,N_15338);
and U15722 (N_15722,N_15005,N_15239);
nor U15723 (N_15723,N_15399,N_15391);
nor U15724 (N_15724,N_15169,N_15151);
xor U15725 (N_15725,N_15373,N_15114);
xor U15726 (N_15726,N_15113,N_15422);
and U15727 (N_15727,N_15434,N_15345);
or U15728 (N_15728,N_15070,N_15464);
nand U15729 (N_15729,N_15098,N_15454);
and U15730 (N_15730,N_15357,N_15064);
or U15731 (N_15731,N_15435,N_15418);
nand U15732 (N_15732,N_15289,N_15386);
nand U15733 (N_15733,N_15021,N_15342);
xor U15734 (N_15734,N_15167,N_15083);
and U15735 (N_15735,N_15057,N_15296);
xnor U15736 (N_15736,N_15089,N_15029);
and U15737 (N_15737,N_15325,N_15275);
nor U15738 (N_15738,N_15001,N_15245);
or U15739 (N_15739,N_15249,N_15126);
or U15740 (N_15740,N_15018,N_15262);
nor U15741 (N_15741,N_15333,N_15493);
nand U15742 (N_15742,N_15231,N_15305);
and U15743 (N_15743,N_15071,N_15075);
xor U15744 (N_15744,N_15217,N_15404);
nor U15745 (N_15745,N_15401,N_15286);
and U15746 (N_15746,N_15331,N_15389);
nor U15747 (N_15747,N_15393,N_15407);
nor U15748 (N_15748,N_15313,N_15463);
nand U15749 (N_15749,N_15017,N_15485);
xnor U15750 (N_15750,N_15398,N_15482);
xor U15751 (N_15751,N_15412,N_15346);
nor U15752 (N_15752,N_15459,N_15437);
or U15753 (N_15753,N_15486,N_15233);
and U15754 (N_15754,N_15195,N_15097);
nor U15755 (N_15755,N_15318,N_15476);
and U15756 (N_15756,N_15387,N_15171);
or U15757 (N_15757,N_15064,N_15009);
xor U15758 (N_15758,N_15078,N_15139);
and U15759 (N_15759,N_15318,N_15221);
xor U15760 (N_15760,N_15311,N_15199);
and U15761 (N_15761,N_15089,N_15428);
nand U15762 (N_15762,N_15333,N_15208);
or U15763 (N_15763,N_15139,N_15099);
and U15764 (N_15764,N_15285,N_15460);
or U15765 (N_15765,N_15462,N_15328);
or U15766 (N_15766,N_15418,N_15143);
or U15767 (N_15767,N_15201,N_15325);
xor U15768 (N_15768,N_15092,N_15213);
or U15769 (N_15769,N_15026,N_15188);
nor U15770 (N_15770,N_15086,N_15186);
and U15771 (N_15771,N_15171,N_15274);
xor U15772 (N_15772,N_15133,N_15473);
nand U15773 (N_15773,N_15472,N_15393);
xnor U15774 (N_15774,N_15201,N_15313);
nor U15775 (N_15775,N_15060,N_15181);
nand U15776 (N_15776,N_15239,N_15043);
nand U15777 (N_15777,N_15106,N_15034);
nand U15778 (N_15778,N_15188,N_15033);
and U15779 (N_15779,N_15161,N_15154);
xnor U15780 (N_15780,N_15221,N_15287);
nand U15781 (N_15781,N_15449,N_15099);
nand U15782 (N_15782,N_15106,N_15340);
or U15783 (N_15783,N_15105,N_15245);
xnor U15784 (N_15784,N_15023,N_15302);
or U15785 (N_15785,N_15335,N_15202);
and U15786 (N_15786,N_15219,N_15130);
xor U15787 (N_15787,N_15280,N_15165);
xor U15788 (N_15788,N_15442,N_15076);
nor U15789 (N_15789,N_15055,N_15377);
or U15790 (N_15790,N_15370,N_15334);
nand U15791 (N_15791,N_15356,N_15449);
or U15792 (N_15792,N_15131,N_15273);
or U15793 (N_15793,N_15080,N_15251);
nand U15794 (N_15794,N_15397,N_15270);
or U15795 (N_15795,N_15484,N_15438);
xor U15796 (N_15796,N_15170,N_15485);
and U15797 (N_15797,N_15121,N_15109);
or U15798 (N_15798,N_15393,N_15228);
or U15799 (N_15799,N_15260,N_15334);
xnor U15800 (N_15800,N_15239,N_15202);
nand U15801 (N_15801,N_15467,N_15296);
nor U15802 (N_15802,N_15337,N_15451);
nor U15803 (N_15803,N_15320,N_15156);
or U15804 (N_15804,N_15072,N_15391);
xnor U15805 (N_15805,N_15352,N_15432);
and U15806 (N_15806,N_15258,N_15335);
or U15807 (N_15807,N_15215,N_15231);
xor U15808 (N_15808,N_15190,N_15482);
xor U15809 (N_15809,N_15408,N_15073);
and U15810 (N_15810,N_15254,N_15499);
xor U15811 (N_15811,N_15348,N_15060);
xnor U15812 (N_15812,N_15304,N_15480);
nand U15813 (N_15813,N_15429,N_15482);
nor U15814 (N_15814,N_15371,N_15251);
and U15815 (N_15815,N_15246,N_15416);
nor U15816 (N_15816,N_15488,N_15388);
and U15817 (N_15817,N_15232,N_15494);
xor U15818 (N_15818,N_15475,N_15366);
or U15819 (N_15819,N_15281,N_15346);
and U15820 (N_15820,N_15031,N_15318);
or U15821 (N_15821,N_15301,N_15376);
nor U15822 (N_15822,N_15436,N_15246);
nor U15823 (N_15823,N_15477,N_15175);
or U15824 (N_15824,N_15421,N_15185);
xor U15825 (N_15825,N_15079,N_15229);
xor U15826 (N_15826,N_15110,N_15396);
xor U15827 (N_15827,N_15406,N_15281);
or U15828 (N_15828,N_15042,N_15356);
xnor U15829 (N_15829,N_15005,N_15038);
xor U15830 (N_15830,N_15207,N_15402);
nor U15831 (N_15831,N_15334,N_15171);
or U15832 (N_15832,N_15103,N_15412);
nor U15833 (N_15833,N_15458,N_15083);
and U15834 (N_15834,N_15466,N_15004);
xnor U15835 (N_15835,N_15343,N_15454);
nand U15836 (N_15836,N_15394,N_15136);
xor U15837 (N_15837,N_15286,N_15449);
and U15838 (N_15838,N_15350,N_15338);
xnor U15839 (N_15839,N_15414,N_15272);
nor U15840 (N_15840,N_15130,N_15054);
nor U15841 (N_15841,N_15248,N_15019);
xnor U15842 (N_15842,N_15317,N_15335);
and U15843 (N_15843,N_15217,N_15036);
xor U15844 (N_15844,N_15420,N_15171);
or U15845 (N_15845,N_15118,N_15335);
nor U15846 (N_15846,N_15232,N_15340);
and U15847 (N_15847,N_15147,N_15180);
and U15848 (N_15848,N_15366,N_15446);
nor U15849 (N_15849,N_15326,N_15161);
nand U15850 (N_15850,N_15315,N_15000);
and U15851 (N_15851,N_15097,N_15450);
or U15852 (N_15852,N_15353,N_15365);
and U15853 (N_15853,N_15222,N_15314);
or U15854 (N_15854,N_15385,N_15456);
xnor U15855 (N_15855,N_15255,N_15336);
or U15856 (N_15856,N_15247,N_15148);
nand U15857 (N_15857,N_15494,N_15103);
nand U15858 (N_15858,N_15115,N_15161);
xor U15859 (N_15859,N_15195,N_15015);
and U15860 (N_15860,N_15341,N_15387);
or U15861 (N_15861,N_15255,N_15116);
and U15862 (N_15862,N_15348,N_15487);
nor U15863 (N_15863,N_15268,N_15286);
nor U15864 (N_15864,N_15253,N_15233);
nand U15865 (N_15865,N_15050,N_15005);
xor U15866 (N_15866,N_15383,N_15266);
and U15867 (N_15867,N_15042,N_15434);
or U15868 (N_15868,N_15146,N_15350);
nor U15869 (N_15869,N_15482,N_15395);
or U15870 (N_15870,N_15119,N_15145);
xnor U15871 (N_15871,N_15218,N_15160);
xnor U15872 (N_15872,N_15056,N_15149);
or U15873 (N_15873,N_15405,N_15257);
nand U15874 (N_15874,N_15102,N_15353);
and U15875 (N_15875,N_15048,N_15102);
and U15876 (N_15876,N_15198,N_15168);
or U15877 (N_15877,N_15440,N_15151);
nand U15878 (N_15878,N_15266,N_15430);
or U15879 (N_15879,N_15211,N_15305);
or U15880 (N_15880,N_15071,N_15201);
xnor U15881 (N_15881,N_15209,N_15178);
and U15882 (N_15882,N_15308,N_15420);
or U15883 (N_15883,N_15387,N_15153);
nor U15884 (N_15884,N_15436,N_15014);
xnor U15885 (N_15885,N_15224,N_15453);
nor U15886 (N_15886,N_15024,N_15363);
or U15887 (N_15887,N_15068,N_15049);
or U15888 (N_15888,N_15193,N_15089);
nor U15889 (N_15889,N_15376,N_15426);
and U15890 (N_15890,N_15494,N_15312);
xnor U15891 (N_15891,N_15010,N_15272);
nand U15892 (N_15892,N_15388,N_15274);
nand U15893 (N_15893,N_15396,N_15398);
nor U15894 (N_15894,N_15329,N_15150);
xnor U15895 (N_15895,N_15126,N_15180);
or U15896 (N_15896,N_15238,N_15221);
or U15897 (N_15897,N_15226,N_15252);
and U15898 (N_15898,N_15375,N_15494);
nand U15899 (N_15899,N_15156,N_15134);
and U15900 (N_15900,N_15204,N_15064);
and U15901 (N_15901,N_15029,N_15291);
nand U15902 (N_15902,N_15347,N_15465);
or U15903 (N_15903,N_15284,N_15467);
nor U15904 (N_15904,N_15365,N_15303);
nor U15905 (N_15905,N_15184,N_15155);
nand U15906 (N_15906,N_15406,N_15136);
xor U15907 (N_15907,N_15169,N_15327);
xor U15908 (N_15908,N_15467,N_15308);
nand U15909 (N_15909,N_15098,N_15245);
nand U15910 (N_15910,N_15447,N_15150);
xnor U15911 (N_15911,N_15195,N_15100);
nor U15912 (N_15912,N_15326,N_15201);
nand U15913 (N_15913,N_15010,N_15452);
or U15914 (N_15914,N_15181,N_15292);
or U15915 (N_15915,N_15160,N_15288);
nor U15916 (N_15916,N_15475,N_15264);
nor U15917 (N_15917,N_15250,N_15465);
nand U15918 (N_15918,N_15480,N_15013);
or U15919 (N_15919,N_15265,N_15070);
xor U15920 (N_15920,N_15390,N_15275);
or U15921 (N_15921,N_15427,N_15348);
and U15922 (N_15922,N_15277,N_15194);
nand U15923 (N_15923,N_15407,N_15191);
nor U15924 (N_15924,N_15197,N_15490);
or U15925 (N_15925,N_15136,N_15238);
nand U15926 (N_15926,N_15488,N_15069);
or U15927 (N_15927,N_15471,N_15321);
xnor U15928 (N_15928,N_15356,N_15417);
and U15929 (N_15929,N_15311,N_15212);
nand U15930 (N_15930,N_15033,N_15205);
or U15931 (N_15931,N_15425,N_15285);
or U15932 (N_15932,N_15417,N_15334);
or U15933 (N_15933,N_15164,N_15414);
nor U15934 (N_15934,N_15127,N_15024);
or U15935 (N_15935,N_15256,N_15389);
xnor U15936 (N_15936,N_15041,N_15203);
nor U15937 (N_15937,N_15345,N_15379);
nand U15938 (N_15938,N_15336,N_15481);
xnor U15939 (N_15939,N_15259,N_15009);
and U15940 (N_15940,N_15266,N_15406);
nor U15941 (N_15941,N_15360,N_15488);
and U15942 (N_15942,N_15491,N_15351);
nand U15943 (N_15943,N_15213,N_15266);
nor U15944 (N_15944,N_15010,N_15177);
xnor U15945 (N_15945,N_15321,N_15104);
xnor U15946 (N_15946,N_15102,N_15041);
xnor U15947 (N_15947,N_15014,N_15235);
nor U15948 (N_15948,N_15319,N_15253);
nand U15949 (N_15949,N_15471,N_15272);
nor U15950 (N_15950,N_15080,N_15204);
xor U15951 (N_15951,N_15344,N_15469);
or U15952 (N_15952,N_15496,N_15152);
or U15953 (N_15953,N_15342,N_15068);
nand U15954 (N_15954,N_15142,N_15316);
and U15955 (N_15955,N_15208,N_15338);
xnor U15956 (N_15956,N_15326,N_15451);
or U15957 (N_15957,N_15146,N_15438);
or U15958 (N_15958,N_15457,N_15487);
xor U15959 (N_15959,N_15141,N_15271);
nor U15960 (N_15960,N_15002,N_15317);
and U15961 (N_15961,N_15009,N_15287);
and U15962 (N_15962,N_15121,N_15150);
xnor U15963 (N_15963,N_15406,N_15342);
and U15964 (N_15964,N_15398,N_15456);
nor U15965 (N_15965,N_15383,N_15355);
xnor U15966 (N_15966,N_15473,N_15356);
or U15967 (N_15967,N_15321,N_15116);
and U15968 (N_15968,N_15330,N_15487);
nor U15969 (N_15969,N_15339,N_15023);
or U15970 (N_15970,N_15189,N_15304);
and U15971 (N_15971,N_15473,N_15286);
xnor U15972 (N_15972,N_15053,N_15172);
nor U15973 (N_15973,N_15061,N_15317);
xnor U15974 (N_15974,N_15226,N_15253);
nand U15975 (N_15975,N_15287,N_15405);
nor U15976 (N_15976,N_15210,N_15003);
and U15977 (N_15977,N_15397,N_15398);
nand U15978 (N_15978,N_15014,N_15191);
xnor U15979 (N_15979,N_15269,N_15219);
or U15980 (N_15980,N_15286,N_15290);
and U15981 (N_15981,N_15149,N_15323);
nand U15982 (N_15982,N_15405,N_15052);
xor U15983 (N_15983,N_15312,N_15300);
or U15984 (N_15984,N_15185,N_15134);
xor U15985 (N_15985,N_15011,N_15295);
nor U15986 (N_15986,N_15442,N_15191);
and U15987 (N_15987,N_15186,N_15317);
nor U15988 (N_15988,N_15073,N_15366);
nand U15989 (N_15989,N_15187,N_15455);
nor U15990 (N_15990,N_15299,N_15146);
nand U15991 (N_15991,N_15354,N_15088);
nor U15992 (N_15992,N_15415,N_15204);
and U15993 (N_15993,N_15217,N_15435);
nor U15994 (N_15994,N_15094,N_15042);
nor U15995 (N_15995,N_15007,N_15110);
and U15996 (N_15996,N_15307,N_15484);
nand U15997 (N_15997,N_15458,N_15360);
nand U15998 (N_15998,N_15442,N_15423);
nor U15999 (N_15999,N_15242,N_15237);
nand U16000 (N_16000,N_15726,N_15687);
nand U16001 (N_16001,N_15772,N_15601);
nand U16002 (N_16002,N_15525,N_15786);
nand U16003 (N_16003,N_15784,N_15551);
nor U16004 (N_16004,N_15899,N_15560);
nand U16005 (N_16005,N_15521,N_15925);
xnor U16006 (N_16006,N_15651,N_15892);
xor U16007 (N_16007,N_15556,N_15978);
xor U16008 (N_16008,N_15540,N_15608);
nor U16009 (N_16009,N_15904,N_15590);
and U16010 (N_16010,N_15977,N_15815);
and U16011 (N_16011,N_15811,N_15634);
xor U16012 (N_16012,N_15652,N_15759);
and U16013 (N_16013,N_15727,N_15664);
nand U16014 (N_16014,N_15967,N_15822);
nor U16015 (N_16015,N_15663,N_15854);
xor U16016 (N_16016,N_15890,N_15922);
and U16017 (N_16017,N_15610,N_15713);
or U16018 (N_16018,N_15564,N_15975);
and U16019 (N_16019,N_15565,N_15505);
nor U16020 (N_16020,N_15766,N_15791);
xor U16021 (N_16021,N_15558,N_15607);
and U16022 (N_16022,N_15718,N_15573);
xor U16023 (N_16023,N_15912,N_15535);
nor U16024 (N_16024,N_15554,N_15571);
and U16025 (N_16025,N_15699,N_15548);
nand U16026 (N_16026,N_15753,N_15812);
xor U16027 (N_16027,N_15657,N_15983);
xor U16028 (N_16028,N_15690,N_15576);
xnor U16029 (N_16029,N_15679,N_15761);
or U16030 (N_16030,N_15821,N_15902);
and U16031 (N_16031,N_15751,N_15875);
or U16032 (N_16032,N_15804,N_15613);
xnor U16033 (N_16033,N_15650,N_15592);
or U16034 (N_16034,N_15619,N_15817);
nand U16035 (N_16035,N_15883,N_15867);
or U16036 (N_16036,N_15615,N_15711);
xnor U16037 (N_16037,N_15924,N_15893);
xor U16038 (N_16038,N_15783,N_15585);
xnor U16039 (N_16039,N_15796,N_15896);
nand U16040 (N_16040,N_15670,N_15760);
nor U16041 (N_16041,N_15536,N_15935);
or U16042 (N_16042,N_15838,N_15996);
or U16043 (N_16043,N_15717,N_15513);
nand U16044 (N_16044,N_15980,N_15775);
and U16045 (N_16045,N_15595,N_15919);
nor U16046 (N_16046,N_15524,N_15943);
or U16047 (N_16047,N_15530,N_15877);
or U16048 (N_16048,N_15516,N_15597);
nand U16049 (N_16049,N_15981,N_15827);
and U16050 (N_16050,N_15777,N_15633);
or U16051 (N_16051,N_15654,N_15839);
nand U16052 (N_16052,N_15616,N_15689);
nor U16053 (N_16053,N_15695,N_15872);
nand U16054 (N_16054,N_15829,N_15742);
nand U16055 (N_16055,N_15789,N_15873);
and U16056 (N_16056,N_15820,N_15696);
xor U16057 (N_16057,N_15646,N_15933);
nand U16058 (N_16058,N_15721,N_15724);
or U16059 (N_16059,N_15602,N_15675);
and U16060 (N_16060,N_15735,N_15946);
nand U16061 (N_16061,N_15984,N_15553);
and U16062 (N_16062,N_15641,N_15862);
or U16063 (N_16063,N_15624,N_15769);
nor U16064 (N_16064,N_15940,N_15776);
nand U16065 (N_16065,N_15974,N_15710);
nor U16066 (N_16066,N_15959,N_15806);
and U16067 (N_16067,N_15858,N_15611);
and U16068 (N_16068,N_15855,N_15744);
nor U16069 (N_16069,N_15960,N_15596);
xor U16070 (N_16070,N_15620,N_15734);
xor U16071 (N_16071,N_15931,N_15770);
nor U16072 (N_16072,N_15517,N_15562);
or U16073 (N_16073,N_15808,N_15968);
nor U16074 (N_16074,N_15880,N_15637);
nand U16075 (N_16075,N_15847,N_15965);
or U16076 (N_16076,N_15976,N_15934);
nor U16077 (N_16077,N_15681,N_15503);
nor U16078 (N_16078,N_15966,N_15972);
nand U16079 (N_16079,N_15989,N_15510);
or U16080 (N_16080,N_15501,N_15843);
and U16081 (N_16081,N_15835,N_15743);
and U16082 (N_16082,N_15531,N_15544);
nand U16083 (N_16083,N_15589,N_15988);
and U16084 (N_16084,N_15701,N_15903);
nand U16085 (N_16085,N_15627,N_15840);
or U16086 (N_16086,N_15618,N_15956);
nor U16087 (N_16087,N_15732,N_15778);
nand U16088 (N_16088,N_15962,N_15938);
and U16089 (N_16089,N_15583,N_15889);
or U16090 (N_16090,N_15771,N_15950);
or U16091 (N_16091,N_15706,N_15729);
and U16092 (N_16092,N_15694,N_15999);
and U16093 (N_16093,N_15522,N_15969);
and U16094 (N_16094,N_15716,N_15911);
or U16095 (N_16095,N_15799,N_15916);
nor U16096 (N_16096,N_15667,N_15685);
nand U16097 (N_16097,N_15655,N_15936);
nand U16098 (N_16098,N_15942,N_15870);
nor U16099 (N_16099,N_15591,N_15567);
and U16100 (N_16100,N_15901,N_15692);
and U16101 (N_16101,N_15550,N_15745);
or U16102 (N_16102,N_15795,N_15702);
xor U16103 (N_16103,N_15863,N_15756);
or U16104 (N_16104,N_15508,N_15955);
nand U16105 (N_16105,N_15635,N_15686);
nor U16106 (N_16106,N_15569,N_15539);
nand U16107 (N_16107,N_15683,N_15780);
xor U16108 (N_16108,N_15794,N_15851);
xor U16109 (N_16109,N_15866,N_15906);
xnor U16110 (N_16110,N_15871,N_15845);
or U16111 (N_16111,N_15653,N_15793);
or U16112 (N_16112,N_15814,N_15830);
xnor U16113 (N_16113,N_15599,N_15606);
xor U16114 (N_16114,N_15684,N_15825);
or U16115 (N_16115,N_15882,N_15700);
nor U16116 (N_16116,N_15671,N_15884);
and U16117 (N_16117,N_15909,N_15860);
nor U16118 (N_16118,N_15659,N_15574);
nand U16119 (N_16119,N_15537,N_15774);
or U16120 (N_16120,N_15810,N_15737);
nor U16121 (N_16121,N_15970,N_15861);
nor U16122 (N_16122,N_15844,N_15728);
nand U16123 (N_16123,N_15639,N_15951);
nor U16124 (N_16124,N_15688,N_15779);
or U16125 (N_16125,N_15673,N_15660);
and U16126 (N_16126,N_15869,N_15908);
or U16127 (N_16127,N_15868,N_15905);
xnor U16128 (N_16128,N_15813,N_15939);
or U16129 (N_16129,N_15894,N_15763);
and U16130 (N_16130,N_15676,N_15831);
xnor U16131 (N_16131,N_15586,N_15807);
and U16132 (N_16132,N_15865,N_15898);
nor U16133 (N_16133,N_15523,N_15948);
or U16134 (N_16134,N_15617,N_15581);
nor U16135 (N_16135,N_15693,N_15926);
or U16136 (N_16136,N_15632,N_15929);
or U16137 (N_16137,N_15719,N_15707);
xor U16138 (N_16138,N_15588,N_15768);
and U16139 (N_16139,N_15644,N_15832);
or U16140 (N_16140,N_15973,N_15656);
xnor U16141 (N_16141,N_15614,N_15918);
and U16142 (N_16142,N_15964,N_15750);
and U16143 (N_16143,N_15913,N_15991);
or U16144 (N_16144,N_15714,N_15559);
xor U16145 (N_16145,N_15547,N_15900);
and U16146 (N_16146,N_15947,N_15785);
nor U16147 (N_16147,N_15930,N_15605);
nand U16148 (N_16148,N_15949,N_15527);
or U16149 (N_16149,N_15740,N_15878);
nor U16150 (N_16150,N_15698,N_15720);
or U16151 (N_16151,N_15741,N_15953);
and U16152 (N_16152,N_15647,N_15837);
nor U16153 (N_16153,N_15738,N_15502);
nand U16154 (N_16154,N_15764,N_15715);
nor U16155 (N_16155,N_15538,N_15891);
nor U16156 (N_16156,N_15542,N_15986);
nor U16157 (N_16157,N_15885,N_15534);
and U16158 (N_16158,N_15747,N_15669);
and U16159 (N_16159,N_15985,N_15665);
and U16160 (N_16160,N_15625,N_15642);
and U16161 (N_16161,N_15703,N_15823);
and U16162 (N_16162,N_15834,N_15725);
nand U16163 (N_16163,N_15612,N_15662);
or U16164 (N_16164,N_15963,N_15888);
or U16165 (N_16165,N_15582,N_15680);
or U16166 (N_16166,N_15677,N_15636);
nand U16167 (N_16167,N_15752,N_15575);
or U16168 (N_16168,N_15824,N_15526);
or U16169 (N_16169,N_15736,N_15897);
or U16170 (N_16170,N_15598,N_15819);
nand U16171 (N_16171,N_15570,N_15923);
nor U16172 (N_16172,N_15971,N_15626);
nor U16173 (N_16173,N_15500,N_15631);
or U16174 (N_16174,N_15767,N_15874);
nor U16175 (N_16175,N_15666,N_15773);
or U16176 (N_16176,N_15826,N_15557);
or U16177 (N_16177,N_15992,N_15762);
or U16178 (N_16178,N_15731,N_15708);
xor U16179 (N_16179,N_15887,N_15543);
nand U16180 (N_16180,N_15842,N_15928);
nor U16181 (N_16181,N_15579,N_15803);
or U16182 (N_16182,N_15957,N_15623);
or U16183 (N_16183,N_15998,N_15781);
nor U16184 (N_16184,N_15529,N_15661);
or U16185 (N_16185,N_15746,N_15853);
and U16186 (N_16186,N_15798,N_15805);
or U16187 (N_16187,N_15649,N_15850);
nand U16188 (N_16188,N_15628,N_15739);
xnor U16189 (N_16189,N_15915,N_15881);
xnor U16190 (N_16190,N_15697,N_15857);
xor U16191 (N_16191,N_15859,N_15994);
and U16192 (N_16192,N_15507,N_15528);
nor U16193 (N_16193,N_15952,N_15841);
xor U16194 (N_16194,N_15809,N_15563);
and U16195 (N_16195,N_15682,N_15648);
and U16196 (N_16196,N_15987,N_15566);
nand U16197 (N_16197,N_15621,N_15638);
nor U16198 (N_16198,N_15712,N_15722);
or U16199 (N_16199,N_15577,N_15552);
xnor U16200 (N_16200,N_15580,N_15997);
nor U16201 (N_16201,N_15749,N_15568);
or U16202 (N_16202,N_15849,N_15800);
nand U16203 (N_16203,N_15758,N_15917);
and U16204 (N_16204,N_15604,N_15630);
nand U16205 (N_16205,N_15937,N_15578);
nor U16206 (N_16206,N_15886,N_15546);
nand U16207 (N_16207,N_15941,N_15895);
or U16208 (N_16208,N_15828,N_15788);
nand U16209 (N_16209,N_15782,N_15512);
nor U16210 (N_16210,N_15982,N_15765);
nand U16211 (N_16211,N_15643,N_15852);
nor U16212 (N_16212,N_15757,N_15914);
and U16213 (N_16213,N_15790,N_15755);
nor U16214 (N_16214,N_15848,N_15518);
xnor U16215 (N_16215,N_15674,N_15593);
nand U16216 (N_16216,N_15920,N_15515);
nand U16217 (N_16217,N_15549,N_15555);
nor U16218 (N_16218,N_15704,N_15532);
nor U16219 (N_16219,N_15910,N_15678);
nand U16220 (N_16220,N_15561,N_15691);
nor U16221 (N_16221,N_15705,N_15545);
nand U16222 (N_16222,N_15907,N_15954);
nand U16223 (N_16223,N_15792,N_15879);
nand U16224 (N_16224,N_15730,N_15801);
xnor U16225 (N_16225,N_15519,N_15645);
or U16226 (N_16226,N_15833,N_15995);
nand U16227 (N_16227,N_15609,N_15603);
xnor U16228 (N_16228,N_15511,N_15709);
xor U16229 (N_16229,N_15864,N_15672);
nor U16230 (N_16230,N_15629,N_15818);
or U16231 (N_16231,N_15927,N_15600);
nor U16232 (N_16232,N_15668,N_15723);
nand U16233 (N_16233,N_15958,N_15640);
or U16234 (N_16234,N_15514,N_15797);
and U16235 (N_16235,N_15594,N_15961);
nand U16236 (N_16236,N_15993,N_15509);
nor U16237 (N_16237,N_15787,N_15856);
xnor U16238 (N_16238,N_15846,N_15572);
xnor U16239 (N_16239,N_15754,N_15944);
nor U16240 (N_16240,N_15945,N_15584);
xnor U16241 (N_16241,N_15533,N_15990);
nor U16242 (N_16242,N_15748,N_15622);
or U16243 (N_16243,N_15587,N_15520);
xor U16244 (N_16244,N_15816,N_15921);
xnor U16245 (N_16245,N_15802,N_15504);
and U16246 (N_16246,N_15876,N_15979);
nor U16247 (N_16247,N_15541,N_15733);
and U16248 (N_16248,N_15932,N_15836);
nor U16249 (N_16249,N_15658,N_15506);
nor U16250 (N_16250,N_15958,N_15642);
nand U16251 (N_16251,N_15699,N_15847);
nor U16252 (N_16252,N_15984,N_15761);
and U16253 (N_16253,N_15691,N_15807);
nor U16254 (N_16254,N_15568,N_15614);
or U16255 (N_16255,N_15737,N_15820);
xnor U16256 (N_16256,N_15873,N_15889);
nor U16257 (N_16257,N_15604,N_15995);
or U16258 (N_16258,N_15964,N_15939);
and U16259 (N_16259,N_15620,N_15765);
nor U16260 (N_16260,N_15755,N_15602);
xor U16261 (N_16261,N_15827,N_15914);
nand U16262 (N_16262,N_15847,N_15653);
or U16263 (N_16263,N_15928,N_15611);
xor U16264 (N_16264,N_15839,N_15553);
nor U16265 (N_16265,N_15872,N_15669);
nand U16266 (N_16266,N_15726,N_15869);
and U16267 (N_16267,N_15646,N_15716);
nor U16268 (N_16268,N_15916,N_15962);
and U16269 (N_16269,N_15638,N_15695);
nor U16270 (N_16270,N_15995,N_15506);
xnor U16271 (N_16271,N_15793,N_15547);
nand U16272 (N_16272,N_15868,N_15691);
and U16273 (N_16273,N_15606,N_15865);
nor U16274 (N_16274,N_15692,N_15760);
and U16275 (N_16275,N_15934,N_15799);
nor U16276 (N_16276,N_15723,N_15730);
nand U16277 (N_16277,N_15536,N_15597);
xnor U16278 (N_16278,N_15628,N_15854);
nor U16279 (N_16279,N_15678,N_15792);
nand U16280 (N_16280,N_15884,N_15666);
nand U16281 (N_16281,N_15623,N_15643);
nand U16282 (N_16282,N_15712,N_15871);
or U16283 (N_16283,N_15583,N_15898);
xnor U16284 (N_16284,N_15884,N_15716);
nor U16285 (N_16285,N_15733,N_15583);
or U16286 (N_16286,N_15638,N_15927);
xnor U16287 (N_16287,N_15635,N_15691);
and U16288 (N_16288,N_15894,N_15968);
nor U16289 (N_16289,N_15793,N_15640);
and U16290 (N_16290,N_15666,N_15688);
and U16291 (N_16291,N_15516,N_15764);
or U16292 (N_16292,N_15554,N_15619);
or U16293 (N_16293,N_15957,N_15526);
or U16294 (N_16294,N_15600,N_15674);
and U16295 (N_16295,N_15611,N_15827);
xnor U16296 (N_16296,N_15794,N_15657);
nand U16297 (N_16297,N_15763,N_15971);
or U16298 (N_16298,N_15679,N_15817);
nor U16299 (N_16299,N_15615,N_15953);
or U16300 (N_16300,N_15681,N_15847);
or U16301 (N_16301,N_15732,N_15862);
or U16302 (N_16302,N_15884,N_15737);
xor U16303 (N_16303,N_15676,N_15843);
nor U16304 (N_16304,N_15724,N_15563);
or U16305 (N_16305,N_15889,N_15681);
or U16306 (N_16306,N_15942,N_15793);
xor U16307 (N_16307,N_15673,N_15966);
nand U16308 (N_16308,N_15671,N_15792);
or U16309 (N_16309,N_15566,N_15889);
xor U16310 (N_16310,N_15834,N_15692);
and U16311 (N_16311,N_15876,N_15917);
or U16312 (N_16312,N_15606,N_15680);
xor U16313 (N_16313,N_15594,N_15911);
nor U16314 (N_16314,N_15622,N_15590);
and U16315 (N_16315,N_15677,N_15767);
nand U16316 (N_16316,N_15903,N_15646);
or U16317 (N_16317,N_15901,N_15762);
nor U16318 (N_16318,N_15782,N_15874);
nor U16319 (N_16319,N_15865,N_15934);
nand U16320 (N_16320,N_15576,N_15993);
nor U16321 (N_16321,N_15832,N_15720);
nor U16322 (N_16322,N_15720,N_15870);
nor U16323 (N_16323,N_15779,N_15519);
xnor U16324 (N_16324,N_15942,N_15523);
and U16325 (N_16325,N_15525,N_15507);
or U16326 (N_16326,N_15502,N_15755);
and U16327 (N_16327,N_15903,N_15920);
and U16328 (N_16328,N_15875,N_15729);
nor U16329 (N_16329,N_15580,N_15736);
nor U16330 (N_16330,N_15889,N_15617);
nor U16331 (N_16331,N_15537,N_15779);
or U16332 (N_16332,N_15965,N_15616);
nor U16333 (N_16333,N_15623,N_15641);
nor U16334 (N_16334,N_15898,N_15984);
xnor U16335 (N_16335,N_15708,N_15586);
xnor U16336 (N_16336,N_15659,N_15642);
and U16337 (N_16337,N_15502,N_15557);
or U16338 (N_16338,N_15864,N_15794);
nor U16339 (N_16339,N_15977,N_15651);
and U16340 (N_16340,N_15961,N_15540);
and U16341 (N_16341,N_15881,N_15577);
nand U16342 (N_16342,N_15636,N_15786);
nor U16343 (N_16343,N_15753,N_15939);
xnor U16344 (N_16344,N_15858,N_15748);
nor U16345 (N_16345,N_15609,N_15926);
or U16346 (N_16346,N_15984,N_15812);
xor U16347 (N_16347,N_15519,N_15869);
or U16348 (N_16348,N_15920,N_15513);
nor U16349 (N_16349,N_15743,N_15605);
or U16350 (N_16350,N_15885,N_15560);
nand U16351 (N_16351,N_15514,N_15747);
or U16352 (N_16352,N_15662,N_15521);
nand U16353 (N_16353,N_15958,N_15593);
or U16354 (N_16354,N_15724,N_15616);
or U16355 (N_16355,N_15754,N_15551);
nand U16356 (N_16356,N_15816,N_15632);
nor U16357 (N_16357,N_15897,N_15516);
and U16358 (N_16358,N_15673,N_15899);
or U16359 (N_16359,N_15895,N_15767);
xor U16360 (N_16360,N_15749,N_15919);
xnor U16361 (N_16361,N_15714,N_15537);
or U16362 (N_16362,N_15666,N_15633);
nor U16363 (N_16363,N_15617,N_15728);
xnor U16364 (N_16364,N_15669,N_15610);
xor U16365 (N_16365,N_15700,N_15974);
and U16366 (N_16366,N_15668,N_15934);
xor U16367 (N_16367,N_15789,N_15900);
or U16368 (N_16368,N_15584,N_15998);
and U16369 (N_16369,N_15650,N_15850);
nor U16370 (N_16370,N_15625,N_15502);
nand U16371 (N_16371,N_15962,N_15641);
and U16372 (N_16372,N_15835,N_15995);
or U16373 (N_16373,N_15775,N_15716);
xnor U16374 (N_16374,N_15827,N_15791);
nand U16375 (N_16375,N_15823,N_15582);
and U16376 (N_16376,N_15792,N_15896);
nor U16377 (N_16377,N_15612,N_15946);
nor U16378 (N_16378,N_15947,N_15961);
nand U16379 (N_16379,N_15686,N_15519);
nand U16380 (N_16380,N_15934,N_15962);
nor U16381 (N_16381,N_15790,N_15652);
nor U16382 (N_16382,N_15901,N_15510);
and U16383 (N_16383,N_15727,N_15879);
or U16384 (N_16384,N_15790,N_15741);
and U16385 (N_16385,N_15629,N_15795);
nand U16386 (N_16386,N_15953,N_15649);
nor U16387 (N_16387,N_15975,N_15576);
nand U16388 (N_16388,N_15742,N_15554);
xnor U16389 (N_16389,N_15744,N_15579);
and U16390 (N_16390,N_15764,N_15684);
xor U16391 (N_16391,N_15643,N_15991);
nand U16392 (N_16392,N_15678,N_15800);
xnor U16393 (N_16393,N_15807,N_15995);
or U16394 (N_16394,N_15678,N_15770);
nand U16395 (N_16395,N_15643,N_15618);
nor U16396 (N_16396,N_15956,N_15732);
and U16397 (N_16397,N_15802,N_15850);
xnor U16398 (N_16398,N_15979,N_15633);
nand U16399 (N_16399,N_15535,N_15915);
or U16400 (N_16400,N_15977,N_15712);
xor U16401 (N_16401,N_15908,N_15532);
and U16402 (N_16402,N_15523,N_15575);
nand U16403 (N_16403,N_15542,N_15540);
and U16404 (N_16404,N_15657,N_15807);
and U16405 (N_16405,N_15549,N_15584);
nor U16406 (N_16406,N_15838,N_15621);
xnor U16407 (N_16407,N_15643,N_15533);
and U16408 (N_16408,N_15959,N_15650);
or U16409 (N_16409,N_15653,N_15928);
xor U16410 (N_16410,N_15774,N_15582);
or U16411 (N_16411,N_15902,N_15627);
xnor U16412 (N_16412,N_15941,N_15911);
nor U16413 (N_16413,N_15972,N_15600);
nand U16414 (N_16414,N_15591,N_15535);
and U16415 (N_16415,N_15835,N_15891);
nor U16416 (N_16416,N_15966,N_15958);
nand U16417 (N_16417,N_15662,N_15807);
nand U16418 (N_16418,N_15712,N_15642);
nor U16419 (N_16419,N_15648,N_15533);
xnor U16420 (N_16420,N_15917,N_15508);
nor U16421 (N_16421,N_15784,N_15968);
nand U16422 (N_16422,N_15674,N_15888);
or U16423 (N_16423,N_15830,N_15954);
nand U16424 (N_16424,N_15572,N_15797);
or U16425 (N_16425,N_15551,N_15741);
nand U16426 (N_16426,N_15938,N_15891);
nor U16427 (N_16427,N_15508,N_15768);
and U16428 (N_16428,N_15896,N_15649);
xor U16429 (N_16429,N_15921,N_15809);
and U16430 (N_16430,N_15621,N_15702);
or U16431 (N_16431,N_15887,N_15717);
and U16432 (N_16432,N_15517,N_15779);
or U16433 (N_16433,N_15637,N_15958);
or U16434 (N_16434,N_15904,N_15793);
or U16435 (N_16435,N_15781,N_15579);
or U16436 (N_16436,N_15947,N_15953);
nand U16437 (N_16437,N_15724,N_15631);
nor U16438 (N_16438,N_15725,N_15545);
and U16439 (N_16439,N_15740,N_15874);
and U16440 (N_16440,N_15746,N_15560);
nor U16441 (N_16441,N_15637,N_15629);
and U16442 (N_16442,N_15901,N_15750);
nand U16443 (N_16443,N_15712,N_15936);
nand U16444 (N_16444,N_15895,N_15608);
nor U16445 (N_16445,N_15701,N_15858);
or U16446 (N_16446,N_15675,N_15899);
nor U16447 (N_16447,N_15544,N_15859);
and U16448 (N_16448,N_15524,N_15582);
xnor U16449 (N_16449,N_15575,N_15545);
xor U16450 (N_16450,N_15611,N_15865);
xor U16451 (N_16451,N_15916,N_15541);
or U16452 (N_16452,N_15679,N_15844);
nand U16453 (N_16453,N_15964,N_15815);
or U16454 (N_16454,N_15887,N_15929);
nor U16455 (N_16455,N_15908,N_15627);
or U16456 (N_16456,N_15514,N_15691);
xnor U16457 (N_16457,N_15772,N_15867);
xnor U16458 (N_16458,N_15589,N_15614);
or U16459 (N_16459,N_15972,N_15920);
and U16460 (N_16460,N_15507,N_15980);
or U16461 (N_16461,N_15515,N_15857);
and U16462 (N_16462,N_15598,N_15748);
nand U16463 (N_16463,N_15970,N_15841);
and U16464 (N_16464,N_15892,N_15652);
nor U16465 (N_16465,N_15753,N_15960);
nor U16466 (N_16466,N_15613,N_15547);
nand U16467 (N_16467,N_15687,N_15819);
or U16468 (N_16468,N_15784,N_15509);
or U16469 (N_16469,N_15653,N_15599);
xor U16470 (N_16470,N_15685,N_15811);
and U16471 (N_16471,N_15814,N_15730);
xnor U16472 (N_16472,N_15807,N_15503);
and U16473 (N_16473,N_15901,N_15764);
nor U16474 (N_16474,N_15809,N_15958);
nand U16475 (N_16475,N_15505,N_15562);
or U16476 (N_16476,N_15525,N_15503);
xor U16477 (N_16477,N_15507,N_15913);
nand U16478 (N_16478,N_15837,N_15783);
or U16479 (N_16479,N_15609,N_15519);
or U16480 (N_16480,N_15981,N_15644);
xnor U16481 (N_16481,N_15721,N_15738);
and U16482 (N_16482,N_15956,N_15559);
or U16483 (N_16483,N_15593,N_15717);
nand U16484 (N_16484,N_15766,N_15511);
and U16485 (N_16485,N_15629,N_15622);
and U16486 (N_16486,N_15697,N_15745);
nand U16487 (N_16487,N_15675,N_15590);
or U16488 (N_16488,N_15577,N_15592);
xor U16489 (N_16489,N_15557,N_15699);
and U16490 (N_16490,N_15851,N_15693);
nor U16491 (N_16491,N_15581,N_15751);
and U16492 (N_16492,N_15564,N_15873);
or U16493 (N_16493,N_15711,N_15647);
nand U16494 (N_16494,N_15745,N_15825);
nor U16495 (N_16495,N_15846,N_15731);
or U16496 (N_16496,N_15995,N_15857);
and U16497 (N_16497,N_15659,N_15645);
nand U16498 (N_16498,N_15938,N_15564);
and U16499 (N_16499,N_15781,N_15804);
nand U16500 (N_16500,N_16497,N_16102);
and U16501 (N_16501,N_16397,N_16007);
nand U16502 (N_16502,N_16110,N_16354);
nand U16503 (N_16503,N_16273,N_16100);
xor U16504 (N_16504,N_16186,N_16219);
or U16505 (N_16505,N_16068,N_16154);
nand U16506 (N_16506,N_16293,N_16173);
and U16507 (N_16507,N_16349,N_16369);
nor U16508 (N_16508,N_16194,N_16137);
xor U16509 (N_16509,N_16227,N_16367);
nor U16510 (N_16510,N_16198,N_16190);
xor U16511 (N_16511,N_16305,N_16380);
or U16512 (N_16512,N_16114,N_16343);
nor U16513 (N_16513,N_16237,N_16012);
nand U16514 (N_16514,N_16252,N_16001);
or U16515 (N_16515,N_16127,N_16083);
nor U16516 (N_16516,N_16040,N_16314);
and U16517 (N_16517,N_16213,N_16030);
nand U16518 (N_16518,N_16467,N_16357);
xor U16519 (N_16519,N_16148,N_16181);
or U16520 (N_16520,N_16346,N_16233);
nand U16521 (N_16521,N_16441,N_16429);
or U16522 (N_16522,N_16300,N_16447);
and U16523 (N_16523,N_16091,N_16368);
xor U16524 (N_16524,N_16076,N_16161);
nor U16525 (N_16525,N_16430,N_16182);
xor U16526 (N_16526,N_16200,N_16426);
nor U16527 (N_16527,N_16218,N_16432);
nor U16528 (N_16528,N_16440,N_16321);
or U16529 (N_16529,N_16010,N_16095);
xor U16530 (N_16530,N_16257,N_16224);
and U16531 (N_16531,N_16312,N_16371);
nand U16532 (N_16532,N_16490,N_16223);
nor U16533 (N_16533,N_16470,N_16058);
nor U16534 (N_16534,N_16342,N_16311);
nor U16535 (N_16535,N_16020,N_16494);
and U16536 (N_16536,N_16269,N_16096);
or U16537 (N_16537,N_16277,N_16128);
nor U16538 (N_16538,N_16370,N_16438);
nand U16539 (N_16539,N_16489,N_16319);
nor U16540 (N_16540,N_16139,N_16283);
and U16541 (N_16541,N_16225,N_16156);
nor U16542 (N_16542,N_16162,N_16138);
nand U16543 (N_16543,N_16451,N_16407);
nor U16544 (N_16544,N_16105,N_16459);
nand U16545 (N_16545,N_16492,N_16104);
or U16546 (N_16546,N_16013,N_16329);
and U16547 (N_16547,N_16498,N_16042);
nand U16548 (N_16548,N_16038,N_16392);
nor U16549 (N_16549,N_16315,N_16109);
nor U16550 (N_16550,N_16199,N_16016);
nor U16551 (N_16551,N_16092,N_16031);
and U16552 (N_16552,N_16131,N_16331);
xor U16553 (N_16553,N_16328,N_16405);
and U16554 (N_16554,N_16072,N_16398);
nor U16555 (N_16555,N_16056,N_16334);
or U16556 (N_16556,N_16340,N_16289);
nor U16557 (N_16557,N_16268,N_16290);
or U16558 (N_16558,N_16093,N_16485);
or U16559 (N_16559,N_16052,N_16070);
and U16560 (N_16560,N_16338,N_16453);
nand U16561 (N_16561,N_16140,N_16471);
or U16562 (N_16562,N_16081,N_16416);
nand U16563 (N_16563,N_16463,N_16055);
xor U16564 (N_16564,N_16390,N_16330);
xor U16565 (N_16565,N_16133,N_16496);
nand U16566 (N_16566,N_16421,N_16391);
and U16567 (N_16567,N_16420,N_16080);
nor U16568 (N_16568,N_16226,N_16043);
nor U16569 (N_16569,N_16255,N_16253);
nor U16570 (N_16570,N_16084,N_16067);
xor U16571 (N_16571,N_16065,N_16073);
xnor U16572 (N_16572,N_16413,N_16151);
nor U16573 (N_16573,N_16347,N_16077);
xnor U16574 (N_16574,N_16166,N_16216);
xor U16575 (N_16575,N_16172,N_16027);
nand U16576 (N_16576,N_16499,N_16383);
xnor U16577 (N_16577,N_16130,N_16442);
or U16578 (N_16578,N_16260,N_16431);
or U16579 (N_16579,N_16170,N_16240);
and U16580 (N_16580,N_16458,N_16248);
nand U16581 (N_16581,N_16404,N_16288);
nand U16582 (N_16582,N_16317,N_16215);
nor U16583 (N_16583,N_16477,N_16455);
nor U16584 (N_16584,N_16469,N_16393);
nand U16585 (N_16585,N_16386,N_16297);
and U16586 (N_16586,N_16122,N_16351);
or U16587 (N_16587,N_16473,N_16256);
or U16588 (N_16588,N_16158,N_16064);
nor U16589 (N_16589,N_16493,N_16488);
and U16590 (N_16590,N_16419,N_16387);
xor U16591 (N_16591,N_16448,N_16206);
nor U16592 (N_16592,N_16232,N_16359);
xnor U16593 (N_16593,N_16125,N_16023);
xor U16594 (N_16594,N_16450,N_16202);
xnor U16595 (N_16595,N_16119,N_16344);
xor U16596 (N_16596,N_16054,N_16204);
nor U16597 (N_16597,N_16082,N_16281);
or U16598 (N_16598,N_16401,N_16481);
nand U16599 (N_16599,N_16325,N_16059);
nand U16600 (N_16600,N_16002,N_16303);
nor U16601 (N_16601,N_16074,N_16090);
or U16602 (N_16602,N_16444,N_16307);
xor U16603 (N_16603,N_16231,N_16124);
and U16604 (N_16604,N_16478,N_16278);
xnor U16605 (N_16605,N_16341,N_16372);
nand U16606 (N_16606,N_16089,N_16376);
and U16607 (N_16607,N_16003,N_16417);
nor U16608 (N_16608,N_16408,N_16403);
and U16609 (N_16609,N_16318,N_16048);
nand U16610 (N_16610,N_16365,N_16388);
nor U16611 (N_16611,N_16142,N_16034);
xnor U16612 (N_16612,N_16456,N_16286);
or U16613 (N_16613,N_16466,N_16272);
or U16614 (N_16614,N_16045,N_16000);
and U16615 (N_16615,N_16422,N_16250);
nor U16616 (N_16616,N_16189,N_16275);
nand U16617 (N_16617,N_16465,N_16150);
nor U16618 (N_16618,N_16239,N_16057);
or U16619 (N_16619,N_16299,N_16284);
xnor U16620 (N_16620,N_16157,N_16350);
and U16621 (N_16621,N_16220,N_16254);
nand U16622 (N_16622,N_16411,N_16271);
and U16623 (N_16623,N_16460,N_16247);
nor U16624 (N_16624,N_16362,N_16461);
xor U16625 (N_16625,N_16021,N_16004);
xor U16626 (N_16626,N_16209,N_16373);
and U16627 (N_16627,N_16258,N_16212);
and U16628 (N_16628,N_16207,N_16160);
nand U16629 (N_16629,N_16101,N_16332);
xnor U16630 (N_16630,N_16075,N_16475);
and U16631 (N_16631,N_16014,N_16452);
nor U16632 (N_16632,N_16188,N_16306);
xnor U16633 (N_16633,N_16366,N_16111);
nand U16634 (N_16634,N_16264,N_16482);
and U16635 (N_16635,N_16434,N_16472);
or U16636 (N_16636,N_16267,N_16241);
nand U16637 (N_16637,N_16017,N_16484);
nand U16638 (N_16638,N_16406,N_16136);
or U16639 (N_16639,N_16086,N_16015);
or U16640 (N_16640,N_16062,N_16320);
xor U16641 (N_16641,N_16063,N_16282);
nor U16642 (N_16642,N_16418,N_16396);
nor U16643 (N_16643,N_16230,N_16153);
or U16644 (N_16644,N_16295,N_16165);
or U16645 (N_16645,N_16108,N_16191);
xnor U16646 (N_16646,N_16279,N_16029);
and U16647 (N_16647,N_16134,N_16280);
or U16648 (N_16648,N_16381,N_16050);
nand U16649 (N_16649,N_16480,N_16353);
nor U16650 (N_16650,N_16266,N_16302);
nor U16651 (N_16651,N_16487,N_16292);
or U16652 (N_16652,N_16177,N_16339);
and U16653 (N_16653,N_16155,N_16201);
xor U16654 (N_16654,N_16246,N_16261);
xor U16655 (N_16655,N_16176,N_16146);
and U16656 (N_16656,N_16423,N_16385);
and U16657 (N_16657,N_16025,N_16159);
nor U16658 (N_16658,N_16106,N_16457);
nand U16659 (N_16659,N_16022,N_16169);
nor U16660 (N_16660,N_16309,N_16141);
nor U16661 (N_16661,N_16298,N_16287);
or U16662 (N_16662,N_16454,N_16196);
nor U16663 (N_16663,N_16363,N_16116);
and U16664 (N_16664,N_16024,N_16235);
xnor U16665 (N_16665,N_16236,N_16414);
and U16666 (N_16666,N_16301,N_16143);
xnor U16667 (N_16667,N_16193,N_16439);
nand U16668 (N_16668,N_16011,N_16449);
or U16669 (N_16669,N_16039,N_16129);
and U16670 (N_16670,N_16427,N_16026);
or U16671 (N_16671,N_16049,N_16375);
nand U16672 (N_16672,N_16117,N_16356);
xor U16673 (N_16673,N_16433,N_16384);
and U16674 (N_16674,N_16036,N_16037);
xnor U16675 (N_16675,N_16121,N_16395);
or U16676 (N_16676,N_16164,N_16047);
xnor U16677 (N_16677,N_16006,N_16175);
nor U16678 (N_16678,N_16364,N_16333);
nand U16679 (N_16679,N_16483,N_16476);
or U16680 (N_16680,N_16069,N_16337);
nor U16681 (N_16681,N_16087,N_16060);
xnor U16682 (N_16682,N_16326,N_16210);
xnor U16683 (N_16683,N_16400,N_16079);
or U16684 (N_16684,N_16491,N_16327);
nor U16685 (N_16685,N_16358,N_16234);
or U16686 (N_16686,N_16051,N_16251);
xnor U16687 (N_16687,N_16208,N_16098);
nor U16688 (N_16688,N_16308,N_16409);
and U16689 (N_16689,N_16115,N_16028);
nand U16690 (N_16690,N_16053,N_16008);
nor U16691 (N_16691,N_16265,N_16399);
xnor U16692 (N_16692,N_16377,N_16018);
and U16693 (N_16693,N_16468,N_16378);
nor U16694 (N_16694,N_16228,N_16382);
nor U16695 (N_16695,N_16291,N_16323);
xnor U16696 (N_16696,N_16183,N_16032);
xnor U16697 (N_16697,N_16379,N_16249);
and U16698 (N_16698,N_16195,N_16044);
nor U16699 (N_16699,N_16187,N_16238);
or U16700 (N_16700,N_16135,N_16035);
nor U16701 (N_16701,N_16197,N_16163);
nor U16702 (N_16702,N_16041,N_16088);
nand U16703 (N_16703,N_16099,N_16174);
or U16704 (N_16704,N_16214,N_16046);
nor U16705 (N_16705,N_16263,N_16242);
nand U16706 (N_16706,N_16474,N_16243);
nor U16707 (N_16707,N_16126,N_16322);
nand U16708 (N_16708,N_16412,N_16374);
nand U16709 (N_16709,N_16147,N_16360);
nor U16710 (N_16710,N_16066,N_16178);
nand U16711 (N_16711,N_16294,N_16203);
or U16712 (N_16712,N_16345,N_16118);
nor U16713 (N_16713,N_16336,N_16410);
or U16714 (N_16714,N_16424,N_16120);
or U16715 (N_16715,N_16192,N_16184);
xor U16716 (N_16716,N_16149,N_16316);
and U16717 (N_16717,N_16436,N_16276);
nor U16718 (N_16718,N_16078,N_16486);
nand U16719 (N_16719,N_16352,N_16107);
and U16720 (N_16720,N_16103,N_16179);
nand U16721 (N_16721,N_16221,N_16145);
nand U16722 (N_16722,N_16185,N_16168);
or U16723 (N_16723,N_16324,N_16152);
nor U16724 (N_16724,N_16304,N_16259);
or U16725 (N_16725,N_16097,N_16171);
and U16726 (N_16726,N_16245,N_16085);
nor U16727 (N_16727,N_16019,N_16389);
and U16728 (N_16728,N_16123,N_16402);
nand U16729 (N_16729,N_16445,N_16094);
nor U16730 (N_16730,N_16005,N_16113);
nand U16731 (N_16731,N_16009,N_16313);
nor U16732 (N_16732,N_16361,N_16211);
nor U16733 (N_16733,N_16180,N_16435);
nor U16734 (N_16734,N_16167,N_16112);
nor U16735 (N_16735,N_16296,N_16415);
and U16736 (N_16736,N_16479,N_16132);
or U16737 (N_16737,N_16443,N_16310);
xor U16738 (N_16738,N_16335,N_16205);
xnor U16739 (N_16739,N_16285,N_16394);
and U16740 (N_16740,N_16446,N_16061);
or U16741 (N_16741,N_16462,N_16222);
xnor U16742 (N_16742,N_16495,N_16428);
xor U16743 (N_16743,N_16348,N_16274);
xor U16744 (N_16744,N_16425,N_16262);
nand U16745 (N_16745,N_16144,N_16270);
xor U16746 (N_16746,N_16355,N_16244);
nand U16747 (N_16747,N_16033,N_16071);
and U16748 (N_16748,N_16229,N_16437);
xnor U16749 (N_16749,N_16217,N_16464);
nand U16750 (N_16750,N_16114,N_16035);
or U16751 (N_16751,N_16423,N_16207);
nand U16752 (N_16752,N_16105,N_16194);
nor U16753 (N_16753,N_16260,N_16103);
and U16754 (N_16754,N_16167,N_16422);
and U16755 (N_16755,N_16244,N_16434);
or U16756 (N_16756,N_16315,N_16067);
nand U16757 (N_16757,N_16292,N_16140);
or U16758 (N_16758,N_16051,N_16165);
nand U16759 (N_16759,N_16348,N_16393);
xnor U16760 (N_16760,N_16432,N_16359);
nand U16761 (N_16761,N_16283,N_16392);
and U16762 (N_16762,N_16045,N_16258);
or U16763 (N_16763,N_16416,N_16073);
nor U16764 (N_16764,N_16128,N_16255);
and U16765 (N_16765,N_16156,N_16323);
and U16766 (N_16766,N_16366,N_16346);
and U16767 (N_16767,N_16309,N_16051);
or U16768 (N_16768,N_16458,N_16328);
nand U16769 (N_16769,N_16388,N_16042);
nor U16770 (N_16770,N_16179,N_16049);
nor U16771 (N_16771,N_16009,N_16459);
or U16772 (N_16772,N_16438,N_16195);
and U16773 (N_16773,N_16124,N_16200);
or U16774 (N_16774,N_16127,N_16206);
or U16775 (N_16775,N_16067,N_16072);
nand U16776 (N_16776,N_16068,N_16273);
nor U16777 (N_16777,N_16225,N_16381);
nand U16778 (N_16778,N_16095,N_16042);
nand U16779 (N_16779,N_16409,N_16264);
nor U16780 (N_16780,N_16385,N_16356);
or U16781 (N_16781,N_16451,N_16008);
xnor U16782 (N_16782,N_16000,N_16123);
nor U16783 (N_16783,N_16058,N_16416);
nor U16784 (N_16784,N_16471,N_16005);
xnor U16785 (N_16785,N_16328,N_16106);
or U16786 (N_16786,N_16227,N_16261);
xor U16787 (N_16787,N_16374,N_16125);
xor U16788 (N_16788,N_16169,N_16463);
xor U16789 (N_16789,N_16243,N_16089);
nor U16790 (N_16790,N_16080,N_16371);
xnor U16791 (N_16791,N_16026,N_16044);
and U16792 (N_16792,N_16150,N_16059);
and U16793 (N_16793,N_16127,N_16147);
nand U16794 (N_16794,N_16154,N_16394);
or U16795 (N_16795,N_16224,N_16000);
xor U16796 (N_16796,N_16194,N_16444);
nand U16797 (N_16797,N_16176,N_16160);
and U16798 (N_16798,N_16285,N_16220);
xnor U16799 (N_16799,N_16352,N_16465);
xnor U16800 (N_16800,N_16396,N_16444);
xnor U16801 (N_16801,N_16044,N_16133);
and U16802 (N_16802,N_16172,N_16018);
or U16803 (N_16803,N_16129,N_16419);
nor U16804 (N_16804,N_16372,N_16302);
and U16805 (N_16805,N_16250,N_16212);
nor U16806 (N_16806,N_16369,N_16375);
xnor U16807 (N_16807,N_16330,N_16425);
nand U16808 (N_16808,N_16124,N_16300);
xnor U16809 (N_16809,N_16111,N_16358);
nor U16810 (N_16810,N_16240,N_16348);
xnor U16811 (N_16811,N_16210,N_16382);
xnor U16812 (N_16812,N_16457,N_16291);
nand U16813 (N_16813,N_16256,N_16207);
nand U16814 (N_16814,N_16178,N_16455);
nor U16815 (N_16815,N_16274,N_16375);
xor U16816 (N_16816,N_16145,N_16236);
xnor U16817 (N_16817,N_16021,N_16070);
or U16818 (N_16818,N_16430,N_16483);
nor U16819 (N_16819,N_16110,N_16419);
and U16820 (N_16820,N_16107,N_16345);
or U16821 (N_16821,N_16100,N_16089);
or U16822 (N_16822,N_16045,N_16222);
xor U16823 (N_16823,N_16132,N_16421);
or U16824 (N_16824,N_16313,N_16368);
nor U16825 (N_16825,N_16135,N_16421);
nor U16826 (N_16826,N_16300,N_16091);
xor U16827 (N_16827,N_16010,N_16190);
nand U16828 (N_16828,N_16221,N_16007);
nand U16829 (N_16829,N_16105,N_16482);
nand U16830 (N_16830,N_16108,N_16315);
or U16831 (N_16831,N_16484,N_16121);
nand U16832 (N_16832,N_16487,N_16009);
or U16833 (N_16833,N_16340,N_16002);
or U16834 (N_16834,N_16169,N_16110);
nor U16835 (N_16835,N_16491,N_16325);
nand U16836 (N_16836,N_16141,N_16028);
nand U16837 (N_16837,N_16087,N_16055);
and U16838 (N_16838,N_16279,N_16130);
nor U16839 (N_16839,N_16215,N_16461);
nor U16840 (N_16840,N_16326,N_16360);
nor U16841 (N_16841,N_16494,N_16443);
xnor U16842 (N_16842,N_16337,N_16312);
or U16843 (N_16843,N_16465,N_16231);
nor U16844 (N_16844,N_16394,N_16489);
nand U16845 (N_16845,N_16377,N_16232);
nor U16846 (N_16846,N_16309,N_16120);
nor U16847 (N_16847,N_16216,N_16109);
nand U16848 (N_16848,N_16003,N_16284);
and U16849 (N_16849,N_16355,N_16120);
and U16850 (N_16850,N_16310,N_16394);
or U16851 (N_16851,N_16258,N_16149);
or U16852 (N_16852,N_16240,N_16105);
nor U16853 (N_16853,N_16208,N_16459);
or U16854 (N_16854,N_16165,N_16344);
xnor U16855 (N_16855,N_16363,N_16247);
or U16856 (N_16856,N_16353,N_16497);
nor U16857 (N_16857,N_16126,N_16018);
xor U16858 (N_16858,N_16488,N_16331);
nor U16859 (N_16859,N_16086,N_16117);
nor U16860 (N_16860,N_16340,N_16324);
nand U16861 (N_16861,N_16328,N_16065);
xnor U16862 (N_16862,N_16445,N_16427);
xnor U16863 (N_16863,N_16416,N_16141);
xnor U16864 (N_16864,N_16185,N_16183);
or U16865 (N_16865,N_16178,N_16132);
nor U16866 (N_16866,N_16343,N_16249);
and U16867 (N_16867,N_16441,N_16332);
and U16868 (N_16868,N_16320,N_16061);
nor U16869 (N_16869,N_16100,N_16458);
xnor U16870 (N_16870,N_16453,N_16216);
xor U16871 (N_16871,N_16053,N_16421);
nand U16872 (N_16872,N_16154,N_16323);
nand U16873 (N_16873,N_16103,N_16466);
xnor U16874 (N_16874,N_16283,N_16091);
nor U16875 (N_16875,N_16258,N_16286);
and U16876 (N_16876,N_16298,N_16490);
and U16877 (N_16877,N_16248,N_16097);
or U16878 (N_16878,N_16233,N_16487);
and U16879 (N_16879,N_16064,N_16033);
nor U16880 (N_16880,N_16151,N_16245);
xnor U16881 (N_16881,N_16395,N_16431);
or U16882 (N_16882,N_16257,N_16351);
nand U16883 (N_16883,N_16308,N_16085);
xor U16884 (N_16884,N_16264,N_16128);
nor U16885 (N_16885,N_16359,N_16327);
nor U16886 (N_16886,N_16288,N_16344);
nand U16887 (N_16887,N_16258,N_16422);
nor U16888 (N_16888,N_16113,N_16468);
xnor U16889 (N_16889,N_16392,N_16126);
nand U16890 (N_16890,N_16031,N_16368);
and U16891 (N_16891,N_16487,N_16464);
nand U16892 (N_16892,N_16219,N_16343);
nor U16893 (N_16893,N_16191,N_16137);
xnor U16894 (N_16894,N_16096,N_16384);
or U16895 (N_16895,N_16165,N_16316);
or U16896 (N_16896,N_16241,N_16380);
nand U16897 (N_16897,N_16135,N_16063);
nand U16898 (N_16898,N_16370,N_16409);
or U16899 (N_16899,N_16310,N_16081);
xnor U16900 (N_16900,N_16305,N_16451);
nor U16901 (N_16901,N_16079,N_16491);
and U16902 (N_16902,N_16149,N_16253);
nand U16903 (N_16903,N_16205,N_16109);
nor U16904 (N_16904,N_16033,N_16010);
nor U16905 (N_16905,N_16489,N_16186);
xor U16906 (N_16906,N_16255,N_16085);
and U16907 (N_16907,N_16060,N_16022);
or U16908 (N_16908,N_16499,N_16033);
and U16909 (N_16909,N_16063,N_16209);
nand U16910 (N_16910,N_16230,N_16324);
or U16911 (N_16911,N_16300,N_16339);
or U16912 (N_16912,N_16194,N_16300);
nor U16913 (N_16913,N_16004,N_16236);
xnor U16914 (N_16914,N_16158,N_16357);
nand U16915 (N_16915,N_16160,N_16416);
nor U16916 (N_16916,N_16108,N_16216);
nor U16917 (N_16917,N_16350,N_16231);
or U16918 (N_16918,N_16210,N_16463);
xnor U16919 (N_16919,N_16492,N_16076);
nand U16920 (N_16920,N_16470,N_16337);
nand U16921 (N_16921,N_16097,N_16096);
nand U16922 (N_16922,N_16270,N_16406);
and U16923 (N_16923,N_16004,N_16417);
and U16924 (N_16924,N_16238,N_16437);
nor U16925 (N_16925,N_16138,N_16337);
or U16926 (N_16926,N_16359,N_16219);
xnor U16927 (N_16927,N_16241,N_16204);
nand U16928 (N_16928,N_16453,N_16267);
nand U16929 (N_16929,N_16168,N_16430);
or U16930 (N_16930,N_16160,N_16340);
and U16931 (N_16931,N_16443,N_16472);
and U16932 (N_16932,N_16036,N_16058);
and U16933 (N_16933,N_16322,N_16475);
and U16934 (N_16934,N_16473,N_16293);
or U16935 (N_16935,N_16494,N_16099);
nor U16936 (N_16936,N_16056,N_16276);
nor U16937 (N_16937,N_16150,N_16475);
xnor U16938 (N_16938,N_16448,N_16060);
and U16939 (N_16939,N_16338,N_16022);
and U16940 (N_16940,N_16276,N_16103);
and U16941 (N_16941,N_16194,N_16067);
nand U16942 (N_16942,N_16455,N_16302);
xnor U16943 (N_16943,N_16326,N_16351);
xor U16944 (N_16944,N_16272,N_16219);
nand U16945 (N_16945,N_16269,N_16199);
or U16946 (N_16946,N_16165,N_16169);
or U16947 (N_16947,N_16247,N_16359);
nand U16948 (N_16948,N_16281,N_16151);
nor U16949 (N_16949,N_16027,N_16012);
nand U16950 (N_16950,N_16113,N_16081);
nand U16951 (N_16951,N_16176,N_16200);
nand U16952 (N_16952,N_16175,N_16377);
or U16953 (N_16953,N_16240,N_16013);
and U16954 (N_16954,N_16330,N_16417);
xor U16955 (N_16955,N_16182,N_16482);
or U16956 (N_16956,N_16093,N_16425);
and U16957 (N_16957,N_16050,N_16098);
nor U16958 (N_16958,N_16273,N_16381);
and U16959 (N_16959,N_16018,N_16088);
nor U16960 (N_16960,N_16115,N_16037);
nand U16961 (N_16961,N_16423,N_16420);
nor U16962 (N_16962,N_16406,N_16380);
nor U16963 (N_16963,N_16104,N_16131);
and U16964 (N_16964,N_16272,N_16460);
or U16965 (N_16965,N_16078,N_16101);
or U16966 (N_16966,N_16497,N_16234);
or U16967 (N_16967,N_16330,N_16331);
or U16968 (N_16968,N_16373,N_16449);
or U16969 (N_16969,N_16331,N_16059);
nand U16970 (N_16970,N_16261,N_16126);
xnor U16971 (N_16971,N_16394,N_16053);
and U16972 (N_16972,N_16021,N_16213);
nand U16973 (N_16973,N_16298,N_16293);
and U16974 (N_16974,N_16388,N_16273);
nor U16975 (N_16975,N_16376,N_16470);
nor U16976 (N_16976,N_16130,N_16033);
nor U16977 (N_16977,N_16003,N_16242);
and U16978 (N_16978,N_16441,N_16350);
nand U16979 (N_16979,N_16481,N_16255);
nor U16980 (N_16980,N_16371,N_16483);
xor U16981 (N_16981,N_16426,N_16119);
nor U16982 (N_16982,N_16266,N_16166);
and U16983 (N_16983,N_16062,N_16167);
and U16984 (N_16984,N_16116,N_16465);
or U16985 (N_16985,N_16148,N_16092);
and U16986 (N_16986,N_16397,N_16330);
or U16987 (N_16987,N_16005,N_16128);
xnor U16988 (N_16988,N_16410,N_16469);
and U16989 (N_16989,N_16047,N_16027);
xor U16990 (N_16990,N_16095,N_16406);
or U16991 (N_16991,N_16206,N_16401);
and U16992 (N_16992,N_16465,N_16232);
nor U16993 (N_16993,N_16328,N_16427);
nand U16994 (N_16994,N_16241,N_16432);
nand U16995 (N_16995,N_16199,N_16352);
xnor U16996 (N_16996,N_16007,N_16429);
nand U16997 (N_16997,N_16098,N_16370);
and U16998 (N_16998,N_16279,N_16252);
nand U16999 (N_16999,N_16192,N_16194);
xnor U17000 (N_17000,N_16680,N_16844);
and U17001 (N_17001,N_16622,N_16849);
nand U17002 (N_17002,N_16576,N_16878);
nor U17003 (N_17003,N_16563,N_16547);
and U17004 (N_17004,N_16664,N_16609);
xor U17005 (N_17005,N_16774,N_16917);
and U17006 (N_17006,N_16566,N_16720);
or U17007 (N_17007,N_16630,N_16751);
or U17008 (N_17008,N_16772,N_16733);
and U17009 (N_17009,N_16560,N_16520);
nand U17010 (N_17010,N_16946,N_16667);
or U17011 (N_17011,N_16603,N_16512);
or U17012 (N_17012,N_16781,N_16871);
nor U17013 (N_17013,N_16658,N_16921);
nor U17014 (N_17014,N_16662,N_16588);
or U17015 (N_17015,N_16968,N_16901);
xor U17016 (N_17016,N_16596,N_16942);
nor U17017 (N_17017,N_16550,N_16686);
xor U17018 (N_17018,N_16952,N_16863);
xnor U17019 (N_17019,N_16979,N_16809);
nand U17020 (N_17020,N_16734,N_16816);
xor U17021 (N_17021,N_16557,N_16530);
nor U17022 (N_17022,N_16922,N_16915);
nand U17023 (N_17023,N_16782,N_16639);
and U17024 (N_17024,N_16534,N_16780);
or U17025 (N_17025,N_16848,N_16999);
xor U17026 (N_17026,N_16784,N_16766);
nor U17027 (N_17027,N_16691,N_16870);
nand U17028 (N_17028,N_16607,N_16793);
nand U17029 (N_17029,N_16642,N_16974);
or U17030 (N_17030,N_16841,N_16684);
nand U17031 (N_17031,N_16626,N_16567);
and U17032 (N_17032,N_16593,N_16888);
and U17033 (N_17033,N_16825,N_16874);
nor U17034 (N_17034,N_16770,N_16624);
and U17035 (N_17035,N_16821,N_16722);
nand U17036 (N_17036,N_16589,N_16716);
nor U17037 (N_17037,N_16523,N_16597);
and U17038 (N_17038,N_16723,N_16862);
or U17039 (N_17039,N_16677,N_16598);
or U17040 (N_17040,N_16570,N_16838);
or U17041 (N_17041,N_16806,N_16859);
and U17042 (N_17042,N_16898,N_16865);
nor U17043 (N_17043,N_16846,N_16771);
or U17044 (N_17044,N_16978,N_16561);
nor U17045 (N_17045,N_16889,N_16619);
xor U17046 (N_17046,N_16829,N_16867);
nor U17047 (N_17047,N_16736,N_16507);
nand U17048 (N_17048,N_16617,N_16540);
and U17049 (N_17049,N_16916,N_16702);
and U17050 (N_17050,N_16805,N_16564);
and U17051 (N_17051,N_16725,N_16698);
nand U17052 (N_17052,N_16590,N_16535);
or U17053 (N_17053,N_16852,N_16818);
and U17054 (N_17054,N_16511,N_16730);
or U17055 (N_17055,N_16802,N_16890);
or U17056 (N_17056,N_16541,N_16940);
and U17057 (N_17057,N_16553,N_16824);
or U17058 (N_17058,N_16972,N_16532);
nor U17059 (N_17059,N_16971,N_16537);
nor U17060 (N_17060,N_16502,N_16804);
and U17061 (N_17061,N_16504,N_16708);
nor U17062 (N_17062,N_16600,N_16932);
and U17063 (N_17063,N_16599,N_16615);
nor U17064 (N_17064,N_16646,N_16672);
nor U17065 (N_17065,N_16761,N_16735);
or U17066 (N_17066,N_16914,N_16980);
or U17067 (N_17067,N_16709,N_16912);
or U17068 (N_17068,N_16933,N_16713);
or U17069 (N_17069,N_16941,N_16591);
and U17070 (N_17070,N_16650,N_16703);
xnor U17071 (N_17071,N_16500,N_16954);
or U17072 (N_17072,N_16756,N_16582);
and U17073 (N_17073,N_16970,N_16690);
nand U17074 (N_17074,N_16528,N_16652);
nand U17075 (N_17075,N_16649,N_16827);
or U17076 (N_17076,N_16855,N_16538);
nand U17077 (N_17077,N_16585,N_16645);
nand U17078 (N_17078,N_16551,N_16747);
nand U17079 (N_17079,N_16765,N_16939);
nand U17080 (N_17080,N_16629,N_16812);
xnor U17081 (N_17081,N_16868,N_16976);
nor U17082 (N_17082,N_16657,N_16760);
nand U17083 (N_17083,N_16907,N_16727);
nor U17084 (N_17084,N_16834,N_16910);
and U17085 (N_17085,N_16923,N_16938);
nor U17086 (N_17086,N_16605,N_16688);
and U17087 (N_17087,N_16982,N_16671);
xor U17088 (N_17088,N_16886,N_16611);
and U17089 (N_17089,N_16643,N_16826);
nor U17090 (N_17090,N_16957,N_16799);
and U17091 (N_17091,N_16842,N_16505);
xnor U17092 (N_17092,N_16847,N_16572);
and U17093 (N_17093,N_16704,N_16992);
and U17094 (N_17094,N_16899,N_16666);
and U17095 (N_17095,N_16819,N_16944);
and U17096 (N_17096,N_16683,N_16800);
nor U17097 (N_17097,N_16858,N_16696);
or U17098 (N_17098,N_16632,N_16955);
xnor U17099 (N_17099,N_16724,N_16920);
and U17100 (N_17100,N_16911,N_16715);
nand U17101 (N_17101,N_16518,N_16533);
nand U17102 (N_17102,N_16909,N_16641);
or U17103 (N_17103,N_16902,N_16988);
nand U17104 (N_17104,N_16559,N_16851);
and U17105 (N_17105,N_16803,N_16794);
or U17106 (N_17106,N_16545,N_16718);
nand U17107 (N_17107,N_16757,N_16670);
xnor U17108 (N_17108,N_16668,N_16750);
xor U17109 (N_17109,N_16953,N_16549);
nand U17110 (N_17110,N_16685,N_16763);
and U17111 (N_17111,N_16701,N_16861);
and U17112 (N_17112,N_16789,N_16711);
nand U17113 (N_17113,N_16513,N_16675);
nor U17114 (N_17114,N_16748,N_16885);
nor U17115 (N_17115,N_16991,N_16694);
and U17116 (N_17116,N_16602,N_16854);
or U17117 (N_17117,N_16501,N_16737);
nor U17118 (N_17118,N_16879,N_16714);
xnor U17119 (N_17119,N_16787,N_16973);
or U17120 (N_17120,N_16571,N_16962);
nand U17121 (N_17121,N_16539,N_16797);
xor U17122 (N_17122,N_16673,N_16731);
or U17123 (N_17123,N_16997,N_16776);
xnor U17124 (N_17124,N_16845,N_16759);
nor U17125 (N_17125,N_16665,N_16964);
xnor U17126 (N_17126,N_16604,N_16949);
or U17127 (N_17127,N_16618,N_16790);
or U17128 (N_17128,N_16613,N_16935);
nand U17129 (N_17129,N_16904,N_16903);
nor U17130 (N_17130,N_16753,N_16929);
or U17131 (N_17131,N_16791,N_16891);
nor U17132 (N_17132,N_16801,N_16638);
nor U17133 (N_17133,N_16882,N_16739);
xor U17134 (N_17134,N_16595,N_16965);
nand U17135 (N_17135,N_16850,N_16640);
nand U17136 (N_17136,N_16936,N_16745);
nand U17137 (N_17137,N_16584,N_16798);
and U17138 (N_17138,N_16749,N_16699);
and U17139 (N_17139,N_16627,N_16987);
and U17140 (N_17140,N_16764,N_16788);
xnor U17141 (N_17141,N_16633,N_16975);
or U17142 (N_17142,N_16959,N_16743);
nand U17143 (N_17143,N_16707,N_16837);
and U17144 (N_17144,N_16578,N_16526);
nand U17145 (N_17145,N_16919,N_16860);
nand U17146 (N_17146,N_16514,N_16918);
nor U17147 (N_17147,N_16913,N_16682);
or U17148 (N_17148,N_16755,N_16767);
and U17149 (N_17149,N_16994,N_16881);
nor U17150 (N_17150,N_16958,N_16637);
or U17151 (N_17151,N_16543,N_16710);
and U17152 (N_17152,N_16717,N_16778);
nor U17153 (N_17153,N_16663,N_16884);
and U17154 (N_17154,N_16529,N_16981);
or U17155 (N_17155,N_16527,N_16823);
or U17156 (N_17156,N_16620,N_16857);
nor U17157 (N_17157,N_16986,N_16897);
or U17158 (N_17158,N_16839,N_16687);
xnor U17159 (N_17159,N_16754,N_16831);
nand U17160 (N_17160,N_16956,N_16947);
xor U17161 (N_17161,N_16817,N_16610);
or U17162 (N_17162,N_16542,N_16741);
and U17163 (N_17163,N_16647,N_16606);
nor U17164 (N_17164,N_16746,N_16833);
xnor U17165 (N_17165,N_16531,N_16556);
nor U17166 (N_17166,N_16517,N_16693);
nor U17167 (N_17167,N_16906,N_16524);
xor U17168 (N_17168,N_16655,N_16586);
or U17169 (N_17169,N_16659,N_16644);
nand U17170 (N_17170,N_16628,N_16742);
xor U17171 (N_17171,N_16726,N_16963);
and U17172 (N_17172,N_16651,N_16840);
and U17173 (N_17173,N_16807,N_16777);
and U17174 (N_17174,N_16892,N_16503);
nor U17175 (N_17175,N_16653,N_16587);
nor U17176 (N_17176,N_16961,N_16575);
nor U17177 (N_17177,N_16506,N_16546);
nand U17178 (N_17178,N_16810,N_16625);
xnor U17179 (N_17179,N_16796,N_16728);
xnor U17180 (N_17180,N_16934,N_16924);
or U17181 (N_17181,N_16752,N_16508);
or U17182 (N_17182,N_16631,N_16768);
or U17183 (N_17183,N_16623,N_16573);
nand U17184 (N_17184,N_16516,N_16555);
xnor U17185 (N_17185,N_16950,N_16983);
nand U17186 (N_17186,N_16880,N_16565);
and U17187 (N_17187,N_16744,N_16943);
xor U17188 (N_17188,N_16905,N_16601);
and U17189 (N_17189,N_16783,N_16592);
xnor U17190 (N_17190,N_16522,N_16896);
and U17191 (N_17191,N_16552,N_16872);
and U17192 (N_17192,N_16729,N_16873);
nor U17193 (N_17193,N_16996,N_16681);
xor U17194 (N_17194,N_16678,N_16967);
xor U17195 (N_17195,N_16758,N_16822);
xor U17196 (N_17196,N_16843,N_16893);
or U17197 (N_17197,N_16554,N_16875);
and U17198 (N_17198,N_16985,N_16654);
and U17199 (N_17199,N_16762,N_16738);
xnor U17200 (N_17200,N_16815,N_16926);
and U17201 (N_17201,N_16521,N_16580);
and U17202 (N_17202,N_16908,N_16960);
xor U17203 (N_17203,N_16695,N_16519);
and U17204 (N_17204,N_16989,N_16864);
and U17205 (N_17205,N_16856,N_16656);
nor U17206 (N_17206,N_16562,N_16674);
or U17207 (N_17207,N_16995,N_16877);
or U17208 (N_17208,N_16883,N_16808);
and U17209 (N_17209,N_16697,N_16583);
nor U17210 (N_17210,N_16568,N_16689);
nand U17211 (N_17211,N_16928,N_16636);
and U17212 (N_17212,N_16869,N_16515);
xor U17213 (N_17213,N_16993,N_16779);
and U17214 (N_17214,N_16925,N_16577);
nand U17215 (N_17215,N_16525,N_16990);
and U17216 (N_17216,N_16951,N_16594);
or U17217 (N_17217,N_16574,N_16814);
nor U17218 (N_17218,N_16692,N_16634);
and U17219 (N_17219,N_16706,N_16966);
xor U17220 (N_17220,N_16785,N_16931);
or U17221 (N_17221,N_16969,N_16828);
and U17222 (N_17222,N_16635,N_16558);
or U17223 (N_17223,N_16719,N_16866);
or U17224 (N_17224,N_16740,N_16876);
and U17225 (N_17225,N_16661,N_16830);
or U17226 (N_17226,N_16579,N_16614);
nand U17227 (N_17227,N_16887,N_16569);
xnor U17228 (N_17228,N_16648,N_16853);
xor U17229 (N_17229,N_16930,N_16732);
nand U17230 (N_17230,N_16548,N_16544);
xor U17231 (N_17231,N_16811,N_16937);
nand U17232 (N_17232,N_16612,N_16832);
nor U17233 (N_17233,N_16792,N_16769);
nor U17234 (N_17234,N_16669,N_16894);
xnor U17235 (N_17235,N_16895,N_16660);
nor U17236 (N_17236,N_16820,N_16509);
or U17237 (N_17237,N_16536,N_16998);
or U17238 (N_17238,N_16948,N_16795);
xnor U17239 (N_17239,N_16945,N_16984);
or U17240 (N_17240,N_16581,N_16836);
nor U17241 (N_17241,N_16608,N_16773);
and U17242 (N_17242,N_16676,N_16712);
or U17243 (N_17243,N_16621,N_16927);
xnor U17244 (N_17244,N_16616,N_16835);
nand U17245 (N_17245,N_16510,N_16775);
nand U17246 (N_17246,N_16679,N_16700);
nand U17247 (N_17247,N_16786,N_16705);
and U17248 (N_17248,N_16977,N_16900);
or U17249 (N_17249,N_16721,N_16813);
and U17250 (N_17250,N_16570,N_16844);
xnor U17251 (N_17251,N_16521,N_16770);
nand U17252 (N_17252,N_16880,N_16806);
or U17253 (N_17253,N_16549,N_16902);
and U17254 (N_17254,N_16640,N_16751);
and U17255 (N_17255,N_16996,N_16563);
nor U17256 (N_17256,N_16867,N_16516);
or U17257 (N_17257,N_16808,N_16615);
nand U17258 (N_17258,N_16511,N_16543);
nand U17259 (N_17259,N_16817,N_16696);
xor U17260 (N_17260,N_16560,N_16744);
xnor U17261 (N_17261,N_16667,N_16541);
nand U17262 (N_17262,N_16731,N_16997);
nand U17263 (N_17263,N_16855,N_16764);
or U17264 (N_17264,N_16893,N_16605);
nor U17265 (N_17265,N_16963,N_16921);
and U17266 (N_17266,N_16700,N_16535);
and U17267 (N_17267,N_16598,N_16951);
nand U17268 (N_17268,N_16559,N_16993);
nand U17269 (N_17269,N_16911,N_16708);
and U17270 (N_17270,N_16733,N_16759);
nand U17271 (N_17271,N_16858,N_16584);
or U17272 (N_17272,N_16948,N_16982);
and U17273 (N_17273,N_16639,N_16775);
xor U17274 (N_17274,N_16600,N_16820);
or U17275 (N_17275,N_16690,N_16953);
xnor U17276 (N_17276,N_16748,N_16916);
nor U17277 (N_17277,N_16917,N_16857);
and U17278 (N_17278,N_16524,N_16722);
nand U17279 (N_17279,N_16643,N_16982);
xor U17280 (N_17280,N_16922,N_16575);
xor U17281 (N_17281,N_16578,N_16891);
nand U17282 (N_17282,N_16563,N_16716);
xnor U17283 (N_17283,N_16644,N_16554);
or U17284 (N_17284,N_16914,N_16664);
nand U17285 (N_17285,N_16607,N_16871);
xnor U17286 (N_17286,N_16907,N_16536);
xnor U17287 (N_17287,N_16849,N_16558);
nor U17288 (N_17288,N_16867,N_16624);
nor U17289 (N_17289,N_16899,N_16776);
nor U17290 (N_17290,N_16685,N_16955);
and U17291 (N_17291,N_16723,N_16595);
and U17292 (N_17292,N_16641,N_16839);
nand U17293 (N_17293,N_16661,N_16767);
nor U17294 (N_17294,N_16645,N_16723);
nor U17295 (N_17295,N_16661,N_16966);
and U17296 (N_17296,N_16743,N_16662);
or U17297 (N_17297,N_16999,N_16876);
xnor U17298 (N_17298,N_16605,N_16574);
nand U17299 (N_17299,N_16982,N_16820);
nor U17300 (N_17300,N_16637,N_16785);
or U17301 (N_17301,N_16621,N_16926);
nand U17302 (N_17302,N_16614,N_16978);
and U17303 (N_17303,N_16903,N_16566);
xor U17304 (N_17304,N_16548,N_16837);
nand U17305 (N_17305,N_16882,N_16602);
or U17306 (N_17306,N_16789,N_16904);
xor U17307 (N_17307,N_16690,N_16750);
and U17308 (N_17308,N_16514,N_16814);
nor U17309 (N_17309,N_16703,N_16503);
or U17310 (N_17310,N_16657,N_16786);
xnor U17311 (N_17311,N_16809,N_16500);
and U17312 (N_17312,N_16913,N_16790);
xnor U17313 (N_17313,N_16625,N_16986);
and U17314 (N_17314,N_16522,N_16621);
and U17315 (N_17315,N_16664,N_16503);
or U17316 (N_17316,N_16702,N_16972);
or U17317 (N_17317,N_16683,N_16991);
xnor U17318 (N_17318,N_16943,N_16938);
nor U17319 (N_17319,N_16824,N_16866);
and U17320 (N_17320,N_16557,N_16894);
nor U17321 (N_17321,N_16882,N_16999);
and U17322 (N_17322,N_16722,N_16766);
nand U17323 (N_17323,N_16570,N_16851);
or U17324 (N_17324,N_16933,N_16682);
nand U17325 (N_17325,N_16757,N_16925);
and U17326 (N_17326,N_16991,N_16671);
nand U17327 (N_17327,N_16791,N_16826);
and U17328 (N_17328,N_16943,N_16823);
nand U17329 (N_17329,N_16652,N_16741);
or U17330 (N_17330,N_16763,N_16640);
nand U17331 (N_17331,N_16787,N_16795);
xor U17332 (N_17332,N_16615,N_16592);
xnor U17333 (N_17333,N_16921,N_16622);
and U17334 (N_17334,N_16612,N_16597);
nor U17335 (N_17335,N_16676,N_16897);
nand U17336 (N_17336,N_16761,N_16678);
xor U17337 (N_17337,N_16699,N_16985);
nand U17338 (N_17338,N_16656,N_16967);
nor U17339 (N_17339,N_16720,N_16710);
and U17340 (N_17340,N_16939,N_16729);
nor U17341 (N_17341,N_16851,N_16978);
nand U17342 (N_17342,N_16519,N_16752);
and U17343 (N_17343,N_16872,N_16695);
nand U17344 (N_17344,N_16964,N_16707);
and U17345 (N_17345,N_16722,N_16569);
nand U17346 (N_17346,N_16906,N_16985);
and U17347 (N_17347,N_16657,N_16925);
xor U17348 (N_17348,N_16836,N_16675);
xnor U17349 (N_17349,N_16889,N_16994);
nand U17350 (N_17350,N_16666,N_16989);
xor U17351 (N_17351,N_16770,N_16536);
and U17352 (N_17352,N_16860,N_16697);
nand U17353 (N_17353,N_16877,N_16774);
and U17354 (N_17354,N_16914,N_16903);
xor U17355 (N_17355,N_16883,N_16713);
xnor U17356 (N_17356,N_16874,N_16767);
or U17357 (N_17357,N_16785,N_16524);
or U17358 (N_17358,N_16699,N_16882);
nor U17359 (N_17359,N_16791,N_16775);
or U17360 (N_17360,N_16839,N_16837);
nor U17361 (N_17361,N_16815,N_16515);
xor U17362 (N_17362,N_16938,N_16574);
or U17363 (N_17363,N_16844,N_16873);
xor U17364 (N_17364,N_16830,N_16814);
nor U17365 (N_17365,N_16698,N_16682);
nand U17366 (N_17366,N_16730,N_16624);
and U17367 (N_17367,N_16731,N_16914);
and U17368 (N_17368,N_16588,N_16767);
xor U17369 (N_17369,N_16881,N_16945);
xor U17370 (N_17370,N_16861,N_16976);
xor U17371 (N_17371,N_16875,N_16649);
nor U17372 (N_17372,N_16648,N_16543);
nand U17373 (N_17373,N_16502,N_16632);
xnor U17374 (N_17374,N_16645,N_16602);
and U17375 (N_17375,N_16561,N_16505);
nand U17376 (N_17376,N_16717,N_16970);
and U17377 (N_17377,N_16921,N_16877);
xor U17378 (N_17378,N_16684,N_16606);
or U17379 (N_17379,N_16996,N_16832);
xnor U17380 (N_17380,N_16773,N_16538);
nand U17381 (N_17381,N_16759,N_16589);
nand U17382 (N_17382,N_16868,N_16872);
xnor U17383 (N_17383,N_16772,N_16746);
nor U17384 (N_17384,N_16685,N_16942);
or U17385 (N_17385,N_16958,N_16724);
and U17386 (N_17386,N_16681,N_16586);
nand U17387 (N_17387,N_16816,N_16740);
nand U17388 (N_17388,N_16636,N_16568);
and U17389 (N_17389,N_16727,N_16560);
nor U17390 (N_17390,N_16649,N_16761);
and U17391 (N_17391,N_16722,N_16853);
and U17392 (N_17392,N_16952,N_16971);
or U17393 (N_17393,N_16778,N_16590);
and U17394 (N_17394,N_16996,N_16561);
and U17395 (N_17395,N_16817,N_16716);
and U17396 (N_17396,N_16627,N_16948);
and U17397 (N_17397,N_16860,N_16810);
and U17398 (N_17398,N_16693,N_16698);
nor U17399 (N_17399,N_16883,N_16626);
and U17400 (N_17400,N_16532,N_16909);
or U17401 (N_17401,N_16820,N_16876);
nor U17402 (N_17402,N_16802,N_16810);
nand U17403 (N_17403,N_16933,N_16749);
nor U17404 (N_17404,N_16582,N_16627);
nor U17405 (N_17405,N_16924,N_16740);
or U17406 (N_17406,N_16589,N_16872);
and U17407 (N_17407,N_16816,N_16533);
nor U17408 (N_17408,N_16505,N_16694);
and U17409 (N_17409,N_16879,N_16982);
and U17410 (N_17410,N_16768,N_16590);
or U17411 (N_17411,N_16948,N_16717);
and U17412 (N_17412,N_16862,N_16801);
xnor U17413 (N_17413,N_16759,N_16717);
and U17414 (N_17414,N_16505,N_16830);
and U17415 (N_17415,N_16963,N_16644);
nor U17416 (N_17416,N_16877,N_16654);
or U17417 (N_17417,N_16546,N_16549);
and U17418 (N_17418,N_16966,N_16777);
xor U17419 (N_17419,N_16641,N_16640);
and U17420 (N_17420,N_16857,N_16527);
and U17421 (N_17421,N_16839,N_16990);
or U17422 (N_17422,N_16833,N_16636);
or U17423 (N_17423,N_16944,N_16726);
nand U17424 (N_17424,N_16964,N_16853);
and U17425 (N_17425,N_16965,N_16554);
nand U17426 (N_17426,N_16658,N_16828);
nand U17427 (N_17427,N_16908,N_16903);
nand U17428 (N_17428,N_16780,N_16913);
nor U17429 (N_17429,N_16921,N_16518);
and U17430 (N_17430,N_16777,N_16936);
nor U17431 (N_17431,N_16822,N_16917);
xnor U17432 (N_17432,N_16518,N_16993);
or U17433 (N_17433,N_16692,N_16566);
nor U17434 (N_17434,N_16753,N_16756);
xor U17435 (N_17435,N_16742,N_16943);
and U17436 (N_17436,N_16594,N_16898);
or U17437 (N_17437,N_16969,N_16761);
xnor U17438 (N_17438,N_16551,N_16954);
nand U17439 (N_17439,N_16661,N_16651);
nor U17440 (N_17440,N_16635,N_16783);
or U17441 (N_17441,N_16631,N_16553);
nor U17442 (N_17442,N_16502,N_16595);
nand U17443 (N_17443,N_16937,N_16847);
xnor U17444 (N_17444,N_16650,N_16926);
nor U17445 (N_17445,N_16959,N_16500);
nand U17446 (N_17446,N_16540,N_16648);
or U17447 (N_17447,N_16878,N_16621);
xor U17448 (N_17448,N_16942,N_16660);
or U17449 (N_17449,N_16547,N_16564);
nor U17450 (N_17450,N_16820,N_16682);
xor U17451 (N_17451,N_16591,N_16573);
nand U17452 (N_17452,N_16912,N_16600);
xnor U17453 (N_17453,N_16804,N_16609);
nand U17454 (N_17454,N_16564,N_16766);
nor U17455 (N_17455,N_16884,N_16534);
xnor U17456 (N_17456,N_16602,N_16528);
nand U17457 (N_17457,N_16620,N_16536);
and U17458 (N_17458,N_16819,N_16928);
and U17459 (N_17459,N_16863,N_16601);
nor U17460 (N_17460,N_16914,N_16602);
nand U17461 (N_17461,N_16775,N_16650);
xnor U17462 (N_17462,N_16500,N_16581);
nand U17463 (N_17463,N_16890,N_16620);
nor U17464 (N_17464,N_16873,N_16769);
or U17465 (N_17465,N_16993,N_16578);
xnor U17466 (N_17466,N_16902,N_16746);
nand U17467 (N_17467,N_16962,N_16835);
xnor U17468 (N_17468,N_16675,N_16611);
and U17469 (N_17469,N_16828,N_16886);
and U17470 (N_17470,N_16900,N_16972);
xnor U17471 (N_17471,N_16938,N_16637);
xor U17472 (N_17472,N_16771,N_16522);
and U17473 (N_17473,N_16582,N_16510);
nand U17474 (N_17474,N_16993,N_16736);
nor U17475 (N_17475,N_16594,N_16820);
xnor U17476 (N_17476,N_16954,N_16942);
xor U17477 (N_17477,N_16963,N_16849);
or U17478 (N_17478,N_16546,N_16690);
or U17479 (N_17479,N_16525,N_16974);
nand U17480 (N_17480,N_16523,N_16844);
or U17481 (N_17481,N_16958,N_16944);
or U17482 (N_17482,N_16542,N_16907);
nor U17483 (N_17483,N_16516,N_16858);
nor U17484 (N_17484,N_16809,N_16629);
and U17485 (N_17485,N_16538,N_16885);
nand U17486 (N_17486,N_16508,N_16519);
or U17487 (N_17487,N_16767,N_16609);
and U17488 (N_17488,N_16618,N_16712);
xnor U17489 (N_17489,N_16666,N_16756);
nand U17490 (N_17490,N_16862,N_16704);
xor U17491 (N_17491,N_16518,N_16535);
or U17492 (N_17492,N_16848,N_16878);
nand U17493 (N_17493,N_16909,N_16940);
or U17494 (N_17494,N_16644,N_16890);
nand U17495 (N_17495,N_16816,N_16955);
xor U17496 (N_17496,N_16767,N_16832);
nand U17497 (N_17497,N_16750,N_16707);
nor U17498 (N_17498,N_16870,N_16810);
and U17499 (N_17499,N_16935,N_16589);
or U17500 (N_17500,N_17493,N_17335);
nor U17501 (N_17501,N_17038,N_17101);
or U17502 (N_17502,N_17011,N_17491);
and U17503 (N_17503,N_17019,N_17466);
xnor U17504 (N_17504,N_17043,N_17482);
nor U17505 (N_17505,N_17305,N_17331);
nand U17506 (N_17506,N_17201,N_17162);
and U17507 (N_17507,N_17248,N_17033);
nand U17508 (N_17508,N_17408,N_17261);
xnor U17509 (N_17509,N_17383,N_17358);
nand U17510 (N_17510,N_17287,N_17231);
or U17511 (N_17511,N_17353,N_17197);
nor U17512 (N_17512,N_17362,N_17403);
xor U17513 (N_17513,N_17181,N_17254);
nor U17514 (N_17514,N_17208,N_17166);
nor U17515 (N_17515,N_17332,N_17303);
nand U17516 (N_17516,N_17456,N_17045);
and U17517 (N_17517,N_17329,N_17235);
nand U17518 (N_17518,N_17334,N_17199);
and U17519 (N_17519,N_17360,N_17202);
nor U17520 (N_17520,N_17020,N_17125);
xnor U17521 (N_17521,N_17176,N_17333);
or U17522 (N_17522,N_17017,N_17191);
or U17523 (N_17523,N_17128,N_17355);
nand U17524 (N_17524,N_17015,N_17008);
or U17525 (N_17525,N_17130,N_17185);
xor U17526 (N_17526,N_17268,N_17463);
nor U17527 (N_17527,N_17114,N_17047);
xnor U17528 (N_17528,N_17279,N_17243);
or U17529 (N_17529,N_17304,N_17432);
or U17530 (N_17530,N_17222,N_17212);
nand U17531 (N_17531,N_17296,N_17413);
nor U17532 (N_17532,N_17242,N_17350);
nand U17533 (N_17533,N_17266,N_17108);
xnor U17534 (N_17534,N_17085,N_17079);
xor U17535 (N_17535,N_17368,N_17445);
xnor U17536 (N_17536,N_17000,N_17451);
or U17537 (N_17537,N_17116,N_17006);
xnor U17538 (N_17538,N_17310,N_17213);
xor U17539 (N_17539,N_17430,N_17071);
or U17540 (N_17540,N_17168,N_17169);
or U17541 (N_17541,N_17431,N_17300);
nor U17542 (N_17542,N_17321,N_17061);
or U17543 (N_17543,N_17215,N_17400);
and U17544 (N_17544,N_17464,N_17091);
nand U17545 (N_17545,N_17029,N_17060);
nand U17546 (N_17546,N_17005,N_17067);
nand U17547 (N_17547,N_17453,N_17066);
or U17548 (N_17548,N_17419,N_17416);
nand U17549 (N_17549,N_17339,N_17050);
nand U17550 (N_17550,N_17399,N_17136);
and U17551 (N_17551,N_17080,N_17224);
and U17552 (N_17552,N_17426,N_17255);
nand U17553 (N_17553,N_17088,N_17188);
and U17554 (N_17554,N_17349,N_17144);
nor U17555 (N_17555,N_17278,N_17264);
and U17556 (N_17556,N_17328,N_17301);
nand U17557 (N_17557,N_17122,N_17238);
or U17558 (N_17558,N_17338,N_17103);
and U17559 (N_17559,N_17113,N_17145);
nor U17560 (N_17560,N_17083,N_17387);
and U17561 (N_17561,N_17455,N_17234);
nor U17562 (N_17562,N_17381,N_17316);
nor U17563 (N_17563,N_17135,N_17433);
xor U17564 (N_17564,N_17452,N_17193);
xor U17565 (N_17565,N_17393,N_17078);
xnor U17566 (N_17566,N_17023,N_17249);
nand U17567 (N_17567,N_17063,N_17485);
nor U17568 (N_17568,N_17072,N_17096);
and U17569 (N_17569,N_17290,N_17121);
nor U17570 (N_17570,N_17076,N_17318);
xnor U17571 (N_17571,N_17271,N_17376);
nor U17572 (N_17572,N_17428,N_17312);
and U17573 (N_17573,N_17173,N_17158);
nand U17574 (N_17574,N_17373,N_17280);
or U17575 (N_17575,N_17089,N_17467);
xor U17576 (N_17576,N_17468,N_17298);
and U17577 (N_17577,N_17094,N_17274);
nand U17578 (N_17578,N_17102,N_17186);
xor U17579 (N_17579,N_17031,N_17109);
and U17580 (N_17580,N_17371,N_17257);
xnor U17581 (N_17581,N_17032,N_17306);
nor U17582 (N_17582,N_17205,N_17471);
and U17583 (N_17583,N_17037,N_17126);
nand U17584 (N_17584,N_17115,N_17036);
nand U17585 (N_17585,N_17475,N_17459);
nor U17586 (N_17586,N_17359,N_17284);
xnor U17587 (N_17587,N_17164,N_17377);
xnor U17588 (N_17588,N_17069,N_17314);
and U17589 (N_17589,N_17337,N_17171);
nand U17590 (N_17590,N_17256,N_17497);
and U17591 (N_17591,N_17175,N_17273);
nand U17592 (N_17592,N_17270,N_17177);
xor U17593 (N_17593,N_17372,N_17039);
xor U17594 (N_17594,N_17075,N_17297);
nor U17595 (N_17595,N_17203,N_17444);
nand U17596 (N_17596,N_17182,N_17093);
nand U17597 (N_17597,N_17095,N_17390);
and U17598 (N_17598,N_17457,N_17228);
or U17599 (N_17599,N_17086,N_17165);
nand U17600 (N_17600,N_17367,N_17178);
nand U17601 (N_17601,N_17288,N_17289);
nand U17602 (N_17602,N_17336,N_17214);
and U17603 (N_17603,N_17356,N_17439);
xor U17604 (N_17604,N_17313,N_17327);
nor U17605 (N_17605,N_17187,N_17219);
nor U17606 (N_17606,N_17041,N_17404);
or U17607 (N_17607,N_17411,N_17395);
or U17608 (N_17608,N_17134,N_17232);
or U17609 (N_17609,N_17216,N_17267);
nand U17610 (N_17610,N_17097,N_17065);
or U17611 (N_17611,N_17237,N_17410);
or U17612 (N_17612,N_17263,N_17105);
xor U17613 (N_17613,N_17340,N_17230);
nor U17614 (N_17614,N_17397,N_17200);
and U17615 (N_17615,N_17450,N_17406);
or U17616 (N_17616,N_17409,N_17281);
xnor U17617 (N_17617,N_17149,N_17379);
xor U17618 (N_17618,N_17272,N_17241);
xnor U17619 (N_17619,N_17365,N_17405);
or U17620 (N_17620,N_17495,N_17448);
nor U17621 (N_17621,N_17309,N_17351);
nand U17622 (N_17622,N_17401,N_17117);
and U17623 (N_17623,N_17124,N_17153);
nor U17624 (N_17624,N_17172,N_17198);
and U17625 (N_17625,N_17221,N_17150);
xnor U17626 (N_17626,N_17488,N_17375);
xnor U17627 (N_17627,N_17291,N_17441);
and U17628 (N_17628,N_17477,N_17174);
or U17629 (N_17629,N_17402,N_17286);
nand U17630 (N_17630,N_17218,N_17276);
and U17631 (N_17631,N_17319,N_17481);
xor U17632 (N_17632,N_17380,N_17293);
nor U17633 (N_17633,N_17081,N_17084);
or U17634 (N_17634,N_17059,N_17077);
xor U17635 (N_17635,N_17342,N_17057);
and U17636 (N_17636,N_17478,N_17167);
or U17637 (N_17637,N_17386,N_17123);
or U17638 (N_17638,N_17308,N_17207);
nand U17639 (N_17639,N_17012,N_17354);
xnor U17640 (N_17640,N_17425,N_17382);
nor U17641 (N_17641,N_17027,N_17460);
nand U17642 (N_17642,N_17100,N_17496);
xor U17643 (N_17643,N_17325,N_17138);
and U17644 (N_17644,N_17447,N_17446);
nand U17645 (N_17645,N_17236,N_17423);
nor U17646 (N_17646,N_17424,N_17152);
xor U17647 (N_17647,N_17090,N_17127);
xnor U17648 (N_17648,N_17398,N_17420);
nand U17649 (N_17649,N_17389,N_17311);
nor U17650 (N_17650,N_17132,N_17357);
nor U17651 (N_17651,N_17192,N_17148);
nand U17652 (N_17652,N_17053,N_17044);
xnor U17653 (N_17653,N_17131,N_17240);
nor U17654 (N_17654,N_17470,N_17010);
or U17655 (N_17655,N_17156,N_17392);
nand U17656 (N_17656,N_17473,N_17396);
or U17657 (N_17657,N_17021,N_17258);
and U17658 (N_17658,N_17087,N_17004);
nor U17659 (N_17659,N_17064,N_17140);
xor U17660 (N_17660,N_17479,N_17474);
and U17661 (N_17661,N_17499,N_17220);
nor U17662 (N_17662,N_17239,N_17210);
xor U17663 (N_17663,N_17322,N_17026);
or U17664 (N_17664,N_17364,N_17442);
xor U17665 (N_17665,N_17143,N_17034);
nand U17666 (N_17666,N_17003,N_17055);
nor U17667 (N_17667,N_17007,N_17363);
or U17668 (N_17668,N_17252,N_17056);
and U17669 (N_17669,N_17412,N_17111);
nand U17670 (N_17670,N_17112,N_17469);
nor U17671 (N_17671,N_17369,N_17217);
and U17672 (N_17672,N_17110,N_17227);
nor U17673 (N_17673,N_17330,N_17407);
nand U17674 (N_17674,N_17299,N_17492);
xor U17675 (N_17675,N_17154,N_17347);
or U17676 (N_17676,N_17099,N_17120);
xnor U17677 (N_17677,N_17098,N_17163);
xnor U17678 (N_17678,N_17253,N_17480);
and U17679 (N_17679,N_17461,N_17265);
xor U17680 (N_17680,N_17048,N_17294);
xnor U17681 (N_17681,N_17344,N_17196);
nand U17682 (N_17682,N_17104,N_17269);
or U17683 (N_17683,N_17370,N_17352);
nand U17684 (N_17684,N_17320,N_17245);
or U17685 (N_17685,N_17250,N_17179);
nor U17686 (N_17686,N_17315,N_17052);
nor U17687 (N_17687,N_17378,N_17106);
nor U17688 (N_17688,N_17429,N_17051);
or U17689 (N_17689,N_17030,N_17229);
or U17690 (N_17690,N_17498,N_17206);
xnor U17691 (N_17691,N_17414,N_17262);
nor U17692 (N_17692,N_17092,N_17194);
or U17693 (N_17693,N_17049,N_17223);
or U17694 (N_17694,N_17494,N_17366);
nand U17695 (N_17695,N_17388,N_17151);
and U17696 (N_17696,N_17462,N_17119);
or U17697 (N_17697,N_17438,N_17183);
xnor U17698 (N_17698,N_17024,N_17141);
and U17699 (N_17699,N_17326,N_17487);
nand U17700 (N_17700,N_17275,N_17082);
and U17701 (N_17701,N_17427,N_17443);
xnor U17702 (N_17702,N_17385,N_17159);
nand U17703 (N_17703,N_17465,N_17483);
and U17704 (N_17704,N_17013,N_17391);
nor U17705 (N_17705,N_17018,N_17345);
xor U17706 (N_17706,N_17054,N_17346);
xor U17707 (N_17707,N_17035,N_17118);
or U17708 (N_17708,N_17454,N_17436);
or U17709 (N_17709,N_17009,N_17180);
or U17710 (N_17710,N_17068,N_17246);
nand U17711 (N_17711,N_17184,N_17014);
or U17712 (N_17712,N_17421,N_17285);
xor U17713 (N_17713,N_17001,N_17062);
nand U17714 (N_17714,N_17283,N_17440);
xnor U17715 (N_17715,N_17259,N_17484);
and U17716 (N_17716,N_17348,N_17139);
or U17717 (N_17717,N_17040,N_17251);
and U17718 (N_17718,N_17307,N_17317);
xnor U17719 (N_17719,N_17324,N_17282);
nand U17720 (N_17720,N_17260,N_17422);
nor U17721 (N_17721,N_17129,N_17155);
nand U17722 (N_17722,N_17341,N_17016);
nand U17723 (N_17723,N_17190,N_17394);
nor U17724 (N_17724,N_17486,N_17449);
nor U17725 (N_17725,N_17490,N_17476);
nand U17726 (N_17726,N_17002,N_17022);
nor U17727 (N_17727,N_17225,N_17157);
nand U17728 (N_17728,N_17434,N_17247);
nor U17729 (N_17729,N_17489,N_17437);
and U17730 (N_17730,N_17374,N_17384);
nand U17731 (N_17731,N_17211,N_17417);
nor U17732 (N_17732,N_17137,N_17142);
nor U17733 (N_17733,N_17295,N_17226);
or U17734 (N_17734,N_17133,N_17028);
and U17735 (N_17735,N_17160,N_17209);
or U17736 (N_17736,N_17189,N_17204);
or U17737 (N_17737,N_17472,N_17418);
and U17738 (N_17738,N_17107,N_17233);
nor U17739 (N_17739,N_17244,N_17302);
or U17740 (N_17740,N_17161,N_17361);
and U17741 (N_17741,N_17323,N_17277);
or U17742 (N_17742,N_17025,N_17435);
and U17743 (N_17743,N_17146,N_17458);
nand U17744 (N_17744,N_17195,N_17415);
or U17745 (N_17745,N_17147,N_17042);
nand U17746 (N_17746,N_17073,N_17070);
nor U17747 (N_17747,N_17292,N_17170);
nor U17748 (N_17748,N_17046,N_17074);
xnor U17749 (N_17749,N_17058,N_17343);
nor U17750 (N_17750,N_17163,N_17168);
nor U17751 (N_17751,N_17315,N_17277);
nor U17752 (N_17752,N_17181,N_17172);
xnor U17753 (N_17753,N_17000,N_17335);
xnor U17754 (N_17754,N_17284,N_17400);
xor U17755 (N_17755,N_17338,N_17287);
and U17756 (N_17756,N_17310,N_17412);
nor U17757 (N_17757,N_17194,N_17043);
xnor U17758 (N_17758,N_17380,N_17115);
xor U17759 (N_17759,N_17059,N_17268);
nor U17760 (N_17760,N_17481,N_17096);
nand U17761 (N_17761,N_17268,N_17452);
xor U17762 (N_17762,N_17206,N_17372);
and U17763 (N_17763,N_17149,N_17040);
nor U17764 (N_17764,N_17376,N_17343);
and U17765 (N_17765,N_17445,N_17490);
or U17766 (N_17766,N_17180,N_17291);
xor U17767 (N_17767,N_17388,N_17270);
and U17768 (N_17768,N_17206,N_17097);
and U17769 (N_17769,N_17121,N_17011);
xor U17770 (N_17770,N_17145,N_17049);
nor U17771 (N_17771,N_17197,N_17312);
nand U17772 (N_17772,N_17374,N_17049);
or U17773 (N_17773,N_17159,N_17017);
nand U17774 (N_17774,N_17478,N_17441);
nor U17775 (N_17775,N_17099,N_17204);
nor U17776 (N_17776,N_17302,N_17026);
or U17777 (N_17777,N_17066,N_17402);
or U17778 (N_17778,N_17411,N_17168);
or U17779 (N_17779,N_17298,N_17285);
xnor U17780 (N_17780,N_17166,N_17013);
nand U17781 (N_17781,N_17088,N_17126);
and U17782 (N_17782,N_17211,N_17115);
or U17783 (N_17783,N_17121,N_17268);
nand U17784 (N_17784,N_17298,N_17175);
nor U17785 (N_17785,N_17066,N_17382);
or U17786 (N_17786,N_17442,N_17037);
and U17787 (N_17787,N_17295,N_17339);
or U17788 (N_17788,N_17157,N_17003);
nand U17789 (N_17789,N_17173,N_17087);
nand U17790 (N_17790,N_17438,N_17452);
nand U17791 (N_17791,N_17373,N_17207);
nor U17792 (N_17792,N_17446,N_17047);
xnor U17793 (N_17793,N_17025,N_17425);
xor U17794 (N_17794,N_17243,N_17312);
xor U17795 (N_17795,N_17162,N_17384);
and U17796 (N_17796,N_17381,N_17265);
nor U17797 (N_17797,N_17291,N_17221);
and U17798 (N_17798,N_17435,N_17257);
and U17799 (N_17799,N_17074,N_17327);
nand U17800 (N_17800,N_17096,N_17105);
nor U17801 (N_17801,N_17324,N_17254);
or U17802 (N_17802,N_17372,N_17486);
and U17803 (N_17803,N_17150,N_17092);
xnor U17804 (N_17804,N_17362,N_17113);
and U17805 (N_17805,N_17196,N_17326);
xnor U17806 (N_17806,N_17379,N_17192);
or U17807 (N_17807,N_17445,N_17046);
nor U17808 (N_17808,N_17426,N_17098);
nand U17809 (N_17809,N_17077,N_17361);
nand U17810 (N_17810,N_17434,N_17228);
nor U17811 (N_17811,N_17183,N_17259);
and U17812 (N_17812,N_17302,N_17044);
nor U17813 (N_17813,N_17300,N_17147);
and U17814 (N_17814,N_17193,N_17379);
xnor U17815 (N_17815,N_17121,N_17144);
nor U17816 (N_17816,N_17168,N_17157);
nor U17817 (N_17817,N_17404,N_17146);
xor U17818 (N_17818,N_17477,N_17235);
nand U17819 (N_17819,N_17264,N_17471);
xor U17820 (N_17820,N_17266,N_17289);
nand U17821 (N_17821,N_17127,N_17467);
nor U17822 (N_17822,N_17242,N_17289);
or U17823 (N_17823,N_17399,N_17342);
xnor U17824 (N_17824,N_17123,N_17479);
nand U17825 (N_17825,N_17204,N_17001);
or U17826 (N_17826,N_17069,N_17483);
nand U17827 (N_17827,N_17307,N_17190);
nor U17828 (N_17828,N_17180,N_17264);
nand U17829 (N_17829,N_17259,N_17434);
xnor U17830 (N_17830,N_17351,N_17406);
or U17831 (N_17831,N_17450,N_17240);
nand U17832 (N_17832,N_17134,N_17034);
and U17833 (N_17833,N_17365,N_17156);
and U17834 (N_17834,N_17107,N_17358);
and U17835 (N_17835,N_17154,N_17064);
and U17836 (N_17836,N_17119,N_17151);
xor U17837 (N_17837,N_17227,N_17344);
xor U17838 (N_17838,N_17167,N_17059);
nor U17839 (N_17839,N_17054,N_17260);
nand U17840 (N_17840,N_17165,N_17463);
xor U17841 (N_17841,N_17491,N_17286);
nand U17842 (N_17842,N_17243,N_17304);
xor U17843 (N_17843,N_17314,N_17496);
or U17844 (N_17844,N_17241,N_17310);
xnor U17845 (N_17845,N_17170,N_17192);
nor U17846 (N_17846,N_17117,N_17275);
and U17847 (N_17847,N_17150,N_17477);
xor U17848 (N_17848,N_17427,N_17024);
nand U17849 (N_17849,N_17101,N_17359);
nor U17850 (N_17850,N_17357,N_17004);
nand U17851 (N_17851,N_17331,N_17149);
and U17852 (N_17852,N_17031,N_17286);
xnor U17853 (N_17853,N_17328,N_17256);
xnor U17854 (N_17854,N_17477,N_17123);
or U17855 (N_17855,N_17078,N_17201);
or U17856 (N_17856,N_17212,N_17250);
or U17857 (N_17857,N_17491,N_17371);
nor U17858 (N_17858,N_17293,N_17146);
or U17859 (N_17859,N_17359,N_17217);
and U17860 (N_17860,N_17047,N_17266);
nor U17861 (N_17861,N_17310,N_17302);
and U17862 (N_17862,N_17425,N_17224);
xnor U17863 (N_17863,N_17459,N_17097);
and U17864 (N_17864,N_17174,N_17362);
nand U17865 (N_17865,N_17376,N_17234);
nand U17866 (N_17866,N_17350,N_17491);
xnor U17867 (N_17867,N_17292,N_17431);
and U17868 (N_17868,N_17238,N_17456);
and U17869 (N_17869,N_17185,N_17038);
xnor U17870 (N_17870,N_17333,N_17396);
and U17871 (N_17871,N_17369,N_17063);
and U17872 (N_17872,N_17401,N_17243);
nand U17873 (N_17873,N_17389,N_17015);
xor U17874 (N_17874,N_17052,N_17278);
nor U17875 (N_17875,N_17099,N_17269);
or U17876 (N_17876,N_17317,N_17108);
xor U17877 (N_17877,N_17021,N_17098);
and U17878 (N_17878,N_17393,N_17372);
and U17879 (N_17879,N_17063,N_17173);
xnor U17880 (N_17880,N_17042,N_17123);
xnor U17881 (N_17881,N_17226,N_17455);
xor U17882 (N_17882,N_17270,N_17421);
nand U17883 (N_17883,N_17242,N_17077);
or U17884 (N_17884,N_17055,N_17006);
nand U17885 (N_17885,N_17386,N_17291);
nor U17886 (N_17886,N_17234,N_17166);
nand U17887 (N_17887,N_17242,N_17104);
xnor U17888 (N_17888,N_17127,N_17457);
or U17889 (N_17889,N_17277,N_17444);
nor U17890 (N_17890,N_17201,N_17236);
or U17891 (N_17891,N_17016,N_17441);
xnor U17892 (N_17892,N_17443,N_17187);
xnor U17893 (N_17893,N_17160,N_17331);
or U17894 (N_17894,N_17220,N_17076);
xnor U17895 (N_17895,N_17301,N_17444);
nand U17896 (N_17896,N_17315,N_17031);
xnor U17897 (N_17897,N_17132,N_17120);
nor U17898 (N_17898,N_17251,N_17190);
and U17899 (N_17899,N_17108,N_17064);
or U17900 (N_17900,N_17169,N_17291);
xor U17901 (N_17901,N_17087,N_17099);
or U17902 (N_17902,N_17472,N_17362);
and U17903 (N_17903,N_17384,N_17302);
xor U17904 (N_17904,N_17287,N_17143);
xor U17905 (N_17905,N_17234,N_17356);
nand U17906 (N_17906,N_17017,N_17123);
and U17907 (N_17907,N_17248,N_17170);
xor U17908 (N_17908,N_17231,N_17455);
nand U17909 (N_17909,N_17440,N_17247);
nand U17910 (N_17910,N_17493,N_17400);
xnor U17911 (N_17911,N_17212,N_17260);
xor U17912 (N_17912,N_17117,N_17111);
xor U17913 (N_17913,N_17062,N_17260);
xnor U17914 (N_17914,N_17052,N_17256);
nand U17915 (N_17915,N_17039,N_17357);
xor U17916 (N_17916,N_17140,N_17419);
xor U17917 (N_17917,N_17272,N_17020);
and U17918 (N_17918,N_17034,N_17212);
and U17919 (N_17919,N_17021,N_17230);
xor U17920 (N_17920,N_17043,N_17129);
and U17921 (N_17921,N_17491,N_17141);
nand U17922 (N_17922,N_17401,N_17175);
nor U17923 (N_17923,N_17006,N_17042);
or U17924 (N_17924,N_17069,N_17460);
xnor U17925 (N_17925,N_17027,N_17233);
nor U17926 (N_17926,N_17191,N_17286);
xnor U17927 (N_17927,N_17189,N_17337);
and U17928 (N_17928,N_17400,N_17259);
xnor U17929 (N_17929,N_17349,N_17417);
nor U17930 (N_17930,N_17230,N_17488);
nand U17931 (N_17931,N_17236,N_17290);
nand U17932 (N_17932,N_17312,N_17172);
and U17933 (N_17933,N_17054,N_17156);
and U17934 (N_17934,N_17450,N_17238);
nor U17935 (N_17935,N_17189,N_17396);
nor U17936 (N_17936,N_17420,N_17278);
and U17937 (N_17937,N_17208,N_17336);
nand U17938 (N_17938,N_17420,N_17378);
and U17939 (N_17939,N_17101,N_17453);
nor U17940 (N_17940,N_17062,N_17470);
nand U17941 (N_17941,N_17340,N_17292);
or U17942 (N_17942,N_17193,N_17355);
or U17943 (N_17943,N_17487,N_17223);
nand U17944 (N_17944,N_17273,N_17154);
or U17945 (N_17945,N_17458,N_17460);
or U17946 (N_17946,N_17277,N_17177);
or U17947 (N_17947,N_17250,N_17176);
xnor U17948 (N_17948,N_17084,N_17481);
nor U17949 (N_17949,N_17371,N_17180);
or U17950 (N_17950,N_17345,N_17349);
nor U17951 (N_17951,N_17282,N_17157);
nor U17952 (N_17952,N_17130,N_17368);
and U17953 (N_17953,N_17302,N_17128);
xnor U17954 (N_17954,N_17118,N_17438);
nand U17955 (N_17955,N_17290,N_17067);
and U17956 (N_17956,N_17078,N_17230);
and U17957 (N_17957,N_17396,N_17382);
or U17958 (N_17958,N_17384,N_17340);
or U17959 (N_17959,N_17336,N_17034);
or U17960 (N_17960,N_17113,N_17485);
or U17961 (N_17961,N_17193,N_17013);
nor U17962 (N_17962,N_17177,N_17426);
nand U17963 (N_17963,N_17011,N_17385);
nor U17964 (N_17964,N_17497,N_17252);
nor U17965 (N_17965,N_17022,N_17052);
nor U17966 (N_17966,N_17395,N_17271);
xnor U17967 (N_17967,N_17481,N_17077);
nor U17968 (N_17968,N_17091,N_17457);
nor U17969 (N_17969,N_17400,N_17191);
nand U17970 (N_17970,N_17345,N_17300);
xor U17971 (N_17971,N_17388,N_17207);
xor U17972 (N_17972,N_17331,N_17281);
and U17973 (N_17973,N_17310,N_17454);
xor U17974 (N_17974,N_17144,N_17101);
and U17975 (N_17975,N_17169,N_17298);
and U17976 (N_17976,N_17377,N_17154);
and U17977 (N_17977,N_17186,N_17398);
nor U17978 (N_17978,N_17161,N_17467);
or U17979 (N_17979,N_17291,N_17095);
xor U17980 (N_17980,N_17048,N_17092);
nand U17981 (N_17981,N_17464,N_17117);
or U17982 (N_17982,N_17171,N_17277);
xor U17983 (N_17983,N_17495,N_17033);
and U17984 (N_17984,N_17423,N_17433);
nor U17985 (N_17985,N_17309,N_17165);
xor U17986 (N_17986,N_17459,N_17374);
nand U17987 (N_17987,N_17041,N_17391);
nand U17988 (N_17988,N_17125,N_17406);
nand U17989 (N_17989,N_17153,N_17282);
xor U17990 (N_17990,N_17006,N_17253);
xor U17991 (N_17991,N_17228,N_17259);
nor U17992 (N_17992,N_17262,N_17011);
xor U17993 (N_17993,N_17321,N_17456);
or U17994 (N_17994,N_17217,N_17273);
or U17995 (N_17995,N_17351,N_17449);
and U17996 (N_17996,N_17317,N_17394);
or U17997 (N_17997,N_17378,N_17291);
and U17998 (N_17998,N_17401,N_17297);
nor U17999 (N_17999,N_17184,N_17282);
and U18000 (N_18000,N_17666,N_17628);
nand U18001 (N_18001,N_17815,N_17954);
xor U18002 (N_18002,N_17529,N_17934);
and U18003 (N_18003,N_17899,N_17804);
xnor U18004 (N_18004,N_17589,N_17681);
nand U18005 (N_18005,N_17844,N_17523);
nand U18006 (N_18006,N_17704,N_17709);
or U18007 (N_18007,N_17941,N_17930);
nor U18008 (N_18008,N_17676,N_17514);
nor U18009 (N_18009,N_17999,N_17763);
or U18010 (N_18010,N_17616,N_17621);
nand U18011 (N_18011,N_17670,N_17861);
xnor U18012 (N_18012,N_17719,N_17707);
xnor U18013 (N_18013,N_17793,N_17914);
or U18014 (N_18014,N_17635,N_17721);
nand U18015 (N_18015,N_17504,N_17886);
nor U18016 (N_18016,N_17591,N_17752);
and U18017 (N_18017,N_17827,N_17813);
nor U18018 (N_18018,N_17610,N_17962);
xor U18019 (N_18019,N_17622,N_17913);
nand U18020 (N_18020,N_17694,N_17658);
xor U18021 (N_18021,N_17674,N_17920);
and U18022 (N_18022,N_17774,N_17547);
nor U18023 (N_18023,N_17933,N_17794);
nand U18024 (N_18024,N_17854,N_17895);
and U18025 (N_18025,N_17546,N_17940);
or U18026 (N_18026,N_17502,N_17873);
and U18027 (N_18027,N_17742,N_17571);
or U18028 (N_18028,N_17651,N_17874);
xnor U18029 (N_18029,N_17530,N_17878);
nor U18030 (N_18030,N_17972,N_17626);
xnor U18031 (N_18031,N_17845,N_17749);
nand U18032 (N_18032,N_17743,N_17801);
or U18033 (N_18033,N_17946,N_17517);
or U18034 (N_18034,N_17617,N_17567);
xor U18035 (N_18035,N_17633,N_17805);
and U18036 (N_18036,N_17842,N_17711);
nand U18037 (N_18037,N_17967,N_17561);
or U18038 (N_18038,N_17905,N_17970);
or U18039 (N_18039,N_17764,N_17862);
xnor U18040 (N_18040,N_17692,N_17532);
nand U18041 (N_18041,N_17679,N_17597);
nor U18042 (N_18042,N_17713,N_17748);
xnor U18043 (N_18043,N_17888,N_17548);
nor U18044 (N_18044,N_17516,N_17853);
or U18045 (N_18045,N_17510,N_17593);
nand U18046 (N_18046,N_17852,N_17935);
xor U18047 (N_18047,N_17531,N_17996);
xor U18048 (N_18048,N_17755,N_17579);
or U18049 (N_18049,N_17686,N_17847);
nor U18050 (N_18050,N_17775,N_17700);
nand U18051 (N_18051,N_17963,N_17642);
or U18052 (N_18052,N_17936,N_17612);
and U18053 (N_18053,N_17543,N_17969);
or U18054 (N_18054,N_17585,N_17981);
nor U18055 (N_18055,N_17648,N_17958);
nand U18056 (N_18056,N_17625,N_17608);
nand U18057 (N_18057,N_17644,N_17799);
or U18058 (N_18058,N_17646,N_17909);
nor U18059 (N_18059,N_17678,N_17515);
nor U18060 (N_18060,N_17927,N_17677);
xor U18061 (N_18061,N_17691,N_17654);
or U18062 (N_18062,N_17839,N_17753);
nand U18063 (N_18063,N_17910,N_17906);
xor U18064 (N_18064,N_17916,N_17965);
nand U18065 (N_18065,N_17866,N_17949);
xnor U18066 (N_18066,N_17766,N_17717);
nor U18067 (N_18067,N_17740,N_17551);
xnor U18068 (N_18068,N_17911,N_17838);
nand U18069 (N_18069,N_17695,N_17986);
nand U18070 (N_18070,N_17993,N_17918);
or U18071 (N_18071,N_17840,N_17860);
nor U18072 (N_18072,N_17896,N_17511);
nor U18073 (N_18073,N_17536,N_17762);
xor U18074 (N_18074,N_17525,N_17639);
xnor U18075 (N_18075,N_17500,N_17797);
nor U18076 (N_18076,N_17758,N_17984);
xnor U18077 (N_18077,N_17557,N_17802);
nor U18078 (N_18078,N_17588,N_17641);
nand U18079 (N_18079,N_17792,N_17615);
and U18080 (N_18080,N_17791,N_17535);
xor U18081 (N_18081,N_17959,N_17982);
or U18082 (N_18082,N_17919,N_17994);
and U18083 (N_18083,N_17950,N_17577);
nand U18084 (N_18084,N_17640,N_17777);
and U18085 (N_18085,N_17836,N_17673);
and U18086 (N_18086,N_17575,N_17668);
nand U18087 (N_18087,N_17811,N_17718);
and U18088 (N_18088,N_17533,N_17956);
or U18089 (N_18089,N_17932,N_17636);
or U18090 (N_18090,N_17783,N_17706);
and U18091 (N_18091,N_17826,N_17618);
and U18092 (N_18092,N_17778,N_17680);
or U18093 (N_18093,N_17759,N_17624);
xor U18094 (N_18094,N_17931,N_17524);
nand U18095 (N_18095,N_17767,N_17971);
nand U18096 (N_18096,N_17509,N_17643);
nand U18097 (N_18097,N_17701,N_17841);
nand U18098 (N_18098,N_17894,N_17693);
and U18099 (N_18099,N_17659,N_17870);
and U18100 (N_18100,N_17587,N_17664);
or U18101 (N_18101,N_17849,N_17505);
nand U18102 (N_18102,N_17924,N_17875);
and U18103 (N_18103,N_17560,N_17627);
nor U18104 (N_18104,N_17921,N_17871);
or U18105 (N_18105,N_17771,N_17929);
or U18106 (N_18106,N_17563,N_17902);
and U18107 (N_18107,N_17915,N_17991);
nand U18108 (N_18108,N_17819,N_17653);
nor U18109 (N_18109,N_17983,N_17922);
nor U18110 (N_18110,N_17903,N_17901);
nor U18111 (N_18111,N_17688,N_17776);
xor U18112 (N_18112,N_17582,N_17623);
xor U18113 (N_18113,N_17832,N_17741);
nand U18114 (N_18114,N_17539,N_17945);
nor U18115 (N_18115,N_17599,N_17816);
or U18116 (N_18116,N_17831,N_17980);
nand U18117 (N_18117,N_17672,N_17837);
nor U18118 (N_18118,N_17848,N_17630);
nand U18119 (N_18119,N_17513,N_17785);
nand U18120 (N_18120,N_17689,N_17881);
xor U18121 (N_18121,N_17992,N_17501);
nand U18122 (N_18122,N_17978,N_17897);
and U18123 (N_18123,N_17558,N_17795);
or U18124 (N_18124,N_17883,N_17747);
or U18125 (N_18125,N_17699,N_17820);
nor U18126 (N_18126,N_17773,N_17825);
and U18127 (N_18127,N_17620,N_17738);
nand U18128 (N_18128,N_17846,N_17540);
or U18129 (N_18129,N_17885,N_17655);
xor U18130 (N_18130,N_17702,N_17534);
nand U18131 (N_18131,N_17818,N_17926);
nand U18132 (N_18132,N_17619,N_17607);
nand U18133 (N_18133,N_17732,N_17581);
nand U18134 (N_18134,N_17729,N_17884);
nor U18135 (N_18135,N_17882,N_17850);
and U18136 (N_18136,N_17966,N_17812);
nand U18137 (N_18137,N_17671,N_17863);
and U18138 (N_18138,N_17953,N_17573);
nor U18139 (N_18139,N_17977,N_17865);
and U18140 (N_18140,N_17851,N_17638);
nand U18141 (N_18141,N_17590,N_17684);
nor U18142 (N_18142,N_17735,N_17868);
nand U18143 (N_18143,N_17614,N_17867);
or U18144 (N_18144,N_17879,N_17698);
nand U18145 (N_18145,N_17864,N_17556);
or U18146 (N_18146,N_17781,N_17961);
nor U18147 (N_18147,N_17989,N_17550);
nor U18148 (N_18148,N_17925,N_17520);
nand U18149 (N_18149,N_17988,N_17583);
and U18150 (N_18150,N_17734,N_17872);
xor U18151 (N_18151,N_17828,N_17697);
xnor U18152 (N_18152,N_17955,N_17807);
or U18153 (N_18153,N_17564,N_17632);
nor U18154 (N_18154,N_17652,N_17716);
and U18155 (N_18155,N_17995,N_17606);
xnor U18156 (N_18156,N_17538,N_17754);
nand U18157 (N_18157,N_17765,N_17603);
nor U18158 (N_18158,N_17726,N_17745);
nand U18159 (N_18159,N_17715,N_17506);
xnor U18160 (N_18160,N_17541,N_17856);
or U18161 (N_18161,N_17917,N_17537);
or U18162 (N_18162,N_17545,N_17650);
or U18163 (N_18163,N_17683,N_17968);
xnor U18164 (N_18164,N_17724,N_17542);
xor U18165 (N_18165,N_17710,N_17800);
nor U18166 (N_18166,N_17647,N_17705);
nand U18167 (N_18167,N_17720,N_17817);
nor U18168 (N_18168,N_17788,N_17733);
nor U18169 (N_18169,N_17736,N_17562);
xor U18170 (N_18170,N_17663,N_17998);
xor U18171 (N_18171,N_17938,N_17889);
or U18172 (N_18172,N_17731,N_17730);
or U18173 (N_18173,N_17568,N_17796);
nor U18174 (N_18174,N_17578,N_17544);
nor U18175 (N_18175,N_17645,N_17876);
xor U18176 (N_18176,N_17789,N_17631);
or U18177 (N_18177,N_17908,N_17601);
xor U18178 (N_18178,N_17843,N_17857);
nor U18179 (N_18179,N_17761,N_17553);
xor U18180 (N_18180,N_17629,N_17833);
nand U18181 (N_18181,N_17574,N_17690);
nor U18182 (N_18182,N_17928,N_17829);
and U18183 (N_18183,N_17559,N_17685);
nand U18184 (N_18184,N_17768,N_17787);
nand U18185 (N_18185,N_17737,N_17580);
or U18186 (N_18186,N_17973,N_17974);
or U18187 (N_18187,N_17725,N_17869);
and U18188 (N_18188,N_17527,N_17576);
and U18189 (N_18189,N_17806,N_17703);
and U18190 (N_18190,N_17552,N_17549);
or U18191 (N_18191,N_17572,N_17669);
nor U18192 (N_18192,N_17780,N_17667);
nand U18193 (N_18193,N_17600,N_17769);
and U18194 (N_18194,N_17605,N_17859);
and U18195 (N_18195,N_17512,N_17757);
nor U18196 (N_18196,N_17808,N_17521);
and U18197 (N_18197,N_17675,N_17985);
or U18198 (N_18198,N_17898,N_17891);
nand U18199 (N_18199,N_17595,N_17660);
xnor U18200 (N_18200,N_17656,N_17662);
and U18201 (N_18201,N_17507,N_17803);
nand U18202 (N_18202,N_17822,N_17830);
xor U18203 (N_18203,N_17942,N_17912);
xnor U18204 (N_18204,N_17979,N_17723);
or U18205 (N_18205,N_17760,N_17739);
and U18206 (N_18206,N_17887,N_17746);
and U18207 (N_18207,N_17712,N_17907);
or U18208 (N_18208,N_17637,N_17790);
and U18209 (N_18209,N_17770,N_17604);
and U18210 (N_18210,N_17855,N_17823);
nor U18211 (N_18211,N_17834,N_17528);
and U18212 (N_18212,N_17798,N_17948);
nor U18213 (N_18213,N_17596,N_17728);
or U18214 (N_18214,N_17987,N_17526);
and U18215 (N_18215,N_17696,N_17592);
or U18216 (N_18216,N_17779,N_17824);
nand U18217 (N_18217,N_17708,N_17727);
nand U18218 (N_18218,N_17858,N_17649);
xor U18219 (N_18219,N_17570,N_17503);
nor U18220 (N_18220,N_17687,N_17611);
or U18221 (N_18221,N_17714,N_17877);
nor U18222 (N_18222,N_17722,N_17613);
nor U18223 (N_18223,N_17522,N_17821);
xnor U18224 (N_18224,N_17756,N_17554);
nand U18225 (N_18225,N_17584,N_17634);
nor U18226 (N_18226,N_17602,N_17661);
nand U18227 (N_18227,N_17990,N_17964);
and U18228 (N_18228,N_17814,N_17784);
nor U18229 (N_18229,N_17890,N_17569);
nor U18230 (N_18230,N_17565,N_17937);
or U18231 (N_18231,N_17555,N_17923);
nor U18232 (N_18232,N_17657,N_17893);
or U18233 (N_18233,N_17786,N_17997);
or U18234 (N_18234,N_17880,N_17508);
or U18235 (N_18235,N_17943,N_17750);
and U18236 (N_18236,N_17960,N_17809);
nand U18237 (N_18237,N_17904,N_17782);
nand U18238 (N_18238,N_17951,N_17665);
xnor U18239 (N_18239,N_17518,N_17751);
nor U18240 (N_18240,N_17772,N_17586);
and U18241 (N_18241,N_17835,N_17598);
or U18242 (N_18242,N_17609,N_17976);
xnor U18243 (N_18243,N_17810,N_17744);
nand U18244 (N_18244,N_17892,N_17682);
and U18245 (N_18245,N_17566,N_17952);
and U18246 (N_18246,N_17939,N_17900);
xor U18247 (N_18247,N_17594,N_17947);
xnor U18248 (N_18248,N_17944,N_17519);
nor U18249 (N_18249,N_17975,N_17957);
nor U18250 (N_18250,N_17687,N_17857);
xor U18251 (N_18251,N_17536,N_17861);
or U18252 (N_18252,N_17741,N_17835);
and U18253 (N_18253,N_17592,N_17963);
nand U18254 (N_18254,N_17894,N_17931);
nand U18255 (N_18255,N_17562,N_17926);
and U18256 (N_18256,N_17684,N_17742);
and U18257 (N_18257,N_17665,N_17631);
nand U18258 (N_18258,N_17530,N_17969);
and U18259 (N_18259,N_17821,N_17925);
and U18260 (N_18260,N_17907,N_17900);
and U18261 (N_18261,N_17952,N_17994);
or U18262 (N_18262,N_17851,N_17982);
or U18263 (N_18263,N_17717,N_17866);
nand U18264 (N_18264,N_17637,N_17561);
and U18265 (N_18265,N_17638,N_17538);
and U18266 (N_18266,N_17819,N_17626);
nor U18267 (N_18267,N_17979,N_17605);
and U18268 (N_18268,N_17740,N_17663);
and U18269 (N_18269,N_17589,N_17973);
and U18270 (N_18270,N_17738,N_17646);
nor U18271 (N_18271,N_17521,N_17852);
xor U18272 (N_18272,N_17746,N_17824);
and U18273 (N_18273,N_17891,N_17613);
or U18274 (N_18274,N_17621,N_17815);
nand U18275 (N_18275,N_17530,N_17827);
and U18276 (N_18276,N_17506,N_17963);
and U18277 (N_18277,N_17825,N_17664);
nor U18278 (N_18278,N_17909,N_17697);
xnor U18279 (N_18279,N_17844,N_17971);
nor U18280 (N_18280,N_17621,N_17998);
xor U18281 (N_18281,N_17928,N_17980);
and U18282 (N_18282,N_17927,N_17837);
nand U18283 (N_18283,N_17863,N_17831);
nand U18284 (N_18284,N_17987,N_17654);
nor U18285 (N_18285,N_17630,N_17669);
nor U18286 (N_18286,N_17902,N_17531);
nor U18287 (N_18287,N_17728,N_17973);
or U18288 (N_18288,N_17876,N_17801);
xnor U18289 (N_18289,N_17554,N_17815);
or U18290 (N_18290,N_17958,N_17614);
nand U18291 (N_18291,N_17739,N_17792);
and U18292 (N_18292,N_17924,N_17729);
or U18293 (N_18293,N_17844,N_17828);
xor U18294 (N_18294,N_17737,N_17749);
nand U18295 (N_18295,N_17907,N_17904);
nor U18296 (N_18296,N_17960,N_17979);
xor U18297 (N_18297,N_17669,N_17596);
nand U18298 (N_18298,N_17688,N_17618);
and U18299 (N_18299,N_17517,N_17819);
and U18300 (N_18300,N_17737,N_17614);
or U18301 (N_18301,N_17620,N_17596);
or U18302 (N_18302,N_17917,N_17502);
nor U18303 (N_18303,N_17989,N_17500);
or U18304 (N_18304,N_17756,N_17835);
nor U18305 (N_18305,N_17889,N_17644);
or U18306 (N_18306,N_17703,N_17788);
and U18307 (N_18307,N_17613,N_17669);
xor U18308 (N_18308,N_17533,N_17850);
nor U18309 (N_18309,N_17526,N_17607);
nand U18310 (N_18310,N_17867,N_17935);
xor U18311 (N_18311,N_17768,N_17922);
or U18312 (N_18312,N_17517,N_17977);
and U18313 (N_18313,N_17789,N_17950);
and U18314 (N_18314,N_17869,N_17649);
nand U18315 (N_18315,N_17502,N_17848);
nor U18316 (N_18316,N_17679,N_17590);
xnor U18317 (N_18317,N_17978,N_17793);
xnor U18318 (N_18318,N_17670,N_17998);
or U18319 (N_18319,N_17725,N_17503);
nor U18320 (N_18320,N_17578,N_17947);
or U18321 (N_18321,N_17786,N_17702);
and U18322 (N_18322,N_17823,N_17529);
or U18323 (N_18323,N_17567,N_17557);
xnor U18324 (N_18324,N_17799,N_17790);
or U18325 (N_18325,N_17958,N_17768);
xnor U18326 (N_18326,N_17943,N_17882);
or U18327 (N_18327,N_17625,N_17727);
nand U18328 (N_18328,N_17739,N_17594);
or U18329 (N_18329,N_17685,N_17565);
and U18330 (N_18330,N_17546,N_17527);
and U18331 (N_18331,N_17517,N_17689);
xor U18332 (N_18332,N_17523,N_17893);
or U18333 (N_18333,N_17657,N_17501);
or U18334 (N_18334,N_17818,N_17536);
and U18335 (N_18335,N_17811,N_17873);
nand U18336 (N_18336,N_17517,N_17890);
and U18337 (N_18337,N_17808,N_17809);
nor U18338 (N_18338,N_17801,N_17748);
xnor U18339 (N_18339,N_17590,N_17811);
or U18340 (N_18340,N_17929,N_17625);
nand U18341 (N_18341,N_17605,N_17699);
nand U18342 (N_18342,N_17932,N_17667);
or U18343 (N_18343,N_17928,N_17820);
or U18344 (N_18344,N_17616,N_17853);
nand U18345 (N_18345,N_17937,N_17562);
xnor U18346 (N_18346,N_17684,N_17639);
or U18347 (N_18347,N_17582,N_17618);
nor U18348 (N_18348,N_17755,N_17604);
nor U18349 (N_18349,N_17589,N_17949);
or U18350 (N_18350,N_17809,N_17861);
nand U18351 (N_18351,N_17703,N_17722);
nand U18352 (N_18352,N_17725,N_17557);
and U18353 (N_18353,N_17762,N_17954);
and U18354 (N_18354,N_17703,N_17612);
xor U18355 (N_18355,N_17599,N_17613);
nand U18356 (N_18356,N_17542,N_17653);
and U18357 (N_18357,N_17570,N_17612);
xor U18358 (N_18358,N_17795,N_17539);
nand U18359 (N_18359,N_17601,N_17812);
or U18360 (N_18360,N_17839,N_17956);
and U18361 (N_18361,N_17612,N_17649);
nor U18362 (N_18362,N_17994,N_17531);
and U18363 (N_18363,N_17920,N_17822);
xnor U18364 (N_18364,N_17909,N_17905);
nand U18365 (N_18365,N_17523,N_17833);
nand U18366 (N_18366,N_17509,N_17592);
or U18367 (N_18367,N_17506,N_17527);
nand U18368 (N_18368,N_17694,N_17695);
nor U18369 (N_18369,N_17619,N_17686);
and U18370 (N_18370,N_17702,N_17922);
and U18371 (N_18371,N_17894,N_17749);
nand U18372 (N_18372,N_17844,N_17532);
nor U18373 (N_18373,N_17636,N_17823);
xnor U18374 (N_18374,N_17712,N_17859);
nor U18375 (N_18375,N_17585,N_17776);
nor U18376 (N_18376,N_17559,N_17860);
or U18377 (N_18377,N_17734,N_17842);
or U18378 (N_18378,N_17555,N_17726);
nand U18379 (N_18379,N_17646,N_17562);
nor U18380 (N_18380,N_17664,N_17630);
nor U18381 (N_18381,N_17749,N_17800);
or U18382 (N_18382,N_17938,N_17515);
and U18383 (N_18383,N_17963,N_17914);
or U18384 (N_18384,N_17865,N_17780);
xor U18385 (N_18385,N_17769,N_17558);
or U18386 (N_18386,N_17643,N_17593);
xor U18387 (N_18387,N_17635,N_17854);
nand U18388 (N_18388,N_17951,N_17724);
xnor U18389 (N_18389,N_17982,N_17829);
xnor U18390 (N_18390,N_17854,N_17923);
nor U18391 (N_18391,N_17951,N_17740);
nand U18392 (N_18392,N_17843,N_17573);
nand U18393 (N_18393,N_17854,N_17536);
xnor U18394 (N_18394,N_17522,N_17833);
nand U18395 (N_18395,N_17564,N_17581);
nand U18396 (N_18396,N_17731,N_17966);
and U18397 (N_18397,N_17532,N_17652);
xor U18398 (N_18398,N_17880,N_17638);
nor U18399 (N_18399,N_17654,N_17675);
xor U18400 (N_18400,N_17593,N_17763);
and U18401 (N_18401,N_17952,N_17623);
xnor U18402 (N_18402,N_17723,N_17717);
or U18403 (N_18403,N_17549,N_17735);
and U18404 (N_18404,N_17973,N_17501);
or U18405 (N_18405,N_17811,N_17952);
or U18406 (N_18406,N_17795,N_17538);
xnor U18407 (N_18407,N_17760,N_17545);
nor U18408 (N_18408,N_17921,N_17603);
and U18409 (N_18409,N_17773,N_17697);
xor U18410 (N_18410,N_17965,N_17667);
nand U18411 (N_18411,N_17981,N_17853);
nand U18412 (N_18412,N_17610,N_17558);
or U18413 (N_18413,N_17513,N_17528);
xnor U18414 (N_18414,N_17851,N_17744);
xnor U18415 (N_18415,N_17667,N_17964);
nor U18416 (N_18416,N_17835,N_17871);
or U18417 (N_18417,N_17923,N_17982);
xnor U18418 (N_18418,N_17703,N_17832);
nor U18419 (N_18419,N_17619,N_17874);
xnor U18420 (N_18420,N_17874,N_17998);
and U18421 (N_18421,N_17936,N_17580);
nand U18422 (N_18422,N_17971,N_17865);
nor U18423 (N_18423,N_17986,N_17521);
nand U18424 (N_18424,N_17673,N_17756);
or U18425 (N_18425,N_17942,N_17964);
nor U18426 (N_18426,N_17857,N_17854);
or U18427 (N_18427,N_17632,N_17648);
and U18428 (N_18428,N_17742,N_17550);
nand U18429 (N_18429,N_17829,N_17653);
xor U18430 (N_18430,N_17964,N_17713);
nand U18431 (N_18431,N_17692,N_17678);
or U18432 (N_18432,N_17856,N_17637);
xnor U18433 (N_18433,N_17703,N_17763);
and U18434 (N_18434,N_17515,N_17572);
nor U18435 (N_18435,N_17840,N_17841);
and U18436 (N_18436,N_17558,N_17863);
nor U18437 (N_18437,N_17840,N_17906);
xor U18438 (N_18438,N_17676,N_17673);
xnor U18439 (N_18439,N_17906,N_17705);
or U18440 (N_18440,N_17651,N_17924);
and U18441 (N_18441,N_17524,N_17902);
nor U18442 (N_18442,N_17552,N_17872);
nand U18443 (N_18443,N_17761,N_17578);
nor U18444 (N_18444,N_17953,N_17550);
or U18445 (N_18445,N_17512,N_17629);
nand U18446 (N_18446,N_17896,N_17899);
xor U18447 (N_18447,N_17833,N_17503);
nor U18448 (N_18448,N_17767,N_17589);
nor U18449 (N_18449,N_17572,N_17967);
xor U18450 (N_18450,N_17860,N_17757);
or U18451 (N_18451,N_17815,N_17697);
nor U18452 (N_18452,N_17932,N_17747);
xor U18453 (N_18453,N_17515,N_17628);
or U18454 (N_18454,N_17691,N_17792);
or U18455 (N_18455,N_17786,N_17521);
or U18456 (N_18456,N_17525,N_17872);
or U18457 (N_18457,N_17841,N_17888);
nand U18458 (N_18458,N_17741,N_17593);
nand U18459 (N_18459,N_17953,N_17997);
nand U18460 (N_18460,N_17879,N_17745);
or U18461 (N_18461,N_17585,N_17748);
or U18462 (N_18462,N_17942,N_17660);
nand U18463 (N_18463,N_17992,N_17877);
xor U18464 (N_18464,N_17712,N_17899);
nor U18465 (N_18465,N_17551,N_17842);
nor U18466 (N_18466,N_17736,N_17574);
or U18467 (N_18467,N_17720,N_17580);
nor U18468 (N_18468,N_17730,N_17905);
or U18469 (N_18469,N_17502,N_17836);
and U18470 (N_18470,N_17920,N_17569);
nor U18471 (N_18471,N_17961,N_17787);
nand U18472 (N_18472,N_17997,N_17819);
xnor U18473 (N_18473,N_17746,N_17911);
and U18474 (N_18474,N_17871,N_17679);
nor U18475 (N_18475,N_17736,N_17768);
nand U18476 (N_18476,N_17908,N_17787);
nor U18477 (N_18477,N_17971,N_17815);
nor U18478 (N_18478,N_17712,N_17774);
nand U18479 (N_18479,N_17998,N_17984);
or U18480 (N_18480,N_17510,N_17587);
nor U18481 (N_18481,N_17854,N_17829);
nor U18482 (N_18482,N_17651,N_17949);
xnor U18483 (N_18483,N_17718,N_17881);
and U18484 (N_18484,N_17529,N_17929);
nor U18485 (N_18485,N_17503,N_17804);
nand U18486 (N_18486,N_17653,N_17649);
or U18487 (N_18487,N_17709,N_17757);
xor U18488 (N_18488,N_17786,N_17844);
and U18489 (N_18489,N_17612,N_17964);
or U18490 (N_18490,N_17616,N_17904);
nor U18491 (N_18491,N_17555,N_17849);
xor U18492 (N_18492,N_17844,N_17752);
or U18493 (N_18493,N_17640,N_17763);
xnor U18494 (N_18494,N_17917,N_17717);
nor U18495 (N_18495,N_17736,N_17867);
and U18496 (N_18496,N_17764,N_17630);
or U18497 (N_18497,N_17775,N_17968);
or U18498 (N_18498,N_17911,N_17872);
or U18499 (N_18499,N_17777,N_17555);
and U18500 (N_18500,N_18351,N_18419);
nand U18501 (N_18501,N_18089,N_18068);
and U18502 (N_18502,N_18463,N_18183);
nor U18503 (N_18503,N_18423,N_18178);
nor U18504 (N_18504,N_18413,N_18016);
and U18505 (N_18505,N_18064,N_18202);
xnor U18506 (N_18506,N_18360,N_18163);
nand U18507 (N_18507,N_18253,N_18464);
or U18508 (N_18508,N_18263,N_18076);
nand U18509 (N_18509,N_18218,N_18245);
or U18510 (N_18510,N_18301,N_18036);
and U18511 (N_18511,N_18269,N_18024);
or U18512 (N_18512,N_18346,N_18223);
nor U18513 (N_18513,N_18381,N_18081);
nand U18514 (N_18514,N_18153,N_18000);
and U18515 (N_18515,N_18227,N_18496);
nand U18516 (N_18516,N_18449,N_18330);
nand U18517 (N_18517,N_18112,N_18184);
nor U18518 (N_18518,N_18467,N_18437);
nand U18519 (N_18519,N_18082,N_18242);
xnor U18520 (N_18520,N_18493,N_18047);
and U18521 (N_18521,N_18215,N_18279);
or U18522 (N_18522,N_18239,N_18280);
nor U18523 (N_18523,N_18389,N_18445);
or U18524 (N_18524,N_18088,N_18264);
or U18525 (N_18525,N_18061,N_18241);
nand U18526 (N_18526,N_18188,N_18379);
or U18527 (N_18527,N_18332,N_18075);
nor U18528 (N_18528,N_18203,N_18315);
or U18529 (N_18529,N_18392,N_18087);
nor U18530 (N_18530,N_18080,N_18362);
nor U18531 (N_18531,N_18273,N_18326);
or U18532 (N_18532,N_18294,N_18124);
nand U18533 (N_18533,N_18451,N_18231);
and U18534 (N_18534,N_18265,N_18444);
nand U18535 (N_18535,N_18165,N_18296);
xor U18536 (N_18536,N_18386,N_18155);
nand U18537 (N_18537,N_18149,N_18492);
nor U18538 (N_18538,N_18353,N_18246);
and U18539 (N_18539,N_18143,N_18176);
and U18540 (N_18540,N_18150,N_18342);
nor U18541 (N_18541,N_18491,N_18040);
nor U18542 (N_18542,N_18222,N_18131);
xnor U18543 (N_18543,N_18441,N_18205);
nand U18544 (N_18544,N_18479,N_18219);
and U18545 (N_18545,N_18236,N_18406);
nor U18546 (N_18546,N_18250,N_18104);
nand U18547 (N_18547,N_18105,N_18375);
nand U18548 (N_18548,N_18192,N_18229);
and U18549 (N_18549,N_18038,N_18424);
nor U18550 (N_18550,N_18216,N_18120);
and U18551 (N_18551,N_18430,N_18457);
or U18552 (N_18552,N_18123,N_18001);
nand U18553 (N_18553,N_18255,N_18220);
xnor U18554 (N_18554,N_18349,N_18022);
and U18555 (N_18555,N_18237,N_18262);
or U18556 (N_18556,N_18108,N_18116);
nand U18557 (N_18557,N_18168,N_18233);
nand U18558 (N_18558,N_18478,N_18495);
or U18559 (N_18559,N_18323,N_18235);
and U18560 (N_18560,N_18044,N_18136);
nor U18561 (N_18561,N_18488,N_18110);
nand U18562 (N_18562,N_18133,N_18432);
nor U18563 (N_18563,N_18194,N_18157);
xnor U18564 (N_18564,N_18293,N_18321);
xnor U18565 (N_18565,N_18204,N_18405);
or U18566 (N_18566,N_18361,N_18093);
nor U18567 (N_18567,N_18051,N_18209);
or U18568 (N_18568,N_18435,N_18476);
nor U18569 (N_18569,N_18130,N_18114);
xnor U18570 (N_18570,N_18489,N_18248);
and U18571 (N_18571,N_18308,N_18128);
nor U18572 (N_18572,N_18487,N_18278);
and U18573 (N_18573,N_18207,N_18456);
nand U18574 (N_18574,N_18345,N_18159);
nand U18575 (N_18575,N_18376,N_18055);
nor U18576 (N_18576,N_18244,N_18023);
or U18577 (N_18577,N_18102,N_18228);
nand U18578 (N_18578,N_18063,N_18459);
nor U18579 (N_18579,N_18497,N_18304);
nand U18580 (N_18580,N_18190,N_18365);
or U18581 (N_18581,N_18210,N_18213);
xnor U18582 (N_18582,N_18395,N_18201);
nand U18583 (N_18583,N_18221,N_18206);
or U18584 (N_18584,N_18359,N_18439);
or U18585 (N_18585,N_18170,N_18230);
nand U18586 (N_18586,N_18310,N_18092);
nand U18587 (N_18587,N_18135,N_18005);
nand U18588 (N_18588,N_18226,N_18481);
nand U18589 (N_18589,N_18084,N_18050);
nor U18590 (N_18590,N_18431,N_18167);
nor U18591 (N_18591,N_18098,N_18035);
xor U18592 (N_18592,N_18161,N_18341);
nor U18593 (N_18593,N_18097,N_18461);
xnor U18594 (N_18594,N_18447,N_18101);
nor U18595 (N_18595,N_18391,N_18307);
nor U18596 (N_18596,N_18193,N_18440);
xor U18597 (N_18597,N_18390,N_18402);
or U18598 (N_18598,N_18212,N_18348);
xor U18599 (N_18599,N_18060,N_18407);
nand U18600 (N_18600,N_18470,N_18319);
nor U18601 (N_18601,N_18281,N_18297);
xor U18602 (N_18602,N_18383,N_18275);
xnor U18603 (N_18603,N_18141,N_18287);
nor U18604 (N_18604,N_18090,N_18498);
xor U18605 (N_18605,N_18303,N_18122);
or U18606 (N_18606,N_18003,N_18409);
nand U18607 (N_18607,N_18134,N_18106);
and U18608 (N_18608,N_18288,N_18306);
xnor U18609 (N_18609,N_18340,N_18015);
nand U18610 (N_18610,N_18477,N_18026);
and U18611 (N_18611,N_18354,N_18388);
or U18612 (N_18612,N_18225,N_18350);
nor U18613 (N_18613,N_18410,N_18078);
or U18614 (N_18614,N_18118,N_18454);
and U18615 (N_18615,N_18455,N_18152);
nand U18616 (N_18616,N_18238,N_18267);
nor U18617 (N_18617,N_18010,N_18119);
and U18618 (N_18618,N_18335,N_18300);
nand U18619 (N_18619,N_18347,N_18420);
and U18620 (N_18620,N_18286,N_18327);
nor U18621 (N_18621,N_18305,N_18107);
xor U18622 (N_18622,N_18031,N_18083);
xor U18623 (N_18623,N_18169,N_18313);
nor U18624 (N_18624,N_18352,N_18485);
xor U18625 (N_18625,N_18195,N_18462);
nand U18626 (N_18626,N_18247,N_18385);
xnor U18627 (N_18627,N_18151,N_18382);
nand U18628 (N_18628,N_18387,N_18041);
and U18629 (N_18629,N_18077,N_18298);
nor U18630 (N_18630,N_18109,N_18418);
or U18631 (N_18631,N_18336,N_18232);
and U18632 (N_18632,N_18025,N_18356);
nor U18633 (N_18633,N_18324,N_18028);
or U18634 (N_18634,N_18191,N_18156);
nand U18635 (N_18635,N_18126,N_18458);
and U18636 (N_18636,N_18013,N_18033);
and U18637 (N_18637,N_18261,N_18096);
and U18638 (N_18638,N_18070,N_18343);
nand U18639 (N_18639,N_18021,N_18069);
nor U18640 (N_18640,N_18249,N_18062);
and U18641 (N_18641,N_18309,N_18117);
xnor U18642 (N_18642,N_18311,N_18052);
or U18643 (N_18643,N_18045,N_18364);
and U18644 (N_18644,N_18295,N_18007);
nand U18645 (N_18645,N_18002,N_18370);
nor U18646 (N_18646,N_18282,N_18085);
nor U18647 (N_18647,N_18373,N_18397);
and U18648 (N_18648,N_18322,N_18466);
xor U18649 (N_18649,N_18056,N_18127);
nor U18650 (N_18650,N_18179,N_18270);
nor U18651 (N_18651,N_18317,N_18049);
nor U18652 (N_18652,N_18048,N_18328);
or U18653 (N_18653,N_18144,N_18164);
nor U18654 (N_18654,N_18411,N_18034);
nor U18655 (N_18655,N_18369,N_18039);
nand U18656 (N_18656,N_18436,N_18032);
nand U18657 (N_18657,N_18465,N_18200);
and U18658 (N_18658,N_18393,N_18181);
or U18659 (N_18659,N_18208,N_18234);
and U18660 (N_18660,N_18312,N_18329);
xor U18661 (N_18661,N_18171,N_18029);
nor U18662 (N_18662,N_18214,N_18079);
nand U18663 (N_18663,N_18408,N_18433);
nand U18664 (N_18664,N_18367,N_18443);
xor U18665 (N_18665,N_18429,N_18442);
nand U18666 (N_18666,N_18103,N_18030);
nor U18667 (N_18667,N_18042,N_18158);
xnor U18668 (N_18668,N_18469,N_18318);
nand U18669 (N_18669,N_18499,N_18371);
nand U18670 (N_18670,N_18357,N_18072);
nor U18671 (N_18671,N_18132,N_18425);
and U18672 (N_18672,N_18073,N_18338);
xnor U18673 (N_18673,N_18115,N_18086);
or U18674 (N_18674,N_18285,N_18074);
or U18675 (N_18675,N_18162,N_18276);
nand U18676 (N_18676,N_18434,N_18412);
and U18677 (N_18677,N_18291,N_18460);
nor U18678 (N_18678,N_18139,N_18289);
nand U18679 (N_18679,N_18320,N_18111);
nand U18680 (N_18680,N_18472,N_18018);
nor U18681 (N_18681,N_18421,N_18417);
nor U18682 (N_18682,N_18172,N_18091);
nor U18683 (N_18683,N_18027,N_18254);
and U18684 (N_18684,N_18145,N_18177);
xor U18685 (N_18685,N_18009,N_18438);
xor U18686 (N_18686,N_18416,N_18271);
and U18687 (N_18687,N_18138,N_18266);
xor U18688 (N_18688,N_18358,N_18196);
and U18689 (N_18689,N_18166,N_18012);
xnor U18690 (N_18690,N_18173,N_18428);
and U18691 (N_18691,N_18316,N_18099);
or U18692 (N_18692,N_18125,N_18259);
nand U18693 (N_18693,N_18272,N_18140);
nand U18694 (N_18694,N_18147,N_18475);
or U18695 (N_18695,N_18199,N_18473);
xor U18696 (N_18696,N_18453,N_18059);
nand U18697 (N_18697,N_18331,N_18251);
and U18698 (N_18698,N_18160,N_18004);
and U18699 (N_18699,N_18474,N_18426);
nand U18700 (N_18700,N_18368,N_18121);
nor U18701 (N_18701,N_18014,N_18484);
nand U18702 (N_18702,N_18401,N_18268);
or U18703 (N_18703,N_18019,N_18174);
xnor U18704 (N_18704,N_18008,N_18129);
nand U18705 (N_18705,N_18274,N_18355);
and U18706 (N_18706,N_18483,N_18017);
nand U18707 (N_18707,N_18185,N_18175);
and U18708 (N_18708,N_18053,N_18224);
or U18709 (N_18709,N_18283,N_18258);
nand U18710 (N_18710,N_18187,N_18180);
or U18711 (N_18711,N_18020,N_18384);
or U18712 (N_18712,N_18422,N_18054);
and U18713 (N_18713,N_18011,N_18257);
and U18714 (N_18714,N_18100,N_18414);
and U18715 (N_18715,N_18182,N_18284);
or U18716 (N_18716,N_18066,N_18374);
nand U18717 (N_18717,N_18094,N_18146);
nor U18718 (N_18718,N_18377,N_18067);
and U18719 (N_18719,N_18046,N_18482);
and U18720 (N_18720,N_18366,N_18372);
xor U18721 (N_18721,N_18189,N_18113);
nand U18722 (N_18722,N_18471,N_18243);
nor U18723 (N_18723,N_18142,N_18334);
nand U18724 (N_18724,N_18148,N_18396);
or U18725 (N_18725,N_18333,N_18198);
nand U18726 (N_18726,N_18043,N_18256);
nand U18727 (N_18727,N_18299,N_18065);
nor U18728 (N_18728,N_18314,N_18494);
xor U18729 (N_18729,N_18240,N_18380);
or U18730 (N_18730,N_18337,N_18398);
and U18731 (N_18731,N_18378,N_18137);
or U18732 (N_18732,N_18290,N_18403);
nand U18733 (N_18733,N_18450,N_18427);
and U18734 (N_18734,N_18452,N_18154);
and U18735 (N_18735,N_18490,N_18344);
and U18736 (N_18736,N_18058,N_18260);
nand U18737 (N_18737,N_18071,N_18486);
or U18738 (N_18738,N_18186,N_18448);
xnor U18739 (N_18739,N_18277,N_18006);
and U18740 (N_18740,N_18480,N_18211);
or U18741 (N_18741,N_18292,N_18399);
and U18742 (N_18742,N_18415,N_18197);
and U18743 (N_18743,N_18400,N_18404);
xor U18744 (N_18744,N_18339,N_18057);
xnor U18745 (N_18745,N_18217,N_18095);
and U18746 (N_18746,N_18325,N_18302);
and U18747 (N_18747,N_18468,N_18037);
and U18748 (N_18748,N_18363,N_18446);
or U18749 (N_18749,N_18252,N_18394);
nor U18750 (N_18750,N_18419,N_18305);
or U18751 (N_18751,N_18468,N_18347);
xnor U18752 (N_18752,N_18258,N_18214);
or U18753 (N_18753,N_18114,N_18153);
nor U18754 (N_18754,N_18187,N_18323);
xnor U18755 (N_18755,N_18186,N_18099);
nand U18756 (N_18756,N_18481,N_18401);
nor U18757 (N_18757,N_18146,N_18260);
or U18758 (N_18758,N_18453,N_18171);
nor U18759 (N_18759,N_18289,N_18025);
or U18760 (N_18760,N_18211,N_18360);
xnor U18761 (N_18761,N_18005,N_18057);
and U18762 (N_18762,N_18400,N_18381);
xor U18763 (N_18763,N_18089,N_18041);
nor U18764 (N_18764,N_18036,N_18398);
xnor U18765 (N_18765,N_18094,N_18065);
or U18766 (N_18766,N_18138,N_18176);
or U18767 (N_18767,N_18335,N_18476);
xnor U18768 (N_18768,N_18047,N_18449);
or U18769 (N_18769,N_18370,N_18202);
and U18770 (N_18770,N_18204,N_18358);
or U18771 (N_18771,N_18433,N_18162);
and U18772 (N_18772,N_18461,N_18426);
nor U18773 (N_18773,N_18447,N_18443);
and U18774 (N_18774,N_18033,N_18306);
nor U18775 (N_18775,N_18218,N_18277);
or U18776 (N_18776,N_18470,N_18390);
or U18777 (N_18777,N_18025,N_18140);
nor U18778 (N_18778,N_18049,N_18354);
xnor U18779 (N_18779,N_18411,N_18473);
nor U18780 (N_18780,N_18257,N_18272);
or U18781 (N_18781,N_18360,N_18086);
or U18782 (N_18782,N_18109,N_18176);
nand U18783 (N_18783,N_18411,N_18189);
and U18784 (N_18784,N_18058,N_18178);
nor U18785 (N_18785,N_18091,N_18188);
xnor U18786 (N_18786,N_18072,N_18150);
nand U18787 (N_18787,N_18182,N_18064);
xor U18788 (N_18788,N_18424,N_18440);
nand U18789 (N_18789,N_18288,N_18329);
or U18790 (N_18790,N_18385,N_18258);
nor U18791 (N_18791,N_18153,N_18248);
xor U18792 (N_18792,N_18225,N_18321);
and U18793 (N_18793,N_18278,N_18111);
and U18794 (N_18794,N_18169,N_18219);
nor U18795 (N_18795,N_18498,N_18042);
or U18796 (N_18796,N_18220,N_18310);
nand U18797 (N_18797,N_18148,N_18025);
xor U18798 (N_18798,N_18108,N_18002);
xnor U18799 (N_18799,N_18311,N_18399);
nor U18800 (N_18800,N_18454,N_18408);
nand U18801 (N_18801,N_18454,N_18349);
and U18802 (N_18802,N_18214,N_18397);
or U18803 (N_18803,N_18125,N_18214);
nor U18804 (N_18804,N_18020,N_18006);
xnor U18805 (N_18805,N_18368,N_18486);
nand U18806 (N_18806,N_18416,N_18381);
or U18807 (N_18807,N_18151,N_18059);
or U18808 (N_18808,N_18203,N_18460);
nor U18809 (N_18809,N_18464,N_18002);
and U18810 (N_18810,N_18243,N_18215);
or U18811 (N_18811,N_18077,N_18303);
xnor U18812 (N_18812,N_18147,N_18424);
nor U18813 (N_18813,N_18452,N_18101);
xor U18814 (N_18814,N_18131,N_18265);
or U18815 (N_18815,N_18077,N_18149);
and U18816 (N_18816,N_18105,N_18458);
nand U18817 (N_18817,N_18063,N_18388);
or U18818 (N_18818,N_18025,N_18481);
nand U18819 (N_18819,N_18346,N_18336);
and U18820 (N_18820,N_18360,N_18081);
xor U18821 (N_18821,N_18057,N_18247);
nand U18822 (N_18822,N_18045,N_18279);
nand U18823 (N_18823,N_18131,N_18482);
nand U18824 (N_18824,N_18022,N_18473);
xnor U18825 (N_18825,N_18303,N_18374);
nand U18826 (N_18826,N_18296,N_18287);
or U18827 (N_18827,N_18163,N_18384);
or U18828 (N_18828,N_18170,N_18456);
or U18829 (N_18829,N_18053,N_18357);
nor U18830 (N_18830,N_18248,N_18039);
nand U18831 (N_18831,N_18326,N_18485);
xnor U18832 (N_18832,N_18485,N_18428);
xor U18833 (N_18833,N_18476,N_18280);
xor U18834 (N_18834,N_18458,N_18185);
nor U18835 (N_18835,N_18110,N_18452);
nor U18836 (N_18836,N_18300,N_18034);
and U18837 (N_18837,N_18314,N_18295);
or U18838 (N_18838,N_18455,N_18304);
and U18839 (N_18839,N_18126,N_18177);
xnor U18840 (N_18840,N_18404,N_18017);
nor U18841 (N_18841,N_18206,N_18409);
or U18842 (N_18842,N_18373,N_18154);
xor U18843 (N_18843,N_18430,N_18452);
xnor U18844 (N_18844,N_18357,N_18486);
xor U18845 (N_18845,N_18154,N_18345);
nand U18846 (N_18846,N_18265,N_18297);
or U18847 (N_18847,N_18435,N_18096);
nand U18848 (N_18848,N_18229,N_18291);
and U18849 (N_18849,N_18445,N_18039);
or U18850 (N_18850,N_18247,N_18001);
or U18851 (N_18851,N_18003,N_18052);
and U18852 (N_18852,N_18265,N_18181);
or U18853 (N_18853,N_18216,N_18113);
nand U18854 (N_18854,N_18383,N_18246);
or U18855 (N_18855,N_18448,N_18365);
nor U18856 (N_18856,N_18466,N_18397);
nor U18857 (N_18857,N_18056,N_18081);
xnor U18858 (N_18858,N_18314,N_18457);
nor U18859 (N_18859,N_18463,N_18404);
nand U18860 (N_18860,N_18014,N_18251);
and U18861 (N_18861,N_18076,N_18168);
nor U18862 (N_18862,N_18132,N_18117);
nor U18863 (N_18863,N_18053,N_18103);
or U18864 (N_18864,N_18274,N_18284);
nand U18865 (N_18865,N_18073,N_18225);
and U18866 (N_18866,N_18443,N_18029);
or U18867 (N_18867,N_18026,N_18056);
and U18868 (N_18868,N_18058,N_18111);
and U18869 (N_18869,N_18352,N_18175);
nand U18870 (N_18870,N_18227,N_18163);
and U18871 (N_18871,N_18393,N_18420);
or U18872 (N_18872,N_18458,N_18199);
nand U18873 (N_18873,N_18150,N_18369);
or U18874 (N_18874,N_18078,N_18061);
and U18875 (N_18875,N_18147,N_18458);
nand U18876 (N_18876,N_18212,N_18015);
or U18877 (N_18877,N_18449,N_18043);
nand U18878 (N_18878,N_18371,N_18118);
nand U18879 (N_18879,N_18267,N_18465);
nand U18880 (N_18880,N_18265,N_18461);
or U18881 (N_18881,N_18328,N_18366);
or U18882 (N_18882,N_18415,N_18407);
nand U18883 (N_18883,N_18074,N_18182);
or U18884 (N_18884,N_18020,N_18081);
xnor U18885 (N_18885,N_18311,N_18430);
or U18886 (N_18886,N_18466,N_18437);
nand U18887 (N_18887,N_18203,N_18361);
xnor U18888 (N_18888,N_18466,N_18223);
nand U18889 (N_18889,N_18270,N_18300);
nand U18890 (N_18890,N_18321,N_18077);
or U18891 (N_18891,N_18423,N_18009);
nand U18892 (N_18892,N_18282,N_18161);
nor U18893 (N_18893,N_18322,N_18325);
and U18894 (N_18894,N_18326,N_18328);
xnor U18895 (N_18895,N_18067,N_18450);
nor U18896 (N_18896,N_18307,N_18453);
xnor U18897 (N_18897,N_18296,N_18181);
and U18898 (N_18898,N_18053,N_18047);
nor U18899 (N_18899,N_18044,N_18440);
or U18900 (N_18900,N_18258,N_18121);
and U18901 (N_18901,N_18195,N_18409);
xor U18902 (N_18902,N_18009,N_18462);
nand U18903 (N_18903,N_18082,N_18303);
or U18904 (N_18904,N_18297,N_18017);
and U18905 (N_18905,N_18151,N_18226);
or U18906 (N_18906,N_18093,N_18387);
xnor U18907 (N_18907,N_18083,N_18139);
nand U18908 (N_18908,N_18279,N_18076);
or U18909 (N_18909,N_18361,N_18144);
and U18910 (N_18910,N_18270,N_18417);
or U18911 (N_18911,N_18010,N_18342);
or U18912 (N_18912,N_18422,N_18169);
and U18913 (N_18913,N_18063,N_18300);
xor U18914 (N_18914,N_18360,N_18426);
or U18915 (N_18915,N_18134,N_18146);
or U18916 (N_18916,N_18461,N_18498);
nor U18917 (N_18917,N_18434,N_18214);
and U18918 (N_18918,N_18078,N_18214);
or U18919 (N_18919,N_18152,N_18132);
nand U18920 (N_18920,N_18171,N_18223);
nand U18921 (N_18921,N_18105,N_18484);
nor U18922 (N_18922,N_18172,N_18393);
or U18923 (N_18923,N_18179,N_18001);
and U18924 (N_18924,N_18429,N_18002);
and U18925 (N_18925,N_18178,N_18131);
xor U18926 (N_18926,N_18144,N_18169);
or U18927 (N_18927,N_18430,N_18091);
nand U18928 (N_18928,N_18291,N_18348);
and U18929 (N_18929,N_18390,N_18010);
and U18930 (N_18930,N_18346,N_18448);
or U18931 (N_18931,N_18111,N_18386);
or U18932 (N_18932,N_18209,N_18123);
and U18933 (N_18933,N_18343,N_18215);
and U18934 (N_18934,N_18477,N_18315);
xnor U18935 (N_18935,N_18184,N_18386);
nand U18936 (N_18936,N_18399,N_18070);
xnor U18937 (N_18937,N_18383,N_18292);
or U18938 (N_18938,N_18144,N_18154);
nor U18939 (N_18939,N_18009,N_18366);
or U18940 (N_18940,N_18184,N_18040);
nand U18941 (N_18941,N_18450,N_18162);
and U18942 (N_18942,N_18108,N_18317);
or U18943 (N_18943,N_18328,N_18231);
xor U18944 (N_18944,N_18476,N_18328);
nand U18945 (N_18945,N_18407,N_18091);
and U18946 (N_18946,N_18168,N_18106);
nand U18947 (N_18947,N_18354,N_18164);
nor U18948 (N_18948,N_18312,N_18488);
or U18949 (N_18949,N_18132,N_18131);
nand U18950 (N_18950,N_18355,N_18053);
nand U18951 (N_18951,N_18409,N_18298);
xor U18952 (N_18952,N_18106,N_18469);
and U18953 (N_18953,N_18087,N_18051);
nor U18954 (N_18954,N_18234,N_18199);
nor U18955 (N_18955,N_18111,N_18025);
xnor U18956 (N_18956,N_18463,N_18293);
xor U18957 (N_18957,N_18015,N_18363);
or U18958 (N_18958,N_18277,N_18035);
nand U18959 (N_18959,N_18059,N_18116);
or U18960 (N_18960,N_18416,N_18433);
and U18961 (N_18961,N_18287,N_18076);
nor U18962 (N_18962,N_18022,N_18372);
and U18963 (N_18963,N_18009,N_18005);
or U18964 (N_18964,N_18108,N_18281);
xnor U18965 (N_18965,N_18015,N_18091);
and U18966 (N_18966,N_18189,N_18203);
and U18967 (N_18967,N_18166,N_18242);
nor U18968 (N_18968,N_18024,N_18394);
nand U18969 (N_18969,N_18181,N_18331);
nor U18970 (N_18970,N_18401,N_18149);
and U18971 (N_18971,N_18284,N_18458);
xnor U18972 (N_18972,N_18315,N_18272);
and U18973 (N_18973,N_18085,N_18135);
nand U18974 (N_18974,N_18150,N_18152);
and U18975 (N_18975,N_18285,N_18078);
xor U18976 (N_18976,N_18467,N_18423);
xnor U18977 (N_18977,N_18271,N_18377);
or U18978 (N_18978,N_18451,N_18112);
nor U18979 (N_18979,N_18321,N_18363);
or U18980 (N_18980,N_18494,N_18337);
and U18981 (N_18981,N_18167,N_18152);
and U18982 (N_18982,N_18263,N_18297);
nand U18983 (N_18983,N_18239,N_18259);
and U18984 (N_18984,N_18087,N_18488);
nor U18985 (N_18985,N_18077,N_18486);
and U18986 (N_18986,N_18005,N_18465);
nor U18987 (N_18987,N_18411,N_18423);
or U18988 (N_18988,N_18338,N_18280);
xor U18989 (N_18989,N_18043,N_18275);
and U18990 (N_18990,N_18037,N_18349);
or U18991 (N_18991,N_18271,N_18240);
nor U18992 (N_18992,N_18439,N_18392);
and U18993 (N_18993,N_18274,N_18132);
nand U18994 (N_18994,N_18091,N_18205);
and U18995 (N_18995,N_18270,N_18457);
or U18996 (N_18996,N_18225,N_18472);
or U18997 (N_18997,N_18068,N_18121);
and U18998 (N_18998,N_18162,N_18253);
xnor U18999 (N_18999,N_18064,N_18025);
xnor U19000 (N_19000,N_18551,N_18799);
and U19001 (N_19001,N_18505,N_18969);
and U19002 (N_19002,N_18849,N_18874);
nor U19003 (N_19003,N_18747,N_18939);
nor U19004 (N_19004,N_18982,N_18852);
and U19005 (N_19005,N_18909,N_18952);
xnor U19006 (N_19006,N_18807,N_18640);
nor U19007 (N_19007,N_18834,N_18615);
or U19008 (N_19008,N_18838,N_18641);
nor U19009 (N_19009,N_18608,N_18637);
xor U19010 (N_19010,N_18787,N_18789);
or U19011 (N_19011,N_18703,N_18788);
and U19012 (N_19012,N_18522,N_18652);
nor U19013 (N_19013,N_18835,N_18613);
nand U19014 (N_19014,N_18825,N_18671);
nand U19015 (N_19015,N_18837,N_18970);
nor U19016 (N_19016,N_18604,N_18512);
nor U19017 (N_19017,N_18539,N_18756);
and U19018 (N_19018,N_18688,N_18518);
or U19019 (N_19019,N_18752,N_18962);
nor U19020 (N_19020,N_18980,N_18612);
nand U19021 (N_19021,N_18684,N_18569);
and U19022 (N_19022,N_18951,N_18664);
or U19023 (N_19023,N_18857,N_18651);
nand U19024 (N_19024,N_18721,N_18996);
xnor U19025 (N_19025,N_18646,N_18830);
xor U19026 (N_19026,N_18736,N_18854);
nor U19027 (N_19027,N_18848,N_18986);
nor U19028 (N_19028,N_18773,N_18727);
or U19029 (N_19029,N_18643,N_18546);
or U19030 (N_19030,N_18508,N_18751);
and U19031 (N_19031,N_18618,N_18655);
nand U19032 (N_19032,N_18988,N_18829);
or U19033 (N_19033,N_18626,N_18908);
or U19034 (N_19034,N_18919,N_18631);
nor U19035 (N_19035,N_18913,N_18823);
or U19036 (N_19036,N_18964,N_18845);
xnor U19037 (N_19037,N_18867,N_18621);
and U19038 (N_19038,N_18759,N_18785);
nand U19039 (N_19039,N_18850,N_18740);
nor U19040 (N_19040,N_18905,N_18635);
and U19041 (N_19041,N_18793,N_18696);
xor U19042 (N_19042,N_18766,N_18983);
nand U19043 (N_19043,N_18953,N_18573);
xnor U19044 (N_19044,N_18761,N_18606);
nand U19045 (N_19045,N_18950,N_18550);
nor U19046 (N_19046,N_18956,N_18517);
nand U19047 (N_19047,N_18661,N_18581);
nand U19048 (N_19048,N_18588,N_18519);
nor U19049 (N_19049,N_18610,N_18527);
nand U19050 (N_19050,N_18899,N_18683);
and U19051 (N_19051,N_18995,N_18973);
xor U19052 (N_19052,N_18593,N_18730);
xor U19053 (N_19053,N_18836,N_18790);
nand U19054 (N_19054,N_18680,N_18911);
xnor U19055 (N_19055,N_18630,N_18743);
and U19056 (N_19056,N_18938,N_18731);
or U19057 (N_19057,N_18757,N_18741);
xor U19058 (N_19058,N_18803,N_18622);
nand U19059 (N_19059,N_18528,N_18726);
xor U19060 (N_19060,N_18690,N_18561);
xor U19061 (N_19061,N_18910,N_18563);
nand U19062 (N_19062,N_18673,N_18859);
or U19063 (N_19063,N_18520,N_18885);
nor U19064 (N_19064,N_18697,N_18605);
nand U19065 (N_19065,N_18501,N_18532);
nor U19066 (N_19066,N_18572,N_18587);
nor U19067 (N_19067,N_18877,N_18792);
and U19068 (N_19068,N_18875,N_18868);
nand U19069 (N_19069,N_18500,N_18750);
nand U19070 (N_19070,N_18960,N_18745);
xor U19071 (N_19071,N_18559,N_18709);
nor U19072 (N_19072,N_18904,N_18704);
or U19073 (N_19073,N_18864,N_18639);
nand U19074 (N_19074,N_18556,N_18524);
or U19075 (N_19075,N_18742,N_18663);
xor U19076 (N_19076,N_18974,N_18928);
nor U19077 (N_19077,N_18933,N_18549);
or U19078 (N_19078,N_18544,N_18797);
or U19079 (N_19079,N_18695,N_18841);
and U19080 (N_19080,N_18887,N_18853);
nor U19081 (N_19081,N_18707,N_18659);
nand U19082 (N_19082,N_18883,N_18945);
or U19083 (N_19083,N_18987,N_18708);
nand U19084 (N_19084,N_18821,N_18884);
or U19085 (N_19085,N_18820,N_18774);
nor U19086 (N_19086,N_18669,N_18922);
nand U19087 (N_19087,N_18513,N_18802);
or U19088 (N_19088,N_18576,N_18586);
or U19089 (N_19089,N_18994,N_18819);
nand U19090 (N_19090,N_18916,N_18907);
or U19091 (N_19091,N_18623,N_18882);
nand U19092 (N_19092,N_18968,N_18993);
xor U19093 (N_19093,N_18846,N_18775);
xor U19094 (N_19094,N_18724,N_18914);
nor U19095 (N_19095,N_18794,N_18542);
and U19096 (N_19096,N_18509,N_18831);
nor U19097 (N_19097,N_18634,N_18525);
and U19098 (N_19098,N_18739,N_18676);
or U19099 (N_19099,N_18959,N_18530);
xor U19100 (N_19100,N_18516,N_18729);
or U19101 (N_19101,N_18903,N_18981);
nor U19102 (N_19102,N_18575,N_18511);
nor U19103 (N_19103,N_18538,N_18900);
or U19104 (N_19104,N_18976,N_18732);
and U19105 (N_19105,N_18706,N_18780);
and U19106 (N_19106,N_18737,N_18689);
nand U19107 (N_19107,N_18601,N_18947);
and U19108 (N_19108,N_18814,N_18585);
and U19109 (N_19109,N_18624,N_18584);
and U19110 (N_19110,N_18557,N_18963);
or U19111 (N_19111,N_18578,N_18860);
or U19112 (N_19112,N_18832,N_18934);
and U19113 (N_19113,N_18529,N_18590);
nor U19114 (N_19114,N_18772,N_18515);
nand U19115 (N_19115,N_18598,N_18826);
or U19116 (N_19116,N_18535,N_18504);
nand U19117 (N_19117,N_18712,N_18733);
nor U19118 (N_19118,N_18713,N_18547);
nor U19119 (N_19119,N_18784,N_18582);
nand U19120 (N_19120,N_18560,N_18992);
nor U19121 (N_19121,N_18754,N_18897);
nand U19122 (N_19122,N_18861,N_18863);
xnor U19123 (N_19123,N_18870,N_18924);
nand U19124 (N_19124,N_18923,N_18577);
xnor U19125 (N_19125,N_18796,N_18523);
and U19126 (N_19126,N_18674,N_18991);
xnor U19127 (N_19127,N_18744,N_18906);
and U19128 (N_19128,N_18779,N_18565);
nor U19129 (N_19129,N_18763,N_18891);
and U19130 (N_19130,N_18912,N_18961);
nand U19131 (N_19131,N_18650,N_18878);
nor U19132 (N_19132,N_18989,N_18999);
nand U19133 (N_19133,N_18662,N_18943);
and U19134 (N_19134,N_18510,N_18812);
or U19135 (N_19135,N_18687,N_18958);
nor U19136 (N_19136,N_18722,N_18638);
or U19137 (N_19137,N_18711,N_18665);
nand U19138 (N_19138,N_18701,N_18648);
or U19139 (N_19139,N_18681,N_18816);
or U19140 (N_19140,N_18723,N_18589);
nor U19141 (N_19141,N_18506,N_18815);
xnor U19142 (N_19142,N_18558,N_18771);
or U19143 (N_19143,N_18984,N_18915);
and U19144 (N_19144,N_18918,N_18998);
nand U19145 (N_19145,N_18675,N_18768);
xor U19146 (N_19146,N_18978,N_18795);
nor U19147 (N_19147,N_18791,N_18843);
or U19148 (N_19148,N_18925,N_18948);
and U19149 (N_19149,N_18886,N_18818);
and U19150 (N_19150,N_18869,N_18502);
nand U19151 (N_19151,N_18540,N_18896);
nand U19152 (N_19152,N_18647,N_18902);
nand U19153 (N_19153,N_18720,N_18738);
and U19154 (N_19154,N_18602,N_18536);
or U19155 (N_19155,N_18679,N_18833);
nand U19156 (N_19156,N_18844,N_18746);
and U19157 (N_19157,N_18548,N_18777);
nand U19158 (N_19158,N_18657,N_18654);
or U19159 (N_19159,N_18660,N_18574);
and U19160 (N_19160,N_18804,N_18614);
nor U19161 (N_19161,N_18801,N_18954);
xnor U19162 (N_19162,N_18871,N_18642);
and U19163 (N_19163,N_18965,N_18955);
nand U19164 (N_19164,N_18620,N_18805);
xor U19165 (N_19165,N_18894,N_18977);
nand U19166 (N_19166,N_18936,N_18892);
xor U19167 (N_19167,N_18594,N_18719);
or U19168 (N_19168,N_18786,N_18734);
nand U19169 (N_19169,N_18931,N_18552);
or U19170 (N_19170,N_18949,N_18972);
nand U19171 (N_19171,N_18607,N_18667);
nand U19172 (N_19172,N_18633,N_18595);
and U19173 (N_19173,N_18856,N_18645);
nor U19174 (N_19174,N_18847,N_18876);
and U19175 (N_19175,N_18917,N_18670);
xor U19176 (N_19176,N_18653,N_18699);
or U19177 (N_19177,N_18503,N_18755);
xor U19178 (N_19178,N_18632,N_18758);
and U19179 (N_19179,N_18842,N_18562);
and U19180 (N_19180,N_18851,N_18636);
nor U19181 (N_19181,N_18658,N_18767);
or U19182 (N_19182,N_18990,N_18717);
nand U19183 (N_19183,N_18625,N_18537);
xnor U19184 (N_19184,N_18580,N_18806);
and U19185 (N_19185,N_18702,N_18985);
and U19186 (N_19186,N_18935,N_18554);
and U19187 (N_19187,N_18782,N_18778);
and U19188 (N_19188,N_18596,N_18776);
or U19189 (N_19189,N_18677,N_18898);
xnor U19190 (N_19190,N_18971,N_18692);
xnor U19191 (N_19191,N_18526,N_18541);
and U19192 (N_19192,N_18611,N_18628);
nand U19193 (N_19193,N_18940,N_18808);
or U19194 (N_19194,N_18855,N_18997);
or U19195 (N_19195,N_18666,N_18881);
or U19196 (N_19196,N_18901,N_18809);
nand U19197 (N_19197,N_18694,N_18749);
or U19198 (N_19198,N_18715,N_18770);
and U19199 (N_19199,N_18895,N_18583);
or U19200 (N_19200,N_18858,N_18800);
xor U19201 (N_19201,N_18822,N_18564);
and U19202 (N_19202,N_18543,N_18597);
xor U19203 (N_19203,N_18693,N_18932);
or U19204 (N_19204,N_18592,N_18827);
and U19205 (N_19205,N_18714,N_18567);
nor U19206 (N_19206,N_18591,N_18725);
nand U19207 (N_19207,N_18839,N_18603);
or U19208 (N_19208,N_18568,N_18685);
or U19209 (N_19209,N_18678,N_18533);
and U19210 (N_19210,N_18609,N_18644);
nor U19211 (N_19211,N_18946,N_18765);
nor U19212 (N_19212,N_18672,N_18599);
xor U19213 (N_19213,N_18686,N_18735);
and U19214 (N_19214,N_18798,N_18942);
xor U19215 (N_19215,N_18728,N_18616);
and U19216 (N_19216,N_18781,N_18893);
nor U19217 (N_19217,N_18880,N_18534);
or U19218 (N_19218,N_18553,N_18930);
xor U19219 (N_19219,N_18941,N_18862);
xor U19220 (N_19220,N_18929,N_18698);
and U19221 (N_19221,N_18718,N_18700);
nor U19222 (N_19222,N_18545,N_18967);
xnor U19223 (N_19223,N_18926,N_18810);
xor U19224 (N_19224,N_18617,N_18813);
nand U19225 (N_19225,N_18760,N_18890);
nor U19226 (N_19226,N_18979,N_18921);
nor U19227 (N_19227,N_18764,N_18872);
nor U19228 (N_19228,N_18710,N_18753);
or U19229 (N_19229,N_18975,N_18566);
and U19230 (N_19230,N_18824,N_18762);
or U19231 (N_19231,N_18811,N_18748);
nor U19232 (N_19232,N_18579,N_18705);
nand U19233 (N_19233,N_18873,N_18571);
nand U19234 (N_19234,N_18944,N_18570);
nand U19235 (N_19235,N_18627,N_18691);
nor U19236 (N_19236,N_18828,N_18656);
nand U19237 (N_19237,N_18600,N_18957);
or U19238 (N_19238,N_18531,N_18769);
nand U19239 (N_19239,N_18889,N_18937);
nand U19240 (N_19240,N_18920,N_18629);
nand U19241 (N_19241,N_18682,N_18879);
nor U19242 (N_19242,N_18817,N_18966);
or U19243 (N_19243,N_18783,N_18555);
and U19244 (N_19244,N_18649,N_18927);
and U19245 (N_19245,N_18840,N_18865);
nand U19246 (N_19246,N_18514,N_18521);
nand U19247 (N_19247,N_18716,N_18507);
nand U19248 (N_19248,N_18888,N_18668);
or U19249 (N_19249,N_18866,N_18619);
xor U19250 (N_19250,N_18836,N_18982);
or U19251 (N_19251,N_18652,N_18878);
or U19252 (N_19252,N_18569,N_18696);
nand U19253 (N_19253,N_18879,N_18992);
nor U19254 (N_19254,N_18923,N_18549);
nand U19255 (N_19255,N_18667,N_18986);
or U19256 (N_19256,N_18679,N_18607);
and U19257 (N_19257,N_18719,N_18880);
nand U19258 (N_19258,N_18978,N_18992);
and U19259 (N_19259,N_18954,N_18629);
or U19260 (N_19260,N_18682,N_18552);
nor U19261 (N_19261,N_18712,N_18827);
nor U19262 (N_19262,N_18605,N_18857);
xnor U19263 (N_19263,N_18543,N_18933);
nor U19264 (N_19264,N_18573,N_18764);
or U19265 (N_19265,N_18512,N_18885);
and U19266 (N_19266,N_18885,N_18960);
nor U19267 (N_19267,N_18515,N_18922);
nor U19268 (N_19268,N_18614,N_18918);
and U19269 (N_19269,N_18919,N_18891);
and U19270 (N_19270,N_18937,N_18607);
and U19271 (N_19271,N_18651,N_18884);
nor U19272 (N_19272,N_18742,N_18576);
nand U19273 (N_19273,N_18509,N_18851);
nor U19274 (N_19274,N_18672,N_18968);
or U19275 (N_19275,N_18553,N_18917);
xnor U19276 (N_19276,N_18808,N_18771);
or U19277 (N_19277,N_18898,N_18895);
xnor U19278 (N_19278,N_18991,N_18562);
and U19279 (N_19279,N_18850,N_18590);
nor U19280 (N_19280,N_18874,N_18798);
xnor U19281 (N_19281,N_18651,N_18534);
nor U19282 (N_19282,N_18503,N_18962);
nor U19283 (N_19283,N_18522,N_18686);
xnor U19284 (N_19284,N_18866,N_18593);
xor U19285 (N_19285,N_18521,N_18663);
nor U19286 (N_19286,N_18813,N_18992);
and U19287 (N_19287,N_18541,N_18860);
nand U19288 (N_19288,N_18878,N_18539);
and U19289 (N_19289,N_18756,N_18538);
and U19290 (N_19290,N_18823,N_18577);
xnor U19291 (N_19291,N_18533,N_18597);
xor U19292 (N_19292,N_18505,N_18807);
or U19293 (N_19293,N_18692,N_18848);
or U19294 (N_19294,N_18992,N_18751);
and U19295 (N_19295,N_18959,N_18519);
nand U19296 (N_19296,N_18897,N_18943);
nor U19297 (N_19297,N_18739,N_18959);
nand U19298 (N_19298,N_18603,N_18523);
nand U19299 (N_19299,N_18818,N_18888);
nor U19300 (N_19300,N_18721,N_18797);
and U19301 (N_19301,N_18531,N_18883);
and U19302 (N_19302,N_18763,N_18881);
nor U19303 (N_19303,N_18793,N_18837);
xnor U19304 (N_19304,N_18760,N_18804);
xor U19305 (N_19305,N_18930,N_18501);
nand U19306 (N_19306,N_18750,N_18518);
xnor U19307 (N_19307,N_18802,N_18696);
nor U19308 (N_19308,N_18943,N_18639);
or U19309 (N_19309,N_18951,N_18523);
xnor U19310 (N_19310,N_18803,N_18507);
xnor U19311 (N_19311,N_18550,N_18635);
or U19312 (N_19312,N_18654,N_18895);
and U19313 (N_19313,N_18530,N_18574);
and U19314 (N_19314,N_18600,N_18564);
nand U19315 (N_19315,N_18928,N_18579);
nand U19316 (N_19316,N_18992,N_18537);
or U19317 (N_19317,N_18969,N_18599);
nand U19318 (N_19318,N_18785,N_18639);
xnor U19319 (N_19319,N_18792,N_18559);
nor U19320 (N_19320,N_18959,N_18681);
nor U19321 (N_19321,N_18582,N_18958);
xor U19322 (N_19322,N_18798,N_18969);
and U19323 (N_19323,N_18864,N_18674);
and U19324 (N_19324,N_18551,N_18927);
nand U19325 (N_19325,N_18658,N_18679);
xnor U19326 (N_19326,N_18722,N_18742);
or U19327 (N_19327,N_18879,N_18607);
xnor U19328 (N_19328,N_18936,N_18761);
and U19329 (N_19329,N_18555,N_18861);
xor U19330 (N_19330,N_18791,N_18576);
and U19331 (N_19331,N_18677,N_18964);
xnor U19332 (N_19332,N_18670,N_18955);
and U19333 (N_19333,N_18686,N_18752);
nand U19334 (N_19334,N_18591,N_18553);
nor U19335 (N_19335,N_18770,N_18505);
nor U19336 (N_19336,N_18783,N_18672);
and U19337 (N_19337,N_18705,N_18810);
xor U19338 (N_19338,N_18867,N_18537);
nand U19339 (N_19339,N_18834,N_18723);
and U19340 (N_19340,N_18702,N_18773);
xor U19341 (N_19341,N_18778,N_18620);
nor U19342 (N_19342,N_18510,N_18526);
nor U19343 (N_19343,N_18720,N_18620);
xnor U19344 (N_19344,N_18689,N_18565);
and U19345 (N_19345,N_18625,N_18670);
xor U19346 (N_19346,N_18865,N_18584);
xnor U19347 (N_19347,N_18757,N_18835);
nor U19348 (N_19348,N_18823,N_18878);
nor U19349 (N_19349,N_18988,N_18501);
nor U19350 (N_19350,N_18650,N_18648);
or U19351 (N_19351,N_18722,N_18867);
nor U19352 (N_19352,N_18751,N_18692);
xnor U19353 (N_19353,N_18993,N_18995);
nor U19354 (N_19354,N_18599,N_18829);
or U19355 (N_19355,N_18657,N_18889);
nand U19356 (N_19356,N_18726,N_18796);
nor U19357 (N_19357,N_18597,N_18798);
and U19358 (N_19358,N_18767,N_18651);
xnor U19359 (N_19359,N_18980,N_18508);
nand U19360 (N_19360,N_18662,N_18874);
and U19361 (N_19361,N_18776,N_18507);
and U19362 (N_19362,N_18879,N_18762);
nor U19363 (N_19363,N_18683,N_18990);
nor U19364 (N_19364,N_18600,N_18916);
or U19365 (N_19365,N_18972,N_18965);
or U19366 (N_19366,N_18929,N_18605);
xnor U19367 (N_19367,N_18770,N_18951);
or U19368 (N_19368,N_18787,N_18855);
nand U19369 (N_19369,N_18800,N_18500);
nand U19370 (N_19370,N_18565,N_18954);
and U19371 (N_19371,N_18986,N_18649);
or U19372 (N_19372,N_18525,N_18655);
or U19373 (N_19373,N_18990,N_18975);
nor U19374 (N_19374,N_18524,N_18860);
xor U19375 (N_19375,N_18777,N_18676);
or U19376 (N_19376,N_18937,N_18536);
xnor U19377 (N_19377,N_18561,N_18858);
nor U19378 (N_19378,N_18734,N_18917);
and U19379 (N_19379,N_18800,N_18509);
xnor U19380 (N_19380,N_18978,N_18701);
nor U19381 (N_19381,N_18606,N_18746);
xnor U19382 (N_19382,N_18701,N_18712);
and U19383 (N_19383,N_18961,N_18651);
nor U19384 (N_19384,N_18536,N_18995);
xnor U19385 (N_19385,N_18530,N_18864);
and U19386 (N_19386,N_18624,N_18904);
nand U19387 (N_19387,N_18918,N_18568);
nand U19388 (N_19388,N_18930,N_18809);
or U19389 (N_19389,N_18705,N_18613);
nor U19390 (N_19390,N_18782,N_18949);
and U19391 (N_19391,N_18568,N_18961);
xor U19392 (N_19392,N_18928,N_18953);
or U19393 (N_19393,N_18993,N_18590);
and U19394 (N_19394,N_18874,N_18762);
xor U19395 (N_19395,N_18732,N_18941);
or U19396 (N_19396,N_18715,N_18616);
or U19397 (N_19397,N_18573,N_18639);
xor U19398 (N_19398,N_18875,N_18846);
nand U19399 (N_19399,N_18963,N_18506);
xnor U19400 (N_19400,N_18646,N_18948);
nor U19401 (N_19401,N_18605,N_18763);
or U19402 (N_19402,N_18802,N_18635);
and U19403 (N_19403,N_18959,N_18571);
nor U19404 (N_19404,N_18968,N_18980);
nand U19405 (N_19405,N_18555,N_18845);
or U19406 (N_19406,N_18903,N_18799);
and U19407 (N_19407,N_18617,N_18948);
and U19408 (N_19408,N_18963,N_18792);
xor U19409 (N_19409,N_18628,N_18772);
or U19410 (N_19410,N_18677,N_18652);
or U19411 (N_19411,N_18933,N_18584);
xnor U19412 (N_19412,N_18717,N_18817);
or U19413 (N_19413,N_18640,N_18902);
and U19414 (N_19414,N_18835,N_18969);
xnor U19415 (N_19415,N_18532,N_18734);
nor U19416 (N_19416,N_18758,N_18918);
or U19417 (N_19417,N_18834,N_18579);
nor U19418 (N_19418,N_18574,N_18992);
and U19419 (N_19419,N_18889,N_18778);
and U19420 (N_19420,N_18933,N_18511);
xor U19421 (N_19421,N_18532,N_18835);
or U19422 (N_19422,N_18875,N_18681);
and U19423 (N_19423,N_18791,N_18861);
and U19424 (N_19424,N_18739,N_18837);
nor U19425 (N_19425,N_18635,N_18798);
and U19426 (N_19426,N_18788,N_18597);
or U19427 (N_19427,N_18515,N_18575);
nor U19428 (N_19428,N_18560,N_18665);
and U19429 (N_19429,N_18937,N_18515);
or U19430 (N_19430,N_18895,N_18908);
and U19431 (N_19431,N_18729,N_18902);
or U19432 (N_19432,N_18840,N_18789);
xor U19433 (N_19433,N_18933,N_18643);
xnor U19434 (N_19434,N_18540,N_18930);
nand U19435 (N_19435,N_18569,N_18887);
nor U19436 (N_19436,N_18685,N_18693);
nand U19437 (N_19437,N_18964,N_18914);
or U19438 (N_19438,N_18811,N_18558);
nor U19439 (N_19439,N_18886,N_18710);
xnor U19440 (N_19440,N_18538,N_18962);
nand U19441 (N_19441,N_18562,N_18723);
nor U19442 (N_19442,N_18632,N_18815);
nand U19443 (N_19443,N_18919,N_18690);
nor U19444 (N_19444,N_18748,N_18592);
nand U19445 (N_19445,N_18591,N_18703);
nand U19446 (N_19446,N_18665,N_18641);
or U19447 (N_19447,N_18903,N_18721);
and U19448 (N_19448,N_18832,N_18589);
or U19449 (N_19449,N_18999,N_18985);
and U19450 (N_19450,N_18942,N_18542);
and U19451 (N_19451,N_18541,N_18777);
or U19452 (N_19452,N_18893,N_18896);
and U19453 (N_19453,N_18520,N_18761);
nand U19454 (N_19454,N_18818,N_18645);
nor U19455 (N_19455,N_18924,N_18994);
and U19456 (N_19456,N_18924,N_18546);
nor U19457 (N_19457,N_18873,N_18921);
nor U19458 (N_19458,N_18760,N_18839);
nor U19459 (N_19459,N_18549,N_18890);
nand U19460 (N_19460,N_18773,N_18518);
xnor U19461 (N_19461,N_18781,N_18715);
nor U19462 (N_19462,N_18922,N_18751);
and U19463 (N_19463,N_18579,N_18541);
xor U19464 (N_19464,N_18610,N_18902);
xnor U19465 (N_19465,N_18968,N_18909);
and U19466 (N_19466,N_18903,N_18818);
xor U19467 (N_19467,N_18562,N_18831);
or U19468 (N_19468,N_18740,N_18930);
xor U19469 (N_19469,N_18659,N_18944);
nor U19470 (N_19470,N_18964,N_18588);
xnor U19471 (N_19471,N_18978,N_18781);
xnor U19472 (N_19472,N_18755,N_18812);
or U19473 (N_19473,N_18782,N_18860);
nand U19474 (N_19474,N_18720,N_18868);
nand U19475 (N_19475,N_18866,N_18814);
xor U19476 (N_19476,N_18668,N_18827);
and U19477 (N_19477,N_18644,N_18662);
xor U19478 (N_19478,N_18844,N_18517);
or U19479 (N_19479,N_18706,N_18535);
and U19480 (N_19480,N_18640,N_18782);
xnor U19481 (N_19481,N_18802,N_18516);
xnor U19482 (N_19482,N_18823,N_18969);
and U19483 (N_19483,N_18938,N_18523);
and U19484 (N_19484,N_18848,N_18702);
nand U19485 (N_19485,N_18756,N_18876);
nor U19486 (N_19486,N_18739,N_18720);
nor U19487 (N_19487,N_18758,N_18915);
nand U19488 (N_19488,N_18902,N_18608);
xor U19489 (N_19489,N_18560,N_18503);
xor U19490 (N_19490,N_18854,N_18751);
nor U19491 (N_19491,N_18594,N_18932);
nor U19492 (N_19492,N_18817,N_18844);
nor U19493 (N_19493,N_18934,N_18606);
nand U19494 (N_19494,N_18843,N_18834);
nor U19495 (N_19495,N_18639,N_18817);
xor U19496 (N_19496,N_18850,N_18804);
xnor U19497 (N_19497,N_18667,N_18533);
nor U19498 (N_19498,N_18756,N_18858);
nand U19499 (N_19499,N_18906,N_18897);
or U19500 (N_19500,N_19141,N_19170);
nand U19501 (N_19501,N_19273,N_19244);
nand U19502 (N_19502,N_19453,N_19472);
nor U19503 (N_19503,N_19282,N_19417);
nor U19504 (N_19504,N_19295,N_19080);
nand U19505 (N_19505,N_19002,N_19399);
nand U19506 (N_19506,N_19293,N_19334);
nand U19507 (N_19507,N_19316,N_19427);
nor U19508 (N_19508,N_19154,N_19359);
and U19509 (N_19509,N_19195,N_19264);
nor U19510 (N_19510,N_19183,N_19039);
and U19511 (N_19511,N_19144,N_19078);
xnor U19512 (N_19512,N_19073,N_19258);
xnor U19513 (N_19513,N_19412,N_19118);
nand U19514 (N_19514,N_19132,N_19299);
or U19515 (N_19515,N_19370,N_19307);
and U19516 (N_19516,N_19232,N_19061);
nor U19517 (N_19517,N_19314,N_19011);
nor U19518 (N_19518,N_19190,N_19013);
xor U19519 (N_19519,N_19283,N_19263);
and U19520 (N_19520,N_19348,N_19159);
nor U19521 (N_19521,N_19395,N_19331);
nand U19522 (N_19522,N_19017,N_19292);
nor U19523 (N_19523,N_19217,N_19241);
nor U19524 (N_19524,N_19239,N_19368);
nand U19525 (N_19525,N_19211,N_19092);
xor U19526 (N_19526,N_19425,N_19112);
nand U19527 (N_19527,N_19450,N_19434);
nand U19528 (N_19528,N_19222,N_19477);
nand U19529 (N_19529,N_19345,N_19396);
and U19530 (N_19530,N_19035,N_19349);
and U19531 (N_19531,N_19094,N_19180);
nand U19532 (N_19532,N_19444,N_19267);
and U19533 (N_19533,N_19469,N_19365);
nor U19534 (N_19534,N_19451,N_19247);
nor U19535 (N_19535,N_19488,N_19318);
xor U19536 (N_19536,N_19219,N_19210);
and U19537 (N_19537,N_19145,N_19034);
nand U19538 (N_19538,N_19231,N_19021);
and U19539 (N_19539,N_19315,N_19446);
and U19540 (N_19540,N_19265,N_19485);
or U19541 (N_19541,N_19326,N_19286);
and U19542 (N_19542,N_19029,N_19487);
xnor U19543 (N_19543,N_19464,N_19194);
or U19544 (N_19544,N_19108,N_19025);
or U19545 (N_19545,N_19323,N_19129);
or U19546 (N_19546,N_19379,N_19317);
nor U19547 (N_19547,N_19491,N_19156);
xnor U19548 (N_19548,N_19285,N_19189);
and U19549 (N_19549,N_19483,N_19304);
nand U19550 (N_19550,N_19256,N_19432);
and U19551 (N_19551,N_19216,N_19065);
nor U19552 (N_19552,N_19044,N_19079);
and U19553 (N_19553,N_19478,N_19452);
nor U19554 (N_19554,N_19208,N_19220);
nor U19555 (N_19555,N_19172,N_19130);
xnor U19556 (N_19556,N_19416,N_19235);
or U19557 (N_19557,N_19030,N_19465);
and U19558 (N_19558,N_19049,N_19347);
or U19559 (N_19559,N_19023,N_19437);
xor U19560 (N_19560,N_19071,N_19184);
nand U19561 (N_19561,N_19266,N_19467);
nor U19562 (N_19562,N_19164,N_19271);
nand U19563 (N_19563,N_19423,N_19440);
nand U19564 (N_19564,N_19188,N_19291);
nor U19565 (N_19565,N_19070,N_19093);
nand U19566 (N_19566,N_19087,N_19436);
nand U19567 (N_19567,N_19223,N_19249);
nand U19568 (N_19568,N_19384,N_19245);
nor U19569 (N_19569,N_19207,N_19042);
xor U19570 (N_19570,N_19001,N_19091);
or U19571 (N_19571,N_19109,N_19288);
nor U19572 (N_19572,N_19294,N_19163);
xor U19573 (N_19573,N_19106,N_19123);
nor U19574 (N_19574,N_19102,N_19233);
or U19575 (N_19575,N_19390,N_19343);
and U19576 (N_19576,N_19240,N_19246);
and U19577 (N_19577,N_19429,N_19424);
and U19578 (N_19578,N_19215,N_19124);
xor U19579 (N_19579,N_19400,N_19369);
nand U19580 (N_19580,N_19252,N_19269);
nor U19581 (N_19581,N_19242,N_19146);
and U19582 (N_19582,N_19155,N_19171);
and U19583 (N_19583,N_19075,N_19138);
nand U19584 (N_19584,N_19279,N_19441);
xnor U19585 (N_19585,N_19344,N_19101);
or U19586 (N_19586,N_19378,N_19320);
xnor U19587 (N_19587,N_19019,N_19476);
nor U19588 (N_19588,N_19214,N_19275);
nand U19589 (N_19589,N_19205,N_19063);
or U19590 (N_19590,N_19122,N_19058);
or U19591 (N_19591,N_19460,N_19408);
and U19592 (N_19592,N_19442,N_19193);
or U19593 (N_19593,N_19260,N_19325);
nand U19594 (N_19594,N_19116,N_19237);
xnor U19595 (N_19595,N_19099,N_19227);
and U19596 (N_19596,N_19421,N_19268);
nand U19597 (N_19597,N_19107,N_19168);
or U19598 (N_19598,N_19470,N_19356);
xnor U19599 (N_19599,N_19324,N_19008);
or U19600 (N_19600,N_19248,N_19339);
or U19601 (N_19601,N_19127,N_19391);
or U19602 (N_19602,N_19026,N_19351);
xnor U19603 (N_19603,N_19322,N_19104);
or U19604 (N_19604,N_19173,N_19401);
nand U19605 (N_19605,N_19040,N_19336);
nand U19606 (N_19606,N_19077,N_19158);
or U19607 (N_19607,N_19474,N_19438);
xnor U19608 (N_19608,N_19016,N_19371);
xor U19609 (N_19609,N_19303,N_19358);
nand U19610 (N_19610,N_19489,N_19298);
nand U19611 (N_19611,N_19302,N_19081);
or U19612 (N_19612,N_19153,N_19114);
or U19613 (N_19613,N_19327,N_19095);
nor U19614 (N_19614,N_19036,N_19103);
and U19615 (N_19615,N_19050,N_19262);
and U19616 (N_19616,N_19306,N_19456);
or U19617 (N_19617,N_19468,N_19150);
nand U19618 (N_19618,N_19407,N_19105);
nand U19619 (N_19619,N_19393,N_19046);
nand U19620 (N_19620,N_19006,N_19354);
xor U19621 (N_19621,N_19226,N_19409);
and U19622 (N_19622,N_19096,N_19454);
nand U19623 (N_19623,N_19128,N_19381);
or U19624 (N_19624,N_19387,N_19475);
and U19625 (N_19625,N_19043,N_19490);
nand U19626 (N_19626,N_19461,N_19360);
nor U19627 (N_19627,N_19082,N_19353);
nand U19628 (N_19628,N_19253,N_19236);
nor U19629 (N_19629,N_19086,N_19342);
nand U19630 (N_19630,N_19352,N_19161);
or U19631 (N_19631,N_19495,N_19031);
xnor U19632 (N_19632,N_19426,N_19167);
and U19633 (N_19633,N_19062,N_19069);
or U19634 (N_19634,N_19402,N_19386);
and U19635 (N_19635,N_19165,N_19330);
and U19636 (N_19636,N_19482,N_19018);
xor U19637 (N_19637,N_19312,N_19251);
and U19638 (N_19638,N_19418,N_19435);
nor U19639 (N_19639,N_19033,N_19152);
xnor U19640 (N_19640,N_19433,N_19428);
nand U19641 (N_19641,N_19300,N_19014);
xor U19642 (N_19642,N_19466,N_19383);
or U19643 (N_19643,N_19126,N_19254);
nor U19644 (N_19644,N_19284,N_19085);
or U19645 (N_19645,N_19406,N_19224);
xnor U19646 (N_19646,N_19178,N_19448);
xor U19647 (N_19647,N_19350,N_19097);
xor U19648 (N_19648,N_19024,N_19281);
or U19649 (N_19649,N_19420,N_19136);
nor U19650 (N_19650,N_19278,N_19289);
xnor U19651 (N_19651,N_19403,N_19319);
nor U19652 (N_19652,N_19486,N_19185);
nor U19653 (N_19653,N_19162,N_19120);
nand U19654 (N_19654,N_19414,N_19052);
xnor U19655 (N_19655,N_19497,N_19179);
nand U19656 (N_19656,N_19047,N_19151);
nand U19657 (N_19657,N_19449,N_19119);
nand U19658 (N_19658,N_19012,N_19243);
xnor U19659 (N_19659,N_19133,N_19204);
xnor U19660 (N_19660,N_19362,N_19377);
nand U19661 (N_19661,N_19169,N_19257);
and U19662 (N_19662,N_19005,N_19056);
or U19663 (N_19663,N_19113,N_19038);
nor U19664 (N_19664,N_19480,N_19007);
nand U19665 (N_19665,N_19481,N_19228);
or U19666 (N_19666,N_19255,N_19121);
nor U19667 (N_19667,N_19479,N_19187);
xnor U19668 (N_19668,N_19147,N_19355);
nor U19669 (N_19669,N_19230,N_19067);
nand U19670 (N_19670,N_19422,N_19198);
nor U19671 (N_19671,N_19332,N_19462);
or U19672 (N_19672,N_19221,N_19000);
or U19673 (N_19673,N_19413,N_19276);
or U19674 (N_19674,N_19131,N_19028);
nand U19675 (N_19675,N_19115,N_19089);
and U19676 (N_19676,N_19280,N_19484);
nand U19677 (N_19677,N_19098,N_19084);
and U19678 (N_19678,N_19447,N_19125);
xor U19679 (N_19679,N_19398,N_19009);
xnor U19680 (N_19680,N_19088,N_19439);
nand U19681 (N_19681,N_19498,N_19225);
nor U19682 (N_19682,N_19492,N_19213);
or U19683 (N_19683,N_19149,N_19032);
nor U19684 (N_19684,N_19430,N_19100);
xnor U19685 (N_19685,N_19297,N_19200);
nand U19686 (N_19686,N_19197,N_19054);
nand U19687 (N_19687,N_19083,N_19037);
and U19688 (N_19688,N_19196,N_19191);
nor U19689 (N_19689,N_19212,N_19367);
nor U19690 (N_19690,N_19134,N_19309);
xnor U19691 (N_19691,N_19457,N_19015);
and U19692 (N_19692,N_19229,N_19305);
or U19693 (N_19693,N_19076,N_19139);
and U19694 (N_19694,N_19186,N_19372);
xor U19695 (N_19695,N_19310,N_19174);
xor U19696 (N_19696,N_19287,N_19311);
and U19697 (N_19697,N_19301,N_19335);
or U19698 (N_19698,N_19329,N_19471);
or U19699 (N_19699,N_19202,N_19074);
or U19700 (N_19700,N_19374,N_19055);
xor U19701 (N_19701,N_19431,N_19182);
nor U19702 (N_19702,N_19376,N_19160);
or U19703 (N_19703,N_19027,N_19411);
and U19704 (N_19704,N_19463,N_19166);
or U19705 (N_19705,N_19117,N_19313);
nor U19706 (N_19706,N_19175,N_19111);
nand U19707 (N_19707,N_19135,N_19259);
or U19708 (N_19708,N_19385,N_19203);
nor U19709 (N_19709,N_19051,N_19364);
and U19710 (N_19710,N_19003,N_19066);
xor U19711 (N_19711,N_19022,N_19415);
or U19712 (N_19712,N_19443,N_19375);
nor U19713 (N_19713,N_19234,N_19277);
xnor U19714 (N_19714,N_19382,N_19199);
xor U19715 (N_19715,N_19380,N_19328);
and U19716 (N_19716,N_19048,N_19060);
nand U19717 (N_19717,N_19410,N_19455);
and U19718 (N_19718,N_19192,N_19361);
or U19719 (N_19719,N_19274,N_19110);
and U19720 (N_19720,N_19206,N_19068);
and U19721 (N_19721,N_19143,N_19072);
or U19722 (N_19722,N_19272,N_19201);
nor U19723 (N_19723,N_19404,N_19493);
and U19724 (N_19724,N_19394,N_19494);
xnor U19725 (N_19725,N_19270,N_19057);
nand U19726 (N_19726,N_19041,N_19366);
xor U19727 (N_19727,N_19357,N_19373);
nor U19728 (N_19728,N_19363,N_19261);
or U19729 (N_19729,N_19142,N_19290);
and U19730 (N_19730,N_19157,N_19238);
and U19731 (N_19731,N_19140,N_19346);
nand U19732 (N_19732,N_19308,N_19137);
nor U19733 (N_19733,N_19053,N_19458);
nor U19734 (N_19734,N_19389,N_19337);
xnor U19735 (N_19735,N_19392,N_19250);
nor U19736 (N_19736,N_19321,N_19090);
or U19737 (N_19737,N_19405,N_19499);
and U19738 (N_19738,N_19388,N_19045);
or U19739 (N_19739,N_19064,N_19496);
nor U19740 (N_19740,N_19473,N_19340);
nor U19741 (N_19741,N_19218,N_19020);
nor U19742 (N_19742,N_19148,N_19010);
and U19743 (N_19743,N_19419,N_19177);
or U19744 (N_19744,N_19445,N_19397);
nand U19745 (N_19745,N_19338,N_19181);
nand U19746 (N_19746,N_19176,N_19459);
xor U19747 (N_19747,N_19296,N_19341);
xnor U19748 (N_19748,N_19004,N_19059);
or U19749 (N_19749,N_19209,N_19333);
and U19750 (N_19750,N_19398,N_19334);
xnor U19751 (N_19751,N_19280,N_19147);
nor U19752 (N_19752,N_19118,N_19203);
nor U19753 (N_19753,N_19276,N_19031);
and U19754 (N_19754,N_19173,N_19033);
nand U19755 (N_19755,N_19493,N_19381);
or U19756 (N_19756,N_19054,N_19250);
or U19757 (N_19757,N_19311,N_19106);
xnor U19758 (N_19758,N_19401,N_19047);
and U19759 (N_19759,N_19268,N_19086);
or U19760 (N_19760,N_19109,N_19261);
and U19761 (N_19761,N_19043,N_19264);
nand U19762 (N_19762,N_19434,N_19241);
nand U19763 (N_19763,N_19190,N_19230);
nand U19764 (N_19764,N_19393,N_19135);
or U19765 (N_19765,N_19002,N_19298);
nor U19766 (N_19766,N_19014,N_19346);
nand U19767 (N_19767,N_19101,N_19290);
and U19768 (N_19768,N_19286,N_19195);
nand U19769 (N_19769,N_19290,N_19199);
nor U19770 (N_19770,N_19055,N_19194);
or U19771 (N_19771,N_19177,N_19198);
xnor U19772 (N_19772,N_19199,N_19295);
xor U19773 (N_19773,N_19004,N_19284);
and U19774 (N_19774,N_19280,N_19441);
nor U19775 (N_19775,N_19184,N_19253);
or U19776 (N_19776,N_19233,N_19019);
or U19777 (N_19777,N_19106,N_19287);
nor U19778 (N_19778,N_19022,N_19083);
xnor U19779 (N_19779,N_19247,N_19265);
xnor U19780 (N_19780,N_19427,N_19166);
and U19781 (N_19781,N_19026,N_19401);
or U19782 (N_19782,N_19038,N_19385);
nand U19783 (N_19783,N_19355,N_19112);
xnor U19784 (N_19784,N_19146,N_19238);
or U19785 (N_19785,N_19150,N_19485);
xnor U19786 (N_19786,N_19033,N_19021);
or U19787 (N_19787,N_19458,N_19461);
xnor U19788 (N_19788,N_19183,N_19238);
nand U19789 (N_19789,N_19084,N_19245);
or U19790 (N_19790,N_19351,N_19370);
nor U19791 (N_19791,N_19202,N_19170);
xor U19792 (N_19792,N_19142,N_19369);
and U19793 (N_19793,N_19059,N_19310);
and U19794 (N_19794,N_19413,N_19377);
and U19795 (N_19795,N_19322,N_19378);
nand U19796 (N_19796,N_19477,N_19412);
or U19797 (N_19797,N_19030,N_19475);
xor U19798 (N_19798,N_19278,N_19021);
nand U19799 (N_19799,N_19100,N_19386);
nor U19800 (N_19800,N_19036,N_19043);
nand U19801 (N_19801,N_19134,N_19347);
or U19802 (N_19802,N_19005,N_19259);
and U19803 (N_19803,N_19043,N_19293);
nand U19804 (N_19804,N_19441,N_19296);
xor U19805 (N_19805,N_19098,N_19008);
or U19806 (N_19806,N_19148,N_19480);
or U19807 (N_19807,N_19288,N_19099);
nand U19808 (N_19808,N_19274,N_19162);
or U19809 (N_19809,N_19386,N_19210);
and U19810 (N_19810,N_19462,N_19094);
or U19811 (N_19811,N_19415,N_19332);
or U19812 (N_19812,N_19012,N_19314);
or U19813 (N_19813,N_19479,N_19445);
and U19814 (N_19814,N_19282,N_19360);
or U19815 (N_19815,N_19400,N_19134);
nand U19816 (N_19816,N_19065,N_19002);
nor U19817 (N_19817,N_19099,N_19102);
nand U19818 (N_19818,N_19369,N_19072);
or U19819 (N_19819,N_19152,N_19302);
nor U19820 (N_19820,N_19297,N_19205);
or U19821 (N_19821,N_19393,N_19117);
nand U19822 (N_19822,N_19018,N_19217);
nor U19823 (N_19823,N_19454,N_19024);
nand U19824 (N_19824,N_19386,N_19371);
and U19825 (N_19825,N_19480,N_19224);
xnor U19826 (N_19826,N_19411,N_19239);
or U19827 (N_19827,N_19365,N_19399);
or U19828 (N_19828,N_19116,N_19061);
nor U19829 (N_19829,N_19221,N_19186);
xor U19830 (N_19830,N_19070,N_19266);
nand U19831 (N_19831,N_19171,N_19153);
nor U19832 (N_19832,N_19493,N_19055);
nor U19833 (N_19833,N_19363,N_19407);
and U19834 (N_19834,N_19225,N_19166);
xnor U19835 (N_19835,N_19423,N_19086);
and U19836 (N_19836,N_19025,N_19217);
or U19837 (N_19837,N_19071,N_19131);
nor U19838 (N_19838,N_19197,N_19028);
and U19839 (N_19839,N_19203,N_19389);
or U19840 (N_19840,N_19020,N_19329);
nand U19841 (N_19841,N_19290,N_19124);
nand U19842 (N_19842,N_19004,N_19243);
and U19843 (N_19843,N_19410,N_19398);
or U19844 (N_19844,N_19280,N_19185);
xnor U19845 (N_19845,N_19128,N_19007);
nor U19846 (N_19846,N_19190,N_19394);
nor U19847 (N_19847,N_19038,N_19152);
xor U19848 (N_19848,N_19059,N_19173);
nand U19849 (N_19849,N_19376,N_19013);
nand U19850 (N_19850,N_19363,N_19262);
or U19851 (N_19851,N_19130,N_19348);
and U19852 (N_19852,N_19182,N_19457);
or U19853 (N_19853,N_19298,N_19143);
and U19854 (N_19854,N_19071,N_19103);
nand U19855 (N_19855,N_19429,N_19489);
and U19856 (N_19856,N_19008,N_19288);
or U19857 (N_19857,N_19386,N_19038);
or U19858 (N_19858,N_19355,N_19148);
nand U19859 (N_19859,N_19137,N_19423);
and U19860 (N_19860,N_19370,N_19310);
or U19861 (N_19861,N_19161,N_19241);
or U19862 (N_19862,N_19070,N_19136);
and U19863 (N_19863,N_19361,N_19395);
and U19864 (N_19864,N_19154,N_19343);
or U19865 (N_19865,N_19087,N_19397);
or U19866 (N_19866,N_19153,N_19234);
nor U19867 (N_19867,N_19061,N_19204);
and U19868 (N_19868,N_19376,N_19464);
xor U19869 (N_19869,N_19350,N_19419);
nor U19870 (N_19870,N_19401,N_19109);
nor U19871 (N_19871,N_19271,N_19292);
and U19872 (N_19872,N_19299,N_19477);
or U19873 (N_19873,N_19385,N_19480);
or U19874 (N_19874,N_19238,N_19488);
xnor U19875 (N_19875,N_19382,N_19101);
and U19876 (N_19876,N_19412,N_19222);
nor U19877 (N_19877,N_19022,N_19292);
xnor U19878 (N_19878,N_19471,N_19252);
nor U19879 (N_19879,N_19029,N_19385);
nor U19880 (N_19880,N_19164,N_19042);
and U19881 (N_19881,N_19390,N_19111);
nand U19882 (N_19882,N_19257,N_19346);
nor U19883 (N_19883,N_19340,N_19026);
xnor U19884 (N_19884,N_19010,N_19488);
nand U19885 (N_19885,N_19318,N_19147);
xnor U19886 (N_19886,N_19419,N_19188);
nor U19887 (N_19887,N_19432,N_19030);
nand U19888 (N_19888,N_19195,N_19301);
nand U19889 (N_19889,N_19414,N_19216);
nor U19890 (N_19890,N_19283,N_19204);
and U19891 (N_19891,N_19314,N_19404);
nand U19892 (N_19892,N_19251,N_19040);
and U19893 (N_19893,N_19003,N_19374);
nand U19894 (N_19894,N_19023,N_19249);
xor U19895 (N_19895,N_19192,N_19171);
nor U19896 (N_19896,N_19273,N_19299);
and U19897 (N_19897,N_19214,N_19426);
nand U19898 (N_19898,N_19496,N_19044);
and U19899 (N_19899,N_19083,N_19335);
or U19900 (N_19900,N_19326,N_19275);
xnor U19901 (N_19901,N_19279,N_19169);
nor U19902 (N_19902,N_19190,N_19095);
and U19903 (N_19903,N_19487,N_19390);
nor U19904 (N_19904,N_19398,N_19229);
or U19905 (N_19905,N_19472,N_19031);
or U19906 (N_19906,N_19296,N_19217);
nand U19907 (N_19907,N_19282,N_19188);
xor U19908 (N_19908,N_19322,N_19256);
xor U19909 (N_19909,N_19127,N_19001);
nand U19910 (N_19910,N_19268,N_19214);
or U19911 (N_19911,N_19383,N_19118);
nor U19912 (N_19912,N_19207,N_19151);
nor U19913 (N_19913,N_19262,N_19241);
nor U19914 (N_19914,N_19149,N_19260);
and U19915 (N_19915,N_19497,N_19205);
nand U19916 (N_19916,N_19119,N_19467);
xnor U19917 (N_19917,N_19341,N_19395);
nor U19918 (N_19918,N_19038,N_19448);
nor U19919 (N_19919,N_19475,N_19161);
nand U19920 (N_19920,N_19097,N_19131);
or U19921 (N_19921,N_19279,N_19136);
or U19922 (N_19922,N_19065,N_19325);
xor U19923 (N_19923,N_19170,N_19435);
nand U19924 (N_19924,N_19441,N_19240);
xor U19925 (N_19925,N_19265,N_19217);
xnor U19926 (N_19926,N_19418,N_19204);
or U19927 (N_19927,N_19136,N_19225);
nand U19928 (N_19928,N_19113,N_19303);
and U19929 (N_19929,N_19117,N_19332);
or U19930 (N_19930,N_19449,N_19006);
or U19931 (N_19931,N_19368,N_19298);
and U19932 (N_19932,N_19316,N_19267);
and U19933 (N_19933,N_19194,N_19251);
xnor U19934 (N_19934,N_19233,N_19369);
nand U19935 (N_19935,N_19429,N_19289);
xnor U19936 (N_19936,N_19154,N_19459);
nor U19937 (N_19937,N_19310,N_19443);
or U19938 (N_19938,N_19406,N_19216);
nor U19939 (N_19939,N_19482,N_19227);
nor U19940 (N_19940,N_19242,N_19244);
nor U19941 (N_19941,N_19473,N_19121);
and U19942 (N_19942,N_19308,N_19256);
xnor U19943 (N_19943,N_19191,N_19198);
and U19944 (N_19944,N_19232,N_19006);
nor U19945 (N_19945,N_19271,N_19224);
or U19946 (N_19946,N_19041,N_19349);
and U19947 (N_19947,N_19375,N_19486);
nor U19948 (N_19948,N_19341,N_19466);
nor U19949 (N_19949,N_19029,N_19286);
and U19950 (N_19950,N_19093,N_19298);
and U19951 (N_19951,N_19139,N_19495);
or U19952 (N_19952,N_19295,N_19024);
nand U19953 (N_19953,N_19162,N_19007);
nor U19954 (N_19954,N_19421,N_19154);
and U19955 (N_19955,N_19027,N_19483);
or U19956 (N_19956,N_19064,N_19465);
nand U19957 (N_19957,N_19224,N_19355);
nor U19958 (N_19958,N_19293,N_19324);
or U19959 (N_19959,N_19377,N_19077);
or U19960 (N_19960,N_19279,N_19383);
xor U19961 (N_19961,N_19172,N_19368);
xnor U19962 (N_19962,N_19437,N_19218);
nor U19963 (N_19963,N_19312,N_19148);
or U19964 (N_19964,N_19107,N_19367);
nor U19965 (N_19965,N_19223,N_19484);
or U19966 (N_19966,N_19159,N_19379);
or U19967 (N_19967,N_19126,N_19332);
xor U19968 (N_19968,N_19497,N_19375);
nand U19969 (N_19969,N_19230,N_19130);
nand U19970 (N_19970,N_19447,N_19244);
and U19971 (N_19971,N_19268,N_19175);
nand U19972 (N_19972,N_19356,N_19159);
nor U19973 (N_19973,N_19132,N_19468);
nor U19974 (N_19974,N_19143,N_19437);
xnor U19975 (N_19975,N_19356,N_19352);
nand U19976 (N_19976,N_19052,N_19033);
xor U19977 (N_19977,N_19178,N_19316);
xnor U19978 (N_19978,N_19455,N_19259);
nand U19979 (N_19979,N_19364,N_19447);
and U19980 (N_19980,N_19008,N_19073);
nand U19981 (N_19981,N_19111,N_19102);
xor U19982 (N_19982,N_19310,N_19281);
or U19983 (N_19983,N_19211,N_19259);
nor U19984 (N_19984,N_19231,N_19307);
and U19985 (N_19985,N_19004,N_19356);
nor U19986 (N_19986,N_19034,N_19492);
nand U19987 (N_19987,N_19442,N_19145);
nand U19988 (N_19988,N_19302,N_19189);
xor U19989 (N_19989,N_19098,N_19320);
and U19990 (N_19990,N_19025,N_19221);
xor U19991 (N_19991,N_19074,N_19026);
nand U19992 (N_19992,N_19455,N_19059);
xnor U19993 (N_19993,N_19046,N_19334);
nand U19994 (N_19994,N_19301,N_19076);
and U19995 (N_19995,N_19101,N_19102);
nand U19996 (N_19996,N_19167,N_19392);
xnor U19997 (N_19997,N_19102,N_19455);
nor U19998 (N_19998,N_19075,N_19383);
or U19999 (N_19999,N_19120,N_19003);
nand U20000 (N_20000,N_19929,N_19822);
or U20001 (N_20001,N_19796,N_19762);
and U20002 (N_20002,N_19709,N_19521);
nand U20003 (N_20003,N_19533,N_19932);
xor U20004 (N_20004,N_19676,N_19827);
and U20005 (N_20005,N_19830,N_19814);
nand U20006 (N_20006,N_19904,N_19607);
xor U20007 (N_20007,N_19541,N_19782);
or U20008 (N_20008,N_19724,N_19760);
or U20009 (N_20009,N_19638,N_19515);
xnor U20010 (N_20010,N_19738,N_19764);
xor U20011 (N_20011,N_19522,N_19661);
nor U20012 (N_20012,N_19912,N_19588);
or U20013 (N_20013,N_19772,N_19909);
and U20014 (N_20014,N_19824,N_19718);
nand U20015 (N_20015,N_19649,N_19897);
or U20016 (N_20016,N_19555,N_19906);
xnor U20017 (N_20017,N_19854,N_19789);
nand U20018 (N_20018,N_19702,N_19846);
and U20019 (N_20019,N_19951,N_19659);
xor U20020 (N_20020,N_19965,N_19500);
or U20021 (N_20021,N_19681,N_19976);
nor U20022 (N_20022,N_19777,N_19883);
or U20023 (N_20023,N_19696,N_19921);
and U20024 (N_20024,N_19766,N_19654);
or U20025 (N_20025,N_19773,N_19606);
and U20026 (N_20026,N_19898,N_19594);
xnor U20027 (N_20027,N_19950,N_19903);
xnor U20028 (N_20028,N_19991,N_19885);
and U20029 (N_20029,N_19916,N_19658);
nor U20030 (N_20030,N_19655,N_19502);
xor U20031 (N_20031,N_19562,N_19964);
nor U20032 (N_20032,N_19569,N_19914);
nor U20033 (N_20033,N_19852,N_19534);
nand U20034 (N_20034,N_19902,N_19949);
xor U20035 (N_20035,N_19675,N_19923);
and U20036 (N_20036,N_19715,N_19806);
and U20037 (N_20037,N_19820,N_19962);
or U20038 (N_20038,N_19836,N_19881);
nand U20039 (N_20039,N_19747,N_19779);
nor U20040 (N_20040,N_19920,N_19616);
nand U20041 (N_20041,N_19683,N_19571);
xor U20042 (N_20042,N_19690,N_19670);
xor U20043 (N_20043,N_19563,N_19841);
nor U20044 (N_20044,N_19855,N_19542);
and U20045 (N_20045,N_19937,N_19989);
xnor U20046 (N_20046,N_19943,N_19660);
nor U20047 (N_20047,N_19842,N_19524);
nor U20048 (N_20048,N_19672,N_19511);
or U20049 (N_20049,N_19860,N_19939);
nor U20050 (N_20050,N_19507,N_19578);
and U20051 (N_20051,N_19759,N_19656);
or U20052 (N_20052,N_19609,N_19810);
and U20053 (N_20053,N_19706,N_19719);
or U20054 (N_20054,N_19746,N_19978);
and U20055 (N_20055,N_19960,N_19730);
xor U20056 (N_20056,N_19972,N_19844);
and U20057 (N_20057,N_19784,N_19774);
xor U20058 (N_20058,N_19858,N_19826);
or U20059 (N_20059,N_19543,N_19816);
or U20060 (N_20060,N_19882,N_19832);
and U20061 (N_20061,N_19629,N_19781);
and U20062 (N_20062,N_19665,N_19662);
and U20063 (N_20063,N_19604,N_19592);
nand U20064 (N_20064,N_19870,N_19942);
nand U20065 (N_20065,N_19861,N_19753);
nand U20066 (N_20066,N_19673,N_19838);
xnor U20067 (N_20067,N_19952,N_19769);
or U20068 (N_20068,N_19776,N_19513);
or U20069 (N_20069,N_19639,N_19856);
nand U20070 (N_20070,N_19552,N_19863);
or U20071 (N_20071,N_19565,N_19704);
nor U20072 (N_20072,N_19582,N_19598);
and U20073 (N_20073,N_19917,N_19732);
and U20074 (N_20074,N_19795,N_19710);
nor U20075 (N_20075,N_19620,N_19530);
xor U20076 (N_20076,N_19630,N_19848);
or U20077 (N_20077,N_19787,N_19599);
or U20078 (N_20078,N_19815,N_19786);
or U20079 (N_20079,N_19845,N_19809);
nor U20080 (N_20080,N_19993,N_19913);
xor U20081 (N_20081,N_19901,N_19969);
xnor U20082 (N_20082,N_19899,N_19603);
or U20083 (N_20083,N_19560,N_19705);
nand U20084 (N_20084,N_19612,N_19590);
xor U20085 (N_20085,N_19928,N_19701);
or U20086 (N_20086,N_19802,N_19636);
xor U20087 (N_20087,N_19539,N_19510);
xor U20088 (N_20088,N_19554,N_19581);
nand U20089 (N_20089,N_19677,N_19589);
nand U20090 (N_20090,N_19884,N_19726);
and U20091 (N_20091,N_19973,N_19935);
nor U20092 (N_20092,N_19548,N_19911);
nand U20093 (N_20093,N_19627,N_19867);
and U20094 (N_20094,N_19817,N_19643);
xor U20095 (N_20095,N_19877,N_19872);
nor U20096 (N_20096,N_19859,N_19591);
nor U20097 (N_20097,N_19615,N_19725);
nor U20098 (N_20098,N_19979,N_19741);
or U20099 (N_20099,N_19794,N_19843);
or U20100 (N_20100,N_19775,N_19503);
nor U20101 (N_20101,N_19595,N_19549);
or U20102 (N_20102,N_19663,N_19980);
and U20103 (N_20103,N_19610,N_19646);
nor U20104 (N_20104,N_19700,N_19653);
xnor U20105 (N_20105,N_19587,N_19669);
nand U20106 (N_20106,N_19650,N_19651);
and U20107 (N_20107,N_19823,N_19608);
and U20108 (N_20108,N_19954,N_19955);
nor U20109 (N_20109,N_19692,N_19977);
xor U20110 (N_20110,N_19757,N_19790);
nor U20111 (N_20111,N_19602,N_19517);
nor U20112 (N_20112,N_19873,N_19573);
nand U20113 (N_20113,N_19601,N_19900);
nand U20114 (N_20114,N_19763,N_19934);
xnor U20115 (N_20115,N_19811,N_19750);
xnor U20116 (N_20116,N_19641,N_19698);
nand U20117 (N_20117,N_19839,N_19857);
nand U20118 (N_20118,N_19987,N_19871);
or U20119 (N_20119,N_19736,N_19925);
and U20120 (N_20120,N_19509,N_19633);
xnor U20121 (N_20121,N_19888,N_19990);
or U20122 (N_20122,N_19564,N_19579);
or U20123 (N_20123,N_19765,N_19880);
nor U20124 (N_20124,N_19679,N_19624);
or U20125 (N_20125,N_19528,N_19828);
or U20126 (N_20126,N_19689,N_19508);
or U20127 (N_20127,N_19975,N_19891);
nand U20128 (N_20128,N_19751,N_19514);
and U20129 (N_20129,N_19527,N_19755);
or U20130 (N_20130,N_19878,N_19926);
and U20131 (N_20131,N_19572,N_19547);
nand U20132 (N_20132,N_19632,N_19731);
xnor U20133 (N_20133,N_19771,N_19748);
nor U20134 (N_20134,N_19927,N_19940);
xnor U20135 (N_20135,N_19545,N_19959);
or U20136 (N_20136,N_19821,N_19797);
and U20137 (N_20137,N_19812,N_19749);
nor U20138 (N_20138,N_19529,N_19966);
and U20139 (N_20139,N_19835,N_19933);
nor U20140 (N_20140,N_19551,N_19804);
and U20141 (N_20141,N_19666,N_19894);
and U20142 (N_20142,N_19600,N_19714);
nand U20143 (N_20143,N_19536,N_19918);
or U20144 (N_20144,N_19567,N_19575);
xor U20145 (N_20145,N_19631,N_19813);
or U20146 (N_20146,N_19825,N_19613);
or U20147 (N_20147,N_19970,N_19559);
nor U20148 (N_20148,N_19668,N_19512);
nor U20149 (N_20149,N_19803,N_19621);
or U20150 (N_20150,N_19586,N_19758);
or U20151 (N_20151,N_19944,N_19687);
xnor U20152 (N_20152,N_19945,N_19694);
nor U20153 (N_20153,N_19874,N_19994);
and U20154 (N_20154,N_19707,N_19961);
xnor U20155 (N_20155,N_19819,N_19713);
xor U20156 (N_20156,N_19685,N_19829);
or U20157 (N_20157,N_19622,N_19519);
nor U20158 (N_20158,N_19734,N_19992);
or U20159 (N_20159,N_19840,N_19642);
or U20160 (N_20160,N_19566,N_19862);
nand U20161 (N_20161,N_19788,N_19958);
and U20162 (N_20162,N_19834,N_19890);
nand U20163 (N_20163,N_19879,N_19780);
or U20164 (N_20164,N_19735,N_19570);
nor U20165 (N_20165,N_19866,N_19761);
nand U20166 (N_20166,N_19652,N_19727);
xnor U20167 (N_20167,N_19876,N_19799);
xor U20168 (N_20168,N_19981,N_19506);
or U20169 (N_20169,N_19645,N_19648);
and U20170 (N_20170,N_19986,N_19583);
nor U20171 (N_20171,N_19896,N_19557);
and U20172 (N_20172,N_19580,N_19739);
nor U20173 (N_20173,N_19938,N_19505);
and U20174 (N_20174,N_19712,N_19693);
nand U20175 (N_20175,N_19635,N_19999);
and U20176 (N_20176,N_19785,N_19550);
xnor U20177 (N_20177,N_19628,N_19611);
or U20178 (N_20178,N_19558,N_19720);
nor U20179 (N_20179,N_19996,N_19801);
and U20180 (N_20180,N_19504,N_19956);
nand U20181 (N_20181,N_19742,N_19864);
nor U20182 (N_20182,N_19971,N_19531);
nor U20183 (N_20183,N_19833,N_19831);
and U20184 (N_20184,N_19818,N_19967);
nor U20185 (N_20185,N_19847,N_19728);
and U20186 (N_20186,N_19593,N_19699);
nor U20187 (N_20187,N_19640,N_19745);
xnor U20188 (N_20188,N_19837,N_19664);
nand U20189 (N_20189,N_19783,N_19585);
nor U20190 (N_20190,N_19995,N_19532);
and U20191 (N_20191,N_19657,N_19983);
or U20192 (N_20192,N_19723,N_19907);
and U20193 (N_20193,N_19919,N_19678);
nand U20194 (N_20194,N_19721,N_19792);
xor U20195 (N_20195,N_19537,N_19623);
or U20196 (N_20196,N_19682,N_19540);
nor U20197 (N_20197,N_19988,N_19667);
or U20198 (N_20198,N_19982,N_19853);
or U20199 (N_20199,N_19688,N_19941);
nand U20200 (N_20200,N_19614,N_19584);
and U20201 (N_20201,N_19936,N_19895);
xnor U20202 (N_20202,N_19644,N_19576);
nand U20203 (N_20203,N_19518,N_19800);
and U20204 (N_20204,N_19671,N_19798);
xnor U20205 (N_20205,N_19791,N_19868);
or U20206 (N_20206,N_19691,N_19930);
and U20207 (N_20207,N_19851,N_19674);
nand U20208 (N_20208,N_19740,N_19910);
nand U20209 (N_20209,N_19605,N_19737);
or U20210 (N_20210,N_19717,N_19538);
and U20211 (N_20211,N_19808,N_19535);
and U20212 (N_20212,N_19849,N_19577);
nand U20213 (N_20213,N_19722,N_19793);
nand U20214 (N_20214,N_19596,N_19695);
nand U20215 (N_20215,N_19703,N_19767);
nor U20216 (N_20216,N_19637,N_19647);
and U20217 (N_20217,N_19963,N_19597);
and U20218 (N_20218,N_19574,N_19546);
nor U20219 (N_20219,N_19915,N_19686);
xnor U20220 (N_20220,N_19985,N_19553);
and U20221 (N_20221,N_19875,N_19619);
xnor U20222 (N_20222,N_19708,N_19520);
or U20223 (N_20223,N_19953,N_19711);
xnor U20224 (N_20224,N_19756,N_19525);
and U20225 (N_20225,N_19947,N_19501);
xor U20226 (N_20226,N_19526,N_19625);
or U20227 (N_20227,N_19908,N_19733);
and U20228 (N_20228,N_19754,N_19889);
nor U20229 (N_20229,N_19850,N_19618);
nand U20230 (N_20230,N_19957,N_19805);
xnor U20231 (N_20231,N_19865,N_19768);
xnor U20232 (N_20232,N_19931,N_19544);
xnor U20233 (N_20233,N_19626,N_19680);
nand U20234 (N_20234,N_19516,N_19770);
or U20235 (N_20235,N_19892,N_19744);
xnor U20236 (N_20236,N_19948,N_19697);
and U20237 (N_20237,N_19946,N_19807);
xnor U20238 (N_20238,N_19924,N_19869);
or U20239 (N_20239,N_19716,N_19523);
and U20240 (N_20240,N_19634,N_19997);
and U20241 (N_20241,N_19893,N_19974);
and U20242 (N_20242,N_19561,N_19568);
or U20243 (N_20243,N_19886,N_19752);
nor U20244 (N_20244,N_19984,N_19556);
or U20245 (N_20245,N_19617,N_19729);
and U20246 (N_20246,N_19905,N_19887);
nand U20247 (N_20247,N_19968,N_19684);
or U20248 (N_20248,N_19778,N_19998);
or U20249 (N_20249,N_19922,N_19743);
nand U20250 (N_20250,N_19615,N_19925);
xor U20251 (N_20251,N_19849,N_19748);
nand U20252 (N_20252,N_19817,N_19995);
xnor U20253 (N_20253,N_19616,N_19930);
and U20254 (N_20254,N_19844,N_19634);
nand U20255 (N_20255,N_19685,N_19511);
or U20256 (N_20256,N_19852,N_19541);
and U20257 (N_20257,N_19694,N_19668);
xnor U20258 (N_20258,N_19518,N_19560);
or U20259 (N_20259,N_19965,N_19679);
and U20260 (N_20260,N_19882,N_19509);
nand U20261 (N_20261,N_19661,N_19923);
nand U20262 (N_20262,N_19741,N_19506);
xor U20263 (N_20263,N_19542,N_19702);
or U20264 (N_20264,N_19891,N_19910);
nand U20265 (N_20265,N_19914,N_19660);
and U20266 (N_20266,N_19618,N_19936);
nand U20267 (N_20267,N_19506,N_19983);
nand U20268 (N_20268,N_19761,N_19972);
or U20269 (N_20269,N_19842,N_19939);
or U20270 (N_20270,N_19789,N_19828);
xnor U20271 (N_20271,N_19715,N_19823);
xnor U20272 (N_20272,N_19836,N_19902);
xnor U20273 (N_20273,N_19843,N_19934);
and U20274 (N_20274,N_19537,N_19596);
or U20275 (N_20275,N_19715,N_19718);
or U20276 (N_20276,N_19951,N_19752);
xor U20277 (N_20277,N_19910,N_19895);
xnor U20278 (N_20278,N_19644,N_19580);
nor U20279 (N_20279,N_19907,N_19910);
xnor U20280 (N_20280,N_19569,N_19648);
nor U20281 (N_20281,N_19838,N_19796);
nand U20282 (N_20282,N_19932,N_19696);
xor U20283 (N_20283,N_19820,N_19808);
nor U20284 (N_20284,N_19614,N_19543);
xor U20285 (N_20285,N_19915,N_19790);
nor U20286 (N_20286,N_19570,N_19655);
nor U20287 (N_20287,N_19839,N_19864);
or U20288 (N_20288,N_19500,N_19589);
nor U20289 (N_20289,N_19914,N_19986);
and U20290 (N_20290,N_19951,N_19547);
nand U20291 (N_20291,N_19507,N_19718);
nand U20292 (N_20292,N_19998,N_19848);
nand U20293 (N_20293,N_19885,N_19661);
and U20294 (N_20294,N_19728,N_19558);
nor U20295 (N_20295,N_19677,N_19912);
or U20296 (N_20296,N_19910,N_19877);
nand U20297 (N_20297,N_19532,N_19783);
nor U20298 (N_20298,N_19538,N_19870);
nand U20299 (N_20299,N_19573,N_19730);
and U20300 (N_20300,N_19654,N_19600);
and U20301 (N_20301,N_19944,N_19629);
and U20302 (N_20302,N_19912,N_19972);
nand U20303 (N_20303,N_19773,N_19582);
nand U20304 (N_20304,N_19585,N_19607);
or U20305 (N_20305,N_19687,N_19964);
or U20306 (N_20306,N_19980,N_19570);
nor U20307 (N_20307,N_19504,N_19871);
xor U20308 (N_20308,N_19896,N_19910);
nand U20309 (N_20309,N_19839,N_19805);
or U20310 (N_20310,N_19617,N_19762);
and U20311 (N_20311,N_19619,N_19985);
and U20312 (N_20312,N_19831,N_19746);
nand U20313 (N_20313,N_19902,N_19713);
nand U20314 (N_20314,N_19727,N_19752);
and U20315 (N_20315,N_19634,N_19988);
xnor U20316 (N_20316,N_19931,N_19775);
or U20317 (N_20317,N_19546,N_19691);
nand U20318 (N_20318,N_19646,N_19964);
nand U20319 (N_20319,N_19757,N_19774);
nand U20320 (N_20320,N_19870,N_19674);
nor U20321 (N_20321,N_19523,N_19711);
nor U20322 (N_20322,N_19870,N_19635);
or U20323 (N_20323,N_19567,N_19907);
xor U20324 (N_20324,N_19816,N_19915);
nor U20325 (N_20325,N_19720,N_19825);
nand U20326 (N_20326,N_19624,N_19759);
xnor U20327 (N_20327,N_19737,N_19894);
or U20328 (N_20328,N_19563,N_19705);
nand U20329 (N_20329,N_19529,N_19969);
or U20330 (N_20330,N_19772,N_19815);
or U20331 (N_20331,N_19609,N_19741);
or U20332 (N_20332,N_19815,N_19734);
nor U20333 (N_20333,N_19785,N_19608);
xnor U20334 (N_20334,N_19950,N_19688);
xnor U20335 (N_20335,N_19832,N_19724);
nand U20336 (N_20336,N_19572,N_19953);
xnor U20337 (N_20337,N_19978,N_19643);
nand U20338 (N_20338,N_19973,N_19564);
nand U20339 (N_20339,N_19777,N_19566);
or U20340 (N_20340,N_19883,N_19856);
or U20341 (N_20341,N_19986,N_19951);
or U20342 (N_20342,N_19932,N_19749);
and U20343 (N_20343,N_19833,N_19686);
and U20344 (N_20344,N_19957,N_19770);
nand U20345 (N_20345,N_19875,N_19763);
xnor U20346 (N_20346,N_19554,N_19857);
or U20347 (N_20347,N_19551,N_19704);
xor U20348 (N_20348,N_19733,N_19926);
and U20349 (N_20349,N_19823,N_19541);
xnor U20350 (N_20350,N_19751,N_19920);
and U20351 (N_20351,N_19694,N_19629);
or U20352 (N_20352,N_19977,N_19723);
nand U20353 (N_20353,N_19841,N_19671);
nor U20354 (N_20354,N_19756,N_19568);
nor U20355 (N_20355,N_19655,N_19722);
xor U20356 (N_20356,N_19601,N_19937);
xor U20357 (N_20357,N_19927,N_19596);
nand U20358 (N_20358,N_19870,N_19866);
and U20359 (N_20359,N_19722,N_19955);
and U20360 (N_20360,N_19919,N_19625);
xor U20361 (N_20361,N_19737,N_19816);
xnor U20362 (N_20362,N_19627,N_19774);
nor U20363 (N_20363,N_19561,N_19786);
or U20364 (N_20364,N_19847,N_19595);
nand U20365 (N_20365,N_19542,N_19690);
nand U20366 (N_20366,N_19786,N_19976);
and U20367 (N_20367,N_19659,N_19576);
nor U20368 (N_20368,N_19538,N_19827);
and U20369 (N_20369,N_19506,N_19783);
xnor U20370 (N_20370,N_19613,N_19816);
or U20371 (N_20371,N_19670,N_19579);
xnor U20372 (N_20372,N_19918,N_19966);
or U20373 (N_20373,N_19517,N_19671);
xor U20374 (N_20374,N_19539,N_19566);
nand U20375 (N_20375,N_19927,N_19770);
nand U20376 (N_20376,N_19742,N_19772);
xor U20377 (N_20377,N_19685,N_19582);
nor U20378 (N_20378,N_19929,N_19710);
and U20379 (N_20379,N_19974,N_19543);
xnor U20380 (N_20380,N_19945,N_19675);
and U20381 (N_20381,N_19502,N_19790);
and U20382 (N_20382,N_19510,N_19717);
nor U20383 (N_20383,N_19731,N_19892);
nor U20384 (N_20384,N_19715,N_19743);
and U20385 (N_20385,N_19725,N_19680);
nor U20386 (N_20386,N_19670,N_19664);
nor U20387 (N_20387,N_19641,N_19783);
nor U20388 (N_20388,N_19942,N_19818);
xnor U20389 (N_20389,N_19698,N_19718);
or U20390 (N_20390,N_19866,N_19844);
or U20391 (N_20391,N_19957,N_19811);
xor U20392 (N_20392,N_19611,N_19955);
or U20393 (N_20393,N_19665,N_19863);
nor U20394 (N_20394,N_19594,N_19576);
nand U20395 (N_20395,N_19649,N_19576);
nor U20396 (N_20396,N_19609,N_19854);
nand U20397 (N_20397,N_19512,N_19942);
nand U20398 (N_20398,N_19569,N_19613);
and U20399 (N_20399,N_19649,N_19815);
nor U20400 (N_20400,N_19703,N_19511);
and U20401 (N_20401,N_19682,N_19769);
xnor U20402 (N_20402,N_19973,N_19605);
nand U20403 (N_20403,N_19746,N_19558);
xnor U20404 (N_20404,N_19864,N_19821);
and U20405 (N_20405,N_19936,N_19642);
and U20406 (N_20406,N_19936,N_19800);
nand U20407 (N_20407,N_19676,N_19520);
and U20408 (N_20408,N_19692,N_19952);
nand U20409 (N_20409,N_19661,N_19579);
nor U20410 (N_20410,N_19535,N_19860);
xor U20411 (N_20411,N_19989,N_19871);
nand U20412 (N_20412,N_19715,N_19526);
xor U20413 (N_20413,N_19721,N_19977);
or U20414 (N_20414,N_19745,N_19661);
and U20415 (N_20415,N_19959,N_19633);
xor U20416 (N_20416,N_19816,N_19624);
and U20417 (N_20417,N_19542,N_19597);
nand U20418 (N_20418,N_19834,N_19530);
xor U20419 (N_20419,N_19711,N_19579);
nand U20420 (N_20420,N_19977,N_19766);
or U20421 (N_20421,N_19506,N_19928);
nand U20422 (N_20422,N_19635,N_19708);
nor U20423 (N_20423,N_19791,N_19500);
nand U20424 (N_20424,N_19951,N_19677);
xnor U20425 (N_20425,N_19539,N_19852);
and U20426 (N_20426,N_19936,N_19613);
xnor U20427 (N_20427,N_19564,N_19596);
or U20428 (N_20428,N_19769,N_19515);
nor U20429 (N_20429,N_19619,N_19660);
and U20430 (N_20430,N_19941,N_19753);
nand U20431 (N_20431,N_19610,N_19924);
and U20432 (N_20432,N_19707,N_19791);
xor U20433 (N_20433,N_19723,N_19778);
or U20434 (N_20434,N_19882,N_19508);
xnor U20435 (N_20435,N_19961,N_19515);
or U20436 (N_20436,N_19780,N_19824);
nand U20437 (N_20437,N_19742,N_19964);
nor U20438 (N_20438,N_19730,N_19621);
xnor U20439 (N_20439,N_19863,N_19955);
nor U20440 (N_20440,N_19628,N_19511);
or U20441 (N_20441,N_19516,N_19706);
or U20442 (N_20442,N_19654,N_19817);
nor U20443 (N_20443,N_19732,N_19731);
nor U20444 (N_20444,N_19853,N_19549);
or U20445 (N_20445,N_19916,N_19822);
xnor U20446 (N_20446,N_19706,N_19802);
xnor U20447 (N_20447,N_19615,N_19562);
xor U20448 (N_20448,N_19629,N_19587);
or U20449 (N_20449,N_19954,N_19568);
nor U20450 (N_20450,N_19679,N_19547);
nor U20451 (N_20451,N_19979,N_19913);
nor U20452 (N_20452,N_19642,N_19914);
nand U20453 (N_20453,N_19649,N_19993);
and U20454 (N_20454,N_19987,N_19666);
or U20455 (N_20455,N_19936,N_19587);
and U20456 (N_20456,N_19906,N_19773);
nand U20457 (N_20457,N_19598,N_19940);
nand U20458 (N_20458,N_19500,N_19635);
and U20459 (N_20459,N_19579,N_19841);
and U20460 (N_20460,N_19710,N_19790);
nor U20461 (N_20461,N_19654,N_19992);
nor U20462 (N_20462,N_19746,N_19833);
and U20463 (N_20463,N_19740,N_19701);
and U20464 (N_20464,N_19718,N_19524);
nor U20465 (N_20465,N_19697,N_19660);
xor U20466 (N_20466,N_19506,N_19834);
xnor U20467 (N_20467,N_19710,N_19755);
nor U20468 (N_20468,N_19567,N_19690);
nor U20469 (N_20469,N_19761,N_19646);
and U20470 (N_20470,N_19598,N_19848);
nor U20471 (N_20471,N_19567,N_19806);
nand U20472 (N_20472,N_19503,N_19741);
nor U20473 (N_20473,N_19899,N_19593);
nand U20474 (N_20474,N_19671,N_19530);
nor U20475 (N_20475,N_19614,N_19769);
and U20476 (N_20476,N_19643,N_19608);
and U20477 (N_20477,N_19921,N_19735);
nand U20478 (N_20478,N_19758,N_19891);
nand U20479 (N_20479,N_19637,N_19863);
and U20480 (N_20480,N_19885,N_19864);
nand U20481 (N_20481,N_19959,N_19617);
or U20482 (N_20482,N_19634,N_19707);
or U20483 (N_20483,N_19827,N_19577);
or U20484 (N_20484,N_19576,N_19507);
xnor U20485 (N_20485,N_19619,N_19685);
or U20486 (N_20486,N_19595,N_19874);
nand U20487 (N_20487,N_19917,N_19890);
nor U20488 (N_20488,N_19878,N_19617);
nor U20489 (N_20489,N_19865,N_19894);
or U20490 (N_20490,N_19813,N_19613);
or U20491 (N_20491,N_19611,N_19849);
nor U20492 (N_20492,N_19758,N_19819);
nor U20493 (N_20493,N_19583,N_19984);
or U20494 (N_20494,N_19508,N_19568);
and U20495 (N_20495,N_19949,N_19574);
or U20496 (N_20496,N_19512,N_19658);
nand U20497 (N_20497,N_19677,N_19976);
xor U20498 (N_20498,N_19508,N_19624);
and U20499 (N_20499,N_19691,N_19732);
nor U20500 (N_20500,N_20166,N_20432);
or U20501 (N_20501,N_20460,N_20367);
or U20502 (N_20502,N_20001,N_20279);
nor U20503 (N_20503,N_20236,N_20039);
xor U20504 (N_20504,N_20191,N_20090);
and U20505 (N_20505,N_20246,N_20402);
and U20506 (N_20506,N_20350,N_20054);
nand U20507 (N_20507,N_20456,N_20304);
nor U20508 (N_20508,N_20475,N_20278);
nand U20509 (N_20509,N_20156,N_20442);
and U20510 (N_20510,N_20225,N_20087);
xor U20511 (N_20511,N_20211,N_20307);
xnor U20512 (N_20512,N_20447,N_20496);
or U20513 (N_20513,N_20231,N_20132);
nand U20514 (N_20514,N_20003,N_20199);
nand U20515 (N_20515,N_20014,N_20445);
xor U20516 (N_20516,N_20458,N_20198);
xor U20517 (N_20517,N_20112,N_20466);
or U20518 (N_20518,N_20433,N_20018);
and U20519 (N_20519,N_20143,N_20467);
nor U20520 (N_20520,N_20435,N_20202);
or U20521 (N_20521,N_20033,N_20016);
or U20522 (N_20522,N_20487,N_20069);
nor U20523 (N_20523,N_20275,N_20127);
xor U20524 (N_20524,N_20044,N_20228);
or U20525 (N_20525,N_20420,N_20378);
xor U20526 (N_20526,N_20427,N_20326);
xor U20527 (N_20527,N_20149,N_20124);
and U20528 (N_20528,N_20148,N_20483);
or U20529 (N_20529,N_20129,N_20260);
nand U20530 (N_20530,N_20123,N_20346);
nand U20531 (N_20531,N_20215,N_20426);
or U20532 (N_20532,N_20360,N_20471);
nand U20533 (N_20533,N_20365,N_20415);
xnor U20534 (N_20534,N_20397,N_20219);
or U20535 (N_20535,N_20007,N_20468);
or U20536 (N_20536,N_20291,N_20137);
xor U20537 (N_20537,N_20393,N_20470);
nor U20538 (N_20538,N_20185,N_20197);
or U20539 (N_20539,N_20400,N_20101);
nor U20540 (N_20540,N_20226,N_20196);
xor U20541 (N_20541,N_20205,N_20392);
xnor U20542 (N_20542,N_20072,N_20419);
nor U20543 (N_20543,N_20422,N_20040);
nor U20544 (N_20544,N_20088,N_20213);
or U20545 (N_20545,N_20201,N_20221);
nor U20546 (N_20546,N_20059,N_20151);
xnor U20547 (N_20547,N_20273,N_20128);
or U20548 (N_20548,N_20333,N_20091);
xnor U20549 (N_20549,N_20325,N_20461);
nor U20550 (N_20550,N_20318,N_20116);
xor U20551 (N_20551,N_20109,N_20009);
nand U20552 (N_20552,N_20429,N_20428);
and U20553 (N_20553,N_20280,N_20288);
xnor U20554 (N_20554,N_20080,N_20452);
nand U20555 (N_20555,N_20203,N_20049);
nand U20556 (N_20556,N_20083,N_20062);
nor U20557 (N_20557,N_20386,N_20448);
and U20558 (N_20558,N_20369,N_20262);
xor U20559 (N_20559,N_20321,N_20383);
nor U20560 (N_20560,N_20038,N_20394);
and U20561 (N_20561,N_20243,N_20484);
nand U20562 (N_20562,N_20008,N_20245);
nand U20563 (N_20563,N_20345,N_20254);
and U20564 (N_20564,N_20287,N_20227);
and U20565 (N_20565,N_20440,N_20424);
xnor U20566 (N_20566,N_20331,N_20403);
nor U20567 (N_20567,N_20404,N_20457);
xor U20568 (N_20568,N_20253,N_20028);
nor U20569 (N_20569,N_20247,N_20381);
and U20570 (N_20570,N_20459,N_20037);
xor U20571 (N_20571,N_20067,N_20261);
and U20572 (N_20572,N_20229,N_20242);
nor U20573 (N_20573,N_20004,N_20107);
or U20574 (N_20574,N_20334,N_20017);
xnor U20575 (N_20575,N_20423,N_20041);
or U20576 (N_20576,N_20061,N_20310);
nor U20577 (N_20577,N_20076,N_20138);
or U20578 (N_20578,N_20252,N_20372);
nand U20579 (N_20579,N_20477,N_20497);
and U20580 (N_20580,N_20286,N_20357);
or U20581 (N_20581,N_20042,N_20319);
and U20582 (N_20582,N_20047,N_20478);
or U20583 (N_20583,N_20111,N_20055);
or U20584 (N_20584,N_20363,N_20349);
or U20585 (N_20585,N_20183,N_20232);
xnor U20586 (N_20586,N_20210,N_20034);
xor U20587 (N_20587,N_20160,N_20388);
xnor U20588 (N_20588,N_20265,N_20015);
xor U20589 (N_20589,N_20025,N_20359);
nor U20590 (N_20590,N_20409,N_20465);
and U20591 (N_20591,N_20058,N_20118);
or U20592 (N_20592,N_20084,N_20158);
and U20593 (N_20593,N_20180,N_20011);
nor U20594 (N_20594,N_20421,N_20413);
and U20595 (N_20595,N_20315,N_20120);
nand U20596 (N_20596,N_20159,N_20224);
nand U20597 (N_20597,N_20340,N_20098);
or U20598 (N_20598,N_20027,N_20113);
or U20599 (N_20599,N_20290,N_20165);
or U20600 (N_20600,N_20283,N_20352);
or U20601 (N_20601,N_20235,N_20479);
or U20602 (N_20602,N_20268,N_20293);
and U20603 (N_20603,N_20256,N_20366);
xor U20604 (N_20604,N_20493,N_20259);
nand U20605 (N_20605,N_20115,N_20031);
nor U20606 (N_20606,N_20207,N_20299);
and U20607 (N_20607,N_20241,N_20002);
nor U20608 (N_20608,N_20481,N_20312);
nand U20609 (N_20609,N_20358,N_20106);
xnor U20610 (N_20610,N_20244,N_20269);
nor U20611 (N_20611,N_20100,N_20328);
nand U20612 (N_20612,N_20104,N_20209);
or U20613 (N_20613,N_20338,N_20292);
nor U20614 (N_20614,N_20356,N_20157);
nand U20615 (N_20615,N_20168,N_20013);
xor U20616 (N_20616,N_20302,N_20463);
and U20617 (N_20617,N_20023,N_20250);
nand U20618 (N_20618,N_20074,N_20119);
nand U20619 (N_20619,N_20045,N_20314);
nand U20620 (N_20620,N_20298,N_20294);
and U20621 (N_20621,N_20396,N_20425);
and U20622 (N_20622,N_20125,N_20026);
nor U20623 (N_20623,N_20057,N_20485);
xor U20624 (N_20624,N_20021,N_20152);
or U20625 (N_20625,N_20323,N_20081);
nor U20626 (N_20626,N_20131,N_20284);
xnor U20627 (N_20627,N_20218,N_20239);
nor U20628 (N_20628,N_20078,N_20146);
or U20629 (N_20629,N_20238,N_20171);
or U20630 (N_20630,N_20341,N_20094);
and U20631 (N_20631,N_20208,N_20093);
or U20632 (N_20632,N_20476,N_20355);
and U20633 (N_20633,N_20214,N_20066);
or U20634 (N_20634,N_20177,N_20324);
xnor U20635 (N_20635,N_20095,N_20434);
nand U20636 (N_20636,N_20301,N_20030);
nand U20637 (N_20637,N_20351,N_20189);
nand U20638 (N_20638,N_20220,N_20150);
and U20639 (N_20639,N_20417,N_20443);
and U20640 (N_20640,N_20414,N_20322);
xor U20641 (N_20641,N_20327,N_20142);
and U20642 (N_20642,N_20418,N_20176);
or U20643 (N_20643,N_20401,N_20234);
or U20644 (N_20644,N_20382,N_20408);
and U20645 (N_20645,N_20005,N_20474);
and U20646 (N_20646,N_20070,N_20188);
nor U20647 (N_20647,N_20405,N_20289);
nand U20648 (N_20648,N_20276,N_20248);
xor U20649 (N_20649,N_20469,N_20453);
or U20650 (N_20650,N_20272,N_20195);
nand U20651 (N_20651,N_20082,N_20173);
nor U20652 (N_20652,N_20343,N_20121);
nor U20653 (N_20653,N_20364,N_20193);
xnor U20654 (N_20654,N_20077,N_20172);
and U20655 (N_20655,N_20135,N_20154);
or U20656 (N_20656,N_20348,N_20489);
xor U20657 (N_20657,N_20130,N_20494);
and U20658 (N_20658,N_20416,N_20395);
or U20659 (N_20659,N_20375,N_20139);
nor U20660 (N_20660,N_20053,N_20462);
nor U20661 (N_20661,N_20455,N_20354);
or U20662 (N_20662,N_20473,N_20398);
or U20663 (N_20663,N_20206,N_20412);
and U20664 (N_20664,N_20126,N_20056);
and U20665 (N_20665,N_20251,N_20051);
and U20666 (N_20666,N_20068,N_20187);
or U20667 (N_20667,N_20029,N_20000);
xnor U20668 (N_20668,N_20336,N_20043);
or U20669 (N_20669,N_20303,N_20380);
or U20670 (N_20670,N_20399,N_20464);
nor U20671 (N_20671,N_20108,N_20089);
xor U20672 (N_20672,N_20376,N_20274);
nor U20673 (N_20673,N_20048,N_20071);
or U20674 (N_20674,N_20263,N_20454);
nor U20675 (N_20675,N_20174,N_20147);
nand U20676 (N_20676,N_20486,N_20438);
and U20677 (N_20677,N_20240,N_20296);
or U20678 (N_20678,N_20249,N_20361);
nor U20679 (N_20679,N_20222,N_20313);
and U20680 (N_20680,N_20295,N_20297);
xor U20681 (N_20681,N_20385,N_20406);
xnor U20682 (N_20682,N_20374,N_20255);
and U20683 (N_20683,N_20110,N_20184);
nand U20684 (N_20684,N_20342,N_20437);
xor U20685 (N_20685,N_20337,N_20389);
and U20686 (N_20686,N_20073,N_20140);
or U20687 (N_20687,N_20217,N_20449);
nand U20688 (N_20688,N_20387,N_20311);
or U20689 (N_20689,N_20164,N_20092);
nor U20690 (N_20690,N_20379,N_20320);
or U20691 (N_20691,N_20178,N_20330);
nand U20692 (N_20692,N_20099,N_20281);
xnor U20693 (N_20693,N_20085,N_20212);
and U20694 (N_20694,N_20194,N_20490);
nand U20695 (N_20695,N_20450,N_20169);
or U20696 (N_20696,N_20145,N_20488);
and U20697 (N_20697,N_20431,N_20498);
xnor U20698 (N_20698,N_20204,N_20006);
nor U20699 (N_20699,N_20155,N_20439);
nor U20700 (N_20700,N_20134,N_20200);
or U20701 (N_20701,N_20192,N_20020);
or U20702 (N_20702,N_20153,N_20179);
or U20703 (N_20703,N_20223,N_20141);
nor U20704 (N_20704,N_20114,N_20391);
xnor U20705 (N_20705,N_20144,N_20258);
or U20706 (N_20706,N_20309,N_20032);
nand U20707 (N_20707,N_20495,N_20036);
or U20708 (N_20708,N_20480,N_20411);
nand U20709 (N_20709,N_20035,N_20163);
and U20710 (N_20710,N_20022,N_20371);
or U20711 (N_20711,N_20407,N_20277);
or U20712 (N_20712,N_20430,N_20216);
and U20713 (N_20713,N_20451,N_20282);
or U20714 (N_20714,N_20060,N_20300);
and U20715 (N_20715,N_20064,N_20335);
and U20716 (N_20716,N_20122,N_20117);
and U20717 (N_20717,N_20102,N_20097);
xnor U20718 (N_20718,N_20170,N_20446);
nand U20719 (N_20719,N_20329,N_20264);
and U20720 (N_20720,N_20332,N_20012);
nor U20721 (N_20721,N_20347,N_20133);
or U20722 (N_20722,N_20410,N_20050);
nor U20723 (N_20723,N_20079,N_20103);
nand U20724 (N_20724,N_20362,N_20065);
nor U20725 (N_20725,N_20181,N_20441);
nor U20726 (N_20726,N_20368,N_20230);
and U20727 (N_20727,N_20096,N_20233);
nor U20728 (N_20728,N_20270,N_20237);
xor U20729 (N_20729,N_20105,N_20373);
or U20730 (N_20730,N_20186,N_20266);
nor U20731 (N_20731,N_20052,N_20285);
and U20732 (N_20732,N_20436,N_20316);
nor U20733 (N_20733,N_20472,N_20267);
and U20734 (N_20734,N_20010,N_20086);
or U20735 (N_20735,N_20482,N_20339);
or U20736 (N_20736,N_20182,N_20317);
xnor U20737 (N_20737,N_20075,N_20190);
xnor U20738 (N_20738,N_20353,N_20063);
and U20739 (N_20739,N_20499,N_20271);
nor U20740 (N_20740,N_20046,N_20384);
xor U20741 (N_20741,N_20390,N_20167);
or U20742 (N_20742,N_20491,N_20019);
nand U20743 (N_20743,N_20306,N_20162);
or U20744 (N_20744,N_20377,N_20492);
xnor U20745 (N_20745,N_20444,N_20344);
nand U20746 (N_20746,N_20257,N_20175);
nor U20747 (N_20747,N_20161,N_20305);
and U20748 (N_20748,N_20024,N_20308);
xnor U20749 (N_20749,N_20370,N_20136);
or U20750 (N_20750,N_20131,N_20053);
and U20751 (N_20751,N_20014,N_20016);
nor U20752 (N_20752,N_20013,N_20461);
and U20753 (N_20753,N_20441,N_20036);
xor U20754 (N_20754,N_20283,N_20126);
or U20755 (N_20755,N_20023,N_20124);
nor U20756 (N_20756,N_20252,N_20302);
xnor U20757 (N_20757,N_20069,N_20162);
nor U20758 (N_20758,N_20328,N_20426);
xnor U20759 (N_20759,N_20133,N_20277);
or U20760 (N_20760,N_20111,N_20181);
and U20761 (N_20761,N_20367,N_20410);
or U20762 (N_20762,N_20310,N_20444);
or U20763 (N_20763,N_20281,N_20021);
and U20764 (N_20764,N_20245,N_20053);
nor U20765 (N_20765,N_20088,N_20018);
or U20766 (N_20766,N_20144,N_20065);
xor U20767 (N_20767,N_20383,N_20272);
nor U20768 (N_20768,N_20250,N_20025);
nand U20769 (N_20769,N_20236,N_20146);
nor U20770 (N_20770,N_20455,N_20261);
and U20771 (N_20771,N_20420,N_20100);
nor U20772 (N_20772,N_20110,N_20043);
and U20773 (N_20773,N_20324,N_20425);
nand U20774 (N_20774,N_20472,N_20367);
nor U20775 (N_20775,N_20330,N_20200);
nand U20776 (N_20776,N_20203,N_20121);
nor U20777 (N_20777,N_20238,N_20296);
and U20778 (N_20778,N_20337,N_20324);
nor U20779 (N_20779,N_20120,N_20466);
and U20780 (N_20780,N_20047,N_20289);
or U20781 (N_20781,N_20469,N_20035);
nor U20782 (N_20782,N_20380,N_20173);
nor U20783 (N_20783,N_20496,N_20257);
and U20784 (N_20784,N_20298,N_20209);
or U20785 (N_20785,N_20491,N_20200);
and U20786 (N_20786,N_20472,N_20127);
nand U20787 (N_20787,N_20294,N_20152);
nand U20788 (N_20788,N_20251,N_20154);
or U20789 (N_20789,N_20288,N_20318);
xnor U20790 (N_20790,N_20162,N_20288);
nor U20791 (N_20791,N_20212,N_20478);
xnor U20792 (N_20792,N_20010,N_20453);
or U20793 (N_20793,N_20328,N_20386);
xnor U20794 (N_20794,N_20268,N_20025);
nor U20795 (N_20795,N_20368,N_20437);
xor U20796 (N_20796,N_20257,N_20468);
or U20797 (N_20797,N_20371,N_20175);
and U20798 (N_20798,N_20266,N_20331);
or U20799 (N_20799,N_20456,N_20069);
or U20800 (N_20800,N_20129,N_20347);
or U20801 (N_20801,N_20248,N_20027);
or U20802 (N_20802,N_20300,N_20374);
nand U20803 (N_20803,N_20315,N_20356);
nand U20804 (N_20804,N_20278,N_20188);
nor U20805 (N_20805,N_20078,N_20356);
nor U20806 (N_20806,N_20325,N_20247);
nor U20807 (N_20807,N_20248,N_20139);
nand U20808 (N_20808,N_20349,N_20052);
nor U20809 (N_20809,N_20115,N_20034);
or U20810 (N_20810,N_20475,N_20196);
or U20811 (N_20811,N_20157,N_20273);
nand U20812 (N_20812,N_20425,N_20341);
or U20813 (N_20813,N_20288,N_20025);
and U20814 (N_20814,N_20067,N_20212);
and U20815 (N_20815,N_20084,N_20488);
and U20816 (N_20816,N_20066,N_20426);
xnor U20817 (N_20817,N_20236,N_20460);
and U20818 (N_20818,N_20217,N_20023);
or U20819 (N_20819,N_20212,N_20344);
and U20820 (N_20820,N_20084,N_20083);
or U20821 (N_20821,N_20157,N_20061);
xor U20822 (N_20822,N_20109,N_20445);
nor U20823 (N_20823,N_20387,N_20468);
and U20824 (N_20824,N_20287,N_20115);
nand U20825 (N_20825,N_20427,N_20289);
xor U20826 (N_20826,N_20490,N_20446);
or U20827 (N_20827,N_20266,N_20020);
xnor U20828 (N_20828,N_20353,N_20184);
nor U20829 (N_20829,N_20106,N_20289);
xnor U20830 (N_20830,N_20107,N_20280);
nor U20831 (N_20831,N_20067,N_20475);
and U20832 (N_20832,N_20117,N_20409);
or U20833 (N_20833,N_20490,N_20358);
xnor U20834 (N_20834,N_20264,N_20360);
nor U20835 (N_20835,N_20325,N_20046);
and U20836 (N_20836,N_20089,N_20110);
or U20837 (N_20837,N_20326,N_20375);
xnor U20838 (N_20838,N_20185,N_20491);
or U20839 (N_20839,N_20320,N_20293);
or U20840 (N_20840,N_20280,N_20000);
xnor U20841 (N_20841,N_20200,N_20458);
and U20842 (N_20842,N_20096,N_20000);
or U20843 (N_20843,N_20151,N_20144);
nor U20844 (N_20844,N_20113,N_20447);
xor U20845 (N_20845,N_20249,N_20188);
or U20846 (N_20846,N_20175,N_20408);
and U20847 (N_20847,N_20105,N_20199);
or U20848 (N_20848,N_20250,N_20138);
xnor U20849 (N_20849,N_20304,N_20330);
and U20850 (N_20850,N_20430,N_20166);
nand U20851 (N_20851,N_20156,N_20441);
nor U20852 (N_20852,N_20078,N_20114);
and U20853 (N_20853,N_20172,N_20134);
or U20854 (N_20854,N_20260,N_20171);
nor U20855 (N_20855,N_20430,N_20460);
xnor U20856 (N_20856,N_20494,N_20016);
and U20857 (N_20857,N_20478,N_20486);
nand U20858 (N_20858,N_20138,N_20068);
or U20859 (N_20859,N_20196,N_20474);
and U20860 (N_20860,N_20184,N_20286);
or U20861 (N_20861,N_20281,N_20116);
nor U20862 (N_20862,N_20302,N_20349);
and U20863 (N_20863,N_20267,N_20221);
and U20864 (N_20864,N_20466,N_20377);
and U20865 (N_20865,N_20405,N_20047);
xnor U20866 (N_20866,N_20192,N_20404);
xor U20867 (N_20867,N_20171,N_20317);
nor U20868 (N_20868,N_20350,N_20326);
xor U20869 (N_20869,N_20252,N_20116);
xor U20870 (N_20870,N_20335,N_20237);
and U20871 (N_20871,N_20075,N_20220);
or U20872 (N_20872,N_20292,N_20317);
nor U20873 (N_20873,N_20124,N_20455);
and U20874 (N_20874,N_20364,N_20484);
or U20875 (N_20875,N_20487,N_20431);
nand U20876 (N_20876,N_20324,N_20247);
or U20877 (N_20877,N_20357,N_20374);
nor U20878 (N_20878,N_20045,N_20290);
nor U20879 (N_20879,N_20264,N_20456);
and U20880 (N_20880,N_20217,N_20495);
and U20881 (N_20881,N_20117,N_20402);
nor U20882 (N_20882,N_20215,N_20469);
nand U20883 (N_20883,N_20212,N_20266);
or U20884 (N_20884,N_20280,N_20004);
nor U20885 (N_20885,N_20286,N_20280);
and U20886 (N_20886,N_20386,N_20139);
xnor U20887 (N_20887,N_20226,N_20390);
xor U20888 (N_20888,N_20303,N_20439);
and U20889 (N_20889,N_20030,N_20357);
nor U20890 (N_20890,N_20102,N_20026);
or U20891 (N_20891,N_20124,N_20159);
nor U20892 (N_20892,N_20176,N_20318);
nor U20893 (N_20893,N_20289,N_20397);
nand U20894 (N_20894,N_20386,N_20459);
and U20895 (N_20895,N_20315,N_20228);
nand U20896 (N_20896,N_20382,N_20421);
xor U20897 (N_20897,N_20264,N_20219);
xnor U20898 (N_20898,N_20016,N_20073);
and U20899 (N_20899,N_20122,N_20318);
and U20900 (N_20900,N_20130,N_20170);
nand U20901 (N_20901,N_20308,N_20116);
nand U20902 (N_20902,N_20450,N_20435);
and U20903 (N_20903,N_20103,N_20245);
or U20904 (N_20904,N_20146,N_20112);
nor U20905 (N_20905,N_20135,N_20308);
and U20906 (N_20906,N_20286,N_20268);
nand U20907 (N_20907,N_20035,N_20389);
xor U20908 (N_20908,N_20278,N_20213);
and U20909 (N_20909,N_20214,N_20442);
xor U20910 (N_20910,N_20338,N_20455);
xnor U20911 (N_20911,N_20093,N_20080);
or U20912 (N_20912,N_20446,N_20391);
xnor U20913 (N_20913,N_20028,N_20310);
or U20914 (N_20914,N_20314,N_20390);
nor U20915 (N_20915,N_20390,N_20133);
nor U20916 (N_20916,N_20036,N_20214);
or U20917 (N_20917,N_20110,N_20012);
and U20918 (N_20918,N_20065,N_20328);
nand U20919 (N_20919,N_20173,N_20463);
nor U20920 (N_20920,N_20053,N_20497);
xor U20921 (N_20921,N_20265,N_20126);
nor U20922 (N_20922,N_20193,N_20366);
nor U20923 (N_20923,N_20293,N_20384);
or U20924 (N_20924,N_20402,N_20421);
and U20925 (N_20925,N_20248,N_20416);
xnor U20926 (N_20926,N_20135,N_20304);
xnor U20927 (N_20927,N_20136,N_20350);
or U20928 (N_20928,N_20402,N_20223);
nand U20929 (N_20929,N_20070,N_20228);
nand U20930 (N_20930,N_20243,N_20423);
and U20931 (N_20931,N_20125,N_20318);
nand U20932 (N_20932,N_20369,N_20070);
nor U20933 (N_20933,N_20413,N_20383);
and U20934 (N_20934,N_20267,N_20019);
xor U20935 (N_20935,N_20035,N_20473);
xnor U20936 (N_20936,N_20156,N_20116);
or U20937 (N_20937,N_20156,N_20456);
xor U20938 (N_20938,N_20128,N_20177);
or U20939 (N_20939,N_20394,N_20206);
xor U20940 (N_20940,N_20333,N_20296);
and U20941 (N_20941,N_20373,N_20237);
nor U20942 (N_20942,N_20091,N_20449);
and U20943 (N_20943,N_20163,N_20277);
nand U20944 (N_20944,N_20075,N_20146);
xnor U20945 (N_20945,N_20470,N_20489);
xor U20946 (N_20946,N_20435,N_20060);
or U20947 (N_20947,N_20133,N_20065);
nor U20948 (N_20948,N_20357,N_20213);
or U20949 (N_20949,N_20339,N_20439);
or U20950 (N_20950,N_20035,N_20240);
or U20951 (N_20951,N_20087,N_20062);
nor U20952 (N_20952,N_20001,N_20313);
and U20953 (N_20953,N_20335,N_20104);
nand U20954 (N_20954,N_20332,N_20009);
xor U20955 (N_20955,N_20313,N_20343);
nor U20956 (N_20956,N_20391,N_20204);
xnor U20957 (N_20957,N_20030,N_20243);
nor U20958 (N_20958,N_20137,N_20066);
or U20959 (N_20959,N_20136,N_20064);
or U20960 (N_20960,N_20011,N_20446);
nand U20961 (N_20961,N_20185,N_20126);
and U20962 (N_20962,N_20021,N_20384);
nand U20963 (N_20963,N_20266,N_20432);
nor U20964 (N_20964,N_20132,N_20306);
xnor U20965 (N_20965,N_20329,N_20317);
nor U20966 (N_20966,N_20015,N_20496);
nand U20967 (N_20967,N_20026,N_20313);
nand U20968 (N_20968,N_20406,N_20214);
xnor U20969 (N_20969,N_20308,N_20239);
nand U20970 (N_20970,N_20277,N_20264);
or U20971 (N_20971,N_20389,N_20326);
and U20972 (N_20972,N_20366,N_20380);
nand U20973 (N_20973,N_20493,N_20176);
xor U20974 (N_20974,N_20128,N_20009);
and U20975 (N_20975,N_20434,N_20126);
or U20976 (N_20976,N_20194,N_20239);
or U20977 (N_20977,N_20363,N_20494);
or U20978 (N_20978,N_20086,N_20324);
or U20979 (N_20979,N_20195,N_20377);
or U20980 (N_20980,N_20229,N_20440);
xnor U20981 (N_20981,N_20475,N_20440);
or U20982 (N_20982,N_20042,N_20460);
nor U20983 (N_20983,N_20479,N_20371);
or U20984 (N_20984,N_20020,N_20075);
and U20985 (N_20985,N_20439,N_20287);
xnor U20986 (N_20986,N_20387,N_20345);
xor U20987 (N_20987,N_20415,N_20328);
nand U20988 (N_20988,N_20252,N_20294);
or U20989 (N_20989,N_20491,N_20138);
xor U20990 (N_20990,N_20457,N_20050);
nand U20991 (N_20991,N_20274,N_20109);
nand U20992 (N_20992,N_20240,N_20469);
or U20993 (N_20993,N_20107,N_20400);
xnor U20994 (N_20994,N_20138,N_20237);
and U20995 (N_20995,N_20068,N_20236);
or U20996 (N_20996,N_20177,N_20392);
xnor U20997 (N_20997,N_20328,N_20329);
xnor U20998 (N_20998,N_20256,N_20270);
nor U20999 (N_20999,N_20041,N_20472);
or U21000 (N_21000,N_20979,N_20918);
nor U21001 (N_21001,N_20581,N_20559);
and U21002 (N_21002,N_20947,N_20861);
and U21003 (N_21003,N_20515,N_20545);
and U21004 (N_21004,N_20969,N_20792);
nor U21005 (N_21005,N_20785,N_20552);
and U21006 (N_21006,N_20822,N_20596);
or U21007 (N_21007,N_20595,N_20733);
or U21008 (N_21008,N_20855,N_20982);
xor U21009 (N_21009,N_20864,N_20632);
nor U21010 (N_21010,N_20702,N_20839);
nor U21011 (N_21011,N_20820,N_20578);
nand U21012 (N_21012,N_20699,N_20629);
nand U21013 (N_21013,N_20992,N_20787);
nor U21014 (N_21014,N_20602,N_20797);
xor U21015 (N_21015,N_20741,N_20932);
nand U21016 (N_21016,N_20843,N_20951);
nand U21017 (N_21017,N_20607,N_20728);
and U21018 (N_21018,N_20533,N_20664);
nand U21019 (N_21019,N_20924,N_20724);
xor U21020 (N_21020,N_20916,N_20673);
and U21021 (N_21021,N_20646,N_20663);
or U21022 (N_21022,N_20966,N_20716);
xnor U21023 (N_21023,N_20621,N_20866);
xor U21024 (N_21024,N_20616,N_20972);
xor U21025 (N_21025,N_20833,N_20897);
and U21026 (N_21026,N_20734,N_20524);
and U21027 (N_21027,N_20744,N_20990);
or U21028 (N_21028,N_20676,N_20721);
nand U21029 (N_21029,N_20917,N_20809);
nor U21030 (N_21030,N_20688,N_20960);
and U21031 (N_21031,N_20998,N_20693);
or U21032 (N_21032,N_20510,N_20643);
and U21033 (N_21033,N_20887,N_20853);
xor U21034 (N_21034,N_20574,N_20652);
nor U21035 (N_21035,N_20747,N_20586);
xnor U21036 (N_21036,N_20715,N_20898);
and U21037 (N_21037,N_20900,N_20953);
and U21038 (N_21038,N_20896,N_20889);
and U21039 (N_21039,N_20644,N_20776);
nand U21040 (N_21040,N_20504,N_20692);
or U21041 (N_21041,N_20807,N_20878);
or U21042 (N_21042,N_20931,N_20937);
nor U21043 (N_21043,N_20973,N_20726);
nor U21044 (N_21044,N_20500,N_20869);
or U21045 (N_21045,N_20709,N_20725);
xnor U21046 (N_21046,N_20752,N_20848);
xnor U21047 (N_21047,N_20825,N_20817);
or U21048 (N_21048,N_20534,N_20984);
nand U21049 (N_21049,N_20642,N_20773);
xnor U21050 (N_21050,N_20767,N_20580);
nor U21051 (N_21051,N_20794,N_20899);
nand U21052 (N_21052,N_20712,N_20964);
or U21053 (N_21053,N_20628,N_20711);
and U21054 (N_21054,N_20668,N_20570);
and U21055 (N_21055,N_20610,N_20930);
or U21056 (N_21056,N_20876,N_20557);
or U21057 (N_21057,N_20754,N_20888);
or U21058 (N_21058,N_20637,N_20775);
nand U21059 (N_21059,N_20626,N_20554);
and U21060 (N_21060,N_20701,N_20849);
xor U21061 (N_21061,N_20880,N_20885);
xnor U21062 (N_21062,N_20913,N_20934);
or U21063 (N_21063,N_20708,N_20871);
xnor U21064 (N_21064,N_20983,N_20971);
nor U21065 (N_21065,N_20999,N_20836);
or U21066 (N_21066,N_20751,N_20639);
xor U21067 (N_21067,N_20538,N_20891);
or U21068 (N_21068,N_20868,N_20525);
or U21069 (N_21069,N_20697,N_20567);
or U21070 (N_21070,N_20873,N_20519);
or U21071 (N_21071,N_20894,N_20845);
xor U21072 (N_21072,N_20617,N_20748);
xor U21073 (N_21073,N_20745,N_20682);
xnor U21074 (N_21074,N_20997,N_20834);
xor U21075 (N_21075,N_20638,N_20563);
or U21076 (N_21076,N_20739,N_20656);
nor U21077 (N_21077,N_20771,N_20886);
nor U21078 (N_21078,N_20690,N_20605);
and U21079 (N_21079,N_20687,N_20950);
nor U21080 (N_21080,N_20561,N_20974);
nor U21081 (N_21081,N_20755,N_20929);
xor U21082 (N_21082,N_20842,N_20501);
xor U21083 (N_21083,N_20890,N_20719);
xnor U21084 (N_21084,N_20986,N_20781);
nand U21085 (N_21085,N_20603,N_20933);
or U21086 (N_21086,N_20989,N_20938);
and U21087 (N_21087,N_20981,N_20750);
and U21088 (N_21088,N_20922,N_20592);
nor U21089 (N_21089,N_20641,N_20671);
and U21090 (N_21090,N_20810,N_20847);
or U21091 (N_21091,N_20818,N_20669);
nand U21092 (N_21092,N_20795,N_20939);
and U21093 (N_21093,N_20560,N_20985);
or U21094 (N_21094,N_20650,N_20941);
nor U21095 (N_21095,N_20620,N_20507);
xor U21096 (N_21096,N_20530,N_20689);
nor U21097 (N_21097,N_20505,N_20928);
or U21098 (N_21098,N_20686,N_20920);
and U21099 (N_21099,N_20582,N_20980);
nand U21100 (N_21100,N_20906,N_20838);
nand U21101 (N_21101,N_20753,N_20766);
nand U21102 (N_21102,N_20713,N_20816);
nor U21103 (N_21103,N_20824,N_20837);
nand U21104 (N_21104,N_20800,N_20539);
or U21105 (N_21105,N_20805,N_20779);
xor U21106 (N_21106,N_20511,N_20556);
xor U21107 (N_21107,N_20698,N_20940);
and U21108 (N_21108,N_20593,N_20865);
xnor U21109 (N_21109,N_20529,N_20901);
xor U21110 (N_21110,N_20679,N_20909);
or U21111 (N_21111,N_20618,N_20640);
nand U21112 (N_21112,N_20589,N_20662);
and U21113 (N_21113,N_20881,N_20978);
xnor U21114 (N_21114,N_20604,N_20811);
xnor U21115 (N_21115,N_20700,N_20718);
xor U21116 (N_21116,N_20970,N_20743);
nand U21117 (N_21117,N_20892,N_20919);
xnor U21118 (N_21118,N_20757,N_20536);
or U21119 (N_21119,N_20645,N_20935);
nor U21120 (N_21120,N_20761,N_20846);
nand U21121 (N_21121,N_20942,N_20691);
xor U21122 (N_21122,N_20550,N_20819);
or U21123 (N_21123,N_20995,N_20526);
and U21124 (N_21124,N_20571,N_20841);
and U21125 (N_21125,N_20591,N_20584);
nand U21126 (N_21126,N_20749,N_20553);
or U21127 (N_21127,N_20952,N_20948);
nand U21128 (N_21128,N_20569,N_20936);
nand U21129 (N_21129,N_20636,N_20883);
nor U21130 (N_21130,N_20949,N_20588);
or U21131 (N_21131,N_20742,N_20677);
nor U21132 (N_21132,N_20625,N_20506);
and U21133 (N_21133,N_20562,N_20587);
nor U21134 (N_21134,N_20812,N_20695);
nor U21135 (N_21135,N_20925,N_20655);
or U21136 (N_21136,N_20759,N_20723);
nor U21137 (N_21137,N_20568,N_20532);
or U21138 (N_21138,N_20879,N_20583);
xor U21139 (N_21139,N_20597,N_20903);
xnor U21140 (N_21140,N_20544,N_20905);
nand U21141 (N_21141,N_20826,N_20962);
and U21142 (N_21142,N_20512,N_20672);
nor U21143 (N_21143,N_20904,N_20710);
or U21144 (N_21144,N_20804,N_20793);
or U21145 (N_21145,N_20872,N_20851);
nand U21146 (N_21146,N_20784,N_20543);
or U21147 (N_21147,N_20615,N_20944);
xor U21148 (N_21148,N_20835,N_20914);
and U21149 (N_21149,N_20730,N_20514);
xnor U21150 (N_21150,N_20831,N_20943);
xor U21151 (N_21151,N_20572,N_20762);
nand U21152 (N_21152,N_20778,N_20874);
nor U21153 (N_21153,N_20737,N_20957);
xor U21154 (N_21154,N_20911,N_20675);
or U21155 (N_21155,N_20707,N_20798);
or U21156 (N_21156,N_20653,N_20564);
nor U21157 (N_21157,N_20867,N_20852);
or U21158 (N_21158,N_20738,N_20786);
or U21159 (N_21159,N_20518,N_20746);
nand U21160 (N_21160,N_20956,N_20788);
or U21161 (N_21161,N_20722,N_20624);
xnor U21162 (N_21162,N_20665,N_20594);
xnor U21163 (N_21163,N_20828,N_20893);
and U21164 (N_21164,N_20740,N_20796);
xnor U21165 (N_21165,N_20667,N_20977);
or U21166 (N_21166,N_20736,N_20954);
nand U21167 (N_21167,N_20609,N_20599);
or U21168 (N_21168,N_20627,N_20541);
nand U21169 (N_21169,N_20635,N_20546);
or U21170 (N_21170,N_20806,N_20774);
nand U21171 (N_21171,N_20622,N_20555);
or U21172 (N_21172,N_20558,N_20516);
and U21173 (N_21173,N_20661,N_20996);
xnor U21174 (N_21174,N_20576,N_20912);
xnor U21175 (N_21175,N_20683,N_20613);
nor U21176 (N_21176,N_20821,N_20877);
nor U21177 (N_21177,N_20769,N_20577);
and U21178 (N_21178,N_20651,N_20684);
nor U21179 (N_21179,N_20542,N_20731);
or U21180 (N_21180,N_20907,N_20720);
nand U21181 (N_21181,N_20658,N_20975);
xor U21182 (N_21182,N_20850,N_20991);
xor U21183 (N_21183,N_20703,N_20612);
xnor U21184 (N_21184,N_20783,N_20548);
nand U21185 (N_21185,N_20598,N_20963);
or U21186 (N_21186,N_20670,N_20790);
nand U21187 (N_21187,N_20647,N_20791);
nor U21188 (N_21188,N_20657,N_20801);
or U21189 (N_21189,N_20884,N_20955);
and U21190 (N_21190,N_20517,N_20993);
or U21191 (N_21191,N_20923,N_20858);
and U21192 (N_21192,N_20531,N_20863);
nand U21193 (N_21193,N_20631,N_20648);
nand U21194 (N_21194,N_20927,N_20520);
nor U21195 (N_21195,N_20535,N_20802);
or U21196 (N_21196,N_20777,N_20547);
or U21197 (N_21197,N_20976,N_20813);
and U21198 (N_21198,N_20523,N_20606);
nor U21199 (N_21199,N_20967,N_20573);
xor U21200 (N_21200,N_20674,N_20756);
nor U21201 (N_21201,N_20860,N_20945);
or U21202 (N_21202,N_20854,N_20946);
nor U21203 (N_21203,N_20528,N_20765);
nor U21204 (N_21204,N_20717,N_20857);
xor U21205 (N_21205,N_20910,N_20611);
nor U21206 (N_21206,N_20830,N_20799);
or U21207 (N_21207,N_20988,N_20649);
and U21208 (N_21208,N_20870,N_20882);
and U21209 (N_21209,N_20961,N_20875);
or U21210 (N_21210,N_20782,N_20705);
xnor U21211 (N_21211,N_20590,N_20729);
xnor U21212 (N_21212,N_20522,N_20508);
nand U21213 (N_21213,N_20549,N_20565);
and U21214 (N_21214,N_20566,N_20763);
xor U21215 (N_21215,N_20965,N_20681);
and U21216 (N_21216,N_20823,N_20680);
or U21217 (N_21217,N_20630,N_20908);
and U21218 (N_21218,N_20660,N_20829);
xor U21219 (N_21219,N_20634,N_20768);
xor U21220 (N_21220,N_20994,N_20902);
or U21221 (N_21221,N_20633,N_20732);
and U21222 (N_21222,N_20540,N_20601);
nand U21223 (N_21223,N_20921,N_20770);
and U21224 (N_21224,N_20727,N_20958);
and U21225 (N_21225,N_20502,N_20527);
nand U21226 (N_21226,N_20968,N_20803);
and U21227 (N_21227,N_20959,N_20814);
xnor U21228 (N_21228,N_20862,N_20614);
and U21229 (N_21229,N_20780,N_20513);
or U21230 (N_21230,N_20859,N_20832);
and U21231 (N_21231,N_20600,N_20895);
and U21232 (N_21232,N_20666,N_20503);
nand U21233 (N_21233,N_20579,N_20608);
and U21234 (N_21234,N_20537,N_20808);
nand U21235 (N_21235,N_20619,N_20575);
and U21236 (N_21236,N_20987,N_20704);
nor U21237 (N_21237,N_20714,N_20654);
nand U21238 (N_21238,N_20789,N_20840);
xnor U21239 (N_21239,N_20678,N_20926);
nand U21240 (N_21240,N_20623,N_20706);
and U21241 (N_21241,N_20856,N_20915);
and U21242 (N_21242,N_20735,N_20827);
and U21243 (N_21243,N_20685,N_20521);
xor U21244 (N_21244,N_20551,N_20760);
xnor U21245 (N_21245,N_20585,N_20815);
and U21246 (N_21246,N_20758,N_20696);
nand U21247 (N_21247,N_20694,N_20509);
xor U21248 (N_21248,N_20764,N_20772);
nor U21249 (N_21249,N_20659,N_20844);
nand U21250 (N_21250,N_20684,N_20778);
and U21251 (N_21251,N_20521,N_20625);
or U21252 (N_21252,N_20620,N_20527);
or U21253 (N_21253,N_20821,N_20601);
nor U21254 (N_21254,N_20605,N_20583);
or U21255 (N_21255,N_20840,N_20550);
nand U21256 (N_21256,N_20923,N_20924);
and U21257 (N_21257,N_20568,N_20769);
and U21258 (N_21258,N_20927,N_20739);
or U21259 (N_21259,N_20715,N_20555);
nor U21260 (N_21260,N_20875,N_20731);
nor U21261 (N_21261,N_20835,N_20841);
or U21262 (N_21262,N_20612,N_20737);
nor U21263 (N_21263,N_20993,N_20869);
nor U21264 (N_21264,N_20743,N_20973);
xor U21265 (N_21265,N_20933,N_20822);
nor U21266 (N_21266,N_20676,N_20886);
nor U21267 (N_21267,N_20642,N_20781);
nor U21268 (N_21268,N_20785,N_20856);
xor U21269 (N_21269,N_20713,N_20769);
nand U21270 (N_21270,N_20707,N_20669);
nor U21271 (N_21271,N_20705,N_20548);
or U21272 (N_21272,N_20995,N_20904);
xor U21273 (N_21273,N_20540,N_20738);
nand U21274 (N_21274,N_20659,N_20527);
nor U21275 (N_21275,N_20610,N_20687);
nand U21276 (N_21276,N_20701,N_20746);
xor U21277 (N_21277,N_20574,N_20763);
xnor U21278 (N_21278,N_20730,N_20581);
or U21279 (N_21279,N_20942,N_20804);
and U21280 (N_21280,N_20560,N_20535);
and U21281 (N_21281,N_20813,N_20509);
xnor U21282 (N_21282,N_20917,N_20680);
nor U21283 (N_21283,N_20919,N_20947);
nand U21284 (N_21284,N_20913,N_20816);
nand U21285 (N_21285,N_20708,N_20999);
nand U21286 (N_21286,N_20710,N_20720);
nor U21287 (N_21287,N_20985,N_20960);
and U21288 (N_21288,N_20586,N_20577);
and U21289 (N_21289,N_20640,N_20830);
nand U21290 (N_21290,N_20609,N_20822);
nand U21291 (N_21291,N_20765,N_20667);
xor U21292 (N_21292,N_20865,N_20588);
or U21293 (N_21293,N_20652,N_20849);
or U21294 (N_21294,N_20878,N_20523);
or U21295 (N_21295,N_20809,N_20994);
and U21296 (N_21296,N_20954,N_20993);
nand U21297 (N_21297,N_20896,N_20852);
nand U21298 (N_21298,N_20770,N_20934);
nor U21299 (N_21299,N_20882,N_20510);
xnor U21300 (N_21300,N_20775,N_20928);
nand U21301 (N_21301,N_20731,N_20522);
and U21302 (N_21302,N_20617,N_20971);
or U21303 (N_21303,N_20541,N_20573);
nand U21304 (N_21304,N_20988,N_20658);
nand U21305 (N_21305,N_20528,N_20951);
nor U21306 (N_21306,N_20961,N_20820);
nor U21307 (N_21307,N_20955,N_20928);
nor U21308 (N_21308,N_20794,N_20726);
xnor U21309 (N_21309,N_20903,N_20881);
and U21310 (N_21310,N_20887,N_20985);
nand U21311 (N_21311,N_20587,N_20512);
nor U21312 (N_21312,N_20912,N_20743);
xor U21313 (N_21313,N_20630,N_20673);
nand U21314 (N_21314,N_20807,N_20560);
xor U21315 (N_21315,N_20557,N_20584);
or U21316 (N_21316,N_20812,N_20567);
or U21317 (N_21317,N_20747,N_20598);
nor U21318 (N_21318,N_20993,N_20543);
nor U21319 (N_21319,N_20754,N_20767);
nand U21320 (N_21320,N_20677,N_20724);
or U21321 (N_21321,N_20966,N_20787);
nand U21322 (N_21322,N_20823,N_20827);
xor U21323 (N_21323,N_20726,N_20713);
or U21324 (N_21324,N_20627,N_20649);
nor U21325 (N_21325,N_20799,N_20598);
and U21326 (N_21326,N_20907,N_20705);
or U21327 (N_21327,N_20558,N_20658);
nand U21328 (N_21328,N_20736,N_20925);
and U21329 (N_21329,N_20575,N_20966);
nor U21330 (N_21330,N_20649,N_20859);
xnor U21331 (N_21331,N_20720,N_20958);
nor U21332 (N_21332,N_20600,N_20630);
nand U21333 (N_21333,N_20593,N_20561);
xnor U21334 (N_21334,N_20540,N_20500);
nand U21335 (N_21335,N_20553,N_20600);
or U21336 (N_21336,N_20837,N_20556);
or U21337 (N_21337,N_20714,N_20953);
nand U21338 (N_21338,N_20594,N_20638);
nand U21339 (N_21339,N_20736,N_20865);
xnor U21340 (N_21340,N_20612,N_20877);
or U21341 (N_21341,N_20800,N_20586);
nor U21342 (N_21342,N_20955,N_20604);
nor U21343 (N_21343,N_20956,N_20519);
and U21344 (N_21344,N_20636,N_20606);
nand U21345 (N_21345,N_20644,N_20926);
and U21346 (N_21346,N_20998,N_20931);
nand U21347 (N_21347,N_20790,N_20928);
nor U21348 (N_21348,N_20834,N_20859);
xnor U21349 (N_21349,N_20530,N_20641);
or U21350 (N_21350,N_20927,N_20544);
nand U21351 (N_21351,N_20905,N_20958);
nor U21352 (N_21352,N_20796,N_20938);
xor U21353 (N_21353,N_20830,N_20945);
xor U21354 (N_21354,N_20515,N_20818);
xnor U21355 (N_21355,N_20511,N_20525);
or U21356 (N_21356,N_20997,N_20776);
nand U21357 (N_21357,N_20677,N_20988);
or U21358 (N_21358,N_20993,N_20974);
and U21359 (N_21359,N_20616,N_20925);
and U21360 (N_21360,N_20969,N_20908);
nor U21361 (N_21361,N_20844,N_20895);
or U21362 (N_21362,N_20664,N_20762);
nand U21363 (N_21363,N_20610,N_20646);
nor U21364 (N_21364,N_20539,N_20546);
or U21365 (N_21365,N_20811,N_20715);
nand U21366 (N_21366,N_20652,N_20824);
nor U21367 (N_21367,N_20994,N_20628);
xnor U21368 (N_21368,N_20684,N_20540);
nand U21369 (N_21369,N_20952,N_20978);
nor U21370 (N_21370,N_20830,N_20785);
nor U21371 (N_21371,N_20613,N_20891);
xnor U21372 (N_21372,N_20515,N_20900);
nand U21373 (N_21373,N_20836,N_20712);
nand U21374 (N_21374,N_20716,N_20673);
and U21375 (N_21375,N_20713,N_20746);
xor U21376 (N_21376,N_20633,N_20827);
nand U21377 (N_21377,N_20685,N_20878);
or U21378 (N_21378,N_20863,N_20892);
nand U21379 (N_21379,N_20602,N_20532);
xnor U21380 (N_21380,N_20687,N_20890);
xnor U21381 (N_21381,N_20551,N_20739);
nand U21382 (N_21382,N_20968,N_20821);
nand U21383 (N_21383,N_20972,N_20504);
nor U21384 (N_21384,N_20785,N_20945);
nor U21385 (N_21385,N_20913,N_20907);
and U21386 (N_21386,N_20934,N_20701);
nand U21387 (N_21387,N_20837,N_20580);
nand U21388 (N_21388,N_20870,N_20846);
and U21389 (N_21389,N_20924,N_20863);
nor U21390 (N_21390,N_20976,N_20612);
xor U21391 (N_21391,N_20860,N_20702);
nor U21392 (N_21392,N_20642,N_20981);
nand U21393 (N_21393,N_20529,N_20795);
nand U21394 (N_21394,N_20695,N_20923);
and U21395 (N_21395,N_20877,N_20657);
or U21396 (N_21396,N_20524,N_20553);
nand U21397 (N_21397,N_20865,N_20513);
nor U21398 (N_21398,N_20708,N_20549);
nor U21399 (N_21399,N_20988,N_20640);
xor U21400 (N_21400,N_20922,N_20865);
xnor U21401 (N_21401,N_20934,N_20837);
nor U21402 (N_21402,N_20577,N_20551);
or U21403 (N_21403,N_20980,N_20806);
or U21404 (N_21404,N_20911,N_20592);
nor U21405 (N_21405,N_20971,N_20596);
or U21406 (N_21406,N_20529,N_20567);
xor U21407 (N_21407,N_20766,N_20703);
or U21408 (N_21408,N_20965,N_20774);
xor U21409 (N_21409,N_20857,N_20824);
nor U21410 (N_21410,N_20939,N_20620);
xor U21411 (N_21411,N_20881,N_20854);
xor U21412 (N_21412,N_20849,N_20893);
nor U21413 (N_21413,N_20870,N_20916);
nand U21414 (N_21414,N_20516,N_20723);
xor U21415 (N_21415,N_20680,N_20595);
nand U21416 (N_21416,N_20565,N_20889);
nand U21417 (N_21417,N_20596,N_20542);
nand U21418 (N_21418,N_20567,N_20690);
or U21419 (N_21419,N_20616,N_20613);
xor U21420 (N_21420,N_20768,N_20638);
nor U21421 (N_21421,N_20512,N_20609);
xnor U21422 (N_21422,N_20935,N_20611);
nand U21423 (N_21423,N_20707,N_20916);
and U21424 (N_21424,N_20850,N_20726);
nor U21425 (N_21425,N_20507,N_20568);
xnor U21426 (N_21426,N_20852,N_20897);
xor U21427 (N_21427,N_20967,N_20931);
nand U21428 (N_21428,N_20635,N_20746);
xnor U21429 (N_21429,N_20536,N_20692);
or U21430 (N_21430,N_20791,N_20906);
or U21431 (N_21431,N_20800,N_20929);
nor U21432 (N_21432,N_20737,N_20991);
nand U21433 (N_21433,N_20711,N_20968);
and U21434 (N_21434,N_20743,N_20698);
nor U21435 (N_21435,N_20787,N_20727);
nand U21436 (N_21436,N_20892,N_20965);
and U21437 (N_21437,N_20551,N_20738);
xor U21438 (N_21438,N_20689,N_20824);
and U21439 (N_21439,N_20885,N_20898);
and U21440 (N_21440,N_20507,N_20723);
or U21441 (N_21441,N_20769,N_20704);
nand U21442 (N_21442,N_20702,N_20987);
and U21443 (N_21443,N_20791,N_20767);
or U21444 (N_21444,N_20907,N_20818);
or U21445 (N_21445,N_20658,N_20508);
xor U21446 (N_21446,N_20751,N_20946);
nand U21447 (N_21447,N_20982,N_20682);
or U21448 (N_21448,N_20932,N_20714);
nand U21449 (N_21449,N_20982,N_20546);
nand U21450 (N_21450,N_20663,N_20868);
nand U21451 (N_21451,N_20812,N_20913);
and U21452 (N_21452,N_20891,N_20907);
nand U21453 (N_21453,N_20993,N_20677);
xnor U21454 (N_21454,N_20833,N_20671);
xnor U21455 (N_21455,N_20911,N_20785);
nand U21456 (N_21456,N_20763,N_20719);
xnor U21457 (N_21457,N_20676,N_20713);
and U21458 (N_21458,N_20528,N_20944);
nand U21459 (N_21459,N_20772,N_20530);
xor U21460 (N_21460,N_20845,N_20642);
nand U21461 (N_21461,N_20658,N_20616);
or U21462 (N_21462,N_20753,N_20539);
and U21463 (N_21463,N_20517,N_20891);
and U21464 (N_21464,N_20871,N_20950);
and U21465 (N_21465,N_20552,N_20945);
xor U21466 (N_21466,N_20541,N_20610);
nand U21467 (N_21467,N_20693,N_20931);
xnor U21468 (N_21468,N_20695,N_20869);
or U21469 (N_21469,N_20588,N_20655);
nor U21470 (N_21470,N_20797,N_20812);
nand U21471 (N_21471,N_20593,N_20951);
nor U21472 (N_21472,N_20512,N_20707);
nor U21473 (N_21473,N_20533,N_20819);
xor U21474 (N_21474,N_20921,N_20822);
nor U21475 (N_21475,N_20877,N_20813);
nand U21476 (N_21476,N_20781,N_20853);
and U21477 (N_21477,N_20809,N_20907);
nand U21478 (N_21478,N_20779,N_20776);
or U21479 (N_21479,N_20576,N_20759);
and U21480 (N_21480,N_20788,N_20602);
or U21481 (N_21481,N_20866,N_20676);
nor U21482 (N_21482,N_20845,N_20834);
or U21483 (N_21483,N_20752,N_20791);
and U21484 (N_21484,N_20723,N_20551);
xor U21485 (N_21485,N_20783,N_20610);
or U21486 (N_21486,N_20609,N_20859);
xor U21487 (N_21487,N_20896,N_20724);
nand U21488 (N_21488,N_20568,N_20835);
or U21489 (N_21489,N_20825,N_20928);
xor U21490 (N_21490,N_20751,N_20626);
xor U21491 (N_21491,N_20724,N_20539);
nor U21492 (N_21492,N_20514,N_20710);
and U21493 (N_21493,N_20698,N_20574);
xor U21494 (N_21494,N_20681,N_20785);
or U21495 (N_21495,N_20583,N_20590);
xor U21496 (N_21496,N_20938,N_20647);
nand U21497 (N_21497,N_20959,N_20905);
xor U21498 (N_21498,N_20693,N_20929);
nand U21499 (N_21499,N_20744,N_20545);
xnor U21500 (N_21500,N_21108,N_21272);
and U21501 (N_21501,N_21298,N_21173);
xor U21502 (N_21502,N_21433,N_21090);
or U21503 (N_21503,N_21266,N_21089);
or U21504 (N_21504,N_21444,N_21439);
xor U21505 (N_21505,N_21037,N_21149);
nor U21506 (N_21506,N_21084,N_21366);
and U21507 (N_21507,N_21303,N_21146);
and U21508 (N_21508,N_21152,N_21115);
nor U21509 (N_21509,N_21411,N_21092);
nor U21510 (N_21510,N_21406,N_21436);
or U21511 (N_21511,N_21123,N_21224);
nor U21512 (N_21512,N_21301,N_21496);
xor U21513 (N_21513,N_21273,N_21395);
nor U21514 (N_21514,N_21056,N_21417);
nand U21515 (N_21515,N_21154,N_21157);
nand U21516 (N_21516,N_21486,N_21355);
and U21517 (N_21517,N_21040,N_21275);
and U21518 (N_21518,N_21315,N_21128);
or U21519 (N_21519,N_21357,N_21286);
nor U21520 (N_21520,N_21344,N_21263);
nor U21521 (N_21521,N_21317,N_21445);
xnor U21522 (N_21522,N_21179,N_21426);
nor U21523 (N_21523,N_21093,N_21454);
nor U21524 (N_21524,N_21342,N_21235);
or U21525 (N_21525,N_21484,N_21251);
or U21526 (N_21526,N_21432,N_21180);
nor U21527 (N_21527,N_21213,N_21494);
nor U21528 (N_21528,N_21393,N_21211);
nor U21529 (N_21529,N_21204,N_21374);
and U21530 (N_21530,N_21060,N_21316);
nor U21531 (N_21531,N_21457,N_21214);
and U21532 (N_21532,N_21421,N_21038);
xor U21533 (N_21533,N_21404,N_21088);
or U21534 (N_21534,N_21323,N_21320);
and U21535 (N_21535,N_21247,N_21049);
or U21536 (N_21536,N_21425,N_21442);
or U21537 (N_21537,N_21377,N_21122);
or U21538 (N_21538,N_21493,N_21289);
nor U21539 (N_21539,N_21368,N_21424);
nand U21540 (N_21540,N_21350,N_21232);
nor U21541 (N_21541,N_21171,N_21267);
nand U21542 (N_21542,N_21447,N_21130);
and U21543 (N_21543,N_21483,N_21324);
or U21544 (N_21544,N_21462,N_21032);
nand U21545 (N_21545,N_21262,N_21162);
or U21546 (N_21546,N_21065,N_21113);
nor U21547 (N_21547,N_21443,N_21140);
nand U21548 (N_21548,N_21375,N_21459);
xor U21549 (N_21549,N_21003,N_21437);
nand U21550 (N_21550,N_21481,N_21230);
and U21551 (N_21551,N_21020,N_21446);
or U21552 (N_21552,N_21326,N_21043);
nand U21553 (N_21553,N_21177,N_21278);
or U21554 (N_21554,N_21014,N_21270);
xnor U21555 (N_21555,N_21402,N_21420);
xor U21556 (N_21556,N_21098,N_21384);
nand U21557 (N_21557,N_21063,N_21004);
and U21558 (N_21558,N_21358,N_21238);
xor U21559 (N_21559,N_21467,N_21222);
xnor U21560 (N_21560,N_21452,N_21047);
xor U21561 (N_21561,N_21422,N_21250);
or U21562 (N_21562,N_21290,N_21260);
xor U21563 (N_21563,N_21490,N_21009);
or U21564 (N_21564,N_21135,N_21382);
or U21565 (N_21565,N_21429,N_21259);
nand U21566 (N_21566,N_21480,N_21245);
nor U21567 (N_21567,N_21472,N_21095);
or U21568 (N_21568,N_21455,N_21195);
nand U21569 (N_21569,N_21000,N_21418);
and U21570 (N_21570,N_21376,N_21293);
or U21571 (N_21571,N_21348,N_21151);
or U21572 (N_21572,N_21170,N_21174);
nor U21573 (N_21573,N_21138,N_21110);
or U21574 (N_21574,N_21282,N_21142);
xnor U21575 (N_21575,N_21302,N_21160);
nor U21576 (N_21576,N_21210,N_21136);
and U21577 (N_21577,N_21497,N_21491);
nand U21578 (N_21578,N_21226,N_21386);
or U21579 (N_21579,N_21062,N_21070);
xor U21580 (N_21580,N_21075,N_21061);
or U21581 (N_21581,N_21013,N_21184);
xnor U21582 (N_21582,N_21137,N_21244);
nor U21583 (N_21583,N_21042,N_21082);
xnor U21584 (N_21584,N_21117,N_21304);
nor U21585 (N_21585,N_21073,N_21161);
xor U21586 (N_21586,N_21207,N_21069);
nand U21587 (N_21587,N_21345,N_21456);
xnor U21588 (N_21588,N_21059,N_21362);
nor U21589 (N_21589,N_21391,N_21008);
nor U21590 (N_21590,N_21478,N_21019);
xnor U21591 (N_21591,N_21125,N_21430);
or U21592 (N_21592,N_21387,N_21223);
nand U21593 (N_21593,N_21237,N_21068);
and U21594 (N_21594,N_21005,N_21066);
xnor U21595 (N_21595,N_21373,N_21033);
nand U21596 (N_21596,N_21091,N_21450);
nor U21597 (N_21597,N_21365,N_21434);
nand U21598 (N_21598,N_21072,N_21340);
and U21599 (N_21599,N_21380,N_21129);
nor U21600 (N_21600,N_21141,N_21264);
nor U21601 (N_21601,N_21339,N_21305);
nand U21602 (N_21602,N_21488,N_21354);
and U21603 (N_21603,N_21175,N_21280);
nor U21604 (N_21604,N_21181,N_21319);
nor U21605 (N_21605,N_21217,N_21194);
nor U21606 (N_21606,N_21103,N_21283);
xnor U21607 (N_21607,N_21246,N_21333);
and U21608 (N_21608,N_21415,N_21026);
nand U21609 (N_21609,N_21461,N_21131);
and U21610 (N_21610,N_21347,N_21118);
or U21611 (N_21611,N_21215,N_21101);
or U21612 (N_21612,N_21423,N_21294);
and U21613 (N_21613,N_21186,N_21416);
xnor U21614 (N_21614,N_21076,N_21458);
xnor U21615 (N_21615,N_21334,N_21035);
or U21616 (N_21616,N_21178,N_21067);
nand U21617 (N_21617,N_21189,N_21468);
and U21618 (N_21618,N_21268,N_21254);
xor U21619 (N_21619,N_21389,N_21364);
nand U21620 (N_21620,N_21288,N_21309);
nand U21621 (N_21621,N_21147,N_21405);
or U21622 (N_21622,N_21127,N_21241);
xor U21623 (N_21623,N_21202,N_21322);
or U21624 (N_21624,N_21407,N_21227);
or U21625 (N_21625,N_21205,N_21485);
and U21626 (N_21626,N_21169,N_21216);
and U21627 (N_21627,N_21102,N_21124);
xnor U21628 (N_21628,N_21109,N_21474);
or U21629 (N_21629,N_21440,N_21126);
or U21630 (N_21630,N_21080,N_21025);
nor U21631 (N_21631,N_21381,N_21475);
nand U21632 (N_21632,N_21401,N_21460);
and U21633 (N_21633,N_21281,N_21312);
nand U21634 (N_21634,N_21242,N_21164);
xor U21635 (N_21635,N_21018,N_21428);
xor U21636 (N_21636,N_21153,N_21306);
and U21637 (N_21637,N_21209,N_21248);
or U21638 (N_21638,N_21097,N_21336);
or U21639 (N_21639,N_21412,N_21297);
or U21640 (N_21640,N_21370,N_21258);
xor U21641 (N_21641,N_21015,N_21240);
xnor U21642 (N_21642,N_21074,N_21337);
and U21643 (N_21643,N_21252,N_21006);
nand U21644 (N_21644,N_21220,N_21408);
nor U21645 (N_21645,N_21200,N_21197);
nor U21646 (N_21646,N_21145,N_21051);
nand U21647 (N_21647,N_21291,N_21203);
nor U21648 (N_21648,N_21168,N_21016);
xnor U21649 (N_21649,N_21010,N_21166);
and U21650 (N_21650,N_21012,N_21045);
xnor U21651 (N_21651,N_21031,N_21172);
or U21652 (N_21652,N_21193,N_21464);
xor U21653 (N_21653,N_21218,N_21495);
xnor U21654 (N_21654,N_21311,N_21292);
and U21655 (N_21655,N_21330,N_21431);
nor U21656 (N_21656,N_21071,N_21188);
or U21657 (N_21657,N_21233,N_21192);
xor U21658 (N_21658,N_21024,N_21121);
or U21659 (N_21659,N_21228,N_21078);
nand U21660 (N_21660,N_21451,N_21116);
or U21661 (N_21661,N_21176,N_21329);
xor U21662 (N_21662,N_21287,N_21034);
nor U21663 (N_21663,N_21327,N_21236);
xor U21664 (N_21664,N_21212,N_21079);
nor U21665 (N_21665,N_21285,N_21284);
xnor U21666 (N_21666,N_21119,N_21346);
or U21667 (N_21667,N_21053,N_21441);
nor U21668 (N_21668,N_21325,N_21397);
xor U21669 (N_21669,N_21021,N_21077);
xor U21670 (N_21670,N_21199,N_21054);
nor U21671 (N_21671,N_21338,N_21271);
nand U21672 (N_21672,N_21165,N_21399);
nand U21673 (N_21673,N_21473,N_21349);
nand U21674 (N_21674,N_21229,N_21388);
or U21675 (N_21675,N_21208,N_21096);
or U21676 (N_21676,N_21114,N_21487);
or U21677 (N_21677,N_21265,N_21328);
nand U21678 (N_21678,N_21100,N_21331);
xor U21679 (N_21679,N_21057,N_21277);
nor U21680 (N_21680,N_21107,N_21296);
or U21681 (N_21681,N_21148,N_21086);
xnor U21682 (N_21682,N_21300,N_21219);
or U21683 (N_21683,N_21150,N_21064);
and U21684 (N_21684,N_21378,N_21087);
and U21685 (N_21685,N_21307,N_21085);
nand U21686 (N_21686,N_21036,N_21023);
and U21687 (N_21687,N_21134,N_21321);
or U21688 (N_21688,N_21352,N_21427);
nor U21689 (N_21689,N_21359,N_21372);
and U21690 (N_21690,N_21081,N_21196);
or U21691 (N_21691,N_21027,N_21133);
and U21692 (N_21692,N_21022,N_21167);
and U21693 (N_21693,N_21234,N_21239);
nor U21694 (N_21694,N_21453,N_21435);
nor U21695 (N_21695,N_21198,N_21041);
nor U21696 (N_21696,N_21385,N_21028);
or U21697 (N_21697,N_21449,N_21231);
and U21698 (N_21698,N_21055,N_21030);
or U21699 (N_21699,N_21191,N_21403);
nor U21700 (N_21700,N_21466,N_21111);
xnor U21701 (N_21701,N_21225,N_21185);
nand U21702 (N_21702,N_21144,N_21469);
nand U21703 (N_21703,N_21398,N_21463);
or U21704 (N_21704,N_21253,N_21257);
and U21705 (N_21705,N_21360,N_21269);
nor U21706 (N_21706,N_21361,N_21308);
xor U21707 (N_21707,N_21390,N_21477);
nand U21708 (N_21708,N_21139,N_21314);
and U21709 (N_21709,N_21353,N_21044);
nand U21710 (N_21710,N_21310,N_21470);
and U21711 (N_21711,N_21120,N_21499);
nand U21712 (N_21712,N_21356,N_21295);
xnor U21713 (N_21713,N_21313,N_21201);
or U21714 (N_21714,N_21143,N_21221);
or U21715 (N_21715,N_21371,N_21112);
xor U21716 (N_21716,N_21029,N_21039);
xnor U21717 (N_21717,N_21052,N_21190);
nand U21718 (N_21718,N_21187,N_21335);
and U21719 (N_21719,N_21448,N_21438);
and U21720 (N_21720,N_21094,N_21394);
nand U21721 (N_21721,N_21396,N_21471);
and U21722 (N_21722,N_21383,N_21255);
nor U21723 (N_21723,N_21479,N_21104);
xor U21724 (N_21724,N_21007,N_21206);
or U21725 (N_21725,N_21050,N_21332);
or U21726 (N_21726,N_21476,N_21243);
nand U21727 (N_21727,N_21099,N_21155);
and U21728 (N_21728,N_21279,N_21498);
or U21729 (N_21729,N_21156,N_21410);
or U21730 (N_21730,N_21409,N_21489);
or U21731 (N_21731,N_21318,N_21106);
or U21732 (N_21732,N_21011,N_21158);
and U21733 (N_21733,N_21256,N_21341);
nand U21734 (N_21734,N_21363,N_21392);
xnor U21735 (N_21735,N_21017,N_21058);
xor U21736 (N_21736,N_21343,N_21369);
xnor U21737 (N_21737,N_21400,N_21182);
or U21738 (N_21738,N_21163,N_21183);
nor U21739 (N_21739,N_21001,N_21414);
nand U21740 (N_21740,N_21492,N_21002);
or U21741 (N_21741,N_21482,N_21261);
nand U21742 (N_21742,N_21299,N_21413);
or U21743 (N_21743,N_21465,N_21132);
xor U21744 (N_21744,N_21367,N_21159);
nor U21745 (N_21745,N_21083,N_21419);
nor U21746 (N_21746,N_21048,N_21046);
or U21747 (N_21747,N_21274,N_21379);
and U21748 (N_21748,N_21276,N_21249);
nor U21749 (N_21749,N_21351,N_21105);
or U21750 (N_21750,N_21210,N_21402);
xor U21751 (N_21751,N_21411,N_21323);
xor U21752 (N_21752,N_21422,N_21107);
nor U21753 (N_21753,N_21392,N_21497);
xnor U21754 (N_21754,N_21382,N_21242);
nor U21755 (N_21755,N_21121,N_21219);
and U21756 (N_21756,N_21291,N_21425);
and U21757 (N_21757,N_21145,N_21041);
xnor U21758 (N_21758,N_21148,N_21260);
nor U21759 (N_21759,N_21409,N_21080);
and U21760 (N_21760,N_21173,N_21308);
or U21761 (N_21761,N_21071,N_21110);
and U21762 (N_21762,N_21246,N_21025);
xor U21763 (N_21763,N_21256,N_21348);
nand U21764 (N_21764,N_21385,N_21354);
or U21765 (N_21765,N_21406,N_21056);
and U21766 (N_21766,N_21043,N_21018);
xnor U21767 (N_21767,N_21305,N_21216);
and U21768 (N_21768,N_21400,N_21486);
and U21769 (N_21769,N_21381,N_21184);
xor U21770 (N_21770,N_21498,N_21251);
nor U21771 (N_21771,N_21374,N_21354);
and U21772 (N_21772,N_21062,N_21144);
and U21773 (N_21773,N_21469,N_21114);
nor U21774 (N_21774,N_21245,N_21361);
nand U21775 (N_21775,N_21001,N_21411);
and U21776 (N_21776,N_21462,N_21409);
and U21777 (N_21777,N_21072,N_21474);
and U21778 (N_21778,N_21391,N_21064);
or U21779 (N_21779,N_21067,N_21025);
xor U21780 (N_21780,N_21100,N_21480);
nand U21781 (N_21781,N_21143,N_21456);
and U21782 (N_21782,N_21436,N_21003);
and U21783 (N_21783,N_21020,N_21443);
nand U21784 (N_21784,N_21223,N_21108);
nor U21785 (N_21785,N_21491,N_21097);
nor U21786 (N_21786,N_21084,N_21121);
nor U21787 (N_21787,N_21431,N_21397);
and U21788 (N_21788,N_21333,N_21426);
or U21789 (N_21789,N_21279,N_21363);
nand U21790 (N_21790,N_21398,N_21154);
and U21791 (N_21791,N_21302,N_21321);
and U21792 (N_21792,N_21491,N_21365);
nand U21793 (N_21793,N_21000,N_21496);
nand U21794 (N_21794,N_21480,N_21411);
and U21795 (N_21795,N_21120,N_21447);
xor U21796 (N_21796,N_21489,N_21335);
xor U21797 (N_21797,N_21462,N_21277);
nand U21798 (N_21798,N_21044,N_21050);
or U21799 (N_21799,N_21257,N_21268);
xnor U21800 (N_21800,N_21401,N_21011);
and U21801 (N_21801,N_21475,N_21316);
and U21802 (N_21802,N_21209,N_21425);
xor U21803 (N_21803,N_21418,N_21068);
nand U21804 (N_21804,N_21395,N_21303);
nor U21805 (N_21805,N_21295,N_21400);
nor U21806 (N_21806,N_21444,N_21036);
nor U21807 (N_21807,N_21019,N_21094);
nor U21808 (N_21808,N_21469,N_21409);
nor U21809 (N_21809,N_21350,N_21026);
nor U21810 (N_21810,N_21467,N_21359);
nor U21811 (N_21811,N_21216,N_21084);
and U21812 (N_21812,N_21259,N_21324);
xnor U21813 (N_21813,N_21396,N_21429);
or U21814 (N_21814,N_21295,N_21147);
nand U21815 (N_21815,N_21130,N_21321);
nor U21816 (N_21816,N_21444,N_21162);
or U21817 (N_21817,N_21187,N_21022);
nand U21818 (N_21818,N_21486,N_21431);
or U21819 (N_21819,N_21105,N_21070);
or U21820 (N_21820,N_21302,N_21233);
nand U21821 (N_21821,N_21459,N_21486);
xor U21822 (N_21822,N_21009,N_21203);
or U21823 (N_21823,N_21198,N_21026);
nand U21824 (N_21824,N_21362,N_21067);
and U21825 (N_21825,N_21223,N_21107);
nor U21826 (N_21826,N_21048,N_21363);
and U21827 (N_21827,N_21404,N_21021);
xor U21828 (N_21828,N_21113,N_21457);
and U21829 (N_21829,N_21407,N_21133);
and U21830 (N_21830,N_21028,N_21052);
and U21831 (N_21831,N_21468,N_21203);
xor U21832 (N_21832,N_21007,N_21273);
nand U21833 (N_21833,N_21002,N_21471);
nand U21834 (N_21834,N_21112,N_21026);
xor U21835 (N_21835,N_21208,N_21265);
xor U21836 (N_21836,N_21237,N_21018);
nor U21837 (N_21837,N_21096,N_21424);
or U21838 (N_21838,N_21092,N_21098);
xnor U21839 (N_21839,N_21181,N_21112);
and U21840 (N_21840,N_21248,N_21018);
nor U21841 (N_21841,N_21317,N_21063);
and U21842 (N_21842,N_21192,N_21490);
and U21843 (N_21843,N_21163,N_21458);
and U21844 (N_21844,N_21354,N_21048);
or U21845 (N_21845,N_21152,N_21496);
and U21846 (N_21846,N_21110,N_21155);
or U21847 (N_21847,N_21374,N_21255);
or U21848 (N_21848,N_21150,N_21252);
nand U21849 (N_21849,N_21030,N_21051);
xnor U21850 (N_21850,N_21161,N_21224);
xnor U21851 (N_21851,N_21052,N_21035);
nor U21852 (N_21852,N_21002,N_21284);
nand U21853 (N_21853,N_21076,N_21277);
or U21854 (N_21854,N_21191,N_21284);
and U21855 (N_21855,N_21003,N_21087);
xor U21856 (N_21856,N_21413,N_21111);
or U21857 (N_21857,N_21198,N_21221);
nor U21858 (N_21858,N_21393,N_21022);
xor U21859 (N_21859,N_21440,N_21128);
and U21860 (N_21860,N_21215,N_21125);
xnor U21861 (N_21861,N_21164,N_21262);
nor U21862 (N_21862,N_21494,N_21426);
nor U21863 (N_21863,N_21470,N_21087);
xnor U21864 (N_21864,N_21405,N_21053);
and U21865 (N_21865,N_21211,N_21134);
nand U21866 (N_21866,N_21158,N_21076);
nand U21867 (N_21867,N_21120,N_21085);
nor U21868 (N_21868,N_21497,N_21039);
nand U21869 (N_21869,N_21238,N_21081);
xor U21870 (N_21870,N_21329,N_21132);
or U21871 (N_21871,N_21349,N_21273);
and U21872 (N_21872,N_21294,N_21476);
xor U21873 (N_21873,N_21390,N_21440);
nor U21874 (N_21874,N_21447,N_21154);
or U21875 (N_21875,N_21145,N_21396);
nand U21876 (N_21876,N_21400,N_21056);
nor U21877 (N_21877,N_21065,N_21023);
or U21878 (N_21878,N_21461,N_21074);
nand U21879 (N_21879,N_21187,N_21240);
nand U21880 (N_21880,N_21161,N_21014);
or U21881 (N_21881,N_21290,N_21156);
nor U21882 (N_21882,N_21095,N_21202);
nand U21883 (N_21883,N_21473,N_21229);
or U21884 (N_21884,N_21363,N_21188);
and U21885 (N_21885,N_21269,N_21172);
xor U21886 (N_21886,N_21296,N_21468);
nor U21887 (N_21887,N_21379,N_21001);
nor U21888 (N_21888,N_21442,N_21455);
nand U21889 (N_21889,N_21113,N_21237);
xnor U21890 (N_21890,N_21298,N_21308);
xnor U21891 (N_21891,N_21428,N_21188);
nand U21892 (N_21892,N_21017,N_21034);
and U21893 (N_21893,N_21453,N_21412);
and U21894 (N_21894,N_21025,N_21112);
and U21895 (N_21895,N_21264,N_21193);
xor U21896 (N_21896,N_21160,N_21303);
and U21897 (N_21897,N_21024,N_21083);
nor U21898 (N_21898,N_21103,N_21126);
nor U21899 (N_21899,N_21265,N_21246);
nor U21900 (N_21900,N_21245,N_21094);
or U21901 (N_21901,N_21465,N_21022);
xnor U21902 (N_21902,N_21386,N_21445);
nand U21903 (N_21903,N_21079,N_21340);
or U21904 (N_21904,N_21291,N_21485);
and U21905 (N_21905,N_21233,N_21414);
nand U21906 (N_21906,N_21055,N_21435);
and U21907 (N_21907,N_21124,N_21293);
nor U21908 (N_21908,N_21309,N_21013);
nand U21909 (N_21909,N_21183,N_21392);
and U21910 (N_21910,N_21229,N_21025);
nor U21911 (N_21911,N_21452,N_21167);
nor U21912 (N_21912,N_21069,N_21087);
nor U21913 (N_21913,N_21130,N_21262);
or U21914 (N_21914,N_21471,N_21120);
nand U21915 (N_21915,N_21078,N_21031);
xnor U21916 (N_21916,N_21350,N_21482);
and U21917 (N_21917,N_21160,N_21158);
xnor U21918 (N_21918,N_21202,N_21464);
nor U21919 (N_21919,N_21160,N_21455);
or U21920 (N_21920,N_21480,N_21414);
and U21921 (N_21921,N_21094,N_21434);
xnor U21922 (N_21922,N_21183,N_21065);
nor U21923 (N_21923,N_21333,N_21342);
nor U21924 (N_21924,N_21326,N_21461);
or U21925 (N_21925,N_21400,N_21497);
nand U21926 (N_21926,N_21055,N_21152);
or U21927 (N_21927,N_21349,N_21034);
and U21928 (N_21928,N_21103,N_21181);
nand U21929 (N_21929,N_21003,N_21036);
or U21930 (N_21930,N_21194,N_21458);
nor U21931 (N_21931,N_21329,N_21277);
nor U21932 (N_21932,N_21156,N_21486);
nor U21933 (N_21933,N_21027,N_21158);
or U21934 (N_21934,N_21259,N_21490);
xor U21935 (N_21935,N_21423,N_21166);
nand U21936 (N_21936,N_21168,N_21410);
nand U21937 (N_21937,N_21396,N_21359);
or U21938 (N_21938,N_21346,N_21274);
and U21939 (N_21939,N_21438,N_21372);
and U21940 (N_21940,N_21153,N_21146);
nor U21941 (N_21941,N_21025,N_21045);
and U21942 (N_21942,N_21039,N_21427);
and U21943 (N_21943,N_21497,N_21184);
or U21944 (N_21944,N_21294,N_21358);
and U21945 (N_21945,N_21224,N_21454);
nor U21946 (N_21946,N_21208,N_21261);
nor U21947 (N_21947,N_21137,N_21117);
or U21948 (N_21948,N_21024,N_21050);
and U21949 (N_21949,N_21407,N_21435);
nor U21950 (N_21950,N_21007,N_21243);
nor U21951 (N_21951,N_21349,N_21082);
nor U21952 (N_21952,N_21086,N_21179);
nor U21953 (N_21953,N_21483,N_21004);
and U21954 (N_21954,N_21414,N_21344);
xor U21955 (N_21955,N_21363,N_21059);
xnor U21956 (N_21956,N_21290,N_21119);
nor U21957 (N_21957,N_21223,N_21004);
and U21958 (N_21958,N_21186,N_21038);
nand U21959 (N_21959,N_21323,N_21449);
nor U21960 (N_21960,N_21127,N_21485);
and U21961 (N_21961,N_21400,N_21383);
nand U21962 (N_21962,N_21283,N_21133);
nand U21963 (N_21963,N_21023,N_21188);
nor U21964 (N_21964,N_21092,N_21350);
and U21965 (N_21965,N_21205,N_21302);
nand U21966 (N_21966,N_21249,N_21479);
xor U21967 (N_21967,N_21162,N_21384);
and U21968 (N_21968,N_21282,N_21130);
xnor U21969 (N_21969,N_21215,N_21288);
and U21970 (N_21970,N_21038,N_21341);
nand U21971 (N_21971,N_21422,N_21301);
xor U21972 (N_21972,N_21228,N_21248);
xor U21973 (N_21973,N_21283,N_21343);
nor U21974 (N_21974,N_21377,N_21084);
nand U21975 (N_21975,N_21308,N_21056);
nor U21976 (N_21976,N_21373,N_21345);
nand U21977 (N_21977,N_21270,N_21363);
nand U21978 (N_21978,N_21237,N_21053);
xnor U21979 (N_21979,N_21397,N_21267);
or U21980 (N_21980,N_21266,N_21466);
xor U21981 (N_21981,N_21326,N_21464);
and U21982 (N_21982,N_21043,N_21123);
xnor U21983 (N_21983,N_21276,N_21180);
and U21984 (N_21984,N_21188,N_21411);
and U21985 (N_21985,N_21453,N_21177);
nand U21986 (N_21986,N_21459,N_21307);
or U21987 (N_21987,N_21075,N_21050);
or U21988 (N_21988,N_21133,N_21017);
nor U21989 (N_21989,N_21367,N_21176);
or U21990 (N_21990,N_21117,N_21209);
nand U21991 (N_21991,N_21460,N_21042);
xnor U21992 (N_21992,N_21364,N_21281);
xor U21993 (N_21993,N_21179,N_21048);
or U21994 (N_21994,N_21054,N_21015);
or U21995 (N_21995,N_21021,N_21033);
and U21996 (N_21996,N_21350,N_21332);
or U21997 (N_21997,N_21442,N_21265);
nand U21998 (N_21998,N_21074,N_21124);
xnor U21999 (N_21999,N_21193,N_21180);
nor U22000 (N_22000,N_21584,N_21919);
xnor U22001 (N_22001,N_21863,N_21599);
or U22002 (N_22002,N_21937,N_21893);
or U22003 (N_22003,N_21925,N_21676);
xor U22004 (N_22004,N_21918,N_21732);
xnor U22005 (N_22005,N_21885,N_21833);
and U22006 (N_22006,N_21727,N_21658);
xnor U22007 (N_22007,N_21894,N_21593);
xor U22008 (N_22008,N_21736,N_21502);
xnor U22009 (N_22009,N_21530,N_21694);
xor U22010 (N_22010,N_21668,N_21608);
nor U22011 (N_22011,N_21980,N_21793);
and U22012 (N_22012,N_21843,N_21892);
nand U22013 (N_22013,N_21982,N_21774);
xor U22014 (N_22014,N_21657,N_21590);
and U22015 (N_22015,N_21822,N_21619);
xnor U22016 (N_22016,N_21751,N_21746);
nand U22017 (N_22017,N_21926,N_21724);
or U22018 (N_22018,N_21591,N_21824);
nor U22019 (N_22019,N_21686,N_21795);
nor U22020 (N_22020,N_21614,N_21517);
nand U22021 (N_22021,N_21604,N_21773);
or U22022 (N_22022,N_21979,N_21531);
nand U22023 (N_22023,N_21511,N_21577);
xnor U22024 (N_22024,N_21884,N_21922);
xnor U22025 (N_22025,N_21681,N_21799);
xnor U22026 (N_22026,N_21905,N_21840);
and U22027 (N_22027,N_21698,N_21923);
and U22028 (N_22028,N_21647,N_21508);
nor U22029 (N_22029,N_21914,N_21632);
nand U22030 (N_22030,N_21940,N_21680);
nor U22031 (N_22031,N_21528,N_21756);
and U22032 (N_22032,N_21986,N_21592);
nand U22033 (N_22033,N_21717,N_21667);
nor U22034 (N_22034,N_21790,N_21711);
nor U22035 (N_22035,N_21660,N_21649);
and U22036 (N_22036,N_21930,N_21935);
xnor U22037 (N_22037,N_21804,N_21639);
xor U22038 (N_22038,N_21520,N_21612);
and U22039 (N_22039,N_21920,N_21771);
and U22040 (N_22040,N_21693,N_21769);
or U22041 (N_22041,N_21755,N_21503);
nor U22042 (N_22042,N_21526,N_21626);
nor U22043 (N_22043,N_21998,N_21844);
xor U22044 (N_22044,N_21868,N_21820);
and U22045 (N_22045,N_21789,N_21785);
nor U22046 (N_22046,N_21749,N_21507);
nor U22047 (N_22047,N_21596,N_21996);
xnor U22048 (N_22048,N_21527,N_21514);
and U22049 (N_22049,N_21725,N_21877);
nand U22050 (N_22050,N_21805,N_21541);
nor U22051 (N_22051,N_21617,N_21906);
or U22052 (N_22052,N_21949,N_21703);
xnor U22053 (N_22053,N_21775,N_21858);
nor U22054 (N_22054,N_21889,N_21762);
nor U22055 (N_22055,N_21791,N_21794);
or U22056 (N_22056,N_21948,N_21651);
xor U22057 (N_22057,N_21722,N_21838);
and U22058 (N_22058,N_21829,N_21974);
and U22059 (N_22059,N_21874,N_21888);
xnor U22060 (N_22060,N_21553,N_21609);
nor U22061 (N_22061,N_21802,N_21635);
and U22062 (N_22062,N_21701,N_21772);
nor U22063 (N_22063,N_21588,N_21916);
and U22064 (N_22064,N_21733,N_21610);
xnor U22065 (N_22065,N_21509,N_21897);
nand U22066 (N_22066,N_21947,N_21666);
xnor U22067 (N_22067,N_21677,N_21830);
xor U22068 (N_22068,N_21927,N_21763);
nor U22069 (N_22069,N_21623,N_21636);
xnor U22070 (N_22070,N_21821,N_21960);
nand U22071 (N_22071,N_21961,N_21903);
and U22072 (N_22072,N_21778,N_21784);
or U22073 (N_22073,N_21534,N_21955);
and U22074 (N_22074,N_21696,N_21574);
nor U22075 (N_22075,N_21896,N_21533);
xor U22076 (N_22076,N_21861,N_21987);
and U22077 (N_22077,N_21572,N_21538);
xor U22078 (N_22078,N_21836,N_21796);
or U22079 (N_22079,N_21522,N_21738);
or U22080 (N_22080,N_21631,N_21846);
or U22081 (N_22081,N_21928,N_21643);
nand U22082 (N_22082,N_21862,N_21656);
and U22083 (N_22083,N_21690,N_21662);
or U22084 (N_22084,N_21652,N_21962);
and U22085 (N_22085,N_21924,N_21835);
and U22086 (N_22086,N_21929,N_21723);
or U22087 (N_22087,N_21899,N_21606);
nor U22088 (N_22088,N_21568,N_21559);
xor U22089 (N_22089,N_21752,N_21873);
or U22090 (N_22090,N_21505,N_21860);
or U22091 (N_22091,N_21827,N_21529);
or U22092 (N_22092,N_21523,N_21841);
nor U22093 (N_22093,N_21707,N_21670);
xnor U22094 (N_22094,N_21566,N_21716);
xor U22095 (N_22095,N_21976,N_21547);
nor U22096 (N_22096,N_21910,N_21519);
xnor U22097 (N_22097,N_21544,N_21640);
or U22098 (N_22098,N_21957,N_21545);
nor U22099 (N_22099,N_21720,N_21787);
nor U22100 (N_22100,N_21999,N_21637);
and U22101 (N_22101,N_21811,N_21826);
nor U22102 (N_22102,N_21758,N_21602);
or U22103 (N_22103,N_21550,N_21539);
nand U22104 (N_22104,N_21628,N_21786);
nor U22105 (N_22105,N_21695,N_21882);
xor U22106 (N_22106,N_21579,N_21663);
nand U22107 (N_22107,N_21839,N_21818);
and U22108 (N_22108,N_21561,N_21779);
and U22109 (N_22109,N_21978,N_21869);
and U22110 (N_22110,N_21780,N_21699);
and U22111 (N_22111,N_21646,N_21513);
nand U22112 (N_22112,N_21819,N_21582);
nand U22113 (N_22113,N_21908,N_21712);
nor U22114 (N_22114,N_21714,N_21573);
and U22115 (N_22115,N_21560,N_21942);
nor U22116 (N_22116,N_21965,N_21985);
or U22117 (N_22117,N_21867,N_21558);
nor U22118 (N_22118,N_21600,N_21759);
or U22119 (N_22119,N_21767,N_21966);
nor U22120 (N_22120,N_21575,N_21806);
and U22121 (N_22121,N_21747,N_21870);
and U22122 (N_22122,N_21580,N_21971);
nor U22123 (N_22123,N_21831,N_21589);
nor U22124 (N_22124,N_21682,N_21587);
nor U22125 (N_22125,N_21941,N_21886);
or U22126 (N_22126,N_21809,N_21684);
xor U22127 (N_22127,N_21645,N_21782);
xnor U22128 (N_22128,N_21598,N_21689);
nor U22129 (N_22129,N_21546,N_21750);
xnor U22130 (N_22130,N_21683,N_21854);
nor U22131 (N_22131,N_21764,N_21653);
and U22132 (N_22132,N_21625,N_21969);
nand U22133 (N_22133,N_21567,N_21601);
nor U22134 (N_22134,N_21953,N_21613);
and U22135 (N_22135,N_21586,N_21810);
or U22136 (N_22136,N_21864,N_21944);
and U22137 (N_22137,N_21501,N_21945);
xnor U22138 (N_22138,N_21706,N_21968);
and U22139 (N_22139,N_21512,N_21972);
nor U22140 (N_22140,N_21876,N_21812);
xor U22141 (N_22141,N_21540,N_21963);
and U22142 (N_22142,N_21611,N_21907);
and U22143 (N_22143,N_21983,N_21880);
or U22144 (N_22144,N_21970,N_21524);
xnor U22145 (N_22145,N_21744,N_21605);
nor U22146 (N_22146,N_21902,N_21692);
nor U22147 (N_22147,N_21909,N_21865);
and U22148 (N_22148,N_21921,N_21548);
and U22149 (N_22149,N_21718,N_21837);
nor U22150 (N_22150,N_21768,N_21770);
xor U22151 (N_22151,N_21890,N_21622);
xor U22152 (N_22152,N_21741,N_21815);
nor U22153 (N_22153,N_21518,N_21557);
nand U22154 (N_22154,N_21765,N_21708);
xnor U22155 (N_22155,N_21964,N_21817);
nor U22156 (N_22156,N_21510,N_21912);
nand U22157 (N_22157,N_21845,N_21766);
xor U22158 (N_22158,N_21828,N_21532);
nor U22159 (N_22159,N_21788,N_21850);
xor U22160 (N_22160,N_21536,N_21737);
nor U22161 (N_22161,N_21571,N_21956);
and U22162 (N_22162,N_21989,N_21506);
nand U22163 (N_22163,N_21917,N_21627);
or U22164 (N_22164,N_21875,N_21549);
or U22165 (N_22165,N_21535,N_21616);
or U22166 (N_22166,N_21687,N_21847);
nor U22167 (N_22167,N_21891,N_21671);
nand U22168 (N_22168,N_21866,N_21853);
nand U22169 (N_22169,N_21642,N_21943);
or U22170 (N_22170,N_21995,N_21709);
nand U22171 (N_22171,N_21783,N_21654);
and U22172 (N_22172,N_21800,N_21742);
and U22173 (N_22173,N_21814,N_21797);
or U22174 (N_22174,N_21992,N_21915);
nand U22175 (N_22175,N_21842,N_21881);
nand U22176 (N_22176,N_21537,N_21556);
and U22177 (N_22177,N_21740,N_21621);
or U22178 (N_22178,N_21745,N_21898);
nor U22179 (N_22179,N_21807,N_21761);
and U22180 (N_22180,N_21624,N_21938);
nor U22181 (N_22181,N_21855,N_21515);
nand U22182 (N_22182,N_21792,N_21597);
nand U22183 (N_22183,N_21500,N_21583);
and U22184 (N_22184,N_21729,N_21721);
or U22185 (N_22185,N_21576,N_21641);
or U22186 (N_22186,N_21993,N_21551);
xor U22187 (N_22187,N_21715,N_21991);
and U22188 (N_22188,N_21959,N_21700);
and U22189 (N_22189,N_21521,N_21697);
nor U22190 (N_22190,N_21994,N_21585);
or U22191 (N_22191,N_21705,N_21674);
nor U22192 (N_22192,N_21638,N_21650);
nand U22193 (N_22193,N_21808,N_21618);
nor U22194 (N_22194,N_21859,N_21669);
nor U22195 (N_22195,N_21932,N_21883);
nor U22196 (N_22196,N_21629,N_21757);
or U22197 (N_22197,N_21603,N_21981);
or U22198 (N_22198,N_21973,N_21879);
and U22199 (N_22199,N_21634,N_21730);
or U22200 (N_22200,N_21954,N_21679);
or U22201 (N_22201,N_21849,N_21728);
nand U22202 (N_22202,N_21967,N_21748);
nor U22203 (N_22203,N_21871,N_21562);
xor U22204 (N_22204,N_21984,N_21803);
nand U22205 (N_22205,N_21911,N_21934);
nand U22206 (N_22206,N_21958,N_21901);
xor U22207 (N_22207,N_21713,N_21832);
and U22208 (N_22208,N_21595,N_21975);
and U22209 (N_22209,N_21813,N_21719);
nand U22210 (N_22210,N_21988,N_21977);
nor U22211 (N_22211,N_21939,N_21659);
nor U22212 (N_22212,N_21904,N_21542);
nand U22213 (N_22213,N_21691,N_21726);
nor U22214 (N_22214,N_21816,N_21798);
xor U22215 (N_22215,N_21936,N_21933);
xor U22216 (N_22216,N_21754,N_21664);
xnor U22217 (N_22217,N_21552,N_21554);
and U22218 (N_22218,N_21675,N_21688);
and U22219 (N_22219,N_21739,N_21872);
nand U22220 (N_22220,N_21633,N_21525);
or U22221 (N_22221,N_21900,N_21685);
or U22222 (N_22222,N_21852,N_21570);
and U22223 (N_22223,N_21777,N_21743);
nor U22224 (N_22224,N_21581,N_21857);
or U22225 (N_22225,N_21776,N_21878);
and U22226 (N_22226,N_21615,N_21825);
nand U22227 (N_22227,N_21563,N_21913);
nand U22228 (N_22228,N_21931,N_21672);
nor U22229 (N_22229,N_21555,N_21856);
nand U22230 (N_22230,N_21753,N_21951);
or U22231 (N_22231,N_21851,N_21997);
and U22232 (N_22232,N_21648,N_21665);
nand U22233 (N_22233,N_21702,N_21895);
and U22234 (N_22234,N_21731,N_21565);
or U22235 (N_22235,N_21655,N_21834);
xor U22236 (N_22236,N_21661,N_21848);
nor U22237 (N_22237,N_21620,N_21644);
xor U22238 (N_22238,N_21543,N_21678);
nor U22239 (N_22239,N_21569,N_21735);
and U22240 (N_22240,N_21704,N_21823);
nand U22241 (N_22241,N_21952,N_21630);
xor U22242 (N_22242,N_21950,N_21760);
nor U22243 (N_22243,N_21734,N_21781);
nor U22244 (N_22244,N_21710,N_21504);
or U22245 (N_22245,N_21516,N_21801);
or U22246 (N_22246,N_21578,N_21564);
or U22247 (N_22247,N_21990,N_21887);
and U22248 (N_22248,N_21594,N_21946);
xor U22249 (N_22249,N_21607,N_21673);
nand U22250 (N_22250,N_21728,N_21988);
or U22251 (N_22251,N_21948,N_21768);
nor U22252 (N_22252,N_21688,N_21538);
nand U22253 (N_22253,N_21788,N_21698);
nor U22254 (N_22254,N_21645,N_21585);
xnor U22255 (N_22255,N_21508,N_21701);
nand U22256 (N_22256,N_21681,N_21651);
nand U22257 (N_22257,N_21552,N_21522);
xnor U22258 (N_22258,N_21815,N_21535);
or U22259 (N_22259,N_21580,N_21783);
nor U22260 (N_22260,N_21829,N_21663);
nand U22261 (N_22261,N_21854,N_21588);
or U22262 (N_22262,N_21710,N_21835);
nor U22263 (N_22263,N_21976,N_21994);
xnor U22264 (N_22264,N_21935,N_21829);
and U22265 (N_22265,N_21546,N_21513);
or U22266 (N_22266,N_21822,N_21823);
nand U22267 (N_22267,N_21726,N_21628);
xor U22268 (N_22268,N_21778,N_21754);
or U22269 (N_22269,N_21677,N_21602);
xnor U22270 (N_22270,N_21831,N_21786);
xor U22271 (N_22271,N_21591,N_21848);
and U22272 (N_22272,N_21968,N_21924);
xnor U22273 (N_22273,N_21993,N_21774);
nand U22274 (N_22274,N_21959,N_21778);
nand U22275 (N_22275,N_21739,N_21692);
xor U22276 (N_22276,N_21509,N_21793);
xnor U22277 (N_22277,N_21858,N_21718);
or U22278 (N_22278,N_21524,N_21788);
nor U22279 (N_22279,N_21772,N_21502);
or U22280 (N_22280,N_21805,N_21716);
and U22281 (N_22281,N_21526,N_21659);
nor U22282 (N_22282,N_21755,N_21573);
and U22283 (N_22283,N_21835,N_21509);
nor U22284 (N_22284,N_21791,N_21760);
nor U22285 (N_22285,N_21616,N_21778);
nand U22286 (N_22286,N_21738,N_21619);
nor U22287 (N_22287,N_21588,N_21938);
or U22288 (N_22288,N_21591,N_21707);
or U22289 (N_22289,N_21810,N_21907);
and U22290 (N_22290,N_21757,N_21867);
nor U22291 (N_22291,N_21915,N_21733);
xnor U22292 (N_22292,N_21817,N_21563);
nor U22293 (N_22293,N_21539,N_21580);
nand U22294 (N_22294,N_21610,N_21557);
and U22295 (N_22295,N_21607,N_21897);
and U22296 (N_22296,N_21821,N_21674);
nor U22297 (N_22297,N_21740,N_21727);
nand U22298 (N_22298,N_21897,N_21648);
nor U22299 (N_22299,N_21819,N_21532);
xnor U22300 (N_22300,N_21960,N_21725);
nor U22301 (N_22301,N_21954,N_21649);
nand U22302 (N_22302,N_21508,N_21609);
or U22303 (N_22303,N_21966,N_21539);
or U22304 (N_22304,N_21807,N_21812);
nor U22305 (N_22305,N_21578,N_21705);
or U22306 (N_22306,N_21611,N_21711);
or U22307 (N_22307,N_21889,N_21550);
nor U22308 (N_22308,N_21761,N_21806);
and U22309 (N_22309,N_21979,N_21893);
nor U22310 (N_22310,N_21925,N_21602);
nor U22311 (N_22311,N_21856,N_21909);
and U22312 (N_22312,N_21529,N_21744);
nor U22313 (N_22313,N_21919,N_21903);
or U22314 (N_22314,N_21613,N_21783);
and U22315 (N_22315,N_21891,N_21876);
or U22316 (N_22316,N_21791,N_21920);
or U22317 (N_22317,N_21806,N_21649);
or U22318 (N_22318,N_21656,N_21684);
nor U22319 (N_22319,N_21528,N_21639);
nor U22320 (N_22320,N_21591,N_21985);
nand U22321 (N_22321,N_21596,N_21843);
nor U22322 (N_22322,N_21781,N_21677);
or U22323 (N_22323,N_21644,N_21647);
nand U22324 (N_22324,N_21910,N_21858);
nor U22325 (N_22325,N_21885,N_21566);
nand U22326 (N_22326,N_21982,N_21672);
nor U22327 (N_22327,N_21682,N_21917);
and U22328 (N_22328,N_21689,N_21926);
nor U22329 (N_22329,N_21542,N_21644);
nand U22330 (N_22330,N_21643,N_21582);
and U22331 (N_22331,N_21515,N_21926);
and U22332 (N_22332,N_21945,N_21519);
or U22333 (N_22333,N_21502,N_21767);
nor U22334 (N_22334,N_21515,N_21684);
nand U22335 (N_22335,N_21600,N_21799);
and U22336 (N_22336,N_21815,N_21708);
xnor U22337 (N_22337,N_21771,N_21969);
nand U22338 (N_22338,N_21990,N_21955);
and U22339 (N_22339,N_21925,N_21688);
xor U22340 (N_22340,N_21558,N_21703);
and U22341 (N_22341,N_21990,N_21547);
or U22342 (N_22342,N_21953,N_21806);
nor U22343 (N_22343,N_21745,N_21644);
and U22344 (N_22344,N_21916,N_21665);
or U22345 (N_22345,N_21707,N_21772);
and U22346 (N_22346,N_21947,N_21526);
and U22347 (N_22347,N_21621,N_21513);
nand U22348 (N_22348,N_21516,N_21832);
xnor U22349 (N_22349,N_21541,N_21942);
or U22350 (N_22350,N_21954,N_21601);
or U22351 (N_22351,N_21852,N_21541);
xnor U22352 (N_22352,N_21638,N_21834);
and U22353 (N_22353,N_21711,N_21915);
nor U22354 (N_22354,N_21720,N_21939);
xnor U22355 (N_22355,N_21834,N_21636);
xor U22356 (N_22356,N_21530,N_21662);
nor U22357 (N_22357,N_21986,N_21557);
xnor U22358 (N_22358,N_21943,N_21571);
nor U22359 (N_22359,N_21559,N_21515);
or U22360 (N_22360,N_21981,N_21970);
nor U22361 (N_22361,N_21659,N_21972);
nor U22362 (N_22362,N_21843,N_21538);
nor U22363 (N_22363,N_21999,N_21936);
nor U22364 (N_22364,N_21860,N_21953);
xor U22365 (N_22365,N_21634,N_21842);
and U22366 (N_22366,N_21806,N_21598);
nor U22367 (N_22367,N_21803,N_21778);
xnor U22368 (N_22368,N_21848,N_21714);
xor U22369 (N_22369,N_21703,N_21615);
xnor U22370 (N_22370,N_21984,N_21841);
or U22371 (N_22371,N_21799,N_21874);
or U22372 (N_22372,N_21736,N_21668);
and U22373 (N_22373,N_21832,N_21746);
or U22374 (N_22374,N_21747,N_21781);
or U22375 (N_22375,N_21984,N_21789);
and U22376 (N_22376,N_21586,N_21873);
and U22377 (N_22377,N_21821,N_21781);
xor U22378 (N_22378,N_21823,N_21712);
xnor U22379 (N_22379,N_21804,N_21815);
xnor U22380 (N_22380,N_21662,N_21890);
nor U22381 (N_22381,N_21965,N_21699);
nand U22382 (N_22382,N_21534,N_21599);
nand U22383 (N_22383,N_21703,N_21950);
xnor U22384 (N_22384,N_21889,N_21599);
or U22385 (N_22385,N_21871,N_21539);
xnor U22386 (N_22386,N_21946,N_21565);
nand U22387 (N_22387,N_21948,N_21567);
and U22388 (N_22388,N_21887,N_21614);
and U22389 (N_22389,N_21932,N_21699);
xor U22390 (N_22390,N_21698,N_21753);
nor U22391 (N_22391,N_21751,N_21591);
and U22392 (N_22392,N_21563,N_21713);
nor U22393 (N_22393,N_21867,N_21672);
xor U22394 (N_22394,N_21785,N_21935);
xnor U22395 (N_22395,N_21870,N_21804);
xnor U22396 (N_22396,N_21589,N_21871);
or U22397 (N_22397,N_21804,N_21822);
or U22398 (N_22398,N_21875,N_21945);
nor U22399 (N_22399,N_21592,N_21683);
xor U22400 (N_22400,N_21765,N_21795);
xnor U22401 (N_22401,N_21730,N_21549);
xnor U22402 (N_22402,N_21539,N_21501);
nand U22403 (N_22403,N_21585,N_21545);
nand U22404 (N_22404,N_21589,N_21982);
and U22405 (N_22405,N_21844,N_21906);
nor U22406 (N_22406,N_21922,N_21569);
and U22407 (N_22407,N_21789,N_21823);
and U22408 (N_22408,N_21684,N_21911);
and U22409 (N_22409,N_21582,N_21571);
nor U22410 (N_22410,N_21823,N_21634);
xnor U22411 (N_22411,N_21981,N_21690);
nor U22412 (N_22412,N_21567,N_21847);
or U22413 (N_22413,N_21983,N_21548);
nand U22414 (N_22414,N_21816,N_21832);
nand U22415 (N_22415,N_21924,N_21530);
or U22416 (N_22416,N_21829,N_21879);
nand U22417 (N_22417,N_21611,N_21875);
nor U22418 (N_22418,N_21950,N_21942);
nor U22419 (N_22419,N_21986,N_21587);
nand U22420 (N_22420,N_21890,N_21985);
or U22421 (N_22421,N_21520,N_21985);
and U22422 (N_22422,N_21661,N_21861);
nor U22423 (N_22423,N_21834,N_21584);
or U22424 (N_22424,N_21965,N_21941);
or U22425 (N_22425,N_21616,N_21587);
and U22426 (N_22426,N_21793,N_21847);
nor U22427 (N_22427,N_21590,N_21847);
nor U22428 (N_22428,N_21863,N_21699);
xor U22429 (N_22429,N_21828,N_21523);
nor U22430 (N_22430,N_21982,N_21566);
and U22431 (N_22431,N_21880,N_21676);
nand U22432 (N_22432,N_21783,N_21565);
nor U22433 (N_22433,N_21762,N_21872);
nand U22434 (N_22434,N_21739,N_21864);
and U22435 (N_22435,N_21767,N_21933);
and U22436 (N_22436,N_21933,N_21692);
or U22437 (N_22437,N_21659,N_21503);
nand U22438 (N_22438,N_21754,N_21523);
nand U22439 (N_22439,N_21741,N_21775);
xnor U22440 (N_22440,N_21965,N_21636);
or U22441 (N_22441,N_21536,N_21807);
nor U22442 (N_22442,N_21848,N_21853);
xor U22443 (N_22443,N_21676,N_21765);
or U22444 (N_22444,N_21955,N_21673);
nor U22445 (N_22445,N_21550,N_21954);
and U22446 (N_22446,N_21753,N_21945);
nor U22447 (N_22447,N_21660,N_21646);
nand U22448 (N_22448,N_21768,N_21886);
nand U22449 (N_22449,N_21663,N_21922);
or U22450 (N_22450,N_21898,N_21848);
xor U22451 (N_22451,N_21860,N_21801);
or U22452 (N_22452,N_21548,N_21815);
and U22453 (N_22453,N_21572,N_21589);
xnor U22454 (N_22454,N_21505,N_21686);
or U22455 (N_22455,N_21848,N_21956);
and U22456 (N_22456,N_21732,N_21538);
xor U22457 (N_22457,N_21654,N_21826);
and U22458 (N_22458,N_21960,N_21538);
xor U22459 (N_22459,N_21629,N_21861);
nand U22460 (N_22460,N_21672,N_21922);
or U22461 (N_22461,N_21697,N_21955);
nor U22462 (N_22462,N_21539,N_21729);
and U22463 (N_22463,N_21668,N_21622);
and U22464 (N_22464,N_21866,N_21702);
xnor U22465 (N_22465,N_21808,N_21779);
or U22466 (N_22466,N_21837,N_21889);
nor U22467 (N_22467,N_21943,N_21826);
or U22468 (N_22468,N_21561,N_21823);
and U22469 (N_22469,N_21548,N_21576);
nor U22470 (N_22470,N_21933,N_21894);
and U22471 (N_22471,N_21703,N_21855);
nor U22472 (N_22472,N_21638,N_21941);
and U22473 (N_22473,N_21949,N_21848);
or U22474 (N_22474,N_21908,N_21761);
or U22475 (N_22475,N_21577,N_21534);
and U22476 (N_22476,N_21682,N_21571);
xnor U22477 (N_22477,N_21787,N_21519);
and U22478 (N_22478,N_21593,N_21561);
xor U22479 (N_22479,N_21608,N_21989);
or U22480 (N_22480,N_21879,N_21552);
and U22481 (N_22481,N_21877,N_21554);
nor U22482 (N_22482,N_21704,N_21605);
nand U22483 (N_22483,N_21922,N_21845);
nand U22484 (N_22484,N_21738,N_21860);
xor U22485 (N_22485,N_21561,N_21600);
and U22486 (N_22486,N_21719,N_21685);
nor U22487 (N_22487,N_21944,N_21783);
xor U22488 (N_22488,N_21864,N_21991);
xor U22489 (N_22489,N_21729,N_21574);
nand U22490 (N_22490,N_21539,N_21597);
nor U22491 (N_22491,N_21760,N_21928);
xnor U22492 (N_22492,N_21949,N_21818);
and U22493 (N_22493,N_21761,N_21934);
xnor U22494 (N_22494,N_21596,N_21562);
nand U22495 (N_22495,N_21552,N_21732);
xor U22496 (N_22496,N_21575,N_21848);
xnor U22497 (N_22497,N_21748,N_21564);
or U22498 (N_22498,N_21996,N_21972);
or U22499 (N_22499,N_21776,N_21816);
nor U22500 (N_22500,N_22461,N_22116);
or U22501 (N_22501,N_22339,N_22201);
and U22502 (N_22502,N_22441,N_22053);
and U22503 (N_22503,N_22212,N_22071);
nand U22504 (N_22504,N_22475,N_22153);
or U22505 (N_22505,N_22350,N_22155);
xor U22506 (N_22506,N_22471,N_22296);
nor U22507 (N_22507,N_22323,N_22092);
and U22508 (N_22508,N_22374,N_22217);
nor U22509 (N_22509,N_22268,N_22266);
nand U22510 (N_22510,N_22105,N_22468);
nor U22511 (N_22511,N_22413,N_22177);
xor U22512 (N_22512,N_22451,N_22481);
nor U22513 (N_22513,N_22467,N_22143);
nand U22514 (N_22514,N_22332,N_22037);
xnor U22515 (N_22515,N_22160,N_22348);
xor U22516 (N_22516,N_22084,N_22173);
nor U22517 (N_22517,N_22402,N_22137);
nor U22518 (N_22518,N_22194,N_22474);
xnor U22519 (N_22519,N_22096,N_22134);
or U22520 (N_22520,N_22012,N_22295);
nand U22521 (N_22521,N_22292,N_22126);
and U22522 (N_22522,N_22305,N_22276);
nand U22523 (N_22523,N_22382,N_22139);
or U22524 (N_22524,N_22453,N_22404);
nand U22525 (N_22525,N_22010,N_22498);
and U22526 (N_22526,N_22219,N_22027);
nor U22527 (N_22527,N_22182,N_22338);
xor U22528 (N_22528,N_22324,N_22437);
nand U22529 (N_22529,N_22238,N_22473);
nand U22530 (N_22530,N_22313,N_22389);
xnor U22531 (N_22531,N_22193,N_22401);
or U22532 (N_22532,N_22470,N_22099);
or U22533 (N_22533,N_22163,N_22063);
nand U22534 (N_22534,N_22421,N_22030);
nor U22535 (N_22535,N_22328,N_22482);
nor U22536 (N_22536,N_22431,N_22432);
and U22537 (N_22537,N_22085,N_22000);
and U22538 (N_22538,N_22111,N_22156);
nand U22539 (N_22539,N_22397,N_22426);
nand U22540 (N_22540,N_22108,N_22357);
xor U22541 (N_22541,N_22480,N_22166);
xnor U22542 (N_22542,N_22388,N_22172);
xnor U22543 (N_22543,N_22428,N_22114);
or U22544 (N_22544,N_22079,N_22297);
and U22545 (N_22545,N_22078,N_22094);
xor U22546 (N_22546,N_22447,N_22039);
nand U22547 (N_22547,N_22393,N_22345);
and U22548 (N_22548,N_22244,N_22265);
nor U22549 (N_22549,N_22145,N_22044);
nor U22550 (N_22550,N_22020,N_22396);
xor U22551 (N_22551,N_22368,N_22170);
and U22552 (N_22552,N_22291,N_22277);
or U22553 (N_22553,N_22060,N_22236);
xnor U22554 (N_22554,N_22015,N_22007);
or U22555 (N_22555,N_22259,N_22331);
and U22556 (N_22556,N_22411,N_22255);
and U22557 (N_22557,N_22211,N_22215);
or U22558 (N_22558,N_22130,N_22086);
nor U22559 (N_22559,N_22135,N_22232);
or U22560 (N_22560,N_22463,N_22442);
and U22561 (N_22561,N_22142,N_22390);
nand U22562 (N_22562,N_22090,N_22290);
nor U22563 (N_22563,N_22425,N_22210);
nand U22564 (N_22564,N_22036,N_22147);
and U22565 (N_22565,N_22140,N_22380);
nor U22566 (N_22566,N_22377,N_22069);
and U22567 (N_22567,N_22486,N_22398);
xor U22568 (N_22568,N_22082,N_22479);
or U22569 (N_22569,N_22131,N_22409);
nor U22570 (N_22570,N_22253,N_22024);
and U22571 (N_22571,N_22077,N_22379);
nor U22572 (N_22572,N_22400,N_22408);
nand U22573 (N_22573,N_22146,N_22176);
nand U22574 (N_22574,N_22187,N_22344);
nor U22575 (N_22575,N_22410,N_22430);
and U22576 (N_22576,N_22033,N_22191);
xor U22577 (N_22577,N_22150,N_22218);
nand U22578 (N_22578,N_22394,N_22376);
or U22579 (N_22579,N_22361,N_22222);
xnor U22580 (N_22580,N_22325,N_22308);
and U22581 (N_22581,N_22301,N_22021);
xor U22582 (N_22582,N_22373,N_22165);
xnor U22583 (N_22583,N_22040,N_22275);
and U22584 (N_22584,N_22250,N_22050);
xnor U22585 (N_22585,N_22422,N_22417);
and U22586 (N_22586,N_22386,N_22449);
nor U22587 (N_22587,N_22127,N_22161);
xnor U22588 (N_22588,N_22423,N_22299);
or U22589 (N_22589,N_22102,N_22336);
or U22590 (N_22590,N_22285,N_22186);
nand U22591 (N_22591,N_22496,N_22042);
nand U22592 (N_22592,N_22066,N_22202);
or U22593 (N_22593,N_22452,N_22469);
nand U22594 (N_22594,N_22075,N_22100);
or U22595 (N_22595,N_22207,N_22310);
nand U22596 (N_22596,N_22028,N_22495);
or U22597 (N_22597,N_22013,N_22043);
and U22598 (N_22598,N_22104,N_22228);
and U22599 (N_22599,N_22263,N_22162);
nand U22600 (N_22600,N_22076,N_22444);
and U22601 (N_22601,N_22129,N_22472);
and U22602 (N_22602,N_22144,N_22184);
nor U22603 (N_22603,N_22216,N_22174);
xor U22604 (N_22604,N_22445,N_22089);
nand U22605 (N_22605,N_22334,N_22269);
nor U22606 (N_22606,N_22103,N_22242);
nor U22607 (N_22607,N_22226,N_22062);
and U22608 (N_22608,N_22483,N_22080);
and U22609 (N_22609,N_22347,N_22018);
nor U22610 (N_22610,N_22321,N_22351);
nor U22611 (N_22611,N_22113,N_22169);
nor U22612 (N_22612,N_22175,N_22004);
or U22613 (N_22613,N_22230,N_22017);
xor U22614 (N_22614,N_22298,N_22261);
nand U22615 (N_22615,N_22340,N_22061);
or U22616 (N_22616,N_22198,N_22258);
and U22617 (N_22617,N_22203,N_22485);
nor U22618 (N_22618,N_22048,N_22288);
and U22619 (N_22619,N_22128,N_22151);
nor U22620 (N_22620,N_22330,N_22183);
nand U22621 (N_22621,N_22136,N_22106);
or U22622 (N_22622,N_22234,N_22171);
nand U22623 (N_22623,N_22121,N_22456);
and U22624 (N_22624,N_22093,N_22287);
nor U22625 (N_22625,N_22178,N_22497);
nand U22626 (N_22626,N_22058,N_22337);
and U22627 (N_22627,N_22306,N_22249);
xor U22628 (N_22628,N_22309,N_22003);
nand U22629 (N_22629,N_22059,N_22322);
xnor U22630 (N_22630,N_22446,N_22035);
nor U22631 (N_22631,N_22001,N_22407);
and U22632 (N_22632,N_22110,N_22458);
nand U22633 (N_22633,N_22091,N_22318);
nand U22634 (N_22634,N_22192,N_22205);
nand U22635 (N_22635,N_22272,N_22164);
nand U22636 (N_22636,N_22117,N_22208);
nand U22637 (N_22637,N_22317,N_22493);
or U22638 (N_22638,N_22476,N_22025);
nor U22639 (N_22639,N_22327,N_22335);
nor U22640 (N_22640,N_22118,N_22439);
nand U22641 (N_22641,N_22056,N_22280);
and U22642 (N_22642,N_22148,N_22354);
or U22643 (N_22643,N_22264,N_22149);
nor U22644 (N_22644,N_22055,N_22267);
and U22645 (N_22645,N_22209,N_22074);
nand U22646 (N_22646,N_22316,N_22239);
and U22647 (N_22647,N_22381,N_22181);
nand U22648 (N_22648,N_22281,N_22366);
nor U22649 (N_22649,N_22022,N_22067);
xor U22650 (N_22650,N_22403,N_22477);
and U22651 (N_22651,N_22200,N_22180);
xnor U22652 (N_22652,N_22240,N_22254);
or U22653 (N_22653,N_22199,N_22141);
nand U22654 (N_22654,N_22154,N_22072);
nor U22655 (N_22655,N_22225,N_22274);
nor U22656 (N_22656,N_22349,N_22246);
nand U22657 (N_22657,N_22233,N_22123);
nand U22658 (N_22658,N_22326,N_22011);
xnor U22659 (N_22659,N_22045,N_22329);
nand U22660 (N_22660,N_22237,N_22358);
xor U22661 (N_22661,N_22286,N_22002);
or U22662 (N_22662,N_22168,N_22307);
nor U22663 (N_22663,N_22188,N_22457);
xnor U22664 (N_22664,N_22138,N_22365);
xor U22665 (N_22665,N_22360,N_22424);
or U22666 (N_22666,N_22070,N_22052);
nor U22667 (N_22667,N_22391,N_22418);
nor U22668 (N_22668,N_22443,N_22227);
and U22669 (N_22669,N_22492,N_22352);
xor U22670 (N_22670,N_22491,N_22383);
or U22671 (N_22671,N_22179,N_22252);
and U22672 (N_22672,N_22438,N_22248);
xor U22673 (N_22673,N_22189,N_22300);
nand U22674 (N_22674,N_22167,N_22235);
nor U22675 (N_22675,N_22204,N_22115);
nor U22676 (N_22676,N_22289,N_22311);
nand U22677 (N_22677,N_22448,N_22392);
nand U22678 (N_22678,N_22466,N_22385);
or U22679 (N_22679,N_22429,N_22120);
nor U22680 (N_22680,N_22098,N_22213);
xor U22681 (N_22681,N_22087,N_22245);
and U22682 (N_22682,N_22112,N_22319);
nor U22683 (N_22683,N_22455,N_22158);
xnor U22684 (N_22684,N_22460,N_22256);
or U22685 (N_22685,N_22315,N_22484);
xnor U22686 (N_22686,N_22465,N_22224);
or U22687 (N_22687,N_22023,N_22006);
and U22688 (N_22688,N_22157,N_22363);
xnor U22689 (N_22689,N_22341,N_22293);
or U22690 (N_22690,N_22419,N_22016);
nor U22691 (N_22691,N_22241,N_22333);
and U22692 (N_22692,N_22064,N_22278);
and U22693 (N_22693,N_22262,N_22353);
and U22694 (N_22694,N_22073,N_22251);
nand U22695 (N_22695,N_22247,N_22054);
or U22696 (N_22696,N_22185,N_22231);
xor U22697 (N_22697,N_22420,N_22372);
and U22698 (N_22698,N_22282,N_22370);
nand U22699 (N_22699,N_22260,N_22359);
nand U22700 (N_22700,N_22019,N_22223);
xnor U22701 (N_22701,N_22005,N_22279);
nor U22702 (N_22702,N_22195,N_22049);
and U22703 (N_22703,N_22435,N_22440);
or U22704 (N_22704,N_22302,N_22459);
nor U22705 (N_22705,N_22047,N_22462);
xor U22706 (N_22706,N_22436,N_22283);
or U22707 (N_22707,N_22412,N_22122);
nand U22708 (N_22708,N_22378,N_22229);
nor U22709 (N_22709,N_22273,N_22034);
nand U22710 (N_22710,N_22367,N_22499);
and U22711 (N_22711,N_22081,N_22101);
xnor U22712 (N_22712,N_22487,N_22009);
xnor U22713 (N_22713,N_22454,N_22364);
nand U22714 (N_22714,N_22008,N_22057);
xnor U22715 (N_22715,N_22119,N_22284);
nor U22716 (N_22716,N_22206,N_22387);
or U22717 (N_22717,N_22221,N_22220);
xor U22718 (N_22718,N_22029,N_22395);
or U22719 (N_22719,N_22405,N_22494);
xnor U22720 (N_22720,N_22304,N_22294);
and U22721 (N_22721,N_22051,N_22190);
and U22722 (N_22722,N_22026,N_22125);
nor U22723 (N_22723,N_22095,N_22068);
and U22724 (N_22724,N_22356,N_22343);
xor U22725 (N_22725,N_22107,N_22490);
or U22726 (N_22726,N_22434,N_22270);
nor U22727 (N_22727,N_22342,N_22046);
xnor U22728 (N_22728,N_22271,N_22488);
nor U22729 (N_22729,N_22320,N_22041);
nand U22730 (N_22730,N_22478,N_22375);
nor U22731 (N_22731,N_22014,N_22038);
or U22732 (N_22732,N_22314,N_22371);
and U22733 (N_22733,N_22088,N_22083);
and U22734 (N_22734,N_22243,N_22152);
and U22735 (N_22735,N_22196,N_22031);
and U22736 (N_22736,N_22406,N_22065);
nor U22737 (N_22737,N_22415,N_22159);
xor U22738 (N_22738,N_22257,N_22097);
or U22739 (N_22739,N_22197,N_22355);
xnor U22740 (N_22740,N_22346,N_22384);
nor U22741 (N_22741,N_22312,N_22399);
nor U22742 (N_22742,N_22124,N_22133);
and U22743 (N_22743,N_22109,N_22362);
xnor U22744 (N_22744,N_22433,N_22464);
and U22745 (N_22745,N_22414,N_22427);
nor U22746 (N_22746,N_22132,N_22416);
or U22747 (N_22747,N_22489,N_22214);
nand U22748 (N_22748,N_22450,N_22032);
or U22749 (N_22749,N_22303,N_22369);
nor U22750 (N_22750,N_22048,N_22281);
xor U22751 (N_22751,N_22205,N_22326);
and U22752 (N_22752,N_22161,N_22328);
nand U22753 (N_22753,N_22038,N_22224);
nand U22754 (N_22754,N_22442,N_22204);
nor U22755 (N_22755,N_22149,N_22422);
xor U22756 (N_22756,N_22020,N_22443);
and U22757 (N_22757,N_22283,N_22402);
and U22758 (N_22758,N_22175,N_22227);
nor U22759 (N_22759,N_22218,N_22072);
nor U22760 (N_22760,N_22104,N_22247);
or U22761 (N_22761,N_22448,N_22255);
xnor U22762 (N_22762,N_22044,N_22229);
xor U22763 (N_22763,N_22088,N_22216);
xnor U22764 (N_22764,N_22143,N_22039);
or U22765 (N_22765,N_22494,N_22162);
and U22766 (N_22766,N_22018,N_22132);
nor U22767 (N_22767,N_22379,N_22132);
xnor U22768 (N_22768,N_22238,N_22057);
nand U22769 (N_22769,N_22143,N_22413);
nor U22770 (N_22770,N_22128,N_22396);
xnor U22771 (N_22771,N_22227,N_22012);
nand U22772 (N_22772,N_22473,N_22475);
nand U22773 (N_22773,N_22028,N_22416);
xor U22774 (N_22774,N_22083,N_22346);
and U22775 (N_22775,N_22121,N_22147);
and U22776 (N_22776,N_22250,N_22159);
xnor U22777 (N_22777,N_22405,N_22039);
nor U22778 (N_22778,N_22396,N_22098);
or U22779 (N_22779,N_22055,N_22139);
nand U22780 (N_22780,N_22302,N_22477);
or U22781 (N_22781,N_22010,N_22007);
nor U22782 (N_22782,N_22495,N_22039);
and U22783 (N_22783,N_22011,N_22000);
xnor U22784 (N_22784,N_22441,N_22400);
or U22785 (N_22785,N_22128,N_22004);
nor U22786 (N_22786,N_22122,N_22159);
xnor U22787 (N_22787,N_22193,N_22289);
xor U22788 (N_22788,N_22422,N_22168);
nand U22789 (N_22789,N_22443,N_22499);
nand U22790 (N_22790,N_22072,N_22324);
or U22791 (N_22791,N_22308,N_22494);
or U22792 (N_22792,N_22471,N_22114);
nor U22793 (N_22793,N_22398,N_22119);
xnor U22794 (N_22794,N_22175,N_22078);
and U22795 (N_22795,N_22460,N_22435);
and U22796 (N_22796,N_22234,N_22026);
xor U22797 (N_22797,N_22377,N_22047);
nand U22798 (N_22798,N_22197,N_22053);
or U22799 (N_22799,N_22423,N_22469);
nand U22800 (N_22800,N_22318,N_22170);
nor U22801 (N_22801,N_22133,N_22378);
or U22802 (N_22802,N_22287,N_22236);
nor U22803 (N_22803,N_22073,N_22120);
or U22804 (N_22804,N_22380,N_22126);
nand U22805 (N_22805,N_22224,N_22007);
or U22806 (N_22806,N_22157,N_22139);
or U22807 (N_22807,N_22103,N_22339);
or U22808 (N_22808,N_22353,N_22466);
xor U22809 (N_22809,N_22445,N_22166);
or U22810 (N_22810,N_22444,N_22248);
or U22811 (N_22811,N_22486,N_22122);
and U22812 (N_22812,N_22125,N_22245);
nand U22813 (N_22813,N_22145,N_22455);
xnor U22814 (N_22814,N_22177,N_22054);
and U22815 (N_22815,N_22350,N_22016);
and U22816 (N_22816,N_22308,N_22453);
xnor U22817 (N_22817,N_22330,N_22377);
nor U22818 (N_22818,N_22487,N_22447);
nor U22819 (N_22819,N_22404,N_22393);
nor U22820 (N_22820,N_22497,N_22184);
xor U22821 (N_22821,N_22192,N_22241);
nand U22822 (N_22822,N_22020,N_22123);
nand U22823 (N_22823,N_22149,N_22199);
nand U22824 (N_22824,N_22123,N_22048);
or U22825 (N_22825,N_22175,N_22197);
nor U22826 (N_22826,N_22096,N_22147);
and U22827 (N_22827,N_22490,N_22171);
xnor U22828 (N_22828,N_22062,N_22248);
or U22829 (N_22829,N_22028,N_22240);
nand U22830 (N_22830,N_22276,N_22101);
nor U22831 (N_22831,N_22209,N_22363);
and U22832 (N_22832,N_22194,N_22137);
xnor U22833 (N_22833,N_22101,N_22087);
nand U22834 (N_22834,N_22397,N_22377);
and U22835 (N_22835,N_22198,N_22385);
nor U22836 (N_22836,N_22468,N_22276);
nor U22837 (N_22837,N_22182,N_22246);
and U22838 (N_22838,N_22166,N_22303);
and U22839 (N_22839,N_22316,N_22133);
xor U22840 (N_22840,N_22345,N_22403);
nor U22841 (N_22841,N_22178,N_22383);
nor U22842 (N_22842,N_22439,N_22109);
nand U22843 (N_22843,N_22378,N_22373);
nand U22844 (N_22844,N_22056,N_22227);
or U22845 (N_22845,N_22364,N_22108);
and U22846 (N_22846,N_22266,N_22285);
nor U22847 (N_22847,N_22059,N_22195);
xnor U22848 (N_22848,N_22187,N_22014);
and U22849 (N_22849,N_22016,N_22051);
nand U22850 (N_22850,N_22243,N_22012);
and U22851 (N_22851,N_22193,N_22098);
xnor U22852 (N_22852,N_22283,N_22117);
nand U22853 (N_22853,N_22041,N_22111);
nor U22854 (N_22854,N_22408,N_22325);
or U22855 (N_22855,N_22279,N_22172);
nor U22856 (N_22856,N_22418,N_22035);
and U22857 (N_22857,N_22207,N_22485);
and U22858 (N_22858,N_22425,N_22255);
nand U22859 (N_22859,N_22122,N_22404);
nand U22860 (N_22860,N_22182,N_22420);
nand U22861 (N_22861,N_22020,N_22248);
and U22862 (N_22862,N_22354,N_22428);
xnor U22863 (N_22863,N_22476,N_22031);
nor U22864 (N_22864,N_22182,N_22376);
nor U22865 (N_22865,N_22425,N_22088);
nor U22866 (N_22866,N_22342,N_22234);
or U22867 (N_22867,N_22309,N_22228);
or U22868 (N_22868,N_22028,N_22200);
nand U22869 (N_22869,N_22189,N_22264);
nor U22870 (N_22870,N_22057,N_22027);
xnor U22871 (N_22871,N_22149,N_22139);
nor U22872 (N_22872,N_22208,N_22052);
and U22873 (N_22873,N_22204,N_22310);
nor U22874 (N_22874,N_22487,N_22396);
nor U22875 (N_22875,N_22273,N_22051);
nor U22876 (N_22876,N_22445,N_22124);
and U22877 (N_22877,N_22053,N_22119);
and U22878 (N_22878,N_22121,N_22132);
and U22879 (N_22879,N_22059,N_22119);
xor U22880 (N_22880,N_22324,N_22371);
nand U22881 (N_22881,N_22370,N_22379);
xor U22882 (N_22882,N_22196,N_22475);
and U22883 (N_22883,N_22096,N_22273);
nand U22884 (N_22884,N_22249,N_22115);
nand U22885 (N_22885,N_22418,N_22056);
or U22886 (N_22886,N_22434,N_22412);
xor U22887 (N_22887,N_22300,N_22190);
and U22888 (N_22888,N_22433,N_22266);
nand U22889 (N_22889,N_22390,N_22464);
nor U22890 (N_22890,N_22486,N_22397);
nand U22891 (N_22891,N_22282,N_22040);
nor U22892 (N_22892,N_22480,N_22092);
nand U22893 (N_22893,N_22257,N_22065);
and U22894 (N_22894,N_22408,N_22028);
or U22895 (N_22895,N_22377,N_22491);
nor U22896 (N_22896,N_22284,N_22421);
xor U22897 (N_22897,N_22145,N_22222);
xnor U22898 (N_22898,N_22121,N_22066);
nand U22899 (N_22899,N_22383,N_22357);
xnor U22900 (N_22900,N_22251,N_22108);
and U22901 (N_22901,N_22020,N_22183);
nand U22902 (N_22902,N_22190,N_22197);
nor U22903 (N_22903,N_22483,N_22493);
nor U22904 (N_22904,N_22295,N_22488);
nor U22905 (N_22905,N_22023,N_22442);
and U22906 (N_22906,N_22268,N_22328);
or U22907 (N_22907,N_22315,N_22359);
nor U22908 (N_22908,N_22372,N_22194);
and U22909 (N_22909,N_22119,N_22488);
and U22910 (N_22910,N_22443,N_22228);
nand U22911 (N_22911,N_22466,N_22203);
nand U22912 (N_22912,N_22150,N_22468);
or U22913 (N_22913,N_22112,N_22220);
or U22914 (N_22914,N_22115,N_22120);
xor U22915 (N_22915,N_22317,N_22183);
nor U22916 (N_22916,N_22422,N_22088);
nand U22917 (N_22917,N_22471,N_22270);
nand U22918 (N_22918,N_22244,N_22173);
nand U22919 (N_22919,N_22247,N_22370);
and U22920 (N_22920,N_22434,N_22120);
or U22921 (N_22921,N_22309,N_22225);
nor U22922 (N_22922,N_22421,N_22373);
and U22923 (N_22923,N_22378,N_22164);
nand U22924 (N_22924,N_22405,N_22306);
nor U22925 (N_22925,N_22187,N_22158);
nand U22926 (N_22926,N_22401,N_22366);
or U22927 (N_22927,N_22352,N_22247);
or U22928 (N_22928,N_22070,N_22374);
and U22929 (N_22929,N_22445,N_22107);
nor U22930 (N_22930,N_22075,N_22378);
nor U22931 (N_22931,N_22116,N_22326);
and U22932 (N_22932,N_22000,N_22429);
nor U22933 (N_22933,N_22450,N_22065);
nor U22934 (N_22934,N_22219,N_22226);
nor U22935 (N_22935,N_22271,N_22306);
or U22936 (N_22936,N_22032,N_22360);
or U22937 (N_22937,N_22369,N_22067);
and U22938 (N_22938,N_22277,N_22441);
xor U22939 (N_22939,N_22109,N_22340);
nand U22940 (N_22940,N_22217,N_22426);
and U22941 (N_22941,N_22237,N_22198);
or U22942 (N_22942,N_22376,N_22066);
and U22943 (N_22943,N_22315,N_22032);
or U22944 (N_22944,N_22166,N_22180);
or U22945 (N_22945,N_22259,N_22208);
or U22946 (N_22946,N_22279,N_22083);
and U22947 (N_22947,N_22057,N_22461);
nand U22948 (N_22948,N_22443,N_22042);
and U22949 (N_22949,N_22371,N_22422);
nor U22950 (N_22950,N_22061,N_22321);
xor U22951 (N_22951,N_22454,N_22212);
xnor U22952 (N_22952,N_22380,N_22141);
and U22953 (N_22953,N_22338,N_22071);
nand U22954 (N_22954,N_22134,N_22291);
and U22955 (N_22955,N_22083,N_22099);
xor U22956 (N_22956,N_22110,N_22277);
and U22957 (N_22957,N_22158,N_22080);
nand U22958 (N_22958,N_22010,N_22033);
xor U22959 (N_22959,N_22401,N_22373);
and U22960 (N_22960,N_22262,N_22221);
nand U22961 (N_22961,N_22271,N_22228);
nor U22962 (N_22962,N_22331,N_22099);
and U22963 (N_22963,N_22096,N_22343);
nor U22964 (N_22964,N_22045,N_22286);
nor U22965 (N_22965,N_22194,N_22000);
and U22966 (N_22966,N_22308,N_22409);
nand U22967 (N_22967,N_22155,N_22330);
and U22968 (N_22968,N_22177,N_22121);
nor U22969 (N_22969,N_22117,N_22383);
or U22970 (N_22970,N_22054,N_22465);
or U22971 (N_22971,N_22400,N_22268);
and U22972 (N_22972,N_22026,N_22065);
or U22973 (N_22973,N_22410,N_22461);
xor U22974 (N_22974,N_22030,N_22320);
nor U22975 (N_22975,N_22263,N_22126);
and U22976 (N_22976,N_22342,N_22392);
and U22977 (N_22977,N_22128,N_22197);
or U22978 (N_22978,N_22173,N_22329);
xnor U22979 (N_22979,N_22079,N_22102);
xnor U22980 (N_22980,N_22306,N_22497);
and U22981 (N_22981,N_22023,N_22392);
and U22982 (N_22982,N_22001,N_22426);
nand U22983 (N_22983,N_22335,N_22407);
and U22984 (N_22984,N_22476,N_22060);
and U22985 (N_22985,N_22360,N_22287);
xnor U22986 (N_22986,N_22029,N_22464);
nand U22987 (N_22987,N_22016,N_22497);
nor U22988 (N_22988,N_22027,N_22382);
nor U22989 (N_22989,N_22102,N_22095);
or U22990 (N_22990,N_22361,N_22494);
nor U22991 (N_22991,N_22476,N_22191);
xnor U22992 (N_22992,N_22421,N_22337);
nand U22993 (N_22993,N_22125,N_22116);
nand U22994 (N_22994,N_22410,N_22438);
nor U22995 (N_22995,N_22380,N_22104);
and U22996 (N_22996,N_22007,N_22146);
xnor U22997 (N_22997,N_22390,N_22150);
and U22998 (N_22998,N_22202,N_22020);
and U22999 (N_22999,N_22292,N_22285);
or U23000 (N_23000,N_22998,N_22878);
and U23001 (N_23001,N_22584,N_22853);
xnor U23002 (N_23002,N_22861,N_22784);
nand U23003 (N_23003,N_22920,N_22902);
xnor U23004 (N_23004,N_22780,N_22982);
nand U23005 (N_23005,N_22627,N_22661);
and U23006 (N_23006,N_22806,N_22548);
xor U23007 (N_23007,N_22538,N_22725);
nor U23008 (N_23008,N_22886,N_22951);
nand U23009 (N_23009,N_22821,N_22828);
nand U23010 (N_23010,N_22810,N_22573);
nor U23011 (N_23011,N_22756,N_22767);
nand U23012 (N_23012,N_22874,N_22608);
xnor U23013 (N_23013,N_22818,N_22803);
nor U23014 (N_23014,N_22936,N_22716);
nor U23015 (N_23015,N_22929,N_22642);
and U23016 (N_23016,N_22906,N_22896);
xor U23017 (N_23017,N_22855,N_22536);
or U23018 (N_23018,N_22659,N_22879);
nor U23019 (N_23019,N_22703,N_22743);
nand U23020 (N_23020,N_22993,N_22647);
nand U23021 (N_23021,N_22771,N_22839);
nor U23022 (N_23022,N_22805,N_22822);
and U23023 (N_23023,N_22513,N_22782);
and U23024 (N_23024,N_22612,N_22997);
nand U23025 (N_23025,N_22903,N_22996);
and U23026 (N_23026,N_22507,N_22582);
or U23027 (N_23027,N_22745,N_22624);
nor U23028 (N_23028,N_22798,N_22986);
or U23029 (N_23029,N_22741,N_22918);
nand U23030 (N_23030,N_22824,N_22788);
nand U23031 (N_23031,N_22511,N_22533);
nand U23032 (N_23032,N_22846,N_22712);
and U23033 (N_23033,N_22719,N_22710);
and U23034 (N_23034,N_22552,N_22924);
or U23035 (N_23035,N_22772,N_22877);
xnor U23036 (N_23036,N_22655,N_22530);
nand U23037 (N_23037,N_22962,N_22979);
nor U23038 (N_23038,N_22945,N_22563);
xnor U23039 (N_23039,N_22983,N_22975);
xnor U23040 (N_23040,N_22505,N_22851);
or U23041 (N_23041,N_22750,N_22724);
and U23042 (N_23042,N_22572,N_22518);
or U23043 (N_23043,N_22674,N_22876);
nand U23044 (N_23044,N_22592,N_22885);
nand U23045 (N_23045,N_22680,N_22893);
or U23046 (N_23046,N_22637,N_22907);
and U23047 (N_23047,N_22746,N_22599);
xnor U23048 (N_23048,N_22663,N_22950);
or U23049 (N_23049,N_22978,N_22574);
xor U23050 (N_23050,N_22889,N_22905);
or U23051 (N_23051,N_22706,N_22510);
nand U23052 (N_23052,N_22671,N_22562);
or U23053 (N_23053,N_22525,N_22587);
nand U23054 (N_23054,N_22921,N_22537);
nand U23055 (N_23055,N_22653,N_22890);
nor U23056 (N_23056,N_22568,N_22985);
and U23057 (N_23057,N_22581,N_22755);
nor U23058 (N_23058,N_22974,N_22698);
xnor U23059 (N_23059,N_22808,N_22875);
xnor U23060 (N_23060,N_22911,N_22912);
or U23061 (N_23061,N_22534,N_22652);
nor U23062 (N_23062,N_22901,N_22579);
xnor U23063 (N_23063,N_22789,N_22629);
nor U23064 (N_23064,N_22994,N_22517);
xor U23065 (N_23065,N_22696,N_22664);
xnor U23066 (N_23066,N_22588,N_22832);
or U23067 (N_23067,N_22506,N_22555);
or U23068 (N_23068,N_22923,N_22963);
nor U23069 (N_23069,N_22881,N_22692);
nor U23070 (N_23070,N_22501,N_22880);
xnor U23071 (N_23071,N_22927,N_22954);
nand U23072 (N_23072,N_22988,N_22728);
or U23073 (N_23073,N_22614,N_22977);
or U23074 (N_23074,N_22593,N_22762);
nor U23075 (N_23075,N_22631,N_22633);
xor U23076 (N_23076,N_22842,N_22723);
nor U23077 (N_23077,N_22730,N_22726);
nand U23078 (N_23078,N_22531,N_22705);
nor U23079 (N_23079,N_22969,N_22502);
xor U23080 (N_23080,N_22882,N_22859);
nand U23081 (N_23081,N_22697,N_22623);
nand U23082 (N_23082,N_22535,N_22625);
nor U23083 (N_23083,N_22564,N_22699);
xnor U23084 (N_23084,N_22558,N_22681);
nand U23085 (N_23085,N_22868,N_22672);
and U23086 (N_23086,N_22778,N_22826);
and U23087 (N_23087,N_22595,N_22503);
and U23088 (N_23088,N_22991,N_22686);
and U23089 (N_23089,N_22753,N_22727);
xnor U23090 (N_23090,N_22961,N_22733);
and U23091 (N_23091,N_22662,N_22952);
or U23092 (N_23092,N_22748,N_22613);
and U23093 (N_23093,N_22900,N_22646);
nor U23094 (N_23094,N_22620,N_22643);
xor U23095 (N_23095,N_22688,N_22999);
nand U23096 (N_23096,N_22667,N_22871);
nor U23097 (N_23097,N_22561,N_22636);
nor U23098 (N_23098,N_22640,N_22892);
or U23099 (N_23099,N_22843,N_22591);
or U23100 (N_23100,N_22687,N_22791);
nor U23101 (N_23101,N_22823,N_22834);
nor U23102 (N_23102,N_22779,N_22575);
xor U23103 (N_23103,N_22632,N_22565);
or U23104 (N_23104,N_22870,N_22500);
xnor U23105 (N_23105,N_22934,N_22528);
xor U23106 (N_23106,N_22731,N_22928);
and U23107 (N_23107,N_22601,N_22759);
and U23108 (N_23108,N_22609,N_22628);
xnor U23109 (N_23109,N_22669,N_22713);
nand U23110 (N_23110,N_22957,N_22542);
nor U23111 (N_23111,N_22840,N_22690);
or U23112 (N_23112,N_22630,N_22651);
nor U23113 (N_23113,N_22797,N_22795);
nand U23114 (N_23114,N_22915,N_22816);
and U23115 (N_23115,N_22891,N_22850);
nor U23116 (N_23116,N_22847,N_22639);
nand U23117 (N_23117,N_22958,N_22666);
and U23118 (N_23118,N_22862,N_22953);
nand U23119 (N_23119,N_22682,N_22973);
or U23120 (N_23120,N_22888,N_22761);
xnor U23121 (N_23121,N_22786,N_22960);
and U23122 (N_23122,N_22838,N_22768);
nor U23123 (N_23123,N_22740,N_22649);
or U23124 (N_23124,N_22551,N_22932);
xor U23125 (N_23125,N_22580,N_22645);
xor U23126 (N_23126,N_22971,N_22635);
or U23127 (N_23127,N_22760,N_22689);
nor U23128 (N_23128,N_22829,N_22956);
or U23129 (N_23129,N_22849,N_22781);
nand U23130 (N_23130,N_22955,N_22769);
xor U23131 (N_23131,N_22913,N_22827);
and U23132 (N_23132,N_22775,N_22641);
xor U23133 (N_23133,N_22966,N_22841);
nand U23134 (N_23134,N_22804,N_22813);
or U23135 (N_23135,N_22939,N_22549);
or U23136 (N_23136,N_22700,N_22749);
xor U23137 (N_23137,N_22863,N_22856);
xnor U23138 (N_23138,N_22708,N_22967);
and U23139 (N_23139,N_22830,N_22949);
and U23140 (N_23140,N_22557,N_22658);
xor U23141 (N_23141,N_22774,N_22948);
and U23142 (N_23142,N_22754,N_22544);
nor U23143 (N_23143,N_22519,N_22509);
and U23144 (N_23144,N_22668,N_22981);
nor U23145 (N_23145,N_22770,N_22576);
nand U23146 (N_23146,N_22515,N_22607);
nand U23147 (N_23147,N_22757,N_22873);
or U23148 (N_23148,N_22701,N_22919);
and U23149 (N_23149,N_22898,N_22704);
and U23150 (N_23150,N_22941,N_22590);
nor U23151 (N_23151,N_22908,N_22989);
xor U23152 (N_23152,N_22776,N_22514);
nand U23153 (N_23153,N_22739,N_22732);
or U23154 (N_23154,N_22793,N_22621);
nor U23155 (N_23155,N_22657,N_22540);
nand U23156 (N_23156,N_22578,N_22938);
or U23157 (N_23157,N_22820,N_22566);
or U23158 (N_23158,N_22819,N_22995);
nor U23159 (N_23159,N_22883,N_22765);
nor U23160 (N_23160,N_22512,N_22872);
xnor U23161 (N_23161,N_22600,N_22931);
nor U23162 (N_23162,N_22887,N_22984);
nor U23163 (N_23163,N_22917,N_22683);
nor U23164 (N_23164,N_22935,N_22707);
nor U23165 (N_23165,N_22837,N_22852);
or U23166 (N_23166,N_22812,N_22718);
nand U23167 (N_23167,N_22744,N_22679);
or U23168 (N_23168,N_22532,N_22922);
or U23169 (N_23169,N_22622,N_22583);
or U23170 (N_23170,N_22764,N_22848);
or U23171 (N_23171,N_22735,N_22702);
nand U23172 (N_23172,N_22940,N_22809);
nor U23173 (N_23173,N_22790,N_22670);
and U23174 (N_23174,N_22550,N_22800);
nand U23175 (N_23175,N_22648,N_22794);
xnor U23176 (N_23176,N_22547,N_22617);
or U23177 (N_23177,N_22527,N_22815);
and U23178 (N_23178,N_22529,N_22729);
or U23179 (N_23179,N_22836,N_22626);
or U23180 (N_23180,N_22865,N_22942);
xor U23181 (N_23181,N_22673,N_22844);
nand U23182 (N_23182,N_22654,N_22721);
nor U23183 (N_23183,N_22554,N_22715);
and U23184 (N_23184,N_22560,N_22546);
xnor U23185 (N_23185,N_22904,N_22976);
nor U23186 (N_23186,N_22720,N_22585);
xor U23187 (N_23187,N_22539,N_22763);
nor U23188 (N_23188,N_22615,N_22899);
or U23189 (N_23189,N_22693,N_22691);
nor U23190 (N_23190,N_22526,N_22930);
nand U23191 (N_23191,N_22783,N_22857);
or U23192 (N_23192,N_22677,N_22678);
nand U23193 (N_23193,N_22675,N_22752);
xor U23194 (N_23194,N_22968,N_22990);
and U23195 (N_23195,N_22959,N_22831);
and U23196 (N_23196,N_22965,N_22577);
or U23197 (N_23197,N_22894,N_22944);
and U23198 (N_23198,N_22597,N_22619);
and U23199 (N_23199,N_22773,N_22736);
xor U23200 (N_23200,N_22858,N_22695);
or U23201 (N_23201,N_22970,N_22650);
nand U23202 (N_23202,N_22937,N_22825);
or U23203 (N_23203,N_22711,N_22787);
nand U23204 (N_23204,N_22802,N_22606);
nor U23205 (N_23205,N_22660,N_22508);
nand U23206 (N_23206,N_22709,N_22522);
or U23207 (N_23207,N_22644,N_22604);
or U23208 (N_23208,N_22602,N_22589);
nor U23209 (N_23209,N_22616,N_22925);
and U23210 (N_23210,N_22747,N_22864);
or U23211 (N_23211,N_22559,N_22926);
nor U23212 (N_23212,N_22964,N_22586);
nand U23213 (N_23213,N_22738,N_22634);
and U23214 (N_23214,N_22570,N_22665);
nand U23215 (N_23215,N_22734,N_22553);
or U23216 (N_23216,N_22610,N_22594);
xnor U23217 (N_23217,N_22605,N_22777);
and U23218 (N_23218,N_22909,N_22524);
nand U23219 (N_23219,N_22766,N_22884);
nor U23220 (N_23220,N_22946,N_22751);
nand U23221 (N_23221,N_22916,N_22799);
xnor U23222 (N_23222,N_22676,N_22933);
nand U23223 (N_23223,N_22571,N_22987);
and U23224 (N_23224,N_22980,N_22656);
xor U23225 (N_23225,N_22504,N_22947);
or U23226 (N_23226,N_22541,N_22722);
and U23227 (N_23227,N_22910,N_22556);
and U23228 (N_23228,N_22835,N_22792);
or U23229 (N_23229,N_22618,N_22737);
nor U23230 (N_23230,N_22694,N_22866);
and U23231 (N_23231,N_22914,N_22717);
and U23232 (N_23232,N_22811,N_22972);
or U23233 (N_23233,N_22569,N_22867);
or U23234 (N_23234,N_22603,N_22785);
xnor U23235 (N_23235,N_22807,N_22854);
and U23236 (N_23236,N_22860,N_22543);
nor U23237 (N_23237,N_22638,N_22596);
or U23238 (N_23238,N_22684,N_22742);
or U23239 (N_23239,N_22897,N_22814);
and U23240 (N_23240,N_22567,N_22545);
nand U23241 (N_23241,N_22521,N_22520);
xnor U23242 (N_23242,N_22895,N_22598);
and U23243 (N_23243,N_22992,N_22817);
or U23244 (N_23244,N_22685,N_22758);
and U23245 (N_23245,N_22845,N_22611);
and U23246 (N_23246,N_22516,N_22943);
nor U23247 (N_23247,N_22796,N_22801);
nand U23248 (N_23248,N_22714,N_22523);
and U23249 (N_23249,N_22833,N_22869);
or U23250 (N_23250,N_22647,N_22835);
or U23251 (N_23251,N_22710,N_22624);
nor U23252 (N_23252,N_22823,N_22570);
xnor U23253 (N_23253,N_22621,N_22508);
nand U23254 (N_23254,N_22692,N_22538);
and U23255 (N_23255,N_22938,N_22603);
or U23256 (N_23256,N_22786,N_22836);
or U23257 (N_23257,N_22832,N_22866);
nor U23258 (N_23258,N_22960,N_22699);
nand U23259 (N_23259,N_22940,N_22774);
nand U23260 (N_23260,N_22957,N_22846);
xor U23261 (N_23261,N_22768,N_22869);
xnor U23262 (N_23262,N_22517,N_22690);
and U23263 (N_23263,N_22807,N_22631);
nor U23264 (N_23264,N_22881,N_22521);
or U23265 (N_23265,N_22550,N_22769);
and U23266 (N_23266,N_22553,N_22884);
nor U23267 (N_23267,N_22506,N_22804);
nand U23268 (N_23268,N_22845,N_22883);
and U23269 (N_23269,N_22643,N_22943);
or U23270 (N_23270,N_22574,N_22507);
xnor U23271 (N_23271,N_22575,N_22706);
and U23272 (N_23272,N_22788,N_22503);
xor U23273 (N_23273,N_22874,N_22573);
or U23274 (N_23274,N_22783,N_22669);
nor U23275 (N_23275,N_22914,N_22536);
and U23276 (N_23276,N_22840,N_22873);
and U23277 (N_23277,N_22525,N_22947);
or U23278 (N_23278,N_22669,N_22876);
nor U23279 (N_23279,N_22941,N_22911);
nand U23280 (N_23280,N_22598,N_22761);
and U23281 (N_23281,N_22890,N_22593);
and U23282 (N_23282,N_22739,N_22686);
nand U23283 (N_23283,N_22731,N_22741);
xnor U23284 (N_23284,N_22989,N_22971);
nor U23285 (N_23285,N_22868,N_22548);
or U23286 (N_23286,N_22575,N_22644);
nor U23287 (N_23287,N_22802,N_22765);
nand U23288 (N_23288,N_22657,N_22574);
nor U23289 (N_23289,N_22866,N_22598);
nand U23290 (N_23290,N_22921,N_22623);
xnor U23291 (N_23291,N_22806,N_22656);
or U23292 (N_23292,N_22892,N_22578);
xor U23293 (N_23293,N_22954,N_22845);
nand U23294 (N_23294,N_22526,N_22974);
xor U23295 (N_23295,N_22523,N_22930);
nand U23296 (N_23296,N_22753,N_22849);
xor U23297 (N_23297,N_22644,N_22869);
nand U23298 (N_23298,N_22945,N_22930);
nor U23299 (N_23299,N_22584,N_22972);
nor U23300 (N_23300,N_22865,N_22895);
and U23301 (N_23301,N_22810,N_22764);
xnor U23302 (N_23302,N_22700,N_22683);
nand U23303 (N_23303,N_22894,N_22550);
or U23304 (N_23304,N_22833,N_22701);
nand U23305 (N_23305,N_22957,N_22606);
and U23306 (N_23306,N_22544,N_22988);
xnor U23307 (N_23307,N_22820,N_22782);
xor U23308 (N_23308,N_22598,N_22787);
nand U23309 (N_23309,N_22830,N_22874);
or U23310 (N_23310,N_22966,N_22836);
xor U23311 (N_23311,N_22964,N_22795);
nand U23312 (N_23312,N_22784,N_22578);
nor U23313 (N_23313,N_22969,N_22590);
and U23314 (N_23314,N_22752,N_22639);
xnor U23315 (N_23315,N_22750,N_22924);
nand U23316 (N_23316,N_22947,N_22602);
or U23317 (N_23317,N_22563,N_22606);
nand U23318 (N_23318,N_22758,N_22726);
nor U23319 (N_23319,N_22692,N_22640);
and U23320 (N_23320,N_22521,N_22920);
and U23321 (N_23321,N_22952,N_22727);
xnor U23322 (N_23322,N_22796,N_22560);
and U23323 (N_23323,N_22502,N_22774);
and U23324 (N_23324,N_22806,N_22531);
and U23325 (N_23325,N_22767,N_22657);
and U23326 (N_23326,N_22950,N_22733);
nand U23327 (N_23327,N_22837,N_22971);
nor U23328 (N_23328,N_22524,N_22912);
xnor U23329 (N_23329,N_22868,N_22836);
and U23330 (N_23330,N_22814,N_22500);
xnor U23331 (N_23331,N_22839,N_22607);
and U23332 (N_23332,N_22722,N_22811);
xnor U23333 (N_23333,N_22868,N_22910);
or U23334 (N_23334,N_22749,N_22543);
and U23335 (N_23335,N_22988,N_22877);
nor U23336 (N_23336,N_22548,N_22789);
or U23337 (N_23337,N_22578,N_22949);
or U23338 (N_23338,N_22556,N_22584);
xnor U23339 (N_23339,N_22989,N_22747);
or U23340 (N_23340,N_22640,N_22845);
or U23341 (N_23341,N_22911,N_22840);
nor U23342 (N_23342,N_22799,N_22845);
xnor U23343 (N_23343,N_22718,N_22630);
xnor U23344 (N_23344,N_22629,N_22533);
nand U23345 (N_23345,N_22682,N_22921);
nor U23346 (N_23346,N_22682,N_22501);
and U23347 (N_23347,N_22874,N_22776);
nand U23348 (N_23348,N_22576,N_22853);
or U23349 (N_23349,N_22845,N_22727);
xnor U23350 (N_23350,N_22621,N_22764);
or U23351 (N_23351,N_22518,N_22714);
nor U23352 (N_23352,N_22561,N_22691);
xor U23353 (N_23353,N_22755,N_22871);
xor U23354 (N_23354,N_22998,N_22824);
or U23355 (N_23355,N_22986,N_22763);
nand U23356 (N_23356,N_22606,N_22526);
xor U23357 (N_23357,N_22871,N_22578);
or U23358 (N_23358,N_22891,N_22856);
nand U23359 (N_23359,N_22525,N_22664);
and U23360 (N_23360,N_22521,N_22710);
nor U23361 (N_23361,N_22983,N_22910);
and U23362 (N_23362,N_22582,N_22535);
nand U23363 (N_23363,N_22700,N_22657);
and U23364 (N_23364,N_22649,N_22689);
xor U23365 (N_23365,N_22612,N_22665);
and U23366 (N_23366,N_22591,N_22779);
and U23367 (N_23367,N_22716,N_22655);
xor U23368 (N_23368,N_22679,N_22839);
or U23369 (N_23369,N_22734,N_22994);
and U23370 (N_23370,N_22660,N_22567);
and U23371 (N_23371,N_22680,N_22529);
nand U23372 (N_23372,N_22917,N_22984);
nand U23373 (N_23373,N_22856,N_22963);
and U23374 (N_23374,N_22682,N_22572);
nor U23375 (N_23375,N_22649,N_22669);
or U23376 (N_23376,N_22574,N_22892);
nand U23377 (N_23377,N_22616,N_22729);
or U23378 (N_23378,N_22883,N_22849);
nand U23379 (N_23379,N_22819,N_22962);
xor U23380 (N_23380,N_22845,N_22893);
nor U23381 (N_23381,N_22935,N_22971);
and U23382 (N_23382,N_22982,N_22882);
nand U23383 (N_23383,N_22595,N_22548);
nand U23384 (N_23384,N_22749,N_22722);
nand U23385 (N_23385,N_22931,N_22571);
nand U23386 (N_23386,N_22820,N_22796);
and U23387 (N_23387,N_22753,N_22810);
nand U23388 (N_23388,N_22629,N_22615);
nor U23389 (N_23389,N_22747,N_22954);
or U23390 (N_23390,N_22987,N_22869);
or U23391 (N_23391,N_22766,N_22640);
nand U23392 (N_23392,N_22914,N_22558);
nand U23393 (N_23393,N_22576,N_22559);
or U23394 (N_23394,N_22711,N_22643);
and U23395 (N_23395,N_22660,N_22829);
nand U23396 (N_23396,N_22803,N_22515);
and U23397 (N_23397,N_22828,N_22815);
nand U23398 (N_23398,N_22761,N_22914);
or U23399 (N_23399,N_22730,N_22747);
nand U23400 (N_23400,N_22597,N_22813);
and U23401 (N_23401,N_22824,N_22988);
or U23402 (N_23402,N_22749,N_22662);
nor U23403 (N_23403,N_22581,N_22999);
or U23404 (N_23404,N_22854,N_22887);
nor U23405 (N_23405,N_22669,N_22708);
nand U23406 (N_23406,N_22526,N_22679);
and U23407 (N_23407,N_22802,N_22914);
nor U23408 (N_23408,N_22562,N_22820);
or U23409 (N_23409,N_22877,N_22618);
nand U23410 (N_23410,N_22697,N_22561);
or U23411 (N_23411,N_22554,N_22713);
nand U23412 (N_23412,N_22588,N_22739);
nor U23413 (N_23413,N_22948,N_22509);
and U23414 (N_23414,N_22816,N_22932);
xor U23415 (N_23415,N_22672,N_22816);
nand U23416 (N_23416,N_22980,N_22752);
or U23417 (N_23417,N_22538,N_22717);
nor U23418 (N_23418,N_22576,N_22516);
nand U23419 (N_23419,N_22829,N_22501);
or U23420 (N_23420,N_22810,N_22859);
nand U23421 (N_23421,N_22968,N_22515);
nand U23422 (N_23422,N_22980,N_22619);
nand U23423 (N_23423,N_22700,N_22934);
or U23424 (N_23424,N_22992,N_22871);
xor U23425 (N_23425,N_22803,N_22963);
and U23426 (N_23426,N_22961,N_22778);
or U23427 (N_23427,N_22564,N_22596);
or U23428 (N_23428,N_22974,N_22730);
xnor U23429 (N_23429,N_22700,N_22806);
nor U23430 (N_23430,N_22724,N_22548);
or U23431 (N_23431,N_22689,N_22935);
and U23432 (N_23432,N_22760,N_22742);
and U23433 (N_23433,N_22640,N_22826);
nor U23434 (N_23434,N_22959,N_22889);
nor U23435 (N_23435,N_22662,N_22643);
nand U23436 (N_23436,N_22721,N_22791);
nand U23437 (N_23437,N_22741,N_22728);
nor U23438 (N_23438,N_22602,N_22535);
nor U23439 (N_23439,N_22569,N_22942);
xor U23440 (N_23440,N_22776,N_22872);
and U23441 (N_23441,N_22832,N_22733);
nor U23442 (N_23442,N_22683,N_22711);
xor U23443 (N_23443,N_22726,N_22695);
nor U23444 (N_23444,N_22684,N_22824);
and U23445 (N_23445,N_22750,N_22610);
xnor U23446 (N_23446,N_22704,N_22564);
and U23447 (N_23447,N_22828,N_22552);
and U23448 (N_23448,N_22739,N_22681);
or U23449 (N_23449,N_22617,N_22621);
or U23450 (N_23450,N_22811,N_22612);
and U23451 (N_23451,N_22867,N_22557);
xnor U23452 (N_23452,N_22731,N_22633);
and U23453 (N_23453,N_22802,N_22758);
xor U23454 (N_23454,N_22873,N_22778);
or U23455 (N_23455,N_22503,N_22861);
xnor U23456 (N_23456,N_22703,N_22657);
and U23457 (N_23457,N_22716,N_22878);
and U23458 (N_23458,N_22805,N_22629);
and U23459 (N_23459,N_22839,N_22926);
nor U23460 (N_23460,N_22511,N_22579);
nor U23461 (N_23461,N_22672,N_22930);
xor U23462 (N_23462,N_22702,N_22943);
and U23463 (N_23463,N_22879,N_22715);
xnor U23464 (N_23464,N_22723,N_22819);
xor U23465 (N_23465,N_22984,N_22943);
nor U23466 (N_23466,N_22556,N_22775);
and U23467 (N_23467,N_22784,N_22510);
or U23468 (N_23468,N_22648,N_22888);
nand U23469 (N_23469,N_22815,N_22886);
or U23470 (N_23470,N_22632,N_22508);
nand U23471 (N_23471,N_22887,N_22943);
and U23472 (N_23472,N_22851,N_22794);
nand U23473 (N_23473,N_22541,N_22760);
xor U23474 (N_23474,N_22623,N_22780);
or U23475 (N_23475,N_22633,N_22821);
nor U23476 (N_23476,N_22654,N_22653);
or U23477 (N_23477,N_22707,N_22741);
nor U23478 (N_23478,N_22555,N_22692);
xor U23479 (N_23479,N_22639,N_22803);
or U23480 (N_23480,N_22862,N_22776);
nor U23481 (N_23481,N_22603,N_22880);
and U23482 (N_23482,N_22961,N_22582);
and U23483 (N_23483,N_22949,N_22714);
nand U23484 (N_23484,N_22669,N_22534);
or U23485 (N_23485,N_22660,N_22786);
and U23486 (N_23486,N_22868,N_22510);
xor U23487 (N_23487,N_22881,N_22723);
or U23488 (N_23488,N_22531,N_22653);
xnor U23489 (N_23489,N_22758,N_22774);
nand U23490 (N_23490,N_22710,N_22983);
and U23491 (N_23491,N_22899,N_22516);
nand U23492 (N_23492,N_22723,N_22827);
and U23493 (N_23493,N_22867,N_22762);
nand U23494 (N_23494,N_22586,N_22911);
nor U23495 (N_23495,N_22504,N_22588);
xnor U23496 (N_23496,N_22897,N_22737);
nor U23497 (N_23497,N_22923,N_22546);
or U23498 (N_23498,N_22520,N_22865);
nand U23499 (N_23499,N_22822,N_22817);
nor U23500 (N_23500,N_23138,N_23428);
and U23501 (N_23501,N_23019,N_23416);
nand U23502 (N_23502,N_23192,N_23010);
nand U23503 (N_23503,N_23142,N_23223);
nand U23504 (N_23504,N_23091,N_23444);
nand U23505 (N_23505,N_23017,N_23246);
nor U23506 (N_23506,N_23033,N_23440);
nand U23507 (N_23507,N_23011,N_23035);
nor U23508 (N_23508,N_23002,N_23047);
and U23509 (N_23509,N_23180,N_23059);
nor U23510 (N_23510,N_23158,N_23294);
xor U23511 (N_23511,N_23382,N_23023);
xnor U23512 (N_23512,N_23490,N_23202);
and U23513 (N_23513,N_23208,N_23216);
or U23514 (N_23514,N_23178,N_23042);
xor U23515 (N_23515,N_23092,N_23187);
nand U23516 (N_23516,N_23296,N_23298);
nand U23517 (N_23517,N_23012,N_23140);
nor U23518 (N_23518,N_23212,N_23262);
or U23519 (N_23519,N_23380,N_23329);
xor U23520 (N_23520,N_23280,N_23462);
or U23521 (N_23521,N_23452,N_23018);
and U23522 (N_23522,N_23277,N_23020);
nand U23523 (N_23523,N_23373,N_23321);
and U23524 (N_23524,N_23314,N_23224);
nor U23525 (N_23525,N_23226,N_23170);
nand U23526 (N_23526,N_23176,N_23413);
and U23527 (N_23527,N_23122,N_23328);
nand U23528 (N_23528,N_23356,N_23389);
xor U23529 (N_23529,N_23097,N_23426);
nor U23530 (N_23530,N_23028,N_23473);
nand U23531 (N_23531,N_23293,N_23250);
nor U23532 (N_23532,N_23197,N_23194);
nor U23533 (N_23533,N_23007,N_23434);
or U23534 (N_23534,N_23248,N_23255);
xor U23535 (N_23535,N_23087,N_23311);
and U23536 (N_23536,N_23319,N_23334);
nor U23537 (N_23537,N_23228,N_23244);
nor U23538 (N_23538,N_23268,N_23256);
nand U23539 (N_23539,N_23271,N_23346);
nand U23540 (N_23540,N_23193,N_23129);
nor U23541 (N_23541,N_23366,N_23353);
xnor U23542 (N_23542,N_23415,N_23204);
xnor U23543 (N_23543,N_23046,N_23207);
nand U23544 (N_23544,N_23040,N_23126);
or U23545 (N_23545,N_23370,N_23069);
and U23546 (N_23546,N_23151,N_23326);
xnor U23547 (N_23547,N_23232,N_23340);
nor U23548 (N_23548,N_23190,N_23198);
or U23549 (N_23549,N_23199,N_23461);
nor U23550 (N_23550,N_23390,N_23481);
nand U23551 (N_23551,N_23006,N_23215);
nor U23552 (N_23552,N_23322,N_23359);
nand U23553 (N_23553,N_23082,N_23484);
nand U23554 (N_23554,N_23474,N_23371);
and U23555 (N_23555,N_23300,N_23430);
nor U23556 (N_23556,N_23029,N_23352);
nand U23557 (N_23557,N_23449,N_23072);
and U23558 (N_23558,N_23281,N_23445);
or U23559 (N_23559,N_23374,N_23175);
or U23560 (N_23560,N_23121,N_23275);
xor U23561 (N_23561,N_23339,N_23480);
nor U23562 (N_23562,N_23306,N_23297);
nor U23563 (N_23563,N_23387,N_23458);
nand U23564 (N_23564,N_23213,N_23379);
and U23565 (N_23565,N_23264,N_23009);
and U23566 (N_23566,N_23441,N_23134);
nand U23567 (N_23567,N_23437,N_23320);
and U23568 (N_23568,N_23291,N_23316);
xor U23569 (N_23569,N_23354,N_23229);
xnor U23570 (N_23570,N_23312,N_23357);
nand U23571 (N_23571,N_23478,N_23234);
nor U23572 (N_23572,N_23031,N_23472);
or U23573 (N_23573,N_23102,N_23128);
nand U23574 (N_23574,N_23000,N_23014);
and U23575 (N_23575,N_23108,N_23396);
or U23576 (N_23576,N_23162,N_23499);
nor U23577 (N_23577,N_23496,N_23290);
nand U23578 (N_23578,N_23165,N_23083);
and U23579 (N_23579,N_23049,N_23350);
xnor U23580 (N_23580,N_23355,N_23203);
xor U23581 (N_23581,N_23111,N_23299);
nand U23582 (N_23582,N_23285,N_23343);
or U23583 (N_23583,N_23062,N_23055);
xnor U23584 (N_23584,N_23420,N_23043);
nand U23585 (N_23585,N_23399,N_23471);
nor U23586 (N_23586,N_23136,N_23177);
xor U23587 (N_23587,N_23094,N_23081);
xnor U23588 (N_23588,N_23377,N_23460);
and U23589 (N_23589,N_23022,N_23447);
nor U23590 (N_23590,N_23470,N_23100);
nand U23591 (N_23591,N_23467,N_23362);
or U23592 (N_23592,N_23130,N_23364);
nand U23593 (N_23593,N_23196,N_23107);
and U23594 (N_23594,N_23331,N_23464);
nor U23595 (N_23595,N_23261,N_23150);
xnor U23596 (N_23596,N_23302,N_23409);
xor U23597 (N_23597,N_23372,N_23336);
and U23598 (N_23598,N_23424,N_23394);
nand U23599 (N_23599,N_23034,N_23061);
nand U23600 (N_23600,N_23421,N_23206);
nand U23601 (N_23601,N_23384,N_23013);
xor U23602 (N_23602,N_23227,N_23147);
xor U23603 (N_23603,N_23454,N_23288);
or U23604 (N_23604,N_23123,N_23341);
xor U23605 (N_23605,N_23408,N_23272);
or U23606 (N_23606,N_23221,N_23279);
xor U23607 (N_23607,N_23309,N_23289);
and U23608 (N_23608,N_23103,N_23497);
or U23609 (N_23609,N_23349,N_23383);
xor U23610 (N_23610,N_23404,N_23431);
xor U23611 (N_23611,N_23469,N_23335);
nand U23612 (N_23612,N_23463,N_23105);
nand U23613 (N_23613,N_23425,N_23179);
nand U23614 (N_23614,N_23378,N_23210);
nand U23615 (N_23615,N_23479,N_23418);
and U23616 (N_23616,N_23025,N_23344);
nand U23617 (N_23617,N_23112,N_23144);
xnor U23618 (N_23618,N_23295,N_23239);
nand U23619 (N_23619,N_23395,N_23201);
xor U23620 (N_23620,N_23269,N_23429);
nor U23621 (N_23621,N_23278,N_23422);
and U23622 (N_23622,N_23067,N_23286);
or U23623 (N_23623,N_23361,N_23358);
nand U23624 (N_23624,N_23058,N_23183);
xor U23625 (N_23625,N_23405,N_23171);
nor U23626 (N_23626,N_23037,N_23241);
or U23627 (N_23627,N_23127,N_23044);
nand U23628 (N_23628,N_23071,N_23304);
and U23629 (N_23629,N_23391,N_23117);
and U23630 (N_23630,N_23149,N_23168);
and U23631 (N_23631,N_23410,N_23200);
xor U23632 (N_23632,N_23393,N_23003);
and U23633 (N_23633,N_23257,N_23095);
nor U23634 (N_23634,N_23085,N_23265);
xor U23635 (N_23635,N_23402,N_23001);
xor U23636 (N_23636,N_23411,N_23016);
xnor U23637 (N_23637,N_23315,N_23096);
nor U23638 (N_23638,N_23026,N_23045);
and U23639 (N_23639,N_23266,N_23076);
or U23640 (N_23640,N_23342,N_23351);
and U23641 (N_23641,N_23041,N_23381);
xnor U23642 (N_23642,N_23073,N_23459);
nand U23643 (N_23643,N_23086,N_23439);
and U23644 (N_23644,N_23063,N_23120);
nor U23645 (N_23645,N_23053,N_23222);
nor U23646 (N_23646,N_23348,N_23488);
xnor U23647 (N_23647,N_23154,N_23468);
or U23648 (N_23648,N_23156,N_23475);
nand U23649 (N_23649,N_23466,N_23231);
nor U23650 (N_23650,N_23407,N_23008);
xnor U23651 (N_23651,N_23423,N_23456);
and U23652 (N_23652,N_23174,N_23465);
xor U23653 (N_23653,N_23125,N_23066);
or U23654 (N_23654,N_23401,N_23078);
and U23655 (N_23655,N_23249,N_23038);
nand U23656 (N_23656,N_23317,N_23330);
or U23657 (N_23657,N_23274,N_23104);
xnor U23658 (N_23658,N_23365,N_23432);
or U23659 (N_23659,N_23163,N_23021);
nand U23660 (N_23660,N_23015,N_23027);
nor U23661 (N_23661,N_23030,N_23345);
nor U23662 (N_23662,N_23109,N_23492);
nor U23663 (N_23663,N_23282,N_23400);
or U23664 (N_23664,N_23186,N_23417);
and U23665 (N_23665,N_23077,N_23476);
nand U23666 (N_23666,N_23483,N_23135);
xnor U23667 (N_23667,N_23181,N_23245);
and U23668 (N_23668,N_23435,N_23427);
nor U23669 (N_23669,N_23386,N_23392);
xnor U23670 (N_23670,N_23301,N_23368);
or U23671 (N_23671,N_23133,N_23148);
or U23672 (N_23672,N_23252,N_23273);
nand U23673 (N_23673,N_23448,N_23267);
nor U23674 (N_23674,N_23442,N_23048);
nor U23675 (N_23675,N_23160,N_23233);
nand U23676 (N_23676,N_23446,N_23307);
xnor U23677 (N_23677,N_23116,N_23385);
xnor U23678 (N_23678,N_23005,N_23036);
and U23679 (N_23679,N_23388,N_23495);
and U23680 (N_23680,N_23433,N_23184);
or U23681 (N_23681,N_23369,N_23360);
xor U23682 (N_23682,N_23419,N_23113);
or U23683 (N_23683,N_23220,N_23088);
xnor U23684 (N_23684,N_23276,N_23137);
or U23685 (N_23685,N_23283,N_23406);
nand U23686 (N_23686,N_23098,N_23143);
or U23687 (N_23687,N_23240,N_23453);
or U23688 (N_23688,N_23367,N_23189);
xnor U23689 (N_23689,N_23068,N_23141);
nand U23690 (N_23690,N_23039,N_23324);
or U23691 (N_23691,N_23214,N_23166);
nand U23692 (N_23692,N_23292,N_23139);
xor U23693 (N_23693,N_23251,N_23494);
xnor U23694 (N_23694,N_23243,N_23236);
nor U23695 (N_23695,N_23209,N_23482);
or U23696 (N_23696,N_23074,N_23089);
and U23697 (N_23697,N_23217,N_23211);
or U23698 (N_23698,N_23101,N_23325);
nor U23699 (N_23699,N_23110,N_23318);
or U23700 (N_23700,N_23079,N_23493);
nand U23701 (N_23701,N_23332,N_23414);
and U23702 (N_23702,N_23258,N_23131);
nand U23703 (N_23703,N_23303,N_23004);
and U23704 (N_23704,N_23075,N_23398);
nor U23705 (N_23705,N_23327,N_23114);
and U23706 (N_23706,N_23443,N_23057);
nor U23707 (N_23707,N_23118,N_23498);
or U23708 (N_23708,N_23333,N_23489);
or U23709 (N_23709,N_23485,N_23337);
or U23710 (N_23710,N_23284,N_23253);
xor U23711 (N_23711,N_23313,N_23173);
nand U23712 (N_23712,N_23132,N_23060);
and U23713 (N_23713,N_23169,N_23225);
nor U23714 (N_23714,N_23185,N_23376);
xor U23715 (N_23715,N_23191,N_23164);
xor U23716 (N_23716,N_23338,N_23146);
nor U23717 (N_23717,N_23486,N_23451);
nor U23718 (N_23718,N_23051,N_23235);
and U23719 (N_23719,N_23375,N_23237);
nand U23720 (N_23720,N_23491,N_23093);
and U23721 (N_23721,N_23064,N_23260);
and U23722 (N_23722,N_23182,N_23153);
xor U23723 (N_23723,N_23056,N_23115);
and U23724 (N_23724,N_23450,N_23219);
nor U23725 (N_23725,N_23436,N_23397);
xor U23726 (N_23726,N_23024,N_23195);
or U23727 (N_23727,N_23487,N_23403);
or U23728 (N_23728,N_23106,N_23157);
or U23729 (N_23729,N_23084,N_23188);
xor U23730 (N_23730,N_23218,N_23065);
nor U23731 (N_23731,N_23119,N_23050);
or U23732 (N_23732,N_23099,N_23347);
xnor U23733 (N_23733,N_23305,N_23455);
and U23734 (N_23734,N_23032,N_23070);
and U23735 (N_23735,N_23124,N_23310);
xor U23736 (N_23736,N_23412,N_23238);
nor U23737 (N_23737,N_23054,N_23145);
xnor U23738 (N_23738,N_23172,N_23230);
nor U23739 (N_23739,N_23323,N_23205);
nor U23740 (N_23740,N_23477,N_23080);
and U23741 (N_23741,N_23308,N_23052);
and U23742 (N_23742,N_23167,N_23254);
and U23743 (N_23743,N_23152,N_23457);
xnor U23744 (N_23744,N_23259,N_23155);
xnor U23745 (N_23745,N_23159,N_23247);
or U23746 (N_23746,N_23270,N_23161);
and U23747 (N_23747,N_23438,N_23263);
xor U23748 (N_23748,N_23090,N_23242);
or U23749 (N_23749,N_23287,N_23363);
xnor U23750 (N_23750,N_23032,N_23035);
or U23751 (N_23751,N_23179,N_23499);
or U23752 (N_23752,N_23466,N_23333);
or U23753 (N_23753,N_23171,N_23303);
nor U23754 (N_23754,N_23183,N_23360);
and U23755 (N_23755,N_23314,N_23297);
or U23756 (N_23756,N_23010,N_23073);
and U23757 (N_23757,N_23357,N_23165);
nand U23758 (N_23758,N_23373,N_23082);
or U23759 (N_23759,N_23309,N_23461);
nand U23760 (N_23760,N_23304,N_23060);
xnor U23761 (N_23761,N_23189,N_23091);
or U23762 (N_23762,N_23211,N_23417);
xor U23763 (N_23763,N_23468,N_23264);
nand U23764 (N_23764,N_23235,N_23222);
xnor U23765 (N_23765,N_23479,N_23084);
xor U23766 (N_23766,N_23244,N_23242);
or U23767 (N_23767,N_23379,N_23173);
or U23768 (N_23768,N_23445,N_23159);
nand U23769 (N_23769,N_23329,N_23425);
and U23770 (N_23770,N_23218,N_23316);
or U23771 (N_23771,N_23314,N_23480);
nand U23772 (N_23772,N_23446,N_23195);
nand U23773 (N_23773,N_23265,N_23275);
nor U23774 (N_23774,N_23288,N_23099);
nor U23775 (N_23775,N_23497,N_23030);
or U23776 (N_23776,N_23128,N_23219);
and U23777 (N_23777,N_23017,N_23060);
nor U23778 (N_23778,N_23051,N_23079);
xnor U23779 (N_23779,N_23060,N_23203);
nor U23780 (N_23780,N_23060,N_23143);
or U23781 (N_23781,N_23067,N_23039);
nor U23782 (N_23782,N_23094,N_23238);
or U23783 (N_23783,N_23001,N_23080);
or U23784 (N_23784,N_23025,N_23391);
nand U23785 (N_23785,N_23123,N_23137);
or U23786 (N_23786,N_23328,N_23436);
and U23787 (N_23787,N_23446,N_23247);
and U23788 (N_23788,N_23310,N_23221);
xor U23789 (N_23789,N_23338,N_23317);
xor U23790 (N_23790,N_23240,N_23051);
xnor U23791 (N_23791,N_23263,N_23282);
xor U23792 (N_23792,N_23240,N_23069);
xnor U23793 (N_23793,N_23457,N_23160);
and U23794 (N_23794,N_23059,N_23433);
or U23795 (N_23795,N_23068,N_23051);
nor U23796 (N_23796,N_23403,N_23083);
xnor U23797 (N_23797,N_23038,N_23169);
nor U23798 (N_23798,N_23484,N_23415);
nor U23799 (N_23799,N_23475,N_23106);
and U23800 (N_23800,N_23453,N_23168);
nor U23801 (N_23801,N_23287,N_23010);
nor U23802 (N_23802,N_23405,N_23219);
xor U23803 (N_23803,N_23244,N_23173);
nand U23804 (N_23804,N_23484,N_23241);
nand U23805 (N_23805,N_23148,N_23423);
and U23806 (N_23806,N_23064,N_23281);
nand U23807 (N_23807,N_23102,N_23119);
xor U23808 (N_23808,N_23090,N_23302);
and U23809 (N_23809,N_23315,N_23127);
nand U23810 (N_23810,N_23206,N_23401);
and U23811 (N_23811,N_23123,N_23284);
nand U23812 (N_23812,N_23272,N_23198);
nand U23813 (N_23813,N_23441,N_23275);
and U23814 (N_23814,N_23142,N_23182);
nor U23815 (N_23815,N_23193,N_23073);
nand U23816 (N_23816,N_23267,N_23161);
xor U23817 (N_23817,N_23322,N_23456);
nor U23818 (N_23818,N_23441,N_23305);
and U23819 (N_23819,N_23373,N_23441);
and U23820 (N_23820,N_23114,N_23422);
and U23821 (N_23821,N_23326,N_23119);
nand U23822 (N_23822,N_23434,N_23375);
xnor U23823 (N_23823,N_23344,N_23356);
xor U23824 (N_23824,N_23174,N_23097);
nand U23825 (N_23825,N_23050,N_23150);
nand U23826 (N_23826,N_23074,N_23143);
nand U23827 (N_23827,N_23022,N_23119);
and U23828 (N_23828,N_23296,N_23098);
nor U23829 (N_23829,N_23398,N_23332);
xnor U23830 (N_23830,N_23169,N_23322);
or U23831 (N_23831,N_23369,N_23414);
nand U23832 (N_23832,N_23168,N_23049);
nand U23833 (N_23833,N_23368,N_23447);
nand U23834 (N_23834,N_23244,N_23459);
xnor U23835 (N_23835,N_23391,N_23170);
nand U23836 (N_23836,N_23025,N_23366);
xnor U23837 (N_23837,N_23109,N_23082);
xnor U23838 (N_23838,N_23484,N_23178);
nand U23839 (N_23839,N_23014,N_23473);
and U23840 (N_23840,N_23264,N_23230);
or U23841 (N_23841,N_23445,N_23429);
nand U23842 (N_23842,N_23328,N_23456);
nand U23843 (N_23843,N_23059,N_23146);
xor U23844 (N_23844,N_23361,N_23318);
or U23845 (N_23845,N_23178,N_23171);
or U23846 (N_23846,N_23456,N_23164);
or U23847 (N_23847,N_23007,N_23212);
and U23848 (N_23848,N_23160,N_23328);
nor U23849 (N_23849,N_23436,N_23267);
nor U23850 (N_23850,N_23072,N_23406);
xnor U23851 (N_23851,N_23010,N_23263);
nor U23852 (N_23852,N_23298,N_23014);
nor U23853 (N_23853,N_23326,N_23159);
xnor U23854 (N_23854,N_23047,N_23074);
nand U23855 (N_23855,N_23461,N_23082);
nor U23856 (N_23856,N_23301,N_23213);
or U23857 (N_23857,N_23008,N_23191);
nand U23858 (N_23858,N_23254,N_23050);
xor U23859 (N_23859,N_23490,N_23152);
and U23860 (N_23860,N_23358,N_23184);
or U23861 (N_23861,N_23293,N_23383);
nor U23862 (N_23862,N_23045,N_23469);
nand U23863 (N_23863,N_23175,N_23000);
or U23864 (N_23864,N_23464,N_23429);
nand U23865 (N_23865,N_23030,N_23244);
or U23866 (N_23866,N_23228,N_23146);
nor U23867 (N_23867,N_23456,N_23075);
or U23868 (N_23868,N_23090,N_23122);
or U23869 (N_23869,N_23391,N_23221);
and U23870 (N_23870,N_23057,N_23407);
nand U23871 (N_23871,N_23075,N_23059);
or U23872 (N_23872,N_23252,N_23331);
xor U23873 (N_23873,N_23388,N_23369);
and U23874 (N_23874,N_23394,N_23461);
nor U23875 (N_23875,N_23206,N_23148);
xnor U23876 (N_23876,N_23491,N_23169);
nand U23877 (N_23877,N_23466,N_23163);
and U23878 (N_23878,N_23317,N_23009);
xnor U23879 (N_23879,N_23190,N_23068);
or U23880 (N_23880,N_23378,N_23172);
xor U23881 (N_23881,N_23150,N_23457);
xor U23882 (N_23882,N_23251,N_23395);
or U23883 (N_23883,N_23107,N_23049);
and U23884 (N_23884,N_23326,N_23466);
nor U23885 (N_23885,N_23052,N_23022);
and U23886 (N_23886,N_23102,N_23249);
xor U23887 (N_23887,N_23425,N_23424);
or U23888 (N_23888,N_23161,N_23378);
or U23889 (N_23889,N_23045,N_23260);
and U23890 (N_23890,N_23494,N_23096);
and U23891 (N_23891,N_23146,N_23396);
or U23892 (N_23892,N_23354,N_23457);
or U23893 (N_23893,N_23008,N_23184);
nand U23894 (N_23894,N_23268,N_23112);
xor U23895 (N_23895,N_23401,N_23412);
nor U23896 (N_23896,N_23043,N_23259);
nand U23897 (N_23897,N_23014,N_23177);
xor U23898 (N_23898,N_23326,N_23231);
xnor U23899 (N_23899,N_23432,N_23099);
nand U23900 (N_23900,N_23276,N_23330);
nor U23901 (N_23901,N_23037,N_23056);
nor U23902 (N_23902,N_23152,N_23151);
nor U23903 (N_23903,N_23144,N_23179);
nor U23904 (N_23904,N_23038,N_23463);
xnor U23905 (N_23905,N_23217,N_23256);
and U23906 (N_23906,N_23484,N_23030);
and U23907 (N_23907,N_23343,N_23441);
and U23908 (N_23908,N_23047,N_23475);
xnor U23909 (N_23909,N_23111,N_23421);
or U23910 (N_23910,N_23296,N_23355);
nand U23911 (N_23911,N_23213,N_23236);
nor U23912 (N_23912,N_23160,N_23334);
or U23913 (N_23913,N_23279,N_23133);
xor U23914 (N_23914,N_23275,N_23037);
nor U23915 (N_23915,N_23197,N_23406);
or U23916 (N_23916,N_23135,N_23449);
nand U23917 (N_23917,N_23351,N_23140);
nand U23918 (N_23918,N_23305,N_23116);
and U23919 (N_23919,N_23217,N_23324);
xnor U23920 (N_23920,N_23236,N_23237);
or U23921 (N_23921,N_23015,N_23369);
nand U23922 (N_23922,N_23448,N_23098);
nand U23923 (N_23923,N_23423,N_23194);
nand U23924 (N_23924,N_23359,N_23050);
and U23925 (N_23925,N_23237,N_23113);
nand U23926 (N_23926,N_23326,N_23285);
nor U23927 (N_23927,N_23373,N_23428);
xor U23928 (N_23928,N_23334,N_23348);
nor U23929 (N_23929,N_23352,N_23158);
nor U23930 (N_23930,N_23407,N_23425);
and U23931 (N_23931,N_23273,N_23164);
nand U23932 (N_23932,N_23356,N_23177);
or U23933 (N_23933,N_23045,N_23158);
xnor U23934 (N_23934,N_23171,N_23481);
and U23935 (N_23935,N_23212,N_23348);
or U23936 (N_23936,N_23184,N_23103);
or U23937 (N_23937,N_23177,N_23465);
xnor U23938 (N_23938,N_23457,N_23058);
or U23939 (N_23939,N_23397,N_23377);
nor U23940 (N_23940,N_23456,N_23314);
and U23941 (N_23941,N_23344,N_23158);
nor U23942 (N_23942,N_23348,N_23481);
and U23943 (N_23943,N_23307,N_23369);
nand U23944 (N_23944,N_23328,N_23258);
and U23945 (N_23945,N_23285,N_23320);
or U23946 (N_23946,N_23095,N_23290);
nand U23947 (N_23947,N_23240,N_23242);
nor U23948 (N_23948,N_23070,N_23431);
xor U23949 (N_23949,N_23348,N_23346);
nor U23950 (N_23950,N_23341,N_23156);
nand U23951 (N_23951,N_23340,N_23293);
and U23952 (N_23952,N_23263,N_23072);
xnor U23953 (N_23953,N_23059,N_23238);
and U23954 (N_23954,N_23276,N_23225);
nand U23955 (N_23955,N_23124,N_23087);
or U23956 (N_23956,N_23247,N_23228);
or U23957 (N_23957,N_23483,N_23058);
nand U23958 (N_23958,N_23103,N_23337);
and U23959 (N_23959,N_23497,N_23106);
or U23960 (N_23960,N_23310,N_23473);
nand U23961 (N_23961,N_23404,N_23324);
nor U23962 (N_23962,N_23370,N_23074);
xor U23963 (N_23963,N_23086,N_23264);
xnor U23964 (N_23964,N_23344,N_23387);
and U23965 (N_23965,N_23426,N_23319);
nor U23966 (N_23966,N_23074,N_23398);
or U23967 (N_23967,N_23252,N_23334);
and U23968 (N_23968,N_23044,N_23281);
or U23969 (N_23969,N_23283,N_23261);
xor U23970 (N_23970,N_23015,N_23178);
nand U23971 (N_23971,N_23413,N_23085);
nand U23972 (N_23972,N_23348,N_23065);
and U23973 (N_23973,N_23366,N_23147);
and U23974 (N_23974,N_23384,N_23021);
nand U23975 (N_23975,N_23345,N_23280);
and U23976 (N_23976,N_23046,N_23184);
xor U23977 (N_23977,N_23141,N_23012);
nor U23978 (N_23978,N_23414,N_23183);
nand U23979 (N_23979,N_23388,N_23444);
or U23980 (N_23980,N_23309,N_23265);
or U23981 (N_23981,N_23022,N_23009);
nor U23982 (N_23982,N_23083,N_23247);
or U23983 (N_23983,N_23427,N_23495);
and U23984 (N_23984,N_23249,N_23476);
nor U23985 (N_23985,N_23083,N_23105);
and U23986 (N_23986,N_23009,N_23101);
nor U23987 (N_23987,N_23457,N_23208);
xor U23988 (N_23988,N_23114,N_23168);
and U23989 (N_23989,N_23371,N_23354);
and U23990 (N_23990,N_23381,N_23369);
nor U23991 (N_23991,N_23250,N_23386);
nand U23992 (N_23992,N_23478,N_23142);
or U23993 (N_23993,N_23470,N_23384);
xor U23994 (N_23994,N_23304,N_23349);
nor U23995 (N_23995,N_23271,N_23283);
nor U23996 (N_23996,N_23302,N_23314);
nor U23997 (N_23997,N_23048,N_23223);
nand U23998 (N_23998,N_23260,N_23127);
nor U23999 (N_23999,N_23316,N_23351);
nor U24000 (N_24000,N_23729,N_23525);
xnor U24001 (N_24001,N_23573,N_23712);
nand U24002 (N_24002,N_23545,N_23871);
nor U24003 (N_24003,N_23682,N_23521);
nand U24004 (N_24004,N_23651,N_23632);
nand U24005 (N_24005,N_23526,N_23600);
nand U24006 (N_24006,N_23750,N_23793);
nor U24007 (N_24007,N_23946,N_23810);
or U24008 (N_24008,N_23735,N_23790);
or U24009 (N_24009,N_23921,N_23605);
nor U24010 (N_24010,N_23674,N_23599);
nor U24011 (N_24011,N_23547,N_23542);
or U24012 (N_24012,N_23552,N_23699);
and U24013 (N_24013,N_23747,N_23940);
and U24014 (N_24014,N_23658,N_23701);
xnor U24015 (N_24015,N_23813,N_23849);
and U24016 (N_24016,N_23645,N_23638);
nand U24017 (N_24017,N_23837,N_23914);
and U24018 (N_24018,N_23690,N_23930);
xnor U24019 (N_24019,N_23831,N_23528);
and U24020 (N_24020,N_23587,N_23666);
xor U24021 (N_24021,N_23620,N_23913);
or U24022 (N_24022,N_23959,N_23500);
xnor U24023 (N_24023,N_23886,N_23548);
and U24024 (N_24024,N_23621,N_23901);
and U24025 (N_24025,N_23564,N_23502);
xor U24026 (N_24026,N_23675,N_23743);
nand U24027 (N_24027,N_23734,N_23834);
nand U24028 (N_24028,N_23697,N_23873);
nand U24029 (N_24029,N_23535,N_23618);
or U24030 (N_24030,N_23981,N_23724);
or U24031 (N_24031,N_23988,N_23749);
and U24032 (N_24032,N_23577,N_23748);
and U24033 (N_24033,N_23556,N_23820);
xor U24034 (N_24034,N_23640,N_23978);
nor U24035 (N_24035,N_23776,N_23878);
nor U24036 (N_24036,N_23537,N_23727);
nand U24037 (N_24037,N_23877,N_23660);
xor U24038 (N_24038,N_23597,N_23713);
nor U24039 (N_24039,N_23707,N_23818);
xor U24040 (N_24040,N_23719,N_23677);
and U24041 (N_24041,N_23527,N_23962);
and U24042 (N_24042,N_23504,N_23728);
and U24043 (N_24043,N_23562,N_23967);
and U24044 (N_24044,N_23874,N_23770);
nand U24045 (N_24045,N_23875,N_23926);
or U24046 (N_24046,N_23541,N_23514);
nor U24047 (N_24047,N_23842,N_23601);
xor U24048 (N_24048,N_23627,N_23530);
or U24049 (N_24049,N_23783,N_23784);
or U24050 (N_24050,N_23567,N_23952);
xnor U24051 (N_24051,N_23678,N_23864);
or U24052 (N_24052,N_23538,N_23911);
and U24053 (N_24053,N_23669,N_23533);
nor U24054 (N_24054,N_23523,N_23672);
nor U24055 (N_24055,N_23615,N_23668);
nand U24056 (N_24056,N_23565,N_23680);
nand U24057 (N_24057,N_23593,N_23858);
nor U24058 (N_24058,N_23778,N_23970);
or U24059 (N_24059,N_23809,N_23825);
xor U24060 (N_24060,N_23862,N_23614);
and U24061 (N_24061,N_23854,N_23887);
nor U24062 (N_24062,N_23944,N_23559);
or U24063 (N_24063,N_23982,N_23844);
or U24064 (N_24064,N_23591,N_23738);
xor U24065 (N_24065,N_23969,N_23897);
nand U24066 (N_24066,N_23852,N_23780);
nand U24067 (N_24067,N_23625,N_23976);
and U24068 (N_24068,N_23850,N_23839);
xnor U24069 (N_24069,N_23964,N_23995);
and U24070 (N_24070,N_23739,N_23581);
nor U24071 (N_24071,N_23694,N_23884);
nand U24072 (N_24072,N_23639,N_23808);
xnor U24073 (N_24073,N_23608,N_23765);
or U24074 (N_24074,N_23829,N_23665);
or U24075 (N_24075,N_23635,N_23937);
or U24076 (N_24076,N_23974,N_23576);
nand U24077 (N_24077,N_23650,N_23841);
nor U24078 (N_24078,N_23972,N_23741);
nand U24079 (N_24079,N_23890,N_23549);
xnor U24080 (N_24080,N_23791,N_23711);
nand U24081 (N_24081,N_23927,N_23859);
nor U24082 (N_24082,N_23636,N_23762);
and U24083 (N_24083,N_23800,N_23836);
nand U24084 (N_24084,N_23616,N_23756);
nand U24085 (N_24085,N_23832,N_23782);
nor U24086 (N_24086,N_23994,N_23965);
or U24087 (N_24087,N_23943,N_23916);
or U24088 (N_24088,N_23622,N_23888);
nor U24089 (N_24089,N_23506,N_23708);
and U24090 (N_24090,N_23709,N_23997);
nor U24091 (N_24091,N_23814,N_23612);
and U24092 (N_24092,N_23896,N_23522);
or U24093 (N_24093,N_23604,N_23744);
nand U24094 (N_24094,N_23643,N_23806);
nand U24095 (N_24095,N_23657,N_23772);
xnor U24096 (N_24096,N_23934,N_23557);
or U24097 (N_24097,N_23582,N_23554);
nor U24098 (N_24098,N_23603,N_23691);
xnor U24099 (N_24099,N_23835,N_23802);
nand U24100 (N_24100,N_23929,N_23764);
nor U24101 (N_24101,N_23991,N_23613);
nand U24102 (N_24102,N_23945,N_23954);
xnor U24103 (N_24103,N_23531,N_23763);
nand U24104 (N_24104,N_23700,N_23592);
nand U24105 (N_24105,N_23652,N_23579);
nand U24106 (N_24106,N_23955,N_23771);
nand U24107 (N_24107,N_23794,N_23948);
nand U24108 (N_24108,N_23895,N_23575);
or U24109 (N_24109,N_23915,N_23681);
nor U24110 (N_24110,N_23755,N_23684);
xor U24111 (N_24111,N_23910,N_23827);
and U24112 (N_24112,N_23840,N_23520);
and U24113 (N_24113,N_23510,N_23501);
or U24114 (N_24114,N_23870,N_23847);
nand U24115 (N_24115,N_23879,N_23907);
nor U24116 (N_24116,N_23898,N_23769);
nand U24117 (N_24117,N_23893,N_23555);
or U24118 (N_24118,N_23993,N_23958);
nor U24119 (N_24119,N_23824,N_23950);
nor U24120 (N_24120,N_23722,N_23863);
and U24121 (N_24121,N_23866,N_23536);
or U24122 (N_24122,N_23792,N_23922);
nor U24123 (N_24123,N_23761,N_23596);
nor U24124 (N_24124,N_23610,N_23947);
or U24125 (N_24125,N_23716,N_23752);
nor U24126 (N_24126,N_23894,N_23653);
or U24127 (N_24127,N_23892,N_23990);
xor U24128 (N_24128,N_23698,N_23787);
nor U24129 (N_24129,N_23920,N_23688);
xor U24130 (N_24130,N_23925,N_23957);
and U24131 (N_24131,N_23598,N_23773);
xnor U24132 (N_24132,N_23642,N_23797);
and U24133 (N_24133,N_23686,N_23626);
or U24134 (N_24134,N_23634,N_23572);
and U24135 (N_24135,N_23705,N_23905);
or U24136 (N_24136,N_23933,N_23558);
or U24137 (N_24137,N_23515,N_23785);
and U24138 (N_24138,N_23508,N_23662);
nor U24139 (N_24139,N_23936,N_23595);
and U24140 (N_24140,N_23833,N_23606);
nor U24141 (N_24141,N_23623,N_23819);
xnor U24142 (N_24142,N_23754,N_23519);
or U24143 (N_24143,N_23723,N_23805);
nor U24144 (N_24144,N_23774,N_23903);
xor U24145 (N_24145,N_23628,N_23986);
nor U24146 (N_24146,N_23918,N_23811);
and U24147 (N_24147,N_23872,N_23885);
nand U24148 (N_24148,N_23753,N_23857);
or U24149 (N_24149,N_23586,N_23524);
and U24150 (N_24150,N_23851,N_23737);
or U24151 (N_24151,N_23693,N_23987);
nor U24152 (N_24152,N_23985,N_23828);
or U24153 (N_24153,N_23823,N_23876);
nor U24154 (N_24154,N_23912,N_23803);
nand U24155 (N_24155,N_23881,N_23908);
nand U24156 (N_24156,N_23736,N_23798);
or U24157 (N_24157,N_23509,N_23961);
nor U24158 (N_24158,N_23503,N_23584);
xnor U24159 (N_24159,N_23717,N_23731);
or U24160 (N_24160,N_23801,N_23726);
and U24161 (N_24161,N_23989,N_23821);
nor U24162 (N_24162,N_23924,N_23721);
or U24163 (N_24163,N_23617,N_23781);
or U24164 (N_24164,N_23529,N_23845);
or U24165 (N_24165,N_23941,N_23696);
and U24166 (N_24166,N_23786,N_23868);
or U24167 (N_24167,N_23505,N_23629);
and U24168 (N_24168,N_23732,N_23740);
and U24169 (N_24169,N_23544,N_23661);
xnor U24170 (N_24170,N_23715,N_23553);
and U24171 (N_24171,N_23561,N_23746);
nor U24172 (N_24172,N_23664,N_23899);
nor U24173 (N_24173,N_23676,N_23546);
xor U24174 (N_24174,N_23685,N_23683);
and U24175 (N_24175,N_23960,N_23935);
nand U24176 (N_24176,N_23900,N_23853);
and U24177 (N_24177,N_23702,N_23817);
xnor U24178 (N_24178,N_23760,N_23869);
xor U24179 (N_24179,N_23889,N_23775);
or U24180 (N_24180,N_23532,N_23644);
nand U24181 (N_24181,N_23550,N_23882);
nand U24182 (N_24182,N_23963,N_23860);
xnor U24183 (N_24183,N_23580,N_23996);
nand U24184 (N_24184,N_23671,N_23904);
or U24185 (N_24185,N_23861,N_23706);
or U24186 (N_24186,N_23759,N_23966);
and U24187 (N_24187,N_23999,N_23807);
or U24188 (N_24188,N_23909,N_23646);
or U24189 (N_24189,N_23607,N_23689);
nor U24190 (N_24190,N_23880,N_23516);
xnor U24191 (N_24191,N_23932,N_23687);
nand U24192 (N_24192,N_23804,N_23795);
nand U24193 (N_24193,N_23679,N_23518);
xor U24194 (N_24194,N_23939,N_23695);
xor U24195 (N_24195,N_23511,N_23512);
nand U24196 (N_24196,N_23822,N_23758);
nand U24197 (N_24197,N_23766,N_23513);
nand U24198 (N_24198,N_23998,N_23585);
nor U24199 (N_24199,N_23631,N_23594);
xnor U24200 (N_24200,N_23619,N_23830);
and U24201 (N_24201,N_23624,N_23551);
or U24202 (N_24202,N_23971,N_23590);
nand U24203 (N_24203,N_23745,N_23649);
nand U24204 (N_24204,N_23725,N_23566);
and U24205 (N_24205,N_23714,N_23571);
nand U24206 (N_24206,N_23655,N_23980);
nor U24207 (N_24207,N_23578,N_23751);
or U24208 (N_24208,N_23956,N_23883);
and U24209 (N_24209,N_23977,N_23906);
nor U24210 (N_24210,N_23659,N_23949);
and U24211 (N_24211,N_23968,N_23641);
or U24212 (N_24212,N_23923,N_23654);
nand U24213 (N_24213,N_23733,N_23816);
xnor U24214 (N_24214,N_23838,N_23570);
and U24215 (N_24215,N_23942,N_23673);
xnor U24216 (N_24216,N_23789,N_23647);
and U24217 (N_24217,N_23667,N_23633);
or U24218 (N_24218,N_23796,N_23534);
nand U24219 (N_24219,N_23663,N_23779);
nand U24220 (N_24220,N_23902,N_23848);
or U24221 (N_24221,N_23588,N_23951);
nand U24222 (N_24222,N_23979,N_23856);
nor U24223 (N_24223,N_23992,N_23757);
nor U24224 (N_24224,N_23919,N_23574);
nand U24225 (N_24225,N_23855,N_23843);
and U24226 (N_24226,N_23767,N_23742);
and U24227 (N_24227,N_23730,N_23583);
or U24228 (N_24228,N_23589,N_23815);
xor U24229 (N_24229,N_23692,N_23540);
nor U24230 (N_24230,N_23670,N_23768);
nand U24231 (N_24231,N_23637,N_23812);
nor U24232 (N_24232,N_23984,N_23648);
xnor U24233 (N_24233,N_23826,N_23931);
nor U24234 (N_24234,N_23602,N_23867);
and U24235 (N_24235,N_23777,N_23609);
nand U24236 (N_24236,N_23973,N_23569);
and U24237 (N_24237,N_23560,N_23568);
and U24238 (N_24238,N_23953,N_23539);
nand U24239 (N_24239,N_23975,N_23891);
nand U24240 (N_24240,N_23704,N_23563);
nor U24241 (N_24241,N_23865,N_23718);
nor U24242 (N_24242,N_23917,N_23938);
nand U24243 (N_24243,N_23611,N_23928);
nor U24244 (N_24244,N_23720,N_23710);
nor U24245 (N_24245,N_23846,N_23507);
xnor U24246 (N_24246,N_23983,N_23517);
xor U24247 (N_24247,N_23543,N_23656);
or U24248 (N_24248,N_23630,N_23799);
xnor U24249 (N_24249,N_23703,N_23788);
and U24250 (N_24250,N_23602,N_23804);
and U24251 (N_24251,N_23845,N_23587);
nor U24252 (N_24252,N_23589,N_23947);
or U24253 (N_24253,N_23889,N_23673);
and U24254 (N_24254,N_23516,N_23774);
nor U24255 (N_24255,N_23502,N_23583);
and U24256 (N_24256,N_23563,N_23974);
and U24257 (N_24257,N_23810,N_23914);
xnor U24258 (N_24258,N_23579,N_23858);
nor U24259 (N_24259,N_23841,N_23833);
and U24260 (N_24260,N_23786,N_23909);
xnor U24261 (N_24261,N_23968,N_23797);
nand U24262 (N_24262,N_23752,N_23913);
nand U24263 (N_24263,N_23964,N_23525);
nand U24264 (N_24264,N_23516,N_23738);
or U24265 (N_24265,N_23855,N_23953);
or U24266 (N_24266,N_23502,N_23754);
nor U24267 (N_24267,N_23665,N_23897);
nand U24268 (N_24268,N_23907,N_23644);
nor U24269 (N_24269,N_23848,N_23968);
or U24270 (N_24270,N_23892,N_23894);
xnor U24271 (N_24271,N_23611,N_23633);
nand U24272 (N_24272,N_23750,N_23949);
xor U24273 (N_24273,N_23670,N_23610);
nor U24274 (N_24274,N_23718,N_23617);
xnor U24275 (N_24275,N_23875,N_23515);
nor U24276 (N_24276,N_23504,N_23919);
xnor U24277 (N_24277,N_23629,N_23973);
nor U24278 (N_24278,N_23882,N_23549);
nand U24279 (N_24279,N_23686,N_23908);
or U24280 (N_24280,N_23913,N_23697);
xnor U24281 (N_24281,N_23801,N_23828);
nor U24282 (N_24282,N_23574,N_23812);
nand U24283 (N_24283,N_23850,N_23819);
and U24284 (N_24284,N_23572,N_23839);
xnor U24285 (N_24285,N_23614,N_23816);
nor U24286 (N_24286,N_23721,N_23699);
nor U24287 (N_24287,N_23945,N_23760);
nand U24288 (N_24288,N_23886,N_23577);
and U24289 (N_24289,N_23686,N_23804);
or U24290 (N_24290,N_23885,N_23938);
or U24291 (N_24291,N_23545,N_23740);
nor U24292 (N_24292,N_23809,N_23834);
nand U24293 (N_24293,N_23944,N_23797);
or U24294 (N_24294,N_23869,N_23815);
nor U24295 (N_24295,N_23536,N_23687);
and U24296 (N_24296,N_23732,N_23801);
xor U24297 (N_24297,N_23686,N_23827);
and U24298 (N_24298,N_23680,N_23528);
xnor U24299 (N_24299,N_23972,N_23607);
xor U24300 (N_24300,N_23761,N_23663);
nor U24301 (N_24301,N_23577,N_23966);
and U24302 (N_24302,N_23808,N_23976);
and U24303 (N_24303,N_23935,N_23574);
nand U24304 (N_24304,N_23582,N_23845);
or U24305 (N_24305,N_23990,N_23962);
and U24306 (N_24306,N_23850,N_23518);
xnor U24307 (N_24307,N_23731,N_23845);
xor U24308 (N_24308,N_23822,N_23699);
xnor U24309 (N_24309,N_23689,N_23871);
nor U24310 (N_24310,N_23584,N_23658);
or U24311 (N_24311,N_23713,N_23593);
nor U24312 (N_24312,N_23901,N_23549);
or U24313 (N_24313,N_23544,N_23947);
nor U24314 (N_24314,N_23895,N_23961);
xor U24315 (N_24315,N_23687,N_23573);
or U24316 (N_24316,N_23742,N_23567);
or U24317 (N_24317,N_23757,N_23860);
nor U24318 (N_24318,N_23643,N_23944);
and U24319 (N_24319,N_23738,N_23935);
xnor U24320 (N_24320,N_23766,N_23664);
nand U24321 (N_24321,N_23504,N_23552);
xor U24322 (N_24322,N_23519,N_23694);
xor U24323 (N_24323,N_23730,N_23970);
or U24324 (N_24324,N_23919,N_23892);
or U24325 (N_24325,N_23791,N_23717);
xnor U24326 (N_24326,N_23922,N_23737);
nor U24327 (N_24327,N_23559,N_23802);
nand U24328 (N_24328,N_23532,N_23647);
nand U24329 (N_24329,N_23946,N_23571);
xor U24330 (N_24330,N_23644,N_23651);
xor U24331 (N_24331,N_23554,N_23825);
nand U24332 (N_24332,N_23727,N_23811);
xor U24333 (N_24333,N_23683,N_23669);
and U24334 (N_24334,N_23601,N_23917);
and U24335 (N_24335,N_23555,N_23510);
nand U24336 (N_24336,N_23846,N_23899);
or U24337 (N_24337,N_23807,N_23636);
nor U24338 (N_24338,N_23588,N_23943);
xnor U24339 (N_24339,N_23818,N_23817);
or U24340 (N_24340,N_23909,N_23709);
xor U24341 (N_24341,N_23639,N_23776);
or U24342 (N_24342,N_23916,N_23861);
nand U24343 (N_24343,N_23817,N_23689);
xnor U24344 (N_24344,N_23995,N_23913);
or U24345 (N_24345,N_23888,N_23567);
nand U24346 (N_24346,N_23875,N_23823);
nor U24347 (N_24347,N_23763,N_23593);
nand U24348 (N_24348,N_23843,N_23811);
xnor U24349 (N_24349,N_23547,N_23568);
and U24350 (N_24350,N_23693,N_23772);
or U24351 (N_24351,N_23622,N_23664);
xor U24352 (N_24352,N_23542,N_23800);
or U24353 (N_24353,N_23612,N_23541);
and U24354 (N_24354,N_23998,N_23795);
nor U24355 (N_24355,N_23581,N_23997);
and U24356 (N_24356,N_23747,N_23663);
or U24357 (N_24357,N_23878,N_23696);
or U24358 (N_24358,N_23596,N_23668);
xnor U24359 (N_24359,N_23676,N_23521);
nor U24360 (N_24360,N_23537,N_23774);
and U24361 (N_24361,N_23751,N_23635);
nand U24362 (N_24362,N_23621,N_23674);
nor U24363 (N_24363,N_23936,N_23530);
nand U24364 (N_24364,N_23786,N_23699);
xor U24365 (N_24365,N_23671,N_23663);
xor U24366 (N_24366,N_23738,N_23836);
nor U24367 (N_24367,N_23832,N_23584);
nor U24368 (N_24368,N_23669,N_23801);
xnor U24369 (N_24369,N_23914,N_23660);
xor U24370 (N_24370,N_23794,N_23847);
and U24371 (N_24371,N_23705,N_23897);
xnor U24372 (N_24372,N_23812,N_23925);
xor U24373 (N_24373,N_23649,N_23705);
xnor U24374 (N_24374,N_23807,N_23693);
nor U24375 (N_24375,N_23605,N_23907);
and U24376 (N_24376,N_23874,N_23546);
nor U24377 (N_24377,N_23558,N_23589);
xnor U24378 (N_24378,N_23583,N_23601);
or U24379 (N_24379,N_23570,N_23946);
and U24380 (N_24380,N_23526,N_23562);
and U24381 (N_24381,N_23681,N_23648);
nand U24382 (N_24382,N_23779,N_23747);
or U24383 (N_24383,N_23515,N_23567);
xor U24384 (N_24384,N_23703,N_23895);
nor U24385 (N_24385,N_23968,N_23638);
nand U24386 (N_24386,N_23942,N_23741);
nand U24387 (N_24387,N_23791,N_23745);
xnor U24388 (N_24388,N_23703,N_23614);
nor U24389 (N_24389,N_23643,N_23715);
or U24390 (N_24390,N_23661,N_23930);
and U24391 (N_24391,N_23511,N_23826);
nor U24392 (N_24392,N_23535,N_23630);
and U24393 (N_24393,N_23504,N_23609);
xor U24394 (N_24394,N_23824,N_23745);
and U24395 (N_24395,N_23871,N_23573);
nor U24396 (N_24396,N_23898,N_23512);
and U24397 (N_24397,N_23699,N_23842);
and U24398 (N_24398,N_23916,N_23526);
and U24399 (N_24399,N_23964,N_23822);
xor U24400 (N_24400,N_23537,N_23912);
nand U24401 (N_24401,N_23865,N_23775);
nor U24402 (N_24402,N_23989,N_23984);
nor U24403 (N_24403,N_23943,N_23566);
nand U24404 (N_24404,N_23889,N_23580);
xnor U24405 (N_24405,N_23949,N_23960);
nand U24406 (N_24406,N_23905,N_23679);
nor U24407 (N_24407,N_23562,N_23752);
or U24408 (N_24408,N_23961,N_23604);
or U24409 (N_24409,N_23594,N_23635);
nor U24410 (N_24410,N_23841,N_23958);
and U24411 (N_24411,N_23553,N_23866);
nand U24412 (N_24412,N_23936,N_23522);
xor U24413 (N_24413,N_23617,N_23892);
and U24414 (N_24414,N_23676,N_23584);
nor U24415 (N_24415,N_23680,N_23909);
nand U24416 (N_24416,N_23548,N_23709);
nand U24417 (N_24417,N_23596,N_23601);
and U24418 (N_24418,N_23568,N_23932);
xor U24419 (N_24419,N_23562,N_23845);
xor U24420 (N_24420,N_23749,N_23720);
xnor U24421 (N_24421,N_23853,N_23650);
nand U24422 (N_24422,N_23937,N_23777);
and U24423 (N_24423,N_23833,N_23571);
and U24424 (N_24424,N_23817,N_23779);
nand U24425 (N_24425,N_23807,N_23644);
or U24426 (N_24426,N_23504,N_23927);
nand U24427 (N_24427,N_23851,N_23889);
or U24428 (N_24428,N_23944,N_23714);
xnor U24429 (N_24429,N_23546,N_23581);
nor U24430 (N_24430,N_23963,N_23892);
or U24431 (N_24431,N_23578,N_23772);
nand U24432 (N_24432,N_23736,N_23782);
nand U24433 (N_24433,N_23682,N_23565);
or U24434 (N_24434,N_23802,N_23984);
and U24435 (N_24435,N_23622,N_23885);
nor U24436 (N_24436,N_23752,N_23883);
nor U24437 (N_24437,N_23511,N_23620);
or U24438 (N_24438,N_23926,N_23572);
or U24439 (N_24439,N_23716,N_23648);
nand U24440 (N_24440,N_23786,N_23666);
or U24441 (N_24441,N_23919,N_23664);
nand U24442 (N_24442,N_23750,N_23928);
nor U24443 (N_24443,N_23893,N_23726);
or U24444 (N_24444,N_23656,N_23982);
nand U24445 (N_24445,N_23617,N_23934);
xor U24446 (N_24446,N_23976,N_23610);
nand U24447 (N_24447,N_23933,N_23751);
and U24448 (N_24448,N_23822,N_23716);
nor U24449 (N_24449,N_23790,N_23780);
nand U24450 (N_24450,N_23667,N_23752);
and U24451 (N_24451,N_23828,N_23569);
xnor U24452 (N_24452,N_23628,N_23575);
nand U24453 (N_24453,N_23937,N_23978);
and U24454 (N_24454,N_23671,N_23816);
xnor U24455 (N_24455,N_23767,N_23641);
and U24456 (N_24456,N_23724,N_23603);
and U24457 (N_24457,N_23986,N_23501);
and U24458 (N_24458,N_23977,N_23547);
nor U24459 (N_24459,N_23662,N_23652);
nand U24460 (N_24460,N_23924,N_23603);
xor U24461 (N_24461,N_23993,N_23616);
nor U24462 (N_24462,N_23786,N_23799);
xnor U24463 (N_24463,N_23596,N_23544);
or U24464 (N_24464,N_23869,N_23713);
nand U24465 (N_24465,N_23857,N_23615);
nor U24466 (N_24466,N_23898,N_23966);
nand U24467 (N_24467,N_23585,N_23680);
and U24468 (N_24468,N_23869,N_23894);
xor U24469 (N_24469,N_23884,N_23678);
and U24470 (N_24470,N_23647,N_23686);
and U24471 (N_24471,N_23671,N_23980);
xor U24472 (N_24472,N_23821,N_23735);
xnor U24473 (N_24473,N_23537,N_23566);
nor U24474 (N_24474,N_23921,N_23661);
nand U24475 (N_24475,N_23511,N_23980);
nand U24476 (N_24476,N_23609,N_23533);
nor U24477 (N_24477,N_23537,N_23628);
nand U24478 (N_24478,N_23609,N_23946);
xnor U24479 (N_24479,N_23963,N_23551);
or U24480 (N_24480,N_23842,N_23551);
or U24481 (N_24481,N_23941,N_23955);
nor U24482 (N_24482,N_23917,N_23592);
nand U24483 (N_24483,N_23948,N_23965);
and U24484 (N_24484,N_23671,N_23983);
nor U24485 (N_24485,N_23987,N_23647);
and U24486 (N_24486,N_23654,N_23704);
and U24487 (N_24487,N_23506,N_23680);
or U24488 (N_24488,N_23905,N_23792);
xor U24489 (N_24489,N_23599,N_23867);
and U24490 (N_24490,N_23786,N_23825);
nand U24491 (N_24491,N_23730,N_23966);
xnor U24492 (N_24492,N_23618,N_23933);
xnor U24493 (N_24493,N_23855,N_23556);
nand U24494 (N_24494,N_23877,N_23924);
xor U24495 (N_24495,N_23630,N_23876);
nand U24496 (N_24496,N_23879,N_23967);
nand U24497 (N_24497,N_23722,N_23834);
nand U24498 (N_24498,N_23746,N_23536);
or U24499 (N_24499,N_23707,N_23536);
or U24500 (N_24500,N_24400,N_24220);
xor U24501 (N_24501,N_24321,N_24326);
nand U24502 (N_24502,N_24248,N_24465);
or U24503 (N_24503,N_24215,N_24475);
xor U24504 (N_24504,N_24271,N_24409);
and U24505 (N_24505,N_24083,N_24257);
nor U24506 (N_24506,N_24340,N_24316);
xnor U24507 (N_24507,N_24158,N_24377);
xor U24508 (N_24508,N_24082,N_24286);
nand U24509 (N_24509,N_24206,N_24021);
nor U24510 (N_24510,N_24254,N_24109);
or U24511 (N_24511,N_24136,N_24490);
nor U24512 (N_24512,N_24107,N_24236);
xor U24513 (N_24513,N_24470,N_24046);
xor U24514 (N_24514,N_24239,N_24094);
and U24515 (N_24515,N_24007,N_24250);
nand U24516 (N_24516,N_24054,N_24324);
and U24517 (N_24517,N_24131,N_24277);
nor U24518 (N_24518,N_24259,N_24114);
nor U24519 (N_24519,N_24414,N_24452);
or U24520 (N_24520,N_24485,N_24432);
and U24521 (N_24521,N_24451,N_24438);
nand U24522 (N_24522,N_24351,N_24121);
nand U24523 (N_24523,N_24193,N_24232);
nand U24524 (N_24524,N_24428,N_24356);
nor U24525 (N_24525,N_24478,N_24405);
or U24526 (N_24526,N_24379,N_24395);
or U24527 (N_24527,N_24137,N_24077);
or U24528 (N_24528,N_24123,N_24088);
xor U24529 (N_24529,N_24383,N_24190);
nor U24530 (N_24530,N_24001,N_24191);
or U24531 (N_24531,N_24081,N_24489);
and U24532 (N_24532,N_24020,N_24102);
nand U24533 (N_24533,N_24210,N_24433);
or U24534 (N_24534,N_24065,N_24181);
or U24535 (N_24535,N_24388,N_24084);
or U24536 (N_24536,N_24427,N_24196);
and U24537 (N_24537,N_24174,N_24033);
nor U24538 (N_24538,N_24365,N_24188);
or U24539 (N_24539,N_24039,N_24437);
or U24540 (N_24540,N_24226,N_24059);
or U24541 (N_24541,N_24079,N_24462);
nor U24542 (N_24542,N_24179,N_24178);
nor U24543 (N_24543,N_24278,N_24342);
or U24544 (N_24544,N_24253,N_24036);
nor U24545 (N_24545,N_24175,N_24423);
and U24546 (N_24546,N_24366,N_24052);
nor U24547 (N_24547,N_24412,N_24314);
and U24548 (N_24548,N_24173,N_24029);
nor U24549 (N_24549,N_24463,N_24170);
or U24550 (N_24550,N_24334,N_24195);
nor U24551 (N_24551,N_24197,N_24481);
or U24552 (N_24552,N_24087,N_24375);
xnor U24553 (N_24553,N_24073,N_24417);
and U24554 (N_24554,N_24296,N_24207);
xor U24555 (N_24555,N_24246,N_24142);
and U24556 (N_24556,N_24143,N_24429);
nor U24557 (N_24557,N_24078,N_24013);
nor U24558 (N_24558,N_24076,N_24219);
nand U24559 (N_24559,N_24002,N_24203);
xnor U24560 (N_24560,N_24223,N_24294);
nand U24561 (N_24561,N_24454,N_24180);
nor U24562 (N_24562,N_24224,N_24100);
nand U24563 (N_24563,N_24252,N_24445);
xor U24564 (N_24564,N_24370,N_24066);
xnor U24565 (N_24565,N_24146,N_24242);
nor U24566 (N_24566,N_24298,N_24488);
or U24567 (N_24567,N_24497,N_24049);
nand U24568 (N_24568,N_24213,N_24315);
and U24569 (N_24569,N_24221,N_24095);
and U24570 (N_24570,N_24310,N_24149);
nor U24571 (N_24571,N_24355,N_24362);
nor U24572 (N_24572,N_24004,N_24291);
or U24573 (N_24573,N_24282,N_24055);
xnor U24574 (N_24574,N_24037,N_24098);
nor U24575 (N_24575,N_24041,N_24110);
xnor U24576 (N_24576,N_24067,N_24408);
or U24577 (N_24577,N_24318,N_24230);
xnor U24578 (N_24578,N_24118,N_24208);
nand U24579 (N_24579,N_24165,N_24374);
xnor U24580 (N_24580,N_24487,N_24168);
nand U24581 (N_24581,N_24272,N_24290);
xor U24582 (N_24582,N_24402,N_24430);
and U24583 (N_24583,N_24369,N_24053);
xnor U24584 (N_24584,N_24472,N_24458);
xor U24585 (N_24585,N_24337,N_24456);
nand U24586 (N_24586,N_24008,N_24038);
or U24587 (N_24587,N_24192,N_24161);
or U24588 (N_24588,N_24348,N_24391);
nor U24589 (N_24589,N_24245,N_24435);
nand U24590 (N_24590,N_24313,N_24032);
nor U24591 (N_24591,N_24350,N_24453);
xor U24592 (N_24592,N_24325,N_24167);
nor U24593 (N_24593,N_24473,N_24422);
xnor U24594 (N_24594,N_24235,N_24205);
nor U24595 (N_24595,N_24460,N_24115);
and U24596 (N_24596,N_24469,N_24225);
and U24597 (N_24597,N_24249,N_24071);
xnor U24598 (N_24598,N_24394,N_24096);
xor U24599 (N_24599,N_24306,N_24336);
nand U24600 (N_24600,N_24025,N_24070);
or U24601 (N_24601,N_24390,N_24166);
and U24602 (N_24602,N_24127,N_24012);
nor U24603 (N_24603,N_24339,N_24101);
xor U24604 (N_24604,N_24468,N_24283);
and U24605 (N_24605,N_24153,N_24119);
xnor U24606 (N_24606,N_24163,N_24048);
nand U24607 (N_24607,N_24256,N_24238);
or U24608 (N_24608,N_24479,N_24217);
xnor U24609 (N_24609,N_24367,N_24464);
and U24610 (N_24610,N_24014,N_24466);
nor U24611 (N_24611,N_24156,N_24421);
and U24612 (N_24612,N_24177,N_24035);
and U24613 (N_24613,N_24028,N_24134);
or U24614 (N_24614,N_24393,N_24474);
or U24615 (N_24615,N_24295,N_24425);
nand U24616 (N_24616,N_24103,N_24263);
xnor U24617 (N_24617,N_24016,N_24361);
nor U24618 (N_24618,N_24439,N_24467);
or U24619 (N_24619,N_24011,N_24386);
or U24620 (N_24620,N_24043,N_24284);
and U24621 (N_24621,N_24234,N_24368);
or U24622 (N_24622,N_24328,N_24147);
nor U24623 (N_24623,N_24116,N_24338);
nand U24624 (N_24624,N_24495,N_24183);
xor U24625 (N_24625,N_24269,N_24128);
and U24626 (N_24626,N_24288,N_24214);
nor U24627 (N_24627,N_24381,N_24132);
nor U24628 (N_24628,N_24061,N_24104);
and U24629 (N_24629,N_24420,N_24304);
or U24630 (N_24630,N_24057,N_24126);
xor U24631 (N_24631,N_24093,N_24212);
nand U24632 (N_24632,N_24130,N_24022);
or U24633 (N_24633,N_24241,N_24292);
xnor U24634 (N_24634,N_24152,N_24410);
or U24635 (N_24635,N_24397,N_24160);
xor U24636 (N_24636,N_24281,N_24371);
or U24637 (N_24637,N_24017,N_24133);
and U24638 (N_24638,N_24260,N_24023);
nand U24639 (N_24639,N_24330,N_24005);
xor U24640 (N_24640,N_24446,N_24018);
nor U24641 (N_24641,N_24332,N_24113);
or U24642 (N_24642,N_24448,N_24498);
nand U24643 (N_24643,N_24124,N_24068);
nor U24644 (N_24644,N_24006,N_24044);
and U24645 (N_24645,N_24247,N_24047);
nor U24646 (N_24646,N_24138,N_24092);
xnor U24647 (N_24647,N_24255,N_24237);
xor U24648 (N_24648,N_24396,N_24144);
and U24649 (N_24649,N_24251,N_24185);
and U24650 (N_24650,N_24494,N_24411);
and U24651 (N_24651,N_24003,N_24484);
nand U24652 (N_24652,N_24015,N_24399);
nand U24653 (N_24653,N_24389,N_24301);
and U24654 (N_24654,N_24483,N_24285);
or U24655 (N_24655,N_24346,N_24154);
and U24656 (N_24656,N_24042,N_24135);
and U24657 (N_24657,N_24204,N_24069);
and U24658 (N_24658,N_24216,N_24162);
xnor U24659 (N_24659,N_24099,N_24085);
nand U24660 (N_24660,N_24312,N_24140);
nor U24661 (N_24661,N_24299,N_24373);
and U24662 (N_24662,N_24406,N_24447);
or U24663 (N_24663,N_24145,N_24151);
nor U24664 (N_24664,N_24496,N_24129);
nor U24665 (N_24665,N_24125,N_24352);
or U24666 (N_24666,N_24027,N_24222);
and U24667 (N_24667,N_24000,N_24074);
nor U24668 (N_24668,N_24331,N_24198);
nor U24669 (N_24669,N_24063,N_24171);
xor U24670 (N_24670,N_24303,N_24407);
and U24671 (N_24671,N_24058,N_24097);
or U24672 (N_24672,N_24380,N_24040);
nand U24673 (N_24673,N_24477,N_24106);
nand U24674 (N_24674,N_24056,N_24026);
and U24675 (N_24675,N_24268,N_24218);
or U24676 (N_24676,N_24276,N_24072);
nor U24677 (N_24677,N_24457,N_24364);
and U24678 (N_24678,N_24434,N_24385);
xor U24679 (N_24679,N_24262,N_24289);
nor U24680 (N_24680,N_24442,N_24243);
xnor U24681 (N_24681,N_24075,N_24319);
nand U24682 (N_24682,N_24019,N_24335);
or U24683 (N_24683,N_24302,N_24010);
nand U24684 (N_24684,N_24347,N_24333);
or U24685 (N_24685,N_24117,N_24461);
nand U24686 (N_24686,N_24086,N_24482);
xnor U24687 (N_24687,N_24492,N_24105);
or U24688 (N_24688,N_24436,N_24392);
or U24689 (N_24689,N_24164,N_24349);
or U24690 (N_24690,N_24264,N_24201);
xor U24691 (N_24691,N_24363,N_24440);
nand U24692 (N_24692,N_24297,N_24341);
and U24693 (N_24693,N_24186,N_24089);
or U24694 (N_24694,N_24307,N_24266);
and U24695 (N_24695,N_24441,N_24202);
xor U24696 (N_24696,N_24279,N_24491);
nand U24697 (N_24697,N_24287,N_24357);
and U24698 (N_24698,N_24444,N_24293);
or U24699 (N_24699,N_24155,N_24176);
nand U24700 (N_24700,N_24024,N_24051);
nor U24701 (N_24701,N_24270,N_24141);
xor U24702 (N_24702,N_24353,N_24240);
nor U24703 (N_24703,N_24354,N_24231);
nand U24704 (N_24704,N_24122,N_24211);
nor U24705 (N_24705,N_24309,N_24187);
nor U24706 (N_24706,N_24359,N_24034);
nand U24707 (N_24707,N_24182,N_24060);
and U24708 (N_24708,N_24227,N_24031);
nand U24709 (N_24709,N_24376,N_24273);
nor U24710 (N_24710,N_24344,N_24418);
and U24711 (N_24711,N_24387,N_24476);
and U24712 (N_24712,N_24317,N_24449);
and U24713 (N_24713,N_24120,N_24308);
nor U24714 (N_24714,N_24320,N_24300);
nor U24715 (N_24715,N_24382,N_24343);
and U24716 (N_24716,N_24413,N_24009);
or U24717 (N_24717,N_24189,N_24200);
or U24718 (N_24718,N_24045,N_24148);
and U24719 (N_24719,N_24030,N_24265);
nand U24720 (N_24720,N_24431,N_24384);
or U24721 (N_24721,N_24244,N_24345);
nand U24722 (N_24722,N_24372,N_24139);
or U24723 (N_24723,N_24112,N_24401);
nand U24724 (N_24724,N_24329,N_24459);
nor U24725 (N_24725,N_24493,N_24261);
or U24726 (N_24726,N_24280,N_24194);
and U24727 (N_24727,N_24424,N_24228);
nor U24728 (N_24728,N_24499,N_24480);
and U24729 (N_24729,N_24311,N_24209);
and U24730 (N_24730,N_24169,N_24090);
and U24731 (N_24731,N_24111,N_24450);
and U24732 (N_24732,N_24275,N_24184);
and U24733 (N_24733,N_24404,N_24108);
xnor U24734 (N_24734,N_24426,N_24274);
nand U24735 (N_24735,N_24199,N_24229);
nor U24736 (N_24736,N_24172,N_24415);
nand U24737 (N_24737,N_24233,N_24267);
nor U24738 (N_24738,N_24157,N_24323);
nand U24739 (N_24739,N_24471,N_24091);
nor U24740 (N_24740,N_24416,N_24486);
nand U24741 (N_24741,N_24360,N_24358);
or U24742 (N_24742,N_24443,N_24062);
and U24743 (N_24743,N_24064,N_24378);
nand U24744 (N_24744,N_24258,N_24398);
nor U24745 (N_24745,N_24050,N_24322);
nor U24746 (N_24746,N_24403,N_24159);
nand U24747 (N_24747,N_24419,N_24455);
or U24748 (N_24748,N_24150,N_24305);
or U24749 (N_24749,N_24080,N_24327);
nand U24750 (N_24750,N_24393,N_24183);
and U24751 (N_24751,N_24061,N_24309);
nor U24752 (N_24752,N_24122,N_24020);
nor U24753 (N_24753,N_24108,N_24402);
and U24754 (N_24754,N_24151,N_24362);
nor U24755 (N_24755,N_24360,N_24210);
or U24756 (N_24756,N_24224,N_24427);
nand U24757 (N_24757,N_24373,N_24062);
xnor U24758 (N_24758,N_24428,N_24049);
nand U24759 (N_24759,N_24203,N_24190);
and U24760 (N_24760,N_24071,N_24241);
and U24761 (N_24761,N_24230,N_24393);
or U24762 (N_24762,N_24170,N_24319);
xnor U24763 (N_24763,N_24191,N_24452);
nand U24764 (N_24764,N_24422,N_24210);
nor U24765 (N_24765,N_24332,N_24264);
nor U24766 (N_24766,N_24206,N_24179);
nor U24767 (N_24767,N_24142,N_24458);
nor U24768 (N_24768,N_24424,N_24390);
nor U24769 (N_24769,N_24239,N_24080);
or U24770 (N_24770,N_24427,N_24483);
or U24771 (N_24771,N_24419,N_24410);
and U24772 (N_24772,N_24311,N_24387);
nor U24773 (N_24773,N_24138,N_24210);
and U24774 (N_24774,N_24004,N_24204);
or U24775 (N_24775,N_24042,N_24473);
or U24776 (N_24776,N_24090,N_24121);
nor U24777 (N_24777,N_24316,N_24335);
nand U24778 (N_24778,N_24305,N_24469);
and U24779 (N_24779,N_24440,N_24027);
nand U24780 (N_24780,N_24193,N_24380);
and U24781 (N_24781,N_24003,N_24343);
and U24782 (N_24782,N_24207,N_24490);
nor U24783 (N_24783,N_24059,N_24496);
nand U24784 (N_24784,N_24466,N_24369);
nand U24785 (N_24785,N_24198,N_24340);
and U24786 (N_24786,N_24330,N_24304);
nand U24787 (N_24787,N_24437,N_24446);
nand U24788 (N_24788,N_24381,N_24145);
and U24789 (N_24789,N_24481,N_24265);
or U24790 (N_24790,N_24387,N_24162);
nor U24791 (N_24791,N_24445,N_24217);
nand U24792 (N_24792,N_24204,N_24023);
or U24793 (N_24793,N_24013,N_24047);
nand U24794 (N_24794,N_24173,N_24419);
or U24795 (N_24795,N_24035,N_24025);
nand U24796 (N_24796,N_24078,N_24149);
or U24797 (N_24797,N_24206,N_24190);
nor U24798 (N_24798,N_24047,N_24477);
and U24799 (N_24799,N_24417,N_24282);
nor U24800 (N_24800,N_24489,N_24121);
xor U24801 (N_24801,N_24428,N_24165);
nor U24802 (N_24802,N_24252,N_24310);
or U24803 (N_24803,N_24300,N_24012);
nor U24804 (N_24804,N_24130,N_24118);
xor U24805 (N_24805,N_24009,N_24110);
nand U24806 (N_24806,N_24245,N_24010);
and U24807 (N_24807,N_24372,N_24347);
nor U24808 (N_24808,N_24273,N_24096);
xor U24809 (N_24809,N_24467,N_24218);
nand U24810 (N_24810,N_24200,N_24081);
and U24811 (N_24811,N_24352,N_24346);
xor U24812 (N_24812,N_24135,N_24238);
xor U24813 (N_24813,N_24457,N_24015);
or U24814 (N_24814,N_24439,N_24489);
and U24815 (N_24815,N_24353,N_24459);
xnor U24816 (N_24816,N_24363,N_24457);
xor U24817 (N_24817,N_24288,N_24399);
nor U24818 (N_24818,N_24480,N_24022);
nor U24819 (N_24819,N_24376,N_24343);
nand U24820 (N_24820,N_24459,N_24287);
nand U24821 (N_24821,N_24498,N_24189);
xnor U24822 (N_24822,N_24055,N_24257);
xor U24823 (N_24823,N_24490,N_24046);
nor U24824 (N_24824,N_24449,N_24133);
nor U24825 (N_24825,N_24442,N_24047);
xnor U24826 (N_24826,N_24432,N_24214);
xnor U24827 (N_24827,N_24035,N_24291);
nand U24828 (N_24828,N_24309,N_24283);
nor U24829 (N_24829,N_24101,N_24015);
nor U24830 (N_24830,N_24231,N_24070);
nand U24831 (N_24831,N_24090,N_24164);
nor U24832 (N_24832,N_24071,N_24349);
xnor U24833 (N_24833,N_24358,N_24069);
xor U24834 (N_24834,N_24048,N_24312);
nor U24835 (N_24835,N_24119,N_24227);
or U24836 (N_24836,N_24190,N_24319);
xnor U24837 (N_24837,N_24013,N_24029);
xor U24838 (N_24838,N_24252,N_24266);
or U24839 (N_24839,N_24130,N_24146);
or U24840 (N_24840,N_24206,N_24492);
xor U24841 (N_24841,N_24352,N_24251);
nor U24842 (N_24842,N_24394,N_24058);
or U24843 (N_24843,N_24134,N_24459);
xnor U24844 (N_24844,N_24450,N_24473);
nor U24845 (N_24845,N_24370,N_24307);
or U24846 (N_24846,N_24280,N_24200);
or U24847 (N_24847,N_24305,N_24383);
or U24848 (N_24848,N_24198,N_24016);
xnor U24849 (N_24849,N_24300,N_24145);
and U24850 (N_24850,N_24222,N_24259);
nor U24851 (N_24851,N_24222,N_24446);
nand U24852 (N_24852,N_24016,N_24024);
or U24853 (N_24853,N_24325,N_24010);
nand U24854 (N_24854,N_24272,N_24285);
nand U24855 (N_24855,N_24344,N_24496);
nand U24856 (N_24856,N_24274,N_24408);
nor U24857 (N_24857,N_24154,N_24367);
xnor U24858 (N_24858,N_24198,N_24324);
xor U24859 (N_24859,N_24233,N_24073);
nor U24860 (N_24860,N_24303,N_24158);
xor U24861 (N_24861,N_24231,N_24272);
nor U24862 (N_24862,N_24009,N_24432);
nand U24863 (N_24863,N_24432,N_24334);
or U24864 (N_24864,N_24343,N_24360);
or U24865 (N_24865,N_24347,N_24048);
xor U24866 (N_24866,N_24400,N_24116);
and U24867 (N_24867,N_24098,N_24018);
xnor U24868 (N_24868,N_24164,N_24456);
xnor U24869 (N_24869,N_24262,N_24048);
nand U24870 (N_24870,N_24092,N_24231);
nand U24871 (N_24871,N_24201,N_24402);
xor U24872 (N_24872,N_24426,N_24087);
and U24873 (N_24873,N_24381,N_24267);
nand U24874 (N_24874,N_24343,N_24212);
nor U24875 (N_24875,N_24050,N_24202);
nor U24876 (N_24876,N_24455,N_24279);
nor U24877 (N_24877,N_24330,N_24029);
nand U24878 (N_24878,N_24333,N_24260);
nand U24879 (N_24879,N_24446,N_24300);
nor U24880 (N_24880,N_24128,N_24175);
nor U24881 (N_24881,N_24048,N_24292);
and U24882 (N_24882,N_24013,N_24397);
and U24883 (N_24883,N_24183,N_24416);
nand U24884 (N_24884,N_24274,N_24047);
xor U24885 (N_24885,N_24244,N_24457);
and U24886 (N_24886,N_24114,N_24081);
or U24887 (N_24887,N_24459,N_24074);
xnor U24888 (N_24888,N_24402,N_24377);
xnor U24889 (N_24889,N_24112,N_24047);
and U24890 (N_24890,N_24499,N_24163);
nor U24891 (N_24891,N_24235,N_24490);
xor U24892 (N_24892,N_24245,N_24459);
nand U24893 (N_24893,N_24201,N_24180);
nand U24894 (N_24894,N_24204,N_24080);
xnor U24895 (N_24895,N_24044,N_24232);
nand U24896 (N_24896,N_24481,N_24323);
and U24897 (N_24897,N_24344,N_24000);
nor U24898 (N_24898,N_24318,N_24006);
or U24899 (N_24899,N_24076,N_24135);
nor U24900 (N_24900,N_24272,N_24453);
nand U24901 (N_24901,N_24022,N_24197);
nor U24902 (N_24902,N_24086,N_24420);
nor U24903 (N_24903,N_24357,N_24094);
or U24904 (N_24904,N_24171,N_24424);
nor U24905 (N_24905,N_24327,N_24149);
and U24906 (N_24906,N_24056,N_24073);
or U24907 (N_24907,N_24261,N_24099);
xnor U24908 (N_24908,N_24225,N_24234);
xnor U24909 (N_24909,N_24377,N_24178);
nor U24910 (N_24910,N_24250,N_24400);
or U24911 (N_24911,N_24223,N_24333);
xor U24912 (N_24912,N_24109,N_24393);
or U24913 (N_24913,N_24343,N_24452);
or U24914 (N_24914,N_24015,N_24250);
or U24915 (N_24915,N_24341,N_24090);
nand U24916 (N_24916,N_24455,N_24373);
xor U24917 (N_24917,N_24303,N_24045);
or U24918 (N_24918,N_24289,N_24440);
nand U24919 (N_24919,N_24329,N_24254);
nand U24920 (N_24920,N_24330,N_24160);
xnor U24921 (N_24921,N_24251,N_24326);
and U24922 (N_24922,N_24044,N_24219);
nand U24923 (N_24923,N_24180,N_24326);
nand U24924 (N_24924,N_24134,N_24320);
and U24925 (N_24925,N_24221,N_24410);
and U24926 (N_24926,N_24157,N_24253);
and U24927 (N_24927,N_24371,N_24398);
xnor U24928 (N_24928,N_24465,N_24097);
nand U24929 (N_24929,N_24009,N_24387);
xor U24930 (N_24930,N_24319,N_24250);
xor U24931 (N_24931,N_24051,N_24307);
xnor U24932 (N_24932,N_24496,N_24025);
nand U24933 (N_24933,N_24339,N_24295);
or U24934 (N_24934,N_24329,N_24450);
xor U24935 (N_24935,N_24044,N_24454);
nor U24936 (N_24936,N_24022,N_24170);
nand U24937 (N_24937,N_24362,N_24308);
or U24938 (N_24938,N_24470,N_24137);
and U24939 (N_24939,N_24248,N_24443);
nor U24940 (N_24940,N_24003,N_24048);
xnor U24941 (N_24941,N_24241,N_24411);
and U24942 (N_24942,N_24248,N_24138);
or U24943 (N_24943,N_24357,N_24300);
xnor U24944 (N_24944,N_24046,N_24404);
or U24945 (N_24945,N_24121,N_24173);
nand U24946 (N_24946,N_24048,N_24166);
and U24947 (N_24947,N_24148,N_24164);
or U24948 (N_24948,N_24231,N_24356);
and U24949 (N_24949,N_24266,N_24308);
nand U24950 (N_24950,N_24028,N_24487);
or U24951 (N_24951,N_24132,N_24463);
and U24952 (N_24952,N_24107,N_24049);
nor U24953 (N_24953,N_24308,N_24151);
xnor U24954 (N_24954,N_24352,N_24166);
nand U24955 (N_24955,N_24337,N_24282);
xor U24956 (N_24956,N_24331,N_24269);
xnor U24957 (N_24957,N_24162,N_24340);
and U24958 (N_24958,N_24172,N_24018);
or U24959 (N_24959,N_24054,N_24370);
nor U24960 (N_24960,N_24014,N_24378);
or U24961 (N_24961,N_24013,N_24146);
and U24962 (N_24962,N_24318,N_24408);
nor U24963 (N_24963,N_24432,N_24430);
xor U24964 (N_24964,N_24279,N_24051);
and U24965 (N_24965,N_24140,N_24192);
and U24966 (N_24966,N_24483,N_24310);
or U24967 (N_24967,N_24075,N_24355);
xnor U24968 (N_24968,N_24026,N_24009);
nor U24969 (N_24969,N_24054,N_24129);
or U24970 (N_24970,N_24103,N_24006);
nor U24971 (N_24971,N_24498,N_24343);
or U24972 (N_24972,N_24242,N_24203);
and U24973 (N_24973,N_24344,N_24334);
nand U24974 (N_24974,N_24457,N_24005);
nor U24975 (N_24975,N_24186,N_24057);
nor U24976 (N_24976,N_24023,N_24203);
xnor U24977 (N_24977,N_24334,N_24178);
xor U24978 (N_24978,N_24027,N_24161);
nand U24979 (N_24979,N_24354,N_24159);
nand U24980 (N_24980,N_24453,N_24156);
and U24981 (N_24981,N_24086,N_24240);
and U24982 (N_24982,N_24462,N_24329);
nor U24983 (N_24983,N_24248,N_24330);
and U24984 (N_24984,N_24050,N_24089);
and U24985 (N_24985,N_24149,N_24492);
xnor U24986 (N_24986,N_24126,N_24156);
xnor U24987 (N_24987,N_24133,N_24313);
and U24988 (N_24988,N_24276,N_24349);
and U24989 (N_24989,N_24475,N_24217);
nor U24990 (N_24990,N_24432,N_24057);
or U24991 (N_24991,N_24024,N_24215);
nor U24992 (N_24992,N_24429,N_24489);
xnor U24993 (N_24993,N_24148,N_24135);
nand U24994 (N_24994,N_24293,N_24278);
xnor U24995 (N_24995,N_24024,N_24008);
nand U24996 (N_24996,N_24026,N_24322);
and U24997 (N_24997,N_24327,N_24309);
or U24998 (N_24998,N_24328,N_24249);
xnor U24999 (N_24999,N_24467,N_24280);
nor UO_0 (O_0,N_24718,N_24632);
nor UO_1 (O_1,N_24983,N_24677);
and UO_2 (O_2,N_24848,N_24539);
or UO_3 (O_3,N_24600,N_24523);
xor UO_4 (O_4,N_24574,N_24738);
nor UO_5 (O_5,N_24585,N_24915);
nand UO_6 (O_6,N_24879,N_24587);
nor UO_7 (O_7,N_24912,N_24541);
and UO_8 (O_8,N_24633,N_24979);
and UO_9 (O_9,N_24544,N_24629);
or UO_10 (O_10,N_24615,N_24785);
xnor UO_11 (O_11,N_24681,N_24901);
or UO_12 (O_12,N_24809,N_24531);
or UO_13 (O_13,N_24588,N_24829);
nand UO_14 (O_14,N_24671,N_24898);
and UO_15 (O_15,N_24945,N_24938);
and UO_16 (O_16,N_24869,N_24579);
nand UO_17 (O_17,N_24920,N_24692);
and UO_18 (O_18,N_24576,N_24936);
nor UO_19 (O_19,N_24834,N_24764);
nand UO_20 (O_20,N_24959,N_24552);
nand UO_21 (O_21,N_24926,N_24674);
xnor UO_22 (O_22,N_24769,N_24673);
nor UO_23 (O_23,N_24739,N_24575);
or UO_24 (O_24,N_24737,N_24540);
or UO_25 (O_25,N_24557,N_24950);
nand UO_26 (O_26,N_24561,N_24717);
or UO_27 (O_27,N_24562,N_24756);
and UO_28 (O_28,N_24865,N_24842);
or UO_29 (O_29,N_24986,N_24830);
xor UO_30 (O_30,N_24942,N_24953);
or UO_31 (O_31,N_24981,N_24762);
xnor UO_32 (O_32,N_24644,N_24522);
xor UO_33 (O_33,N_24995,N_24962);
nor UO_34 (O_34,N_24598,N_24690);
nand UO_35 (O_35,N_24759,N_24887);
nand UO_36 (O_36,N_24667,N_24796);
or UO_37 (O_37,N_24768,N_24727);
xnor UO_38 (O_38,N_24560,N_24643);
xnor UO_39 (O_39,N_24777,N_24859);
and UO_40 (O_40,N_24716,N_24812);
xnor UO_41 (O_41,N_24826,N_24696);
and UO_42 (O_42,N_24658,N_24649);
or UO_43 (O_43,N_24925,N_24661);
or UO_44 (O_44,N_24932,N_24614);
nand UO_45 (O_45,N_24928,N_24930);
or UO_46 (O_46,N_24998,N_24849);
and UO_47 (O_47,N_24607,N_24726);
or UO_48 (O_48,N_24967,N_24804);
nor UO_49 (O_49,N_24878,N_24889);
xor UO_50 (O_50,N_24908,N_24518);
nand UO_51 (O_51,N_24511,N_24807);
nor UO_52 (O_52,N_24698,N_24646);
xnor UO_53 (O_53,N_24994,N_24919);
xnor UO_54 (O_54,N_24870,N_24927);
and UO_55 (O_55,N_24874,N_24773);
nand UO_56 (O_56,N_24701,N_24578);
xor UO_57 (O_57,N_24694,N_24987);
and UO_58 (O_58,N_24965,N_24886);
nor UO_59 (O_59,N_24503,N_24907);
nand UO_60 (O_60,N_24728,N_24592);
nor UO_61 (O_61,N_24564,N_24820);
and UO_62 (O_62,N_24894,N_24736);
and UO_63 (O_63,N_24563,N_24982);
nand UO_64 (O_64,N_24897,N_24668);
xor UO_65 (O_65,N_24533,N_24755);
nor UO_66 (O_66,N_24641,N_24631);
and UO_67 (O_67,N_24740,N_24754);
nand UO_68 (O_68,N_24891,N_24570);
nand UO_69 (O_69,N_24850,N_24753);
and UO_70 (O_70,N_24622,N_24551);
xor UO_71 (O_71,N_24628,N_24831);
nor UO_72 (O_72,N_24862,N_24654);
nor UO_73 (O_73,N_24767,N_24731);
xnor UO_74 (O_74,N_24672,N_24597);
or UO_75 (O_75,N_24960,N_24558);
and UO_76 (O_76,N_24937,N_24525);
nand UO_77 (O_77,N_24724,N_24860);
xnor UO_78 (O_78,N_24711,N_24559);
nor UO_79 (O_79,N_24792,N_24515);
xor UO_80 (O_80,N_24864,N_24969);
nand UO_81 (O_81,N_24702,N_24747);
xnor UO_82 (O_82,N_24619,N_24856);
and UO_83 (O_83,N_24506,N_24931);
and UO_84 (O_84,N_24800,N_24660);
nand UO_85 (O_85,N_24903,N_24623);
or UO_86 (O_86,N_24589,N_24722);
xor UO_87 (O_87,N_24803,N_24910);
nor UO_88 (O_88,N_24844,N_24941);
nand UO_89 (O_89,N_24833,N_24914);
and UO_90 (O_90,N_24757,N_24909);
and UO_91 (O_91,N_24710,N_24758);
nor UO_92 (O_92,N_24707,N_24847);
nor UO_93 (O_93,N_24991,N_24837);
and UO_94 (O_94,N_24521,N_24993);
xnor UO_95 (O_95,N_24642,N_24788);
or UO_96 (O_96,N_24999,N_24582);
nand UO_97 (O_97,N_24772,N_24542);
nor UO_98 (O_98,N_24565,N_24682);
xor UO_99 (O_99,N_24851,N_24896);
nor UO_100 (O_100,N_24989,N_24504);
or UO_101 (O_101,N_24958,N_24666);
nand UO_102 (O_102,N_24516,N_24900);
nand UO_103 (O_103,N_24952,N_24881);
and UO_104 (O_104,N_24955,N_24899);
nand UO_105 (O_105,N_24954,N_24584);
or UO_106 (O_106,N_24975,N_24876);
xor UO_107 (O_107,N_24921,N_24923);
and UO_108 (O_108,N_24590,N_24841);
xnor UO_109 (O_109,N_24624,N_24655);
and UO_110 (O_110,N_24935,N_24613);
and UO_111 (O_111,N_24806,N_24693);
nand UO_112 (O_112,N_24729,N_24885);
or UO_113 (O_113,N_24978,N_24517);
nand UO_114 (O_114,N_24853,N_24527);
xnor UO_115 (O_115,N_24605,N_24818);
xnor UO_116 (O_116,N_24752,N_24947);
xnor UO_117 (O_117,N_24595,N_24918);
xor UO_118 (O_118,N_24951,N_24653);
nor UO_119 (O_119,N_24827,N_24770);
xnor UO_120 (O_120,N_24810,N_24948);
xor UO_121 (O_121,N_24713,N_24794);
nand UO_122 (O_122,N_24974,N_24890);
or UO_123 (O_123,N_24502,N_24888);
and UO_124 (O_124,N_24594,N_24581);
or UO_125 (O_125,N_24944,N_24635);
nand UO_126 (O_126,N_24980,N_24700);
or UO_127 (O_127,N_24612,N_24922);
nor UO_128 (O_128,N_24766,N_24811);
nor UO_129 (O_129,N_24520,N_24514);
or UO_130 (O_130,N_24683,N_24873);
xnor UO_131 (O_131,N_24508,N_24882);
and UO_132 (O_132,N_24712,N_24970);
and UO_133 (O_133,N_24573,N_24996);
or UO_134 (O_134,N_24976,N_24904);
xor UO_135 (O_135,N_24745,N_24748);
or UO_136 (O_136,N_24593,N_24943);
and UO_137 (O_137,N_24984,N_24609);
xnor UO_138 (O_138,N_24507,N_24648);
or UO_139 (O_139,N_24824,N_24783);
nand UO_140 (O_140,N_24524,N_24647);
and UO_141 (O_141,N_24709,N_24547);
or UO_142 (O_142,N_24688,N_24610);
and UO_143 (O_143,N_24530,N_24577);
and UO_144 (O_144,N_24966,N_24832);
and UO_145 (O_145,N_24686,N_24815);
xnor UO_146 (O_146,N_24534,N_24793);
or UO_147 (O_147,N_24608,N_24664);
or UO_148 (O_148,N_24538,N_24680);
nand UO_149 (O_149,N_24961,N_24548);
xnor UO_150 (O_150,N_24733,N_24567);
nand UO_151 (O_151,N_24782,N_24821);
xor UO_152 (O_152,N_24705,N_24536);
nor UO_153 (O_153,N_24684,N_24805);
nor UO_154 (O_154,N_24669,N_24699);
xor UO_155 (O_155,N_24637,N_24819);
nand UO_156 (O_156,N_24656,N_24866);
nor UO_157 (O_157,N_24751,N_24621);
xnor UO_158 (O_158,N_24808,N_24781);
xnor UO_159 (O_159,N_24940,N_24670);
and UO_160 (O_160,N_24732,N_24634);
or UO_161 (O_161,N_24638,N_24973);
and UO_162 (O_162,N_24790,N_24857);
nor UO_163 (O_163,N_24846,N_24645);
nor UO_164 (O_164,N_24854,N_24528);
nand UO_165 (O_165,N_24786,N_24549);
xor UO_166 (O_166,N_24550,N_24929);
and UO_167 (O_167,N_24852,N_24687);
and UO_168 (O_168,N_24553,N_24905);
nor UO_169 (O_169,N_24868,N_24985);
nand UO_170 (O_170,N_24741,N_24957);
and UO_171 (O_171,N_24665,N_24675);
and UO_172 (O_172,N_24532,N_24750);
xor UO_173 (O_173,N_24799,N_24743);
nand UO_174 (O_174,N_24529,N_24895);
and UO_175 (O_175,N_24863,N_24586);
nand UO_176 (O_176,N_24840,N_24992);
and UO_177 (O_177,N_24836,N_24893);
nor UO_178 (O_178,N_24744,N_24787);
nand UO_179 (O_179,N_24636,N_24990);
xnor UO_180 (O_180,N_24545,N_24599);
nor UO_181 (O_181,N_24556,N_24580);
nor UO_182 (O_182,N_24780,N_24761);
nor UO_183 (O_183,N_24971,N_24839);
nand UO_184 (O_184,N_24604,N_24679);
nor UO_185 (O_185,N_24946,N_24537);
nor UO_186 (O_186,N_24569,N_24704);
nor UO_187 (O_187,N_24546,N_24509);
or UO_188 (O_188,N_24512,N_24977);
or UO_189 (O_189,N_24639,N_24708);
and UO_190 (O_190,N_24572,N_24640);
and UO_191 (O_191,N_24685,N_24779);
nand UO_192 (O_192,N_24902,N_24798);
or UO_193 (O_193,N_24997,N_24652);
nor UO_194 (O_194,N_24867,N_24775);
nand UO_195 (O_195,N_24568,N_24858);
xor UO_196 (O_196,N_24776,N_24924);
and UO_197 (O_197,N_24723,N_24725);
nor UO_198 (O_198,N_24988,N_24880);
or UO_199 (O_199,N_24855,N_24911);
and UO_200 (O_200,N_24823,N_24676);
and UO_201 (O_201,N_24843,N_24972);
xnor UO_202 (O_202,N_24662,N_24730);
nand UO_203 (O_203,N_24949,N_24917);
nor UO_204 (O_204,N_24765,N_24861);
nand UO_205 (O_205,N_24760,N_24611);
nor UO_206 (O_206,N_24571,N_24956);
and UO_207 (O_207,N_24825,N_24845);
nor UO_208 (O_208,N_24620,N_24715);
nor UO_209 (O_209,N_24519,N_24602);
xor UO_210 (O_210,N_24703,N_24583);
nand UO_211 (O_211,N_24964,N_24746);
and UO_212 (O_212,N_24872,N_24500);
or UO_213 (O_213,N_24513,N_24802);
nor UO_214 (O_214,N_24801,N_24892);
and UO_215 (O_215,N_24828,N_24795);
or UO_216 (O_216,N_24734,N_24596);
nand UO_217 (O_217,N_24616,N_24774);
or UO_218 (O_218,N_24883,N_24939);
and UO_219 (O_219,N_24813,N_24817);
and UO_220 (O_220,N_24933,N_24697);
or UO_221 (O_221,N_24606,N_24625);
and UO_222 (O_222,N_24784,N_24657);
xor UO_223 (O_223,N_24543,N_24913);
xnor UO_224 (O_224,N_24554,N_24797);
and UO_225 (O_225,N_24626,N_24603);
nor UO_226 (O_226,N_24884,N_24721);
xnor UO_227 (O_227,N_24555,N_24789);
xor UO_228 (O_228,N_24618,N_24719);
xnor UO_229 (O_229,N_24535,N_24877);
xnor UO_230 (O_230,N_24875,N_24749);
xnor UO_231 (O_231,N_24526,N_24720);
or UO_232 (O_232,N_24906,N_24630);
or UO_233 (O_233,N_24678,N_24505);
or UO_234 (O_234,N_24822,N_24651);
and UO_235 (O_235,N_24778,N_24659);
nand UO_236 (O_236,N_24742,N_24934);
xnor UO_237 (O_237,N_24706,N_24566);
nor UO_238 (O_238,N_24510,N_24835);
nor UO_239 (O_239,N_24501,N_24689);
and UO_240 (O_240,N_24871,N_24601);
xnor UO_241 (O_241,N_24627,N_24763);
nor UO_242 (O_242,N_24771,N_24650);
xor UO_243 (O_243,N_24695,N_24714);
nand UO_244 (O_244,N_24814,N_24591);
xnor UO_245 (O_245,N_24968,N_24791);
nand UO_246 (O_246,N_24963,N_24916);
and UO_247 (O_247,N_24691,N_24663);
and UO_248 (O_248,N_24816,N_24735);
nand UO_249 (O_249,N_24617,N_24838);
nand UO_250 (O_250,N_24926,N_24825);
nor UO_251 (O_251,N_24819,N_24821);
nor UO_252 (O_252,N_24762,N_24982);
nor UO_253 (O_253,N_24913,N_24867);
and UO_254 (O_254,N_24698,N_24899);
and UO_255 (O_255,N_24723,N_24531);
xor UO_256 (O_256,N_24624,N_24942);
nor UO_257 (O_257,N_24900,N_24901);
nand UO_258 (O_258,N_24764,N_24718);
nor UO_259 (O_259,N_24943,N_24819);
nor UO_260 (O_260,N_24702,N_24761);
nor UO_261 (O_261,N_24822,N_24836);
xor UO_262 (O_262,N_24804,N_24717);
nor UO_263 (O_263,N_24606,N_24653);
or UO_264 (O_264,N_24524,N_24750);
nor UO_265 (O_265,N_24705,N_24673);
or UO_266 (O_266,N_24714,N_24595);
nor UO_267 (O_267,N_24700,N_24945);
nand UO_268 (O_268,N_24560,N_24529);
nand UO_269 (O_269,N_24869,N_24994);
xnor UO_270 (O_270,N_24746,N_24524);
xnor UO_271 (O_271,N_24923,N_24915);
and UO_272 (O_272,N_24956,N_24522);
nor UO_273 (O_273,N_24857,N_24595);
nand UO_274 (O_274,N_24940,N_24522);
nor UO_275 (O_275,N_24767,N_24868);
and UO_276 (O_276,N_24906,N_24759);
or UO_277 (O_277,N_24936,N_24943);
xor UO_278 (O_278,N_24828,N_24898);
nand UO_279 (O_279,N_24780,N_24511);
and UO_280 (O_280,N_24646,N_24558);
nand UO_281 (O_281,N_24995,N_24867);
nor UO_282 (O_282,N_24702,N_24840);
xnor UO_283 (O_283,N_24622,N_24650);
nor UO_284 (O_284,N_24981,N_24864);
xnor UO_285 (O_285,N_24594,N_24650);
or UO_286 (O_286,N_24968,N_24964);
nor UO_287 (O_287,N_24620,N_24768);
or UO_288 (O_288,N_24538,N_24951);
xnor UO_289 (O_289,N_24862,N_24694);
nor UO_290 (O_290,N_24938,N_24795);
nand UO_291 (O_291,N_24573,N_24675);
or UO_292 (O_292,N_24747,N_24530);
or UO_293 (O_293,N_24722,N_24710);
nor UO_294 (O_294,N_24942,N_24932);
or UO_295 (O_295,N_24635,N_24668);
nand UO_296 (O_296,N_24833,N_24705);
or UO_297 (O_297,N_24837,N_24699);
or UO_298 (O_298,N_24947,N_24818);
nand UO_299 (O_299,N_24929,N_24627);
and UO_300 (O_300,N_24728,N_24590);
or UO_301 (O_301,N_24504,N_24756);
nor UO_302 (O_302,N_24575,N_24761);
xnor UO_303 (O_303,N_24989,N_24717);
and UO_304 (O_304,N_24633,N_24962);
and UO_305 (O_305,N_24789,N_24773);
nand UO_306 (O_306,N_24797,N_24547);
and UO_307 (O_307,N_24811,N_24808);
xor UO_308 (O_308,N_24777,N_24696);
xnor UO_309 (O_309,N_24887,N_24634);
nor UO_310 (O_310,N_24898,N_24510);
nor UO_311 (O_311,N_24792,N_24692);
or UO_312 (O_312,N_24597,N_24867);
nor UO_313 (O_313,N_24826,N_24779);
nor UO_314 (O_314,N_24927,N_24608);
xnor UO_315 (O_315,N_24741,N_24754);
nand UO_316 (O_316,N_24819,N_24678);
nand UO_317 (O_317,N_24931,N_24556);
nor UO_318 (O_318,N_24681,N_24896);
nand UO_319 (O_319,N_24666,N_24962);
or UO_320 (O_320,N_24626,N_24665);
and UO_321 (O_321,N_24746,N_24608);
and UO_322 (O_322,N_24873,N_24736);
nor UO_323 (O_323,N_24841,N_24923);
or UO_324 (O_324,N_24708,N_24831);
or UO_325 (O_325,N_24599,N_24783);
nor UO_326 (O_326,N_24653,N_24618);
nand UO_327 (O_327,N_24554,N_24521);
nor UO_328 (O_328,N_24698,N_24523);
nor UO_329 (O_329,N_24883,N_24783);
nor UO_330 (O_330,N_24860,N_24578);
xnor UO_331 (O_331,N_24918,N_24660);
nand UO_332 (O_332,N_24727,N_24879);
xnor UO_333 (O_333,N_24632,N_24614);
and UO_334 (O_334,N_24709,N_24917);
nor UO_335 (O_335,N_24666,N_24775);
or UO_336 (O_336,N_24577,N_24527);
xor UO_337 (O_337,N_24606,N_24929);
and UO_338 (O_338,N_24936,N_24793);
nand UO_339 (O_339,N_24633,N_24670);
or UO_340 (O_340,N_24911,N_24995);
nor UO_341 (O_341,N_24648,N_24526);
nand UO_342 (O_342,N_24807,N_24946);
nand UO_343 (O_343,N_24808,N_24861);
nor UO_344 (O_344,N_24834,N_24566);
or UO_345 (O_345,N_24557,N_24703);
nor UO_346 (O_346,N_24748,N_24906);
nor UO_347 (O_347,N_24608,N_24998);
nand UO_348 (O_348,N_24980,N_24829);
nor UO_349 (O_349,N_24770,N_24573);
nand UO_350 (O_350,N_24700,N_24828);
or UO_351 (O_351,N_24741,N_24630);
nand UO_352 (O_352,N_24819,N_24644);
nor UO_353 (O_353,N_24716,N_24598);
xor UO_354 (O_354,N_24745,N_24531);
xor UO_355 (O_355,N_24600,N_24919);
xnor UO_356 (O_356,N_24633,N_24721);
and UO_357 (O_357,N_24804,N_24909);
or UO_358 (O_358,N_24801,N_24603);
nor UO_359 (O_359,N_24553,N_24528);
xnor UO_360 (O_360,N_24887,N_24637);
and UO_361 (O_361,N_24744,N_24907);
nand UO_362 (O_362,N_24504,N_24591);
or UO_363 (O_363,N_24833,N_24850);
xnor UO_364 (O_364,N_24564,N_24924);
xor UO_365 (O_365,N_24801,N_24831);
and UO_366 (O_366,N_24906,N_24830);
xor UO_367 (O_367,N_24702,N_24815);
xnor UO_368 (O_368,N_24603,N_24813);
nand UO_369 (O_369,N_24900,N_24922);
or UO_370 (O_370,N_24525,N_24668);
nand UO_371 (O_371,N_24504,N_24687);
xnor UO_372 (O_372,N_24990,N_24732);
nand UO_373 (O_373,N_24501,N_24901);
xnor UO_374 (O_374,N_24694,N_24981);
xnor UO_375 (O_375,N_24541,N_24547);
xnor UO_376 (O_376,N_24693,N_24548);
or UO_377 (O_377,N_24998,N_24505);
nand UO_378 (O_378,N_24675,N_24750);
nor UO_379 (O_379,N_24829,N_24653);
nor UO_380 (O_380,N_24738,N_24847);
and UO_381 (O_381,N_24790,N_24718);
and UO_382 (O_382,N_24798,N_24668);
nor UO_383 (O_383,N_24921,N_24501);
nor UO_384 (O_384,N_24712,N_24820);
and UO_385 (O_385,N_24788,N_24776);
nand UO_386 (O_386,N_24728,N_24529);
nor UO_387 (O_387,N_24918,N_24640);
nor UO_388 (O_388,N_24831,N_24672);
or UO_389 (O_389,N_24910,N_24721);
nand UO_390 (O_390,N_24536,N_24631);
nand UO_391 (O_391,N_24976,N_24919);
nor UO_392 (O_392,N_24719,N_24531);
nor UO_393 (O_393,N_24586,N_24624);
nor UO_394 (O_394,N_24550,N_24608);
or UO_395 (O_395,N_24635,N_24675);
nor UO_396 (O_396,N_24824,N_24981);
nor UO_397 (O_397,N_24954,N_24780);
or UO_398 (O_398,N_24571,N_24927);
xor UO_399 (O_399,N_24922,N_24833);
or UO_400 (O_400,N_24680,N_24897);
or UO_401 (O_401,N_24614,N_24671);
or UO_402 (O_402,N_24644,N_24744);
xnor UO_403 (O_403,N_24804,N_24512);
nor UO_404 (O_404,N_24748,N_24813);
xor UO_405 (O_405,N_24557,N_24784);
and UO_406 (O_406,N_24955,N_24631);
nor UO_407 (O_407,N_24784,N_24731);
xor UO_408 (O_408,N_24591,N_24712);
xnor UO_409 (O_409,N_24586,N_24507);
nand UO_410 (O_410,N_24935,N_24516);
xor UO_411 (O_411,N_24899,N_24975);
nor UO_412 (O_412,N_24603,N_24631);
or UO_413 (O_413,N_24501,N_24743);
nand UO_414 (O_414,N_24952,N_24789);
and UO_415 (O_415,N_24962,N_24566);
nand UO_416 (O_416,N_24531,N_24981);
and UO_417 (O_417,N_24677,N_24942);
nor UO_418 (O_418,N_24596,N_24714);
xor UO_419 (O_419,N_24914,N_24528);
xnor UO_420 (O_420,N_24804,N_24718);
or UO_421 (O_421,N_24521,N_24731);
and UO_422 (O_422,N_24819,N_24558);
nand UO_423 (O_423,N_24500,N_24538);
xor UO_424 (O_424,N_24570,N_24846);
nor UO_425 (O_425,N_24878,N_24965);
and UO_426 (O_426,N_24572,N_24573);
or UO_427 (O_427,N_24682,N_24588);
xnor UO_428 (O_428,N_24726,N_24957);
xor UO_429 (O_429,N_24507,N_24630);
and UO_430 (O_430,N_24529,N_24841);
xor UO_431 (O_431,N_24741,N_24666);
and UO_432 (O_432,N_24535,N_24586);
nor UO_433 (O_433,N_24778,N_24624);
nand UO_434 (O_434,N_24521,N_24593);
xnor UO_435 (O_435,N_24886,N_24996);
xor UO_436 (O_436,N_24734,N_24627);
or UO_437 (O_437,N_24930,N_24892);
and UO_438 (O_438,N_24850,N_24765);
nand UO_439 (O_439,N_24965,N_24706);
nand UO_440 (O_440,N_24551,N_24963);
nand UO_441 (O_441,N_24903,N_24683);
or UO_442 (O_442,N_24565,N_24719);
and UO_443 (O_443,N_24747,N_24571);
nand UO_444 (O_444,N_24611,N_24646);
nor UO_445 (O_445,N_24850,N_24774);
and UO_446 (O_446,N_24795,N_24903);
nand UO_447 (O_447,N_24875,N_24798);
xor UO_448 (O_448,N_24666,N_24746);
nand UO_449 (O_449,N_24604,N_24931);
and UO_450 (O_450,N_24739,N_24525);
or UO_451 (O_451,N_24525,N_24918);
nand UO_452 (O_452,N_24878,N_24746);
and UO_453 (O_453,N_24690,N_24707);
nor UO_454 (O_454,N_24677,N_24547);
nor UO_455 (O_455,N_24568,N_24502);
nor UO_456 (O_456,N_24932,N_24701);
and UO_457 (O_457,N_24536,N_24736);
and UO_458 (O_458,N_24881,N_24502);
and UO_459 (O_459,N_24645,N_24895);
nor UO_460 (O_460,N_24682,N_24647);
and UO_461 (O_461,N_24810,N_24914);
xor UO_462 (O_462,N_24874,N_24796);
xnor UO_463 (O_463,N_24805,N_24601);
xnor UO_464 (O_464,N_24693,N_24625);
xnor UO_465 (O_465,N_24780,N_24704);
nand UO_466 (O_466,N_24766,N_24987);
and UO_467 (O_467,N_24882,N_24824);
nand UO_468 (O_468,N_24888,N_24849);
or UO_469 (O_469,N_24652,N_24675);
or UO_470 (O_470,N_24672,N_24702);
and UO_471 (O_471,N_24870,N_24976);
nand UO_472 (O_472,N_24747,N_24801);
nand UO_473 (O_473,N_24621,N_24924);
xor UO_474 (O_474,N_24919,N_24611);
or UO_475 (O_475,N_24896,N_24758);
nand UO_476 (O_476,N_24755,N_24686);
and UO_477 (O_477,N_24593,N_24957);
nand UO_478 (O_478,N_24722,N_24796);
xor UO_479 (O_479,N_24894,N_24799);
and UO_480 (O_480,N_24811,N_24599);
xnor UO_481 (O_481,N_24667,N_24744);
xnor UO_482 (O_482,N_24767,N_24849);
or UO_483 (O_483,N_24734,N_24991);
nor UO_484 (O_484,N_24653,N_24615);
xor UO_485 (O_485,N_24781,N_24784);
or UO_486 (O_486,N_24935,N_24626);
nand UO_487 (O_487,N_24654,N_24780);
nor UO_488 (O_488,N_24505,N_24600);
nand UO_489 (O_489,N_24962,N_24808);
xor UO_490 (O_490,N_24851,N_24526);
or UO_491 (O_491,N_24701,N_24799);
nor UO_492 (O_492,N_24514,N_24553);
xor UO_493 (O_493,N_24504,N_24803);
xor UO_494 (O_494,N_24701,N_24808);
or UO_495 (O_495,N_24521,N_24913);
xor UO_496 (O_496,N_24758,N_24948);
or UO_497 (O_497,N_24565,N_24503);
nor UO_498 (O_498,N_24945,N_24654);
nor UO_499 (O_499,N_24642,N_24847);
and UO_500 (O_500,N_24597,N_24557);
nor UO_501 (O_501,N_24848,N_24881);
nor UO_502 (O_502,N_24518,N_24743);
nand UO_503 (O_503,N_24579,N_24714);
xor UO_504 (O_504,N_24737,N_24790);
or UO_505 (O_505,N_24535,N_24962);
nor UO_506 (O_506,N_24732,N_24630);
nor UO_507 (O_507,N_24973,N_24518);
and UO_508 (O_508,N_24816,N_24794);
nor UO_509 (O_509,N_24673,N_24821);
nand UO_510 (O_510,N_24748,N_24621);
nor UO_511 (O_511,N_24817,N_24995);
nand UO_512 (O_512,N_24947,N_24629);
nor UO_513 (O_513,N_24595,N_24533);
nor UO_514 (O_514,N_24510,N_24628);
nor UO_515 (O_515,N_24826,N_24537);
nor UO_516 (O_516,N_24912,N_24979);
nor UO_517 (O_517,N_24772,N_24571);
nor UO_518 (O_518,N_24694,N_24890);
nor UO_519 (O_519,N_24883,N_24719);
xnor UO_520 (O_520,N_24755,N_24712);
xnor UO_521 (O_521,N_24749,N_24589);
or UO_522 (O_522,N_24759,N_24698);
nor UO_523 (O_523,N_24702,N_24952);
and UO_524 (O_524,N_24624,N_24765);
nand UO_525 (O_525,N_24583,N_24569);
or UO_526 (O_526,N_24910,N_24562);
nor UO_527 (O_527,N_24989,N_24829);
nand UO_528 (O_528,N_24748,N_24738);
and UO_529 (O_529,N_24609,N_24620);
or UO_530 (O_530,N_24769,N_24534);
nor UO_531 (O_531,N_24610,N_24975);
xor UO_532 (O_532,N_24531,N_24657);
and UO_533 (O_533,N_24709,N_24678);
or UO_534 (O_534,N_24834,N_24778);
or UO_535 (O_535,N_24609,N_24890);
nand UO_536 (O_536,N_24640,N_24916);
nor UO_537 (O_537,N_24965,N_24847);
or UO_538 (O_538,N_24704,N_24608);
and UO_539 (O_539,N_24784,N_24889);
xnor UO_540 (O_540,N_24913,N_24746);
and UO_541 (O_541,N_24852,N_24838);
or UO_542 (O_542,N_24782,N_24865);
and UO_543 (O_543,N_24728,N_24873);
xnor UO_544 (O_544,N_24539,N_24750);
or UO_545 (O_545,N_24931,N_24773);
and UO_546 (O_546,N_24553,N_24921);
nand UO_547 (O_547,N_24547,N_24553);
and UO_548 (O_548,N_24645,N_24538);
nand UO_549 (O_549,N_24712,N_24987);
nor UO_550 (O_550,N_24540,N_24735);
or UO_551 (O_551,N_24670,N_24996);
nor UO_552 (O_552,N_24870,N_24539);
nor UO_553 (O_553,N_24768,N_24508);
and UO_554 (O_554,N_24563,N_24747);
and UO_555 (O_555,N_24844,N_24602);
nand UO_556 (O_556,N_24749,N_24784);
nand UO_557 (O_557,N_24592,N_24970);
nand UO_558 (O_558,N_24912,N_24940);
xnor UO_559 (O_559,N_24510,N_24630);
or UO_560 (O_560,N_24752,N_24524);
nor UO_561 (O_561,N_24706,N_24789);
nand UO_562 (O_562,N_24654,N_24786);
or UO_563 (O_563,N_24655,N_24708);
xor UO_564 (O_564,N_24837,N_24563);
nor UO_565 (O_565,N_24892,N_24531);
or UO_566 (O_566,N_24732,N_24711);
nor UO_567 (O_567,N_24840,N_24721);
xor UO_568 (O_568,N_24979,N_24548);
nor UO_569 (O_569,N_24836,N_24767);
and UO_570 (O_570,N_24889,N_24991);
or UO_571 (O_571,N_24524,N_24748);
nor UO_572 (O_572,N_24794,N_24507);
nor UO_573 (O_573,N_24829,N_24791);
and UO_574 (O_574,N_24915,N_24563);
or UO_575 (O_575,N_24934,N_24791);
nor UO_576 (O_576,N_24932,N_24894);
xor UO_577 (O_577,N_24899,N_24863);
or UO_578 (O_578,N_24864,N_24860);
xor UO_579 (O_579,N_24509,N_24994);
nand UO_580 (O_580,N_24790,N_24984);
nor UO_581 (O_581,N_24583,N_24599);
or UO_582 (O_582,N_24531,N_24508);
nor UO_583 (O_583,N_24905,N_24851);
xor UO_584 (O_584,N_24600,N_24816);
xor UO_585 (O_585,N_24916,N_24590);
nand UO_586 (O_586,N_24766,N_24900);
nor UO_587 (O_587,N_24640,N_24963);
and UO_588 (O_588,N_24695,N_24832);
xnor UO_589 (O_589,N_24749,N_24933);
xnor UO_590 (O_590,N_24648,N_24529);
xor UO_591 (O_591,N_24769,N_24724);
nor UO_592 (O_592,N_24709,N_24948);
nor UO_593 (O_593,N_24856,N_24555);
nand UO_594 (O_594,N_24524,N_24804);
xnor UO_595 (O_595,N_24878,N_24824);
nand UO_596 (O_596,N_24943,N_24559);
and UO_597 (O_597,N_24867,N_24848);
nor UO_598 (O_598,N_24844,N_24626);
xor UO_599 (O_599,N_24832,N_24694);
nor UO_600 (O_600,N_24589,N_24797);
nor UO_601 (O_601,N_24793,N_24680);
xnor UO_602 (O_602,N_24768,N_24677);
nand UO_603 (O_603,N_24511,N_24757);
nor UO_604 (O_604,N_24668,N_24795);
and UO_605 (O_605,N_24875,N_24534);
nor UO_606 (O_606,N_24516,N_24994);
nand UO_607 (O_607,N_24691,N_24862);
xnor UO_608 (O_608,N_24506,N_24527);
or UO_609 (O_609,N_24956,N_24714);
nor UO_610 (O_610,N_24636,N_24517);
nand UO_611 (O_611,N_24671,N_24651);
nor UO_612 (O_612,N_24915,N_24673);
nor UO_613 (O_613,N_24521,N_24808);
nand UO_614 (O_614,N_24812,N_24967);
nand UO_615 (O_615,N_24734,N_24960);
nand UO_616 (O_616,N_24596,N_24884);
xnor UO_617 (O_617,N_24652,N_24596);
nand UO_618 (O_618,N_24522,N_24979);
and UO_619 (O_619,N_24791,N_24528);
or UO_620 (O_620,N_24883,N_24506);
and UO_621 (O_621,N_24819,N_24807);
nor UO_622 (O_622,N_24582,N_24589);
or UO_623 (O_623,N_24733,N_24502);
nand UO_624 (O_624,N_24507,N_24707);
xor UO_625 (O_625,N_24896,N_24907);
or UO_626 (O_626,N_24599,N_24748);
and UO_627 (O_627,N_24832,N_24994);
nor UO_628 (O_628,N_24833,N_24770);
or UO_629 (O_629,N_24766,N_24712);
xnor UO_630 (O_630,N_24924,N_24996);
nor UO_631 (O_631,N_24833,N_24793);
xor UO_632 (O_632,N_24829,N_24925);
or UO_633 (O_633,N_24697,N_24918);
xnor UO_634 (O_634,N_24507,N_24721);
nand UO_635 (O_635,N_24566,N_24728);
nand UO_636 (O_636,N_24965,N_24520);
or UO_637 (O_637,N_24777,N_24504);
nor UO_638 (O_638,N_24603,N_24520);
nand UO_639 (O_639,N_24853,N_24542);
nor UO_640 (O_640,N_24991,N_24988);
nor UO_641 (O_641,N_24863,N_24540);
and UO_642 (O_642,N_24985,N_24997);
xnor UO_643 (O_643,N_24827,N_24808);
xnor UO_644 (O_644,N_24708,N_24595);
nor UO_645 (O_645,N_24714,N_24952);
nand UO_646 (O_646,N_24791,N_24874);
and UO_647 (O_647,N_24838,N_24700);
nand UO_648 (O_648,N_24983,N_24518);
nor UO_649 (O_649,N_24688,N_24726);
and UO_650 (O_650,N_24970,N_24515);
and UO_651 (O_651,N_24986,N_24725);
and UO_652 (O_652,N_24750,N_24517);
nand UO_653 (O_653,N_24514,N_24532);
nand UO_654 (O_654,N_24792,N_24604);
nor UO_655 (O_655,N_24732,N_24515);
or UO_656 (O_656,N_24534,N_24654);
xnor UO_657 (O_657,N_24549,N_24948);
xor UO_658 (O_658,N_24767,N_24739);
nand UO_659 (O_659,N_24565,N_24874);
nand UO_660 (O_660,N_24813,N_24799);
nand UO_661 (O_661,N_24808,N_24525);
and UO_662 (O_662,N_24678,N_24742);
or UO_663 (O_663,N_24545,N_24626);
xor UO_664 (O_664,N_24872,N_24617);
xor UO_665 (O_665,N_24857,N_24777);
or UO_666 (O_666,N_24568,N_24864);
nand UO_667 (O_667,N_24683,N_24758);
xnor UO_668 (O_668,N_24936,N_24678);
or UO_669 (O_669,N_24967,N_24581);
xnor UO_670 (O_670,N_24660,N_24595);
and UO_671 (O_671,N_24686,N_24621);
xnor UO_672 (O_672,N_24821,N_24951);
nor UO_673 (O_673,N_24638,N_24632);
nand UO_674 (O_674,N_24575,N_24858);
nand UO_675 (O_675,N_24564,N_24594);
xnor UO_676 (O_676,N_24728,N_24524);
and UO_677 (O_677,N_24964,N_24933);
and UO_678 (O_678,N_24962,N_24678);
and UO_679 (O_679,N_24679,N_24982);
xnor UO_680 (O_680,N_24547,N_24552);
nor UO_681 (O_681,N_24845,N_24957);
and UO_682 (O_682,N_24507,N_24569);
or UO_683 (O_683,N_24635,N_24986);
nand UO_684 (O_684,N_24522,N_24545);
xnor UO_685 (O_685,N_24926,N_24961);
and UO_686 (O_686,N_24974,N_24763);
nor UO_687 (O_687,N_24512,N_24714);
and UO_688 (O_688,N_24666,N_24930);
xor UO_689 (O_689,N_24925,N_24544);
and UO_690 (O_690,N_24536,N_24693);
nor UO_691 (O_691,N_24784,N_24827);
nor UO_692 (O_692,N_24824,N_24818);
or UO_693 (O_693,N_24535,N_24654);
or UO_694 (O_694,N_24552,N_24556);
or UO_695 (O_695,N_24682,N_24907);
or UO_696 (O_696,N_24669,N_24939);
or UO_697 (O_697,N_24558,N_24725);
or UO_698 (O_698,N_24648,N_24811);
nor UO_699 (O_699,N_24654,N_24569);
nor UO_700 (O_700,N_24534,N_24661);
xor UO_701 (O_701,N_24882,N_24619);
nand UO_702 (O_702,N_24840,N_24897);
nor UO_703 (O_703,N_24670,N_24830);
nand UO_704 (O_704,N_24773,N_24953);
nor UO_705 (O_705,N_24865,N_24678);
xnor UO_706 (O_706,N_24526,N_24610);
xnor UO_707 (O_707,N_24814,N_24805);
nor UO_708 (O_708,N_24769,N_24648);
and UO_709 (O_709,N_24988,N_24863);
nand UO_710 (O_710,N_24544,N_24792);
and UO_711 (O_711,N_24916,N_24601);
xnor UO_712 (O_712,N_24665,N_24846);
nor UO_713 (O_713,N_24768,N_24711);
nand UO_714 (O_714,N_24807,N_24665);
nor UO_715 (O_715,N_24908,N_24734);
or UO_716 (O_716,N_24986,N_24671);
or UO_717 (O_717,N_24518,N_24868);
xor UO_718 (O_718,N_24559,N_24502);
and UO_719 (O_719,N_24872,N_24777);
xor UO_720 (O_720,N_24537,N_24755);
nand UO_721 (O_721,N_24651,N_24753);
nand UO_722 (O_722,N_24535,N_24850);
nand UO_723 (O_723,N_24672,N_24752);
and UO_724 (O_724,N_24661,N_24725);
or UO_725 (O_725,N_24823,N_24754);
and UO_726 (O_726,N_24981,N_24955);
nor UO_727 (O_727,N_24879,N_24507);
and UO_728 (O_728,N_24597,N_24623);
xnor UO_729 (O_729,N_24648,N_24661);
nand UO_730 (O_730,N_24787,N_24527);
xor UO_731 (O_731,N_24570,N_24966);
and UO_732 (O_732,N_24860,N_24989);
and UO_733 (O_733,N_24969,N_24705);
nand UO_734 (O_734,N_24976,N_24698);
or UO_735 (O_735,N_24544,N_24654);
and UO_736 (O_736,N_24906,N_24671);
or UO_737 (O_737,N_24558,N_24845);
nand UO_738 (O_738,N_24855,N_24985);
nand UO_739 (O_739,N_24615,N_24503);
nor UO_740 (O_740,N_24541,N_24831);
nand UO_741 (O_741,N_24963,N_24724);
nor UO_742 (O_742,N_24559,N_24909);
nand UO_743 (O_743,N_24605,N_24974);
xor UO_744 (O_744,N_24551,N_24584);
or UO_745 (O_745,N_24904,N_24710);
nand UO_746 (O_746,N_24606,N_24782);
nor UO_747 (O_747,N_24673,N_24641);
nor UO_748 (O_748,N_24613,N_24592);
or UO_749 (O_749,N_24776,N_24725);
nor UO_750 (O_750,N_24775,N_24558);
nor UO_751 (O_751,N_24587,N_24960);
nand UO_752 (O_752,N_24855,N_24701);
or UO_753 (O_753,N_24806,N_24604);
or UO_754 (O_754,N_24605,N_24924);
xnor UO_755 (O_755,N_24812,N_24916);
and UO_756 (O_756,N_24875,N_24768);
and UO_757 (O_757,N_24762,N_24638);
xnor UO_758 (O_758,N_24570,N_24686);
or UO_759 (O_759,N_24741,N_24879);
and UO_760 (O_760,N_24721,N_24906);
nor UO_761 (O_761,N_24666,N_24761);
xor UO_762 (O_762,N_24861,N_24982);
xor UO_763 (O_763,N_24951,N_24896);
or UO_764 (O_764,N_24725,N_24913);
or UO_765 (O_765,N_24830,N_24716);
nor UO_766 (O_766,N_24888,N_24834);
nand UO_767 (O_767,N_24533,N_24935);
xor UO_768 (O_768,N_24622,N_24635);
nor UO_769 (O_769,N_24895,N_24843);
nor UO_770 (O_770,N_24500,N_24795);
nor UO_771 (O_771,N_24813,N_24715);
xnor UO_772 (O_772,N_24988,N_24834);
nor UO_773 (O_773,N_24698,N_24525);
nand UO_774 (O_774,N_24848,N_24989);
and UO_775 (O_775,N_24767,N_24607);
and UO_776 (O_776,N_24856,N_24773);
xnor UO_777 (O_777,N_24599,N_24997);
or UO_778 (O_778,N_24860,N_24654);
or UO_779 (O_779,N_24816,N_24680);
or UO_780 (O_780,N_24503,N_24827);
nand UO_781 (O_781,N_24513,N_24951);
xnor UO_782 (O_782,N_24982,N_24528);
nand UO_783 (O_783,N_24532,N_24542);
nor UO_784 (O_784,N_24737,N_24641);
nand UO_785 (O_785,N_24529,N_24787);
and UO_786 (O_786,N_24751,N_24537);
nand UO_787 (O_787,N_24632,N_24773);
or UO_788 (O_788,N_24911,N_24583);
nor UO_789 (O_789,N_24808,N_24542);
nand UO_790 (O_790,N_24936,N_24555);
and UO_791 (O_791,N_24649,N_24530);
xor UO_792 (O_792,N_24911,N_24648);
xnor UO_793 (O_793,N_24706,N_24601);
nor UO_794 (O_794,N_24623,N_24707);
xor UO_795 (O_795,N_24775,N_24522);
nand UO_796 (O_796,N_24965,N_24569);
xnor UO_797 (O_797,N_24593,N_24605);
and UO_798 (O_798,N_24964,N_24775);
nor UO_799 (O_799,N_24763,N_24506);
or UO_800 (O_800,N_24655,N_24666);
xor UO_801 (O_801,N_24879,N_24646);
and UO_802 (O_802,N_24850,N_24710);
or UO_803 (O_803,N_24550,N_24696);
and UO_804 (O_804,N_24903,N_24688);
nand UO_805 (O_805,N_24928,N_24580);
nand UO_806 (O_806,N_24692,N_24959);
and UO_807 (O_807,N_24885,N_24754);
and UO_808 (O_808,N_24997,N_24505);
nor UO_809 (O_809,N_24938,N_24717);
nor UO_810 (O_810,N_24578,N_24622);
and UO_811 (O_811,N_24942,N_24744);
nand UO_812 (O_812,N_24730,N_24969);
xor UO_813 (O_813,N_24597,N_24669);
nand UO_814 (O_814,N_24697,N_24940);
nand UO_815 (O_815,N_24918,N_24527);
nand UO_816 (O_816,N_24992,N_24550);
or UO_817 (O_817,N_24665,N_24632);
xnor UO_818 (O_818,N_24558,N_24995);
nand UO_819 (O_819,N_24779,N_24756);
nor UO_820 (O_820,N_24718,N_24516);
or UO_821 (O_821,N_24997,N_24639);
nand UO_822 (O_822,N_24820,N_24558);
xnor UO_823 (O_823,N_24529,N_24991);
or UO_824 (O_824,N_24917,N_24551);
nor UO_825 (O_825,N_24927,N_24925);
or UO_826 (O_826,N_24545,N_24759);
or UO_827 (O_827,N_24625,N_24818);
nor UO_828 (O_828,N_24750,N_24644);
and UO_829 (O_829,N_24996,N_24648);
or UO_830 (O_830,N_24736,N_24518);
or UO_831 (O_831,N_24868,N_24641);
or UO_832 (O_832,N_24803,N_24630);
nor UO_833 (O_833,N_24576,N_24533);
xnor UO_834 (O_834,N_24786,N_24849);
nor UO_835 (O_835,N_24753,N_24942);
or UO_836 (O_836,N_24789,N_24566);
and UO_837 (O_837,N_24957,N_24606);
and UO_838 (O_838,N_24657,N_24619);
xnor UO_839 (O_839,N_24523,N_24549);
xnor UO_840 (O_840,N_24693,N_24591);
and UO_841 (O_841,N_24761,N_24944);
nand UO_842 (O_842,N_24818,N_24500);
nor UO_843 (O_843,N_24815,N_24864);
nor UO_844 (O_844,N_24996,N_24551);
nand UO_845 (O_845,N_24544,N_24664);
nand UO_846 (O_846,N_24653,N_24572);
nand UO_847 (O_847,N_24801,N_24918);
and UO_848 (O_848,N_24603,N_24894);
nand UO_849 (O_849,N_24963,N_24891);
xor UO_850 (O_850,N_24655,N_24542);
and UO_851 (O_851,N_24609,N_24903);
nor UO_852 (O_852,N_24942,N_24867);
or UO_853 (O_853,N_24594,N_24525);
nor UO_854 (O_854,N_24765,N_24927);
or UO_855 (O_855,N_24958,N_24610);
or UO_856 (O_856,N_24770,N_24639);
nor UO_857 (O_857,N_24774,N_24820);
and UO_858 (O_858,N_24519,N_24512);
nand UO_859 (O_859,N_24896,N_24528);
nand UO_860 (O_860,N_24766,N_24765);
or UO_861 (O_861,N_24777,N_24632);
or UO_862 (O_862,N_24989,N_24977);
or UO_863 (O_863,N_24509,N_24508);
or UO_864 (O_864,N_24611,N_24675);
nand UO_865 (O_865,N_24812,N_24693);
nor UO_866 (O_866,N_24977,N_24542);
and UO_867 (O_867,N_24872,N_24783);
nor UO_868 (O_868,N_24620,N_24510);
xor UO_869 (O_869,N_24554,N_24689);
xnor UO_870 (O_870,N_24625,N_24655);
nand UO_871 (O_871,N_24517,N_24813);
or UO_872 (O_872,N_24501,N_24600);
nand UO_873 (O_873,N_24752,N_24694);
nand UO_874 (O_874,N_24818,N_24540);
and UO_875 (O_875,N_24565,N_24878);
nand UO_876 (O_876,N_24641,N_24878);
xnor UO_877 (O_877,N_24753,N_24539);
xor UO_878 (O_878,N_24693,N_24934);
nand UO_879 (O_879,N_24759,N_24970);
or UO_880 (O_880,N_24984,N_24898);
nor UO_881 (O_881,N_24661,N_24532);
nand UO_882 (O_882,N_24821,N_24643);
and UO_883 (O_883,N_24632,N_24993);
nor UO_884 (O_884,N_24827,N_24583);
and UO_885 (O_885,N_24810,N_24723);
or UO_886 (O_886,N_24849,N_24775);
nand UO_887 (O_887,N_24829,N_24674);
xnor UO_888 (O_888,N_24791,N_24555);
nor UO_889 (O_889,N_24805,N_24795);
nand UO_890 (O_890,N_24809,N_24544);
nor UO_891 (O_891,N_24872,N_24569);
nand UO_892 (O_892,N_24897,N_24618);
nor UO_893 (O_893,N_24888,N_24525);
nand UO_894 (O_894,N_24533,N_24727);
or UO_895 (O_895,N_24740,N_24704);
and UO_896 (O_896,N_24510,N_24777);
or UO_897 (O_897,N_24977,N_24628);
nand UO_898 (O_898,N_24553,N_24818);
or UO_899 (O_899,N_24672,N_24748);
or UO_900 (O_900,N_24790,N_24933);
nand UO_901 (O_901,N_24710,N_24626);
or UO_902 (O_902,N_24949,N_24728);
and UO_903 (O_903,N_24825,N_24731);
and UO_904 (O_904,N_24838,N_24512);
nand UO_905 (O_905,N_24585,N_24993);
nor UO_906 (O_906,N_24952,N_24614);
nor UO_907 (O_907,N_24755,N_24658);
and UO_908 (O_908,N_24622,N_24869);
and UO_909 (O_909,N_24746,N_24606);
and UO_910 (O_910,N_24503,N_24889);
nor UO_911 (O_911,N_24552,N_24754);
xnor UO_912 (O_912,N_24976,N_24663);
and UO_913 (O_913,N_24993,N_24949);
or UO_914 (O_914,N_24910,N_24819);
nor UO_915 (O_915,N_24611,N_24697);
nand UO_916 (O_916,N_24892,N_24684);
or UO_917 (O_917,N_24649,N_24922);
or UO_918 (O_918,N_24913,N_24884);
xor UO_919 (O_919,N_24913,N_24713);
nor UO_920 (O_920,N_24671,N_24583);
xor UO_921 (O_921,N_24634,N_24658);
xnor UO_922 (O_922,N_24673,N_24913);
or UO_923 (O_923,N_24725,N_24526);
or UO_924 (O_924,N_24794,N_24804);
and UO_925 (O_925,N_24578,N_24658);
nor UO_926 (O_926,N_24652,N_24602);
or UO_927 (O_927,N_24818,N_24849);
xnor UO_928 (O_928,N_24914,N_24611);
nand UO_929 (O_929,N_24783,N_24842);
or UO_930 (O_930,N_24854,N_24735);
nand UO_931 (O_931,N_24673,N_24572);
nand UO_932 (O_932,N_24769,N_24801);
xnor UO_933 (O_933,N_24620,N_24708);
nor UO_934 (O_934,N_24522,N_24882);
or UO_935 (O_935,N_24922,N_24746);
nand UO_936 (O_936,N_24874,N_24806);
nand UO_937 (O_937,N_24743,N_24932);
xnor UO_938 (O_938,N_24735,N_24980);
and UO_939 (O_939,N_24712,N_24693);
xnor UO_940 (O_940,N_24941,N_24870);
nor UO_941 (O_941,N_24817,N_24803);
nor UO_942 (O_942,N_24563,N_24633);
or UO_943 (O_943,N_24588,N_24968);
xnor UO_944 (O_944,N_24912,N_24728);
and UO_945 (O_945,N_24959,N_24554);
xnor UO_946 (O_946,N_24628,N_24651);
and UO_947 (O_947,N_24637,N_24869);
xor UO_948 (O_948,N_24863,N_24943);
or UO_949 (O_949,N_24925,N_24920);
nor UO_950 (O_950,N_24689,N_24663);
nand UO_951 (O_951,N_24850,N_24539);
nor UO_952 (O_952,N_24619,N_24516);
xnor UO_953 (O_953,N_24623,N_24565);
nand UO_954 (O_954,N_24865,N_24800);
xnor UO_955 (O_955,N_24692,N_24514);
or UO_956 (O_956,N_24601,N_24663);
and UO_957 (O_957,N_24751,N_24653);
nor UO_958 (O_958,N_24674,N_24525);
or UO_959 (O_959,N_24573,N_24623);
nand UO_960 (O_960,N_24653,N_24960);
nand UO_961 (O_961,N_24663,N_24749);
nor UO_962 (O_962,N_24894,N_24674);
xor UO_963 (O_963,N_24978,N_24864);
or UO_964 (O_964,N_24750,N_24632);
xor UO_965 (O_965,N_24687,N_24924);
or UO_966 (O_966,N_24908,N_24500);
xnor UO_967 (O_967,N_24895,N_24561);
nor UO_968 (O_968,N_24753,N_24946);
nand UO_969 (O_969,N_24927,N_24977);
xor UO_970 (O_970,N_24914,N_24639);
or UO_971 (O_971,N_24947,N_24843);
or UO_972 (O_972,N_24781,N_24645);
nand UO_973 (O_973,N_24759,N_24971);
or UO_974 (O_974,N_24873,N_24781);
or UO_975 (O_975,N_24743,N_24522);
nor UO_976 (O_976,N_24845,N_24977);
nand UO_977 (O_977,N_24567,N_24500);
or UO_978 (O_978,N_24524,N_24672);
xnor UO_979 (O_979,N_24673,N_24908);
and UO_980 (O_980,N_24708,N_24938);
nor UO_981 (O_981,N_24778,N_24531);
nand UO_982 (O_982,N_24623,N_24516);
and UO_983 (O_983,N_24694,N_24905);
or UO_984 (O_984,N_24978,N_24783);
nand UO_985 (O_985,N_24522,N_24904);
or UO_986 (O_986,N_24631,N_24847);
and UO_987 (O_987,N_24630,N_24924);
and UO_988 (O_988,N_24687,N_24664);
or UO_989 (O_989,N_24511,N_24516);
or UO_990 (O_990,N_24964,N_24747);
nand UO_991 (O_991,N_24747,N_24623);
nand UO_992 (O_992,N_24840,N_24938);
or UO_993 (O_993,N_24903,N_24733);
xnor UO_994 (O_994,N_24676,N_24704);
nand UO_995 (O_995,N_24871,N_24862);
nand UO_996 (O_996,N_24847,N_24880);
and UO_997 (O_997,N_24586,N_24978);
or UO_998 (O_998,N_24567,N_24803);
and UO_999 (O_999,N_24946,N_24727);
and UO_1000 (O_1000,N_24859,N_24999);
or UO_1001 (O_1001,N_24617,N_24776);
or UO_1002 (O_1002,N_24833,N_24727);
xor UO_1003 (O_1003,N_24988,N_24536);
xor UO_1004 (O_1004,N_24602,N_24713);
xor UO_1005 (O_1005,N_24759,N_24627);
or UO_1006 (O_1006,N_24902,N_24916);
xor UO_1007 (O_1007,N_24569,N_24945);
xor UO_1008 (O_1008,N_24611,N_24590);
or UO_1009 (O_1009,N_24622,N_24963);
and UO_1010 (O_1010,N_24583,N_24595);
nor UO_1011 (O_1011,N_24755,N_24701);
and UO_1012 (O_1012,N_24579,N_24751);
or UO_1013 (O_1013,N_24762,N_24533);
xnor UO_1014 (O_1014,N_24541,N_24826);
xor UO_1015 (O_1015,N_24908,N_24881);
or UO_1016 (O_1016,N_24666,N_24909);
nor UO_1017 (O_1017,N_24947,N_24699);
xnor UO_1018 (O_1018,N_24617,N_24942);
nand UO_1019 (O_1019,N_24827,N_24880);
and UO_1020 (O_1020,N_24786,N_24779);
or UO_1021 (O_1021,N_24945,N_24724);
and UO_1022 (O_1022,N_24600,N_24809);
xnor UO_1023 (O_1023,N_24847,N_24639);
or UO_1024 (O_1024,N_24910,N_24965);
or UO_1025 (O_1025,N_24842,N_24524);
nor UO_1026 (O_1026,N_24747,N_24703);
or UO_1027 (O_1027,N_24683,N_24739);
xnor UO_1028 (O_1028,N_24505,N_24745);
xnor UO_1029 (O_1029,N_24634,N_24867);
nand UO_1030 (O_1030,N_24698,N_24526);
xnor UO_1031 (O_1031,N_24735,N_24714);
nor UO_1032 (O_1032,N_24872,N_24638);
or UO_1033 (O_1033,N_24984,N_24721);
xor UO_1034 (O_1034,N_24689,N_24635);
or UO_1035 (O_1035,N_24500,N_24994);
and UO_1036 (O_1036,N_24735,N_24929);
and UO_1037 (O_1037,N_24659,N_24764);
xnor UO_1038 (O_1038,N_24817,N_24710);
nand UO_1039 (O_1039,N_24628,N_24590);
xor UO_1040 (O_1040,N_24510,N_24624);
and UO_1041 (O_1041,N_24826,N_24552);
or UO_1042 (O_1042,N_24957,N_24566);
or UO_1043 (O_1043,N_24696,N_24562);
xnor UO_1044 (O_1044,N_24782,N_24778);
nand UO_1045 (O_1045,N_24849,N_24862);
xor UO_1046 (O_1046,N_24878,N_24662);
nor UO_1047 (O_1047,N_24840,N_24966);
and UO_1048 (O_1048,N_24849,N_24654);
and UO_1049 (O_1049,N_24999,N_24918);
xnor UO_1050 (O_1050,N_24943,N_24562);
nand UO_1051 (O_1051,N_24974,N_24847);
nor UO_1052 (O_1052,N_24795,N_24810);
nor UO_1053 (O_1053,N_24501,N_24913);
or UO_1054 (O_1054,N_24701,N_24828);
and UO_1055 (O_1055,N_24921,N_24982);
nor UO_1056 (O_1056,N_24898,N_24796);
and UO_1057 (O_1057,N_24799,N_24707);
xor UO_1058 (O_1058,N_24583,N_24918);
and UO_1059 (O_1059,N_24962,N_24665);
and UO_1060 (O_1060,N_24891,N_24680);
and UO_1061 (O_1061,N_24890,N_24626);
nor UO_1062 (O_1062,N_24527,N_24741);
and UO_1063 (O_1063,N_24995,N_24697);
xnor UO_1064 (O_1064,N_24999,N_24682);
nand UO_1065 (O_1065,N_24698,N_24551);
nand UO_1066 (O_1066,N_24980,N_24908);
xnor UO_1067 (O_1067,N_24814,N_24969);
or UO_1068 (O_1068,N_24836,N_24768);
and UO_1069 (O_1069,N_24636,N_24647);
nand UO_1070 (O_1070,N_24655,N_24551);
and UO_1071 (O_1071,N_24681,N_24541);
xnor UO_1072 (O_1072,N_24889,N_24616);
and UO_1073 (O_1073,N_24607,N_24787);
nand UO_1074 (O_1074,N_24988,N_24594);
nand UO_1075 (O_1075,N_24690,N_24590);
xnor UO_1076 (O_1076,N_24903,N_24791);
nand UO_1077 (O_1077,N_24671,N_24967);
or UO_1078 (O_1078,N_24796,N_24678);
or UO_1079 (O_1079,N_24721,N_24508);
or UO_1080 (O_1080,N_24871,N_24675);
and UO_1081 (O_1081,N_24754,N_24895);
or UO_1082 (O_1082,N_24957,N_24503);
and UO_1083 (O_1083,N_24766,N_24747);
nand UO_1084 (O_1084,N_24638,N_24500);
or UO_1085 (O_1085,N_24774,N_24957);
or UO_1086 (O_1086,N_24871,N_24850);
nor UO_1087 (O_1087,N_24893,N_24537);
and UO_1088 (O_1088,N_24736,N_24535);
nor UO_1089 (O_1089,N_24839,N_24834);
nor UO_1090 (O_1090,N_24767,N_24784);
nor UO_1091 (O_1091,N_24728,N_24735);
nor UO_1092 (O_1092,N_24838,N_24990);
or UO_1093 (O_1093,N_24791,N_24744);
nor UO_1094 (O_1094,N_24995,N_24847);
nor UO_1095 (O_1095,N_24755,N_24529);
xnor UO_1096 (O_1096,N_24788,N_24912);
and UO_1097 (O_1097,N_24611,N_24670);
and UO_1098 (O_1098,N_24584,N_24850);
or UO_1099 (O_1099,N_24834,N_24961);
xnor UO_1100 (O_1100,N_24918,N_24790);
nand UO_1101 (O_1101,N_24553,N_24906);
nand UO_1102 (O_1102,N_24547,N_24869);
and UO_1103 (O_1103,N_24806,N_24631);
nor UO_1104 (O_1104,N_24588,N_24557);
xor UO_1105 (O_1105,N_24804,N_24797);
xor UO_1106 (O_1106,N_24713,N_24560);
and UO_1107 (O_1107,N_24864,N_24762);
or UO_1108 (O_1108,N_24829,N_24991);
or UO_1109 (O_1109,N_24750,N_24605);
and UO_1110 (O_1110,N_24553,N_24715);
nand UO_1111 (O_1111,N_24568,N_24823);
xnor UO_1112 (O_1112,N_24744,N_24999);
nor UO_1113 (O_1113,N_24598,N_24731);
nand UO_1114 (O_1114,N_24963,N_24590);
nor UO_1115 (O_1115,N_24599,N_24584);
or UO_1116 (O_1116,N_24997,N_24967);
xnor UO_1117 (O_1117,N_24768,N_24600);
and UO_1118 (O_1118,N_24752,N_24982);
or UO_1119 (O_1119,N_24702,N_24598);
nor UO_1120 (O_1120,N_24533,N_24558);
xor UO_1121 (O_1121,N_24650,N_24843);
nand UO_1122 (O_1122,N_24715,N_24799);
nor UO_1123 (O_1123,N_24863,N_24709);
xor UO_1124 (O_1124,N_24931,N_24743);
xor UO_1125 (O_1125,N_24923,N_24514);
xor UO_1126 (O_1126,N_24900,N_24918);
and UO_1127 (O_1127,N_24675,N_24546);
nand UO_1128 (O_1128,N_24702,N_24715);
or UO_1129 (O_1129,N_24541,N_24528);
and UO_1130 (O_1130,N_24515,N_24757);
nand UO_1131 (O_1131,N_24945,N_24807);
xnor UO_1132 (O_1132,N_24670,N_24975);
and UO_1133 (O_1133,N_24548,N_24886);
nand UO_1134 (O_1134,N_24686,N_24759);
or UO_1135 (O_1135,N_24868,N_24531);
nor UO_1136 (O_1136,N_24573,N_24840);
and UO_1137 (O_1137,N_24941,N_24530);
nand UO_1138 (O_1138,N_24593,N_24786);
or UO_1139 (O_1139,N_24787,N_24507);
nand UO_1140 (O_1140,N_24802,N_24500);
nor UO_1141 (O_1141,N_24946,N_24840);
and UO_1142 (O_1142,N_24986,N_24818);
and UO_1143 (O_1143,N_24516,N_24690);
nand UO_1144 (O_1144,N_24949,N_24523);
and UO_1145 (O_1145,N_24524,N_24656);
nand UO_1146 (O_1146,N_24914,N_24934);
or UO_1147 (O_1147,N_24988,N_24813);
xnor UO_1148 (O_1148,N_24779,N_24953);
nor UO_1149 (O_1149,N_24952,N_24510);
or UO_1150 (O_1150,N_24587,N_24853);
and UO_1151 (O_1151,N_24563,N_24655);
nand UO_1152 (O_1152,N_24521,N_24748);
and UO_1153 (O_1153,N_24546,N_24880);
xor UO_1154 (O_1154,N_24798,N_24985);
nor UO_1155 (O_1155,N_24665,N_24735);
and UO_1156 (O_1156,N_24730,N_24986);
and UO_1157 (O_1157,N_24678,N_24909);
and UO_1158 (O_1158,N_24593,N_24822);
xnor UO_1159 (O_1159,N_24900,N_24555);
xnor UO_1160 (O_1160,N_24807,N_24943);
nor UO_1161 (O_1161,N_24770,N_24870);
xnor UO_1162 (O_1162,N_24509,N_24701);
nor UO_1163 (O_1163,N_24758,N_24606);
or UO_1164 (O_1164,N_24906,N_24911);
nor UO_1165 (O_1165,N_24663,N_24523);
and UO_1166 (O_1166,N_24819,N_24534);
and UO_1167 (O_1167,N_24602,N_24975);
or UO_1168 (O_1168,N_24643,N_24878);
nor UO_1169 (O_1169,N_24758,N_24678);
and UO_1170 (O_1170,N_24940,N_24749);
xor UO_1171 (O_1171,N_24688,N_24793);
or UO_1172 (O_1172,N_24653,N_24602);
xnor UO_1173 (O_1173,N_24554,N_24900);
and UO_1174 (O_1174,N_24782,N_24523);
and UO_1175 (O_1175,N_24519,N_24784);
nand UO_1176 (O_1176,N_24857,N_24919);
nand UO_1177 (O_1177,N_24923,N_24761);
nor UO_1178 (O_1178,N_24870,N_24966);
and UO_1179 (O_1179,N_24911,N_24592);
nand UO_1180 (O_1180,N_24564,N_24968);
or UO_1181 (O_1181,N_24958,N_24986);
xnor UO_1182 (O_1182,N_24577,N_24569);
or UO_1183 (O_1183,N_24520,N_24606);
nand UO_1184 (O_1184,N_24867,N_24892);
xor UO_1185 (O_1185,N_24535,N_24839);
or UO_1186 (O_1186,N_24652,N_24544);
nand UO_1187 (O_1187,N_24864,N_24910);
nor UO_1188 (O_1188,N_24709,N_24721);
and UO_1189 (O_1189,N_24565,N_24549);
xor UO_1190 (O_1190,N_24782,N_24570);
xnor UO_1191 (O_1191,N_24561,N_24703);
nand UO_1192 (O_1192,N_24942,N_24573);
and UO_1193 (O_1193,N_24639,N_24794);
and UO_1194 (O_1194,N_24523,N_24592);
nor UO_1195 (O_1195,N_24506,N_24556);
or UO_1196 (O_1196,N_24634,N_24932);
nand UO_1197 (O_1197,N_24923,N_24735);
or UO_1198 (O_1198,N_24918,N_24998);
and UO_1199 (O_1199,N_24936,N_24651);
nand UO_1200 (O_1200,N_24909,N_24658);
xor UO_1201 (O_1201,N_24533,N_24796);
and UO_1202 (O_1202,N_24646,N_24553);
xor UO_1203 (O_1203,N_24661,N_24993);
nor UO_1204 (O_1204,N_24799,N_24919);
nor UO_1205 (O_1205,N_24565,N_24828);
xor UO_1206 (O_1206,N_24725,N_24731);
xnor UO_1207 (O_1207,N_24590,N_24851);
xnor UO_1208 (O_1208,N_24882,N_24983);
nor UO_1209 (O_1209,N_24516,N_24716);
xnor UO_1210 (O_1210,N_24953,N_24676);
and UO_1211 (O_1211,N_24752,N_24951);
or UO_1212 (O_1212,N_24627,N_24881);
and UO_1213 (O_1213,N_24983,N_24610);
or UO_1214 (O_1214,N_24612,N_24926);
or UO_1215 (O_1215,N_24831,N_24535);
and UO_1216 (O_1216,N_24629,N_24853);
and UO_1217 (O_1217,N_24867,N_24677);
nor UO_1218 (O_1218,N_24784,N_24680);
and UO_1219 (O_1219,N_24611,N_24587);
or UO_1220 (O_1220,N_24616,N_24627);
nand UO_1221 (O_1221,N_24690,N_24629);
nor UO_1222 (O_1222,N_24991,N_24591);
and UO_1223 (O_1223,N_24530,N_24783);
and UO_1224 (O_1224,N_24794,N_24801);
nand UO_1225 (O_1225,N_24867,N_24997);
nand UO_1226 (O_1226,N_24508,N_24847);
nor UO_1227 (O_1227,N_24647,N_24657);
or UO_1228 (O_1228,N_24812,N_24939);
xnor UO_1229 (O_1229,N_24826,N_24561);
nor UO_1230 (O_1230,N_24942,N_24725);
or UO_1231 (O_1231,N_24636,N_24582);
nand UO_1232 (O_1232,N_24920,N_24653);
nor UO_1233 (O_1233,N_24518,N_24953);
nand UO_1234 (O_1234,N_24850,N_24793);
and UO_1235 (O_1235,N_24721,N_24786);
nor UO_1236 (O_1236,N_24626,N_24882);
nand UO_1237 (O_1237,N_24963,N_24844);
nand UO_1238 (O_1238,N_24707,N_24684);
nand UO_1239 (O_1239,N_24677,N_24559);
nor UO_1240 (O_1240,N_24920,N_24604);
nor UO_1241 (O_1241,N_24528,N_24581);
nand UO_1242 (O_1242,N_24604,N_24648);
nor UO_1243 (O_1243,N_24754,N_24803);
and UO_1244 (O_1244,N_24796,N_24705);
or UO_1245 (O_1245,N_24538,N_24803);
or UO_1246 (O_1246,N_24651,N_24989);
or UO_1247 (O_1247,N_24678,N_24630);
nand UO_1248 (O_1248,N_24910,N_24674);
and UO_1249 (O_1249,N_24779,N_24828);
or UO_1250 (O_1250,N_24948,N_24825);
nor UO_1251 (O_1251,N_24931,N_24794);
or UO_1252 (O_1252,N_24895,N_24537);
nand UO_1253 (O_1253,N_24689,N_24873);
xor UO_1254 (O_1254,N_24503,N_24534);
nand UO_1255 (O_1255,N_24581,N_24744);
and UO_1256 (O_1256,N_24586,N_24965);
or UO_1257 (O_1257,N_24594,N_24579);
and UO_1258 (O_1258,N_24693,N_24891);
xnor UO_1259 (O_1259,N_24953,N_24559);
or UO_1260 (O_1260,N_24982,N_24834);
xnor UO_1261 (O_1261,N_24580,N_24861);
nand UO_1262 (O_1262,N_24558,N_24929);
nor UO_1263 (O_1263,N_24704,N_24565);
xor UO_1264 (O_1264,N_24639,N_24668);
and UO_1265 (O_1265,N_24792,N_24815);
or UO_1266 (O_1266,N_24662,N_24719);
nor UO_1267 (O_1267,N_24668,N_24596);
nand UO_1268 (O_1268,N_24767,N_24730);
and UO_1269 (O_1269,N_24781,N_24926);
and UO_1270 (O_1270,N_24581,N_24874);
and UO_1271 (O_1271,N_24784,N_24511);
or UO_1272 (O_1272,N_24775,N_24871);
nand UO_1273 (O_1273,N_24866,N_24579);
or UO_1274 (O_1274,N_24668,N_24882);
or UO_1275 (O_1275,N_24726,N_24569);
nand UO_1276 (O_1276,N_24677,N_24554);
and UO_1277 (O_1277,N_24748,N_24573);
or UO_1278 (O_1278,N_24977,N_24913);
or UO_1279 (O_1279,N_24506,N_24734);
or UO_1280 (O_1280,N_24678,N_24932);
xnor UO_1281 (O_1281,N_24871,N_24718);
and UO_1282 (O_1282,N_24876,N_24843);
and UO_1283 (O_1283,N_24667,N_24785);
xnor UO_1284 (O_1284,N_24673,N_24882);
or UO_1285 (O_1285,N_24801,N_24976);
xnor UO_1286 (O_1286,N_24540,N_24557);
nand UO_1287 (O_1287,N_24845,N_24788);
nand UO_1288 (O_1288,N_24940,N_24791);
xnor UO_1289 (O_1289,N_24932,N_24846);
or UO_1290 (O_1290,N_24958,N_24609);
or UO_1291 (O_1291,N_24510,N_24925);
xnor UO_1292 (O_1292,N_24926,N_24573);
nor UO_1293 (O_1293,N_24687,N_24718);
nor UO_1294 (O_1294,N_24785,N_24523);
nor UO_1295 (O_1295,N_24567,N_24715);
xnor UO_1296 (O_1296,N_24819,N_24703);
or UO_1297 (O_1297,N_24936,N_24665);
and UO_1298 (O_1298,N_24690,N_24857);
xor UO_1299 (O_1299,N_24583,N_24863);
or UO_1300 (O_1300,N_24860,N_24592);
or UO_1301 (O_1301,N_24872,N_24719);
xor UO_1302 (O_1302,N_24942,N_24621);
nand UO_1303 (O_1303,N_24749,N_24956);
nor UO_1304 (O_1304,N_24849,N_24730);
nand UO_1305 (O_1305,N_24806,N_24603);
xor UO_1306 (O_1306,N_24990,N_24883);
nand UO_1307 (O_1307,N_24996,N_24665);
and UO_1308 (O_1308,N_24641,N_24680);
or UO_1309 (O_1309,N_24708,N_24935);
xnor UO_1310 (O_1310,N_24535,N_24668);
and UO_1311 (O_1311,N_24598,N_24615);
nand UO_1312 (O_1312,N_24765,N_24520);
nor UO_1313 (O_1313,N_24933,N_24914);
xnor UO_1314 (O_1314,N_24770,N_24512);
nor UO_1315 (O_1315,N_24765,N_24868);
or UO_1316 (O_1316,N_24896,N_24635);
xnor UO_1317 (O_1317,N_24622,N_24696);
xor UO_1318 (O_1318,N_24827,N_24500);
and UO_1319 (O_1319,N_24763,N_24726);
nand UO_1320 (O_1320,N_24806,N_24895);
and UO_1321 (O_1321,N_24783,N_24739);
and UO_1322 (O_1322,N_24832,N_24665);
nand UO_1323 (O_1323,N_24771,N_24817);
xor UO_1324 (O_1324,N_24570,N_24959);
nor UO_1325 (O_1325,N_24652,N_24703);
and UO_1326 (O_1326,N_24602,N_24922);
nor UO_1327 (O_1327,N_24749,N_24685);
nand UO_1328 (O_1328,N_24901,N_24944);
xnor UO_1329 (O_1329,N_24730,N_24994);
xor UO_1330 (O_1330,N_24696,N_24661);
nor UO_1331 (O_1331,N_24730,N_24547);
or UO_1332 (O_1332,N_24582,N_24799);
xnor UO_1333 (O_1333,N_24883,N_24641);
xnor UO_1334 (O_1334,N_24927,N_24726);
xor UO_1335 (O_1335,N_24993,N_24876);
and UO_1336 (O_1336,N_24988,N_24795);
xnor UO_1337 (O_1337,N_24841,N_24830);
nor UO_1338 (O_1338,N_24980,N_24534);
or UO_1339 (O_1339,N_24604,N_24883);
nand UO_1340 (O_1340,N_24552,N_24720);
xnor UO_1341 (O_1341,N_24985,N_24570);
nand UO_1342 (O_1342,N_24707,N_24792);
or UO_1343 (O_1343,N_24661,N_24710);
xnor UO_1344 (O_1344,N_24509,N_24881);
xnor UO_1345 (O_1345,N_24530,N_24960);
nor UO_1346 (O_1346,N_24955,N_24579);
xor UO_1347 (O_1347,N_24763,N_24655);
nor UO_1348 (O_1348,N_24518,N_24674);
and UO_1349 (O_1349,N_24922,N_24628);
and UO_1350 (O_1350,N_24516,N_24653);
nor UO_1351 (O_1351,N_24757,N_24853);
nand UO_1352 (O_1352,N_24670,N_24565);
or UO_1353 (O_1353,N_24817,N_24773);
nand UO_1354 (O_1354,N_24979,N_24689);
and UO_1355 (O_1355,N_24687,N_24520);
xor UO_1356 (O_1356,N_24851,N_24838);
or UO_1357 (O_1357,N_24796,N_24837);
nor UO_1358 (O_1358,N_24815,N_24948);
xor UO_1359 (O_1359,N_24830,N_24854);
or UO_1360 (O_1360,N_24849,N_24671);
nor UO_1361 (O_1361,N_24652,N_24683);
nand UO_1362 (O_1362,N_24988,N_24718);
xnor UO_1363 (O_1363,N_24953,N_24966);
or UO_1364 (O_1364,N_24754,N_24978);
or UO_1365 (O_1365,N_24918,N_24919);
and UO_1366 (O_1366,N_24883,N_24838);
nor UO_1367 (O_1367,N_24933,N_24890);
xnor UO_1368 (O_1368,N_24893,N_24988);
and UO_1369 (O_1369,N_24530,N_24504);
xnor UO_1370 (O_1370,N_24974,N_24972);
nand UO_1371 (O_1371,N_24869,N_24741);
and UO_1372 (O_1372,N_24875,N_24995);
xor UO_1373 (O_1373,N_24558,N_24965);
and UO_1374 (O_1374,N_24826,N_24750);
nor UO_1375 (O_1375,N_24645,N_24663);
nand UO_1376 (O_1376,N_24938,N_24972);
and UO_1377 (O_1377,N_24819,N_24743);
xor UO_1378 (O_1378,N_24655,N_24541);
and UO_1379 (O_1379,N_24652,N_24986);
and UO_1380 (O_1380,N_24620,N_24636);
xnor UO_1381 (O_1381,N_24962,N_24706);
or UO_1382 (O_1382,N_24976,N_24929);
and UO_1383 (O_1383,N_24515,N_24690);
and UO_1384 (O_1384,N_24593,N_24548);
or UO_1385 (O_1385,N_24974,N_24892);
nand UO_1386 (O_1386,N_24822,N_24938);
nor UO_1387 (O_1387,N_24965,N_24508);
nor UO_1388 (O_1388,N_24955,N_24950);
and UO_1389 (O_1389,N_24751,N_24730);
nor UO_1390 (O_1390,N_24973,N_24747);
nand UO_1391 (O_1391,N_24689,N_24924);
xnor UO_1392 (O_1392,N_24702,N_24987);
or UO_1393 (O_1393,N_24652,N_24790);
xor UO_1394 (O_1394,N_24955,N_24883);
nand UO_1395 (O_1395,N_24960,N_24984);
and UO_1396 (O_1396,N_24866,N_24821);
and UO_1397 (O_1397,N_24698,N_24813);
and UO_1398 (O_1398,N_24520,N_24657);
xor UO_1399 (O_1399,N_24938,N_24949);
nand UO_1400 (O_1400,N_24731,N_24625);
nand UO_1401 (O_1401,N_24702,N_24563);
nand UO_1402 (O_1402,N_24666,N_24620);
nor UO_1403 (O_1403,N_24700,N_24555);
and UO_1404 (O_1404,N_24590,N_24927);
nor UO_1405 (O_1405,N_24773,N_24904);
nor UO_1406 (O_1406,N_24854,N_24975);
nand UO_1407 (O_1407,N_24996,N_24730);
nand UO_1408 (O_1408,N_24575,N_24634);
nor UO_1409 (O_1409,N_24646,N_24597);
nand UO_1410 (O_1410,N_24782,N_24909);
or UO_1411 (O_1411,N_24708,N_24625);
xor UO_1412 (O_1412,N_24895,N_24847);
nor UO_1413 (O_1413,N_24525,N_24630);
nor UO_1414 (O_1414,N_24873,N_24611);
nand UO_1415 (O_1415,N_24843,N_24962);
xor UO_1416 (O_1416,N_24657,N_24587);
or UO_1417 (O_1417,N_24754,N_24523);
xor UO_1418 (O_1418,N_24678,N_24701);
nor UO_1419 (O_1419,N_24899,N_24533);
nor UO_1420 (O_1420,N_24872,N_24887);
and UO_1421 (O_1421,N_24734,N_24566);
nand UO_1422 (O_1422,N_24517,N_24652);
or UO_1423 (O_1423,N_24581,N_24991);
or UO_1424 (O_1424,N_24877,N_24775);
nor UO_1425 (O_1425,N_24999,N_24942);
nand UO_1426 (O_1426,N_24881,N_24624);
xor UO_1427 (O_1427,N_24773,N_24569);
nor UO_1428 (O_1428,N_24710,N_24503);
xnor UO_1429 (O_1429,N_24934,N_24838);
and UO_1430 (O_1430,N_24548,N_24562);
nor UO_1431 (O_1431,N_24901,N_24835);
nor UO_1432 (O_1432,N_24823,N_24892);
nor UO_1433 (O_1433,N_24743,N_24995);
and UO_1434 (O_1434,N_24623,N_24962);
xnor UO_1435 (O_1435,N_24512,N_24758);
or UO_1436 (O_1436,N_24610,N_24757);
nand UO_1437 (O_1437,N_24831,N_24926);
xnor UO_1438 (O_1438,N_24756,N_24796);
xor UO_1439 (O_1439,N_24991,N_24646);
xor UO_1440 (O_1440,N_24990,N_24988);
nand UO_1441 (O_1441,N_24688,N_24577);
xnor UO_1442 (O_1442,N_24810,N_24802);
nand UO_1443 (O_1443,N_24552,N_24513);
nand UO_1444 (O_1444,N_24932,N_24750);
xor UO_1445 (O_1445,N_24749,N_24796);
xor UO_1446 (O_1446,N_24710,N_24947);
nor UO_1447 (O_1447,N_24905,N_24602);
nor UO_1448 (O_1448,N_24573,N_24687);
xor UO_1449 (O_1449,N_24691,N_24812);
or UO_1450 (O_1450,N_24658,N_24570);
nand UO_1451 (O_1451,N_24899,N_24927);
and UO_1452 (O_1452,N_24731,N_24607);
xnor UO_1453 (O_1453,N_24702,N_24943);
nand UO_1454 (O_1454,N_24506,N_24518);
or UO_1455 (O_1455,N_24506,N_24769);
nand UO_1456 (O_1456,N_24814,N_24877);
nand UO_1457 (O_1457,N_24634,N_24667);
nor UO_1458 (O_1458,N_24898,N_24896);
or UO_1459 (O_1459,N_24736,N_24875);
xor UO_1460 (O_1460,N_24637,N_24581);
nor UO_1461 (O_1461,N_24628,N_24865);
nor UO_1462 (O_1462,N_24546,N_24682);
or UO_1463 (O_1463,N_24916,N_24592);
nor UO_1464 (O_1464,N_24970,N_24700);
nor UO_1465 (O_1465,N_24841,N_24790);
nand UO_1466 (O_1466,N_24906,N_24973);
nand UO_1467 (O_1467,N_24870,N_24691);
nor UO_1468 (O_1468,N_24884,N_24631);
and UO_1469 (O_1469,N_24991,N_24925);
nor UO_1470 (O_1470,N_24968,N_24928);
nand UO_1471 (O_1471,N_24824,N_24777);
xnor UO_1472 (O_1472,N_24505,N_24629);
and UO_1473 (O_1473,N_24938,N_24942);
xor UO_1474 (O_1474,N_24836,N_24560);
and UO_1475 (O_1475,N_24961,N_24809);
and UO_1476 (O_1476,N_24931,N_24713);
or UO_1477 (O_1477,N_24910,N_24997);
and UO_1478 (O_1478,N_24978,N_24839);
or UO_1479 (O_1479,N_24622,N_24554);
nand UO_1480 (O_1480,N_24960,N_24618);
xor UO_1481 (O_1481,N_24862,N_24623);
nand UO_1482 (O_1482,N_24987,N_24991);
xnor UO_1483 (O_1483,N_24777,N_24763);
or UO_1484 (O_1484,N_24777,N_24998);
and UO_1485 (O_1485,N_24501,N_24927);
nor UO_1486 (O_1486,N_24955,N_24607);
and UO_1487 (O_1487,N_24897,N_24683);
or UO_1488 (O_1488,N_24635,N_24794);
and UO_1489 (O_1489,N_24828,N_24843);
or UO_1490 (O_1490,N_24621,N_24573);
nor UO_1491 (O_1491,N_24966,N_24538);
xor UO_1492 (O_1492,N_24720,N_24902);
xnor UO_1493 (O_1493,N_24629,N_24533);
and UO_1494 (O_1494,N_24895,N_24601);
or UO_1495 (O_1495,N_24975,N_24585);
and UO_1496 (O_1496,N_24624,N_24806);
nand UO_1497 (O_1497,N_24754,N_24994);
or UO_1498 (O_1498,N_24933,N_24912);
and UO_1499 (O_1499,N_24940,N_24692);
and UO_1500 (O_1500,N_24881,N_24751);
xnor UO_1501 (O_1501,N_24842,N_24927);
nand UO_1502 (O_1502,N_24673,N_24559);
xnor UO_1503 (O_1503,N_24587,N_24829);
nor UO_1504 (O_1504,N_24937,N_24623);
nand UO_1505 (O_1505,N_24838,N_24843);
and UO_1506 (O_1506,N_24589,N_24618);
or UO_1507 (O_1507,N_24743,N_24641);
and UO_1508 (O_1508,N_24751,N_24889);
nor UO_1509 (O_1509,N_24892,N_24940);
nor UO_1510 (O_1510,N_24660,N_24523);
or UO_1511 (O_1511,N_24998,N_24732);
nor UO_1512 (O_1512,N_24897,N_24643);
or UO_1513 (O_1513,N_24788,N_24774);
or UO_1514 (O_1514,N_24707,N_24581);
nor UO_1515 (O_1515,N_24942,N_24900);
and UO_1516 (O_1516,N_24952,N_24871);
nand UO_1517 (O_1517,N_24737,N_24880);
and UO_1518 (O_1518,N_24660,N_24751);
nand UO_1519 (O_1519,N_24939,N_24944);
nand UO_1520 (O_1520,N_24902,N_24645);
or UO_1521 (O_1521,N_24806,N_24889);
nor UO_1522 (O_1522,N_24584,N_24575);
nor UO_1523 (O_1523,N_24635,N_24506);
and UO_1524 (O_1524,N_24508,N_24561);
or UO_1525 (O_1525,N_24542,N_24558);
xor UO_1526 (O_1526,N_24920,N_24559);
xnor UO_1527 (O_1527,N_24724,N_24997);
or UO_1528 (O_1528,N_24698,N_24945);
or UO_1529 (O_1529,N_24748,N_24932);
nor UO_1530 (O_1530,N_24568,N_24965);
xor UO_1531 (O_1531,N_24908,N_24862);
nor UO_1532 (O_1532,N_24600,N_24836);
or UO_1533 (O_1533,N_24915,N_24982);
or UO_1534 (O_1534,N_24877,N_24892);
nand UO_1535 (O_1535,N_24537,N_24953);
and UO_1536 (O_1536,N_24806,N_24932);
or UO_1537 (O_1537,N_24588,N_24654);
xor UO_1538 (O_1538,N_24694,N_24755);
nor UO_1539 (O_1539,N_24554,N_24680);
nor UO_1540 (O_1540,N_24898,N_24565);
nor UO_1541 (O_1541,N_24519,N_24690);
xnor UO_1542 (O_1542,N_24939,N_24802);
nor UO_1543 (O_1543,N_24606,N_24971);
nor UO_1544 (O_1544,N_24718,N_24755);
and UO_1545 (O_1545,N_24738,N_24658);
nor UO_1546 (O_1546,N_24590,N_24703);
nand UO_1547 (O_1547,N_24775,N_24715);
nor UO_1548 (O_1548,N_24784,N_24971);
nor UO_1549 (O_1549,N_24825,N_24521);
or UO_1550 (O_1550,N_24604,N_24731);
and UO_1551 (O_1551,N_24772,N_24869);
nor UO_1552 (O_1552,N_24919,N_24909);
nand UO_1553 (O_1553,N_24652,N_24904);
nand UO_1554 (O_1554,N_24602,N_24703);
nor UO_1555 (O_1555,N_24986,N_24881);
and UO_1556 (O_1556,N_24559,N_24941);
or UO_1557 (O_1557,N_24583,N_24941);
and UO_1558 (O_1558,N_24858,N_24506);
or UO_1559 (O_1559,N_24796,N_24775);
or UO_1560 (O_1560,N_24829,N_24567);
nand UO_1561 (O_1561,N_24966,N_24842);
nand UO_1562 (O_1562,N_24841,N_24617);
nor UO_1563 (O_1563,N_24895,N_24932);
nand UO_1564 (O_1564,N_24800,N_24901);
xor UO_1565 (O_1565,N_24651,N_24579);
xor UO_1566 (O_1566,N_24543,N_24822);
and UO_1567 (O_1567,N_24764,N_24608);
xnor UO_1568 (O_1568,N_24588,N_24544);
and UO_1569 (O_1569,N_24704,N_24502);
nor UO_1570 (O_1570,N_24990,N_24997);
nor UO_1571 (O_1571,N_24762,N_24552);
nor UO_1572 (O_1572,N_24998,N_24563);
or UO_1573 (O_1573,N_24558,N_24686);
and UO_1574 (O_1574,N_24782,N_24974);
and UO_1575 (O_1575,N_24850,N_24784);
nor UO_1576 (O_1576,N_24629,N_24572);
xnor UO_1577 (O_1577,N_24531,N_24651);
xnor UO_1578 (O_1578,N_24886,N_24958);
or UO_1579 (O_1579,N_24517,N_24789);
xor UO_1580 (O_1580,N_24842,N_24655);
nand UO_1581 (O_1581,N_24912,N_24610);
and UO_1582 (O_1582,N_24789,N_24536);
or UO_1583 (O_1583,N_24994,N_24768);
nand UO_1584 (O_1584,N_24979,N_24635);
or UO_1585 (O_1585,N_24909,N_24826);
and UO_1586 (O_1586,N_24992,N_24522);
nand UO_1587 (O_1587,N_24895,N_24985);
or UO_1588 (O_1588,N_24652,N_24754);
nand UO_1589 (O_1589,N_24871,N_24838);
xor UO_1590 (O_1590,N_24600,N_24620);
and UO_1591 (O_1591,N_24560,N_24810);
xnor UO_1592 (O_1592,N_24526,N_24764);
nand UO_1593 (O_1593,N_24907,N_24662);
nor UO_1594 (O_1594,N_24735,N_24733);
xor UO_1595 (O_1595,N_24523,N_24826);
xor UO_1596 (O_1596,N_24532,N_24797);
nor UO_1597 (O_1597,N_24820,N_24614);
nand UO_1598 (O_1598,N_24752,N_24561);
nand UO_1599 (O_1599,N_24575,N_24907);
or UO_1600 (O_1600,N_24641,N_24937);
and UO_1601 (O_1601,N_24567,N_24738);
nand UO_1602 (O_1602,N_24938,N_24753);
xor UO_1603 (O_1603,N_24530,N_24552);
nand UO_1604 (O_1604,N_24962,N_24989);
and UO_1605 (O_1605,N_24840,N_24503);
and UO_1606 (O_1606,N_24840,N_24598);
and UO_1607 (O_1607,N_24566,N_24719);
or UO_1608 (O_1608,N_24757,N_24531);
nor UO_1609 (O_1609,N_24669,N_24648);
and UO_1610 (O_1610,N_24772,N_24604);
nor UO_1611 (O_1611,N_24806,N_24683);
or UO_1612 (O_1612,N_24714,N_24996);
or UO_1613 (O_1613,N_24509,N_24915);
and UO_1614 (O_1614,N_24536,N_24975);
and UO_1615 (O_1615,N_24714,N_24916);
xor UO_1616 (O_1616,N_24741,N_24994);
and UO_1617 (O_1617,N_24553,N_24519);
or UO_1618 (O_1618,N_24774,N_24834);
and UO_1619 (O_1619,N_24847,N_24737);
or UO_1620 (O_1620,N_24803,N_24510);
nand UO_1621 (O_1621,N_24816,N_24838);
nand UO_1622 (O_1622,N_24659,N_24587);
nor UO_1623 (O_1623,N_24519,N_24739);
nand UO_1624 (O_1624,N_24983,N_24921);
xor UO_1625 (O_1625,N_24953,N_24978);
and UO_1626 (O_1626,N_24841,N_24963);
xor UO_1627 (O_1627,N_24692,N_24534);
xor UO_1628 (O_1628,N_24597,N_24790);
xor UO_1629 (O_1629,N_24837,N_24634);
nor UO_1630 (O_1630,N_24805,N_24780);
xor UO_1631 (O_1631,N_24507,N_24936);
and UO_1632 (O_1632,N_24536,N_24963);
and UO_1633 (O_1633,N_24696,N_24653);
and UO_1634 (O_1634,N_24994,N_24805);
nand UO_1635 (O_1635,N_24628,N_24557);
nor UO_1636 (O_1636,N_24856,N_24917);
nand UO_1637 (O_1637,N_24553,N_24730);
and UO_1638 (O_1638,N_24895,N_24527);
nor UO_1639 (O_1639,N_24986,N_24763);
or UO_1640 (O_1640,N_24783,N_24710);
or UO_1641 (O_1641,N_24968,N_24627);
and UO_1642 (O_1642,N_24857,N_24969);
or UO_1643 (O_1643,N_24579,N_24785);
nand UO_1644 (O_1644,N_24945,N_24608);
and UO_1645 (O_1645,N_24892,N_24843);
nand UO_1646 (O_1646,N_24763,N_24790);
or UO_1647 (O_1647,N_24588,N_24581);
or UO_1648 (O_1648,N_24699,N_24941);
and UO_1649 (O_1649,N_24815,N_24703);
or UO_1650 (O_1650,N_24555,N_24631);
or UO_1651 (O_1651,N_24848,N_24510);
nand UO_1652 (O_1652,N_24623,N_24811);
or UO_1653 (O_1653,N_24757,N_24683);
nand UO_1654 (O_1654,N_24652,N_24526);
xnor UO_1655 (O_1655,N_24953,N_24972);
and UO_1656 (O_1656,N_24982,N_24667);
xor UO_1657 (O_1657,N_24649,N_24892);
nor UO_1658 (O_1658,N_24747,N_24654);
or UO_1659 (O_1659,N_24786,N_24759);
nand UO_1660 (O_1660,N_24670,N_24788);
nor UO_1661 (O_1661,N_24708,N_24738);
xnor UO_1662 (O_1662,N_24835,N_24888);
nand UO_1663 (O_1663,N_24733,N_24606);
nand UO_1664 (O_1664,N_24548,N_24639);
or UO_1665 (O_1665,N_24908,N_24568);
and UO_1666 (O_1666,N_24863,N_24979);
xor UO_1667 (O_1667,N_24518,N_24662);
and UO_1668 (O_1668,N_24829,N_24594);
nand UO_1669 (O_1669,N_24918,N_24587);
or UO_1670 (O_1670,N_24830,N_24588);
nor UO_1671 (O_1671,N_24579,N_24944);
or UO_1672 (O_1672,N_24609,N_24563);
or UO_1673 (O_1673,N_24735,N_24562);
nand UO_1674 (O_1674,N_24744,N_24719);
nand UO_1675 (O_1675,N_24817,N_24848);
nor UO_1676 (O_1676,N_24633,N_24623);
or UO_1677 (O_1677,N_24991,N_24599);
or UO_1678 (O_1678,N_24571,N_24729);
nand UO_1679 (O_1679,N_24528,N_24657);
xor UO_1680 (O_1680,N_24800,N_24510);
or UO_1681 (O_1681,N_24629,N_24954);
nand UO_1682 (O_1682,N_24539,N_24736);
and UO_1683 (O_1683,N_24571,N_24698);
and UO_1684 (O_1684,N_24829,N_24908);
and UO_1685 (O_1685,N_24651,N_24560);
and UO_1686 (O_1686,N_24511,N_24799);
xor UO_1687 (O_1687,N_24657,N_24565);
nor UO_1688 (O_1688,N_24966,N_24669);
nor UO_1689 (O_1689,N_24623,N_24886);
or UO_1690 (O_1690,N_24814,N_24509);
and UO_1691 (O_1691,N_24585,N_24808);
xor UO_1692 (O_1692,N_24946,N_24979);
and UO_1693 (O_1693,N_24723,N_24800);
or UO_1694 (O_1694,N_24540,N_24942);
or UO_1695 (O_1695,N_24619,N_24797);
nor UO_1696 (O_1696,N_24551,N_24772);
nor UO_1697 (O_1697,N_24946,N_24941);
or UO_1698 (O_1698,N_24578,N_24784);
xnor UO_1699 (O_1699,N_24932,N_24647);
and UO_1700 (O_1700,N_24747,N_24799);
nand UO_1701 (O_1701,N_24759,N_24853);
and UO_1702 (O_1702,N_24669,N_24713);
xnor UO_1703 (O_1703,N_24546,N_24765);
or UO_1704 (O_1704,N_24706,N_24803);
xnor UO_1705 (O_1705,N_24544,N_24737);
nor UO_1706 (O_1706,N_24767,N_24881);
nand UO_1707 (O_1707,N_24968,N_24998);
and UO_1708 (O_1708,N_24511,N_24529);
xnor UO_1709 (O_1709,N_24529,N_24756);
and UO_1710 (O_1710,N_24769,N_24526);
xor UO_1711 (O_1711,N_24702,N_24509);
nand UO_1712 (O_1712,N_24943,N_24778);
xnor UO_1713 (O_1713,N_24597,N_24876);
nand UO_1714 (O_1714,N_24806,N_24804);
and UO_1715 (O_1715,N_24753,N_24812);
xnor UO_1716 (O_1716,N_24731,N_24526);
nor UO_1717 (O_1717,N_24619,N_24501);
nand UO_1718 (O_1718,N_24734,N_24986);
or UO_1719 (O_1719,N_24727,N_24748);
and UO_1720 (O_1720,N_24621,N_24992);
and UO_1721 (O_1721,N_24593,N_24603);
and UO_1722 (O_1722,N_24636,N_24667);
xor UO_1723 (O_1723,N_24974,N_24855);
nand UO_1724 (O_1724,N_24906,N_24905);
nor UO_1725 (O_1725,N_24747,N_24648);
xnor UO_1726 (O_1726,N_24884,N_24679);
nor UO_1727 (O_1727,N_24520,N_24935);
xor UO_1728 (O_1728,N_24944,N_24559);
and UO_1729 (O_1729,N_24514,N_24824);
and UO_1730 (O_1730,N_24891,N_24571);
xor UO_1731 (O_1731,N_24766,N_24913);
and UO_1732 (O_1732,N_24840,N_24670);
or UO_1733 (O_1733,N_24581,N_24751);
and UO_1734 (O_1734,N_24835,N_24928);
xor UO_1735 (O_1735,N_24598,N_24764);
xnor UO_1736 (O_1736,N_24949,N_24721);
nor UO_1737 (O_1737,N_24838,N_24792);
nor UO_1738 (O_1738,N_24869,N_24778);
or UO_1739 (O_1739,N_24777,N_24917);
nand UO_1740 (O_1740,N_24952,N_24602);
xor UO_1741 (O_1741,N_24635,N_24813);
or UO_1742 (O_1742,N_24695,N_24712);
or UO_1743 (O_1743,N_24506,N_24712);
xor UO_1744 (O_1744,N_24653,N_24632);
or UO_1745 (O_1745,N_24931,N_24917);
nand UO_1746 (O_1746,N_24762,N_24538);
or UO_1747 (O_1747,N_24512,N_24628);
or UO_1748 (O_1748,N_24986,N_24857);
and UO_1749 (O_1749,N_24506,N_24966);
and UO_1750 (O_1750,N_24639,N_24596);
nand UO_1751 (O_1751,N_24832,N_24556);
nand UO_1752 (O_1752,N_24815,N_24730);
nor UO_1753 (O_1753,N_24813,N_24738);
and UO_1754 (O_1754,N_24891,N_24744);
and UO_1755 (O_1755,N_24518,N_24837);
or UO_1756 (O_1756,N_24552,N_24846);
nand UO_1757 (O_1757,N_24660,N_24959);
and UO_1758 (O_1758,N_24844,N_24847);
and UO_1759 (O_1759,N_24937,N_24871);
xnor UO_1760 (O_1760,N_24575,N_24513);
or UO_1761 (O_1761,N_24961,N_24566);
or UO_1762 (O_1762,N_24891,N_24955);
nor UO_1763 (O_1763,N_24551,N_24768);
nor UO_1764 (O_1764,N_24528,N_24610);
nor UO_1765 (O_1765,N_24645,N_24869);
and UO_1766 (O_1766,N_24585,N_24857);
and UO_1767 (O_1767,N_24632,N_24899);
nand UO_1768 (O_1768,N_24773,N_24745);
xor UO_1769 (O_1769,N_24949,N_24595);
or UO_1770 (O_1770,N_24589,N_24869);
or UO_1771 (O_1771,N_24665,N_24728);
or UO_1772 (O_1772,N_24827,N_24670);
or UO_1773 (O_1773,N_24543,N_24896);
and UO_1774 (O_1774,N_24743,N_24645);
nand UO_1775 (O_1775,N_24872,N_24678);
nand UO_1776 (O_1776,N_24599,N_24669);
nand UO_1777 (O_1777,N_24577,N_24704);
or UO_1778 (O_1778,N_24917,N_24553);
and UO_1779 (O_1779,N_24641,N_24630);
nand UO_1780 (O_1780,N_24870,N_24764);
nor UO_1781 (O_1781,N_24777,N_24977);
or UO_1782 (O_1782,N_24889,N_24713);
or UO_1783 (O_1783,N_24854,N_24965);
and UO_1784 (O_1784,N_24568,N_24756);
and UO_1785 (O_1785,N_24785,N_24946);
and UO_1786 (O_1786,N_24970,N_24773);
or UO_1787 (O_1787,N_24530,N_24953);
and UO_1788 (O_1788,N_24680,N_24831);
and UO_1789 (O_1789,N_24569,N_24815);
xnor UO_1790 (O_1790,N_24979,N_24805);
xor UO_1791 (O_1791,N_24941,N_24687);
and UO_1792 (O_1792,N_24833,N_24928);
nand UO_1793 (O_1793,N_24919,N_24884);
nor UO_1794 (O_1794,N_24786,N_24853);
or UO_1795 (O_1795,N_24805,N_24872);
or UO_1796 (O_1796,N_24634,N_24709);
nor UO_1797 (O_1797,N_24674,N_24939);
nand UO_1798 (O_1798,N_24905,N_24507);
and UO_1799 (O_1799,N_24808,N_24769);
or UO_1800 (O_1800,N_24718,N_24854);
xor UO_1801 (O_1801,N_24582,N_24613);
nor UO_1802 (O_1802,N_24843,N_24949);
or UO_1803 (O_1803,N_24748,N_24889);
xnor UO_1804 (O_1804,N_24728,N_24525);
xor UO_1805 (O_1805,N_24646,N_24545);
and UO_1806 (O_1806,N_24714,N_24689);
xor UO_1807 (O_1807,N_24945,N_24989);
and UO_1808 (O_1808,N_24822,N_24561);
or UO_1809 (O_1809,N_24676,N_24637);
and UO_1810 (O_1810,N_24523,N_24638);
nand UO_1811 (O_1811,N_24817,N_24593);
nor UO_1812 (O_1812,N_24556,N_24873);
xnor UO_1813 (O_1813,N_24699,N_24876);
nor UO_1814 (O_1814,N_24668,N_24659);
or UO_1815 (O_1815,N_24955,N_24576);
or UO_1816 (O_1816,N_24681,N_24817);
nor UO_1817 (O_1817,N_24581,N_24941);
nor UO_1818 (O_1818,N_24711,N_24537);
and UO_1819 (O_1819,N_24604,N_24675);
xnor UO_1820 (O_1820,N_24613,N_24838);
nand UO_1821 (O_1821,N_24927,N_24961);
nor UO_1822 (O_1822,N_24579,N_24679);
nand UO_1823 (O_1823,N_24843,N_24859);
nand UO_1824 (O_1824,N_24619,N_24620);
xor UO_1825 (O_1825,N_24943,N_24823);
and UO_1826 (O_1826,N_24970,N_24925);
xor UO_1827 (O_1827,N_24835,N_24831);
or UO_1828 (O_1828,N_24797,N_24681);
or UO_1829 (O_1829,N_24893,N_24934);
nor UO_1830 (O_1830,N_24590,N_24770);
xnor UO_1831 (O_1831,N_24843,N_24741);
nor UO_1832 (O_1832,N_24668,N_24651);
and UO_1833 (O_1833,N_24998,N_24936);
nor UO_1834 (O_1834,N_24540,N_24858);
nand UO_1835 (O_1835,N_24522,N_24653);
or UO_1836 (O_1836,N_24724,N_24982);
nand UO_1837 (O_1837,N_24846,N_24626);
nor UO_1838 (O_1838,N_24944,N_24912);
or UO_1839 (O_1839,N_24846,N_24844);
or UO_1840 (O_1840,N_24704,N_24615);
or UO_1841 (O_1841,N_24719,N_24974);
nand UO_1842 (O_1842,N_24686,N_24858);
and UO_1843 (O_1843,N_24601,N_24757);
xor UO_1844 (O_1844,N_24506,N_24702);
nor UO_1845 (O_1845,N_24578,N_24694);
and UO_1846 (O_1846,N_24759,N_24951);
nand UO_1847 (O_1847,N_24944,N_24588);
nand UO_1848 (O_1848,N_24793,N_24589);
or UO_1849 (O_1849,N_24556,N_24517);
xnor UO_1850 (O_1850,N_24894,N_24747);
xor UO_1851 (O_1851,N_24521,N_24832);
xnor UO_1852 (O_1852,N_24524,N_24567);
nand UO_1853 (O_1853,N_24682,N_24572);
and UO_1854 (O_1854,N_24549,N_24928);
and UO_1855 (O_1855,N_24514,N_24864);
xnor UO_1856 (O_1856,N_24757,N_24927);
nand UO_1857 (O_1857,N_24771,N_24656);
xnor UO_1858 (O_1858,N_24726,N_24778);
nand UO_1859 (O_1859,N_24612,N_24597);
and UO_1860 (O_1860,N_24655,N_24644);
xor UO_1861 (O_1861,N_24674,N_24979);
and UO_1862 (O_1862,N_24513,N_24677);
and UO_1863 (O_1863,N_24585,N_24753);
nor UO_1864 (O_1864,N_24835,N_24564);
nand UO_1865 (O_1865,N_24941,N_24557);
nor UO_1866 (O_1866,N_24638,N_24960);
and UO_1867 (O_1867,N_24918,N_24545);
and UO_1868 (O_1868,N_24651,N_24766);
xor UO_1869 (O_1869,N_24971,N_24820);
nand UO_1870 (O_1870,N_24980,N_24752);
nand UO_1871 (O_1871,N_24952,N_24508);
nor UO_1872 (O_1872,N_24748,N_24686);
and UO_1873 (O_1873,N_24644,N_24749);
and UO_1874 (O_1874,N_24614,N_24716);
xnor UO_1875 (O_1875,N_24562,N_24564);
nand UO_1876 (O_1876,N_24900,N_24617);
and UO_1877 (O_1877,N_24725,N_24652);
and UO_1878 (O_1878,N_24807,N_24640);
nor UO_1879 (O_1879,N_24567,N_24981);
and UO_1880 (O_1880,N_24926,N_24921);
and UO_1881 (O_1881,N_24504,N_24968);
nand UO_1882 (O_1882,N_24902,N_24654);
nand UO_1883 (O_1883,N_24727,N_24663);
and UO_1884 (O_1884,N_24682,N_24601);
nor UO_1885 (O_1885,N_24528,N_24544);
and UO_1886 (O_1886,N_24517,N_24738);
and UO_1887 (O_1887,N_24757,N_24607);
xnor UO_1888 (O_1888,N_24879,N_24629);
nor UO_1889 (O_1889,N_24795,N_24700);
or UO_1890 (O_1890,N_24611,N_24729);
nand UO_1891 (O_1891,N_24572,N_24797);
nand UO_1892 (O_1892,N_24609,N_24799);
and UO_1893 (O_1893,N_24608,N_24987);
nand UO_1894 (O_1894,N_24778,N_24574);
nand UO_1895 (O_1895,N_24569,N_24602);
nand UO_1896 (O_1896,N_24581,N_24695);
xor UO_1897 (O_1897,N_24751,N_24909);
nand UO_1898 (O_1898,N_24887,N_24850);
or UO_1899 (O_1899,N_24628,N_24688);
or UO_1900 (O_1900,N_24991,N_24604);
and UO_1901 (O_1901,N_24975,N_24712);
nand UO_1902 (O_1902,N_24941,N_24787);
nor UO_1903 (O_1903,N_24785,N_24713);
or UO_1904 (O_1904,N_24522,N_24911);
xor UO_1905 (O_1905,N_24711,N_24799);
and UO_1906 (O_1906,N_24862,N_24763);
nand UO_1907 (O_1907,N_24683,N_24537);
or UO_1908 (O_1908,N_24656,N_24788);
nor UO_1909 (O_1909,N_24867,N_24668);
nor UO_1910 (O_1910,N_24663,N_24693);
nor UO_1911 (O_1911,N_24888,N_24795);
nor UO_1912 (O_1912,N_24663,N_24742);
nand UO_1913 (O_1913,N_24882,N_24817);
nand UO_1914 (O_1914,N_24558,N_24788);
xor UO_1915 (O_1915,N_24806,N_24535);
and UO_1916 (O_1916,N_24678,N_24527);
nor UO_1917 (O_1917,N_24644,N_24847);
and UO_1918 (O_1918,N_24635,N_24757);
or UO_1919 (O_1919,N_24952,N_24926);
nor UO_1920 (O_1920,N_24919,N_24638);
xor UO_1921 (O_1921,N_24608,N_24943);
or UO_1922 (O_1922,N_24559,N_24791);
and UO_1923 (O_1923,N_24713,N_24671);
nand UO_1924 (O_1924,N_24816,N_24861);
or UO_1925 (O_1925,N_24558,N_24833);
or UO_1926 (O_1926,N_24677,N_24588);
nand UO_1927 (O_1927,N_24555,N_24677);
and UO_1928 (O_1928,N_24530,N_24927);
nand UO_1929 (O_1929,N_24922,N_24891);
xnor UO_1930 (O_1930,N_24948,N_24992);
or UO_1931 (O_1931,N_24936,N_24540);
xor UO_1932 (O_1932,N_24877,N_24961);
xor UO_1933 (O_1933,N_24530,N_24944);
nand UO_1934 (O_1934,N_24724,N_24919);
nor UO_1935 (O_1935,N_24620,N_24888);
nand UO_1936 (O_1936,N_24645,N_24651);
xor UO_1937 (O_1937,N_24734,N_24694);
or UO_1938 (O_1938,N_24696,N_24807);
nor UO_1939 (O_1939,N_24532,N_24957);
nand UO_1940 (O_1940,N_24703,N_24573);
nand UO_1941 (O_1941,N_24820,N_24947);
nor UO_1942 (O_1942,N_24859,N_24564);
or UO_1943 (O_1943,N_24570,N_24949);
nor UO_1944 (O_1944,N_24908,N_24863);
nand UO_1945 (O_1945,N_24942,N_24836);
and UO_1946 (O_1946,N_24829,N_24672);
xnor UO_1947 (O_1947,N_24684,N_24826);
nor UO_1948 (O_1948,N_24899,N_24543);
nor UO_1949 (O_1949,N_24647,N_24865);
nand UO_1950 (O_1950,N_24582,N_24900);
nor UO_1951 (O_1951,N_24598,N_24581);
xnor UO_1952 (O_1952,N_24929,N_24956);
nand UO_1953 (O_1953,N_24920,N_24796);
nand UO_1954 (O_1954,N_24528,N_24852);
or UO_1955 (O_1955,N_24830,N_24508);
and UO_1956 (O_1956,N_24784,N_24880);
and UO_1957 (O_1957,N_24752,N_24512);
xor UO_1958 (O_1958,N_24716,N_24894);
or UO_1959 (O_1959,N_24850,N_24826);
nand UO_1960 (O_1960,N_24520,N_24840);
nor UO_1961 (O_1961,N_24570,N_24621);
nand UO_1962 (O_1962,N_24832,N_24841);
xnor UO_1963 (O_1963,N_24878,N_24789);
or UO_1964 (O_1964,N_24618,N_24772);
and UO_1965 (O_1965,N_24906,N_24728);
nor UO_1966 (O_1966,N_24832,N_24732);
or UO_1967 (O_1967,N_24821,N_24942);
nand UO_1968 (O_1968,N_24641,N_24950);
nand UO_1969 (O_1969,N_24512,N_24999);
nor UO_1970 (O_1970,N_24649,N_24653);
xnor UO_1971 (O_1971,N_24837,N_24964);
and UO_1972 (O_1972,N_24515,N_24774);
nand UO_1973 (O_1973,N_24840,N_24687);
xnor UO_1974 (O_1974,N_24542,N_24616);
nand UO_1975 (O_1975,N_24609,N_24771);
nand UO_1976 (O_1976,N_24663,N_24741);
xor UO_1977 (O_1977,N_24567,N_24594);
nor UO_1978 (O_1978,N_24900,N_24705);
or UO_1979 (O_1979,N_24975,N_24539);
nor UO_1980 (O_1980,N_24658,N_24543);
nor UO_1981 (O_1981,N_24828,N_24860);
nor UO_1982 (O_1982,N_24615,N_24742);
or UO_1983 (O_1983,N_24747,N_24694);
nor UO_1984 (O_1984,N_24635,N_24929);
nor UO_1985 (O_1985,N_24885,N_24743);
nand UO_1986 (O_1986,N_24953,N_24960);
nand UO_1987 (O_1987,N_24896,N_24581);
or UO_1988 (O_1988,N_24772,N_24631);
xor UO_1989 (O_1989,N_24835,N_24613);
nor UO_1990 (O_1990,N_24744,N_24895);
and UO_1991 (O_1991,N_24833,N_24857);
xnor UO_1992 (O_1992,N_24563,N_24526);
nor UO_1993 (O_1993,N_24775,N_24929);
xnor UO_1994 (O_1994,N_24775,N_24668);
nand UO_1995 (O_1995,N_24500,N_24503);
or UO_1996 (O_1996,N_24986,N_24655);
nor UO_1997 (O_1997,N_24907,N_24899);
and UO_1998 (O_1998,N_24501,N_24983);
or UO_1999 (O_1999,N_24796,N_24801);
nor UO_2000 (O_2000,N_24883,N_24599);
nor UO_2001 (O_2001,N_24666,N_24972);
nor UO_2002 (O_2002,N_24775,N_24664);
nor UO_2003 (O_2003,N_24558,N_24816);
nand UO_2004 (O_2004,N_24745,N_24694);
xnor UO_2005 (O_2005,N_24725,N_24667);
nand UO_2006 (O_2006,N_24686,N_24985);
xor UO_2007 (O_2007,N_24883,N_24596);
nand UO_2008 (O_2008,N_24789,N_24997);
or UO_2009 (O_2009,N_24729,N_24531);
or UO_2010 (O_2010,N_24581,N_24856);
nand UO_2011 (O_2011,N_24638,N_24853);
xor UO_2012 (O_2012,N_24975,N_24804);
or UO_2013 (O_2013,N_24818,N_24622);
xor UO_2014 (O_2014,N_24682,N_24880);
nand UO_2015 (O_2015,N_24732,N_24696);
nand UO_2016 (O_2016,N_24838,N_24651);
or UO_2017 (O_2017,N_24562,N_24830);
or UO_2018 (O_2018,N_24734,N_24981);
nor UO_2019 (O_2019,N_24989,N_24878);
nor UO_2020 (O_2020,N_24860,N_24503);
and UO_2021 (O_2021,N_24949,N_24723);
and UO_2022 (O_2022,N_24913,N_24776);
nor UO_2023 (O_2023,N_24999,N_24855);
nand UO_2024 (O_2024,N_24991,N_24903);
and UO_2025 (O_2025,N_24513,N_24999);
or UO_2026 (O_2026,N_24731,N_24529);
nor UO_2027 (O_2027,N_24731,N_24801);
or UO_2028 (O_2028,N_24961,N_24546);
nor UO_2029 (O_2029,N_24677,N_24574);
nand UO_2030 (O_2030,N_24614,N_24541);
nand UO_2031 (O_2031,N_24786,N_24867);
and UO_2032 (O_2032,N_24891,N_24510);
nand UO_2033 (O_2033,N_24820,N_24964);
and UO_2034 (O_2034,N_24806,N_24505);
nor UO_2035 (O_2035,N_24974,N_24608);
and UO_2036 (O_2036,N_24940,N_24747);
nor UO_2037 (O_2037,N_24889,N_24817);
or UO_2038 (O_2038,N_24803,N_24533);
and UO_2039 (O_2039,N_24969,N_24810);
or UO_2040 (O_2040,N_24891,N_24605);
and UO_2041 (O_2041,N_24617,N_24639);
nand UO_2042 (O_2042,N_24732,N_24607);
and UO_2043 (O_2043,N_24942,N_24947);
and UO_2044 (O_2044,N_24656,N_24746);
xor UO_2045 (O_2045,N_24537,N_24971);
and UO_2046 (O_2046,N_24509,N_24851);
nand UO_2047 (O_2047,N_24835,N_24863);
or UO_2048 (O_2048,N_24547,N_24550);
and UO_2049 (O_2049,N_24715,N_24991);
or UO_2050 (O_2050,N_24553,N_24991);
nor UO_2051 (O_2051,N_24887,N_24903);
xor UO_2052 (O_2052,N_24983,N_24607);
nand UO_2053 (O_2053,N_24545,N_24955);
or UO_2054 (O_2054,N_24957,N_24850);
and UO_2055 (O_2055,N_24645,N_24659);
nand UO_2056 (O_2056,N_24668,N_24556);
and UO_2057 (O_2057,N_24619,N_24723);
or UO_2058 (O_2058,N_24575,N_24979);
nand UO_2059 (O_2059,N_24995,N_24560);
or UO_2060 (O_2060,N_24567,N_24947);
and UO_2061 (O_2061,N_24500,N_24640);
and UO_2062 (O_2062,N_24552,N_24635);
or UO_2063 (O_2063,N_24684,N_24872);
xor UO_2064 (O_2064,N_24589,N_24962);
xor UO_2065 (O_2065,N_24640,N_24808);
xor UO_2066 (O_2066,N_24560,N_24965);
nand UO_2067 (O_2067,N_24751,N_24905);
or UO_2068 (O_2068,N_24700,N_24748);
nor UO_2069 (O_2069,N_24522,N_24688);
nor UO_2070 (O_2070,N_24896,N_24593);
xnor UO_2071 (O_2071,N_24858,N_24776);
xor UO_2072 (O_2072,N_24551,N_24676);
and UO_2073 (O_2073,N_24794,N_24942);
nand UO_2074 (O_2074,N_24776,N_24536);
nand UO_2075 (O_2075,N_24584,N_24690);
nor UO_2076 (O_2076,N_24677,N_24918);
xor UO_2077 (O_2077,N_24809,N_24772);
nand UO_2078 (O_2078,N_24686,N_24652);
nand UO_2079 (O_2079,N_24568,N_24541);
and UO_2080 (O_2080,N_24702,N_24921);
xnor UO_2081 (O_2081,N_24805,N_24754);
nand UO_2082 (O_2082,N_24830,N_24767);
or UO_2083 (O_2083,N_24517,N_24741);
and UO_2084 (O_2084,N_24704,N_24912);
or UO_2085 (O_2085,N_24606,N_24689);
nor UO_2086 (O_2086,N_24902,N_24950);
or UO_2087 (O_2087,N_24762,N_24843);
and UO_2088 (O_2088,N_24781,N_24957);
nand UO_2089 (O_2089,N_24893,N_24800);
xnor UO_2090 (O_2090,N_24552,N_24724);
or UO_2091 (O_2091,N_24638,N_24910);
nor UO_2092 (O_2092,N_24897,N_24537);
nor UO_2093 (O_2093,N_24634,N_24861);
xor UO_2094 (O_2094,N_24669,N_24925);
nand UO_2095 (O_2095,N_24798,N_24849);
nor UO_2096 (O_2096,N_24963,N_24532);
and UO_2097 (O_2097,N_24809,N_24975);
xor UO_2098 (O_2098,N_24576,N_24543);
nand UO_2099 (O_2099,N_24976,N_24596);
nand UO_2100 (O_2100,N_24798,N_24608);
and UO_2101 (O_2101,N_24855,N_24656);
nand UO_2102 (O_2102,N_24668,N_24531);
and UO_2103 (O_2103,N_24958,N_24759);
nor UO_2104 (O_2104,N_24934,N_24805);
xor UO_2105 (O_2105,N_24607,N_24763);
or UO_2106 (O_2106,N_24756,N_24911);
nand UO_2107 (O_2107,N_24999,N_24776);
nand UO_2108 (O_2108,N_24509,N_24985);
or UO_2109 (O_2109,N_24900,N_24894);
and UO_2110 (O_2110,N_24803,N_24574);
nor UO_2111 (O_2111,N_24836,N_24864);
or UO_2112 (O_2112,N_24691,N_24821);
nand UO_2113 (O_2113,N_24995,N_24548);
and UO_2114 (O_2114,N_24861,N_24909);
or UO_2115 (O_2115,N_24774,N_24519);
nor UO_2116 (O_2116,N_24520,N_24874);
nand UO_2117 (O_2117,N_24540,N_24830);
and UO_2118 (O_2118,N_24926,N_24917);
and UO_2119 (O_2119,N_24623,N_24519);
nor UO_2120 (O_2120,N_24533,N_24839);
xor UO_2121 (O_2121,N_24647,N_24707);
nor UO_2122 (O_2122,N_24937,N_24515);
nor UO_2123 (O_2123,N_24972,N_24721);
or UO_2124 (O_2124,N_24890,N_24530);
nand UO_2125 (O_2125,N_24748,N_24547);
nor UO_2126 (O_2126,N_24832,N_24855);
xnor UO_2127 (O_2127,N_24636,N_24928);
nand UO_2128 (O_2128,N_24828,N_24695);
nand UO_2129 (O_2129,N_24863,N_24569);
nand UO_2130 (O_2130,N_24778,N_24609);
or UO_2131 (O_2131,N_24820,N_24882);
xnor UO_2132 (O_2132,N_24720,N_24913);
nand UO_2133 (O_2133,N_24551,N_24623);
nor UO_2134 (O_2134,N_24756,N_24563);
or UO_2135 (O_2135,N_24504,N_24940);
or UO_2136 (O_2136,N_24868,N_24840);
xnor UO_2137 (O_2137,N_24649,N_24550);
xnor UO_2138 (O_2138,N_24703,N_24716);
nand UO_2139 (O_2139,N_24588,N_24974);
nand UO_2140 (O_2140,N_24623,N_24798);
and UO_2141 (O_2141,N_24866,N_24574);
nand UO_2142 (O_2142,N_24570,N_24654);
nor UO_2143 (O_2143,N_24501,N_24579);
and UO_2144 (O_2144,N_24754,N_24833);
and UO_2145 (O_2145,N_24782,N_24819);
nand UO_2146 (O_2146,N_24704,N_24945);
nand UO_2147 (O_2147,N_24978,N_24500);
nand UO_2148 (O_2148,N_24891,N_24786);
nor UO_2149 (O_2149,N_24981,N_24676);
or UO_2150 (O_2150,N_24529,N_24505);
nor UO_2151 (O_2151,N_24898,N_24523);
or UO_2152 (O_2152,N_24830,N_24689);
nand UO_2153 (O_2153,N_24581,N_24824);
or UO_2154 (O_2154,N_24507,N_24582);
xor UO_2155 (O_2155,N_24943,N_24601);
xnor UO_2156 (O_2156,N_24768,N_24679);
nor UO_2157 (O_2157,N_24605,N_24791);
nand UO_2158 (O_2158,N_24657,N_24956);
and UO_2159 (O_2159,N_24708,N_24727);
nand UO_2160 (O_2160,N_24507,N_24724);
xor UO_2161 (O_2161,N_24920,N_24615);
and UO_2162 (O_2162,N_24957,N_24988);
nand UO_2163 (O_2163,N_24893,N_24849);
nand UO_2164 (O_2164,N_24790,N_24767);
nor UO_2165 (O_2165,N_24872,N_24931);
xnor UO_2166 (O_2166,N_24820,N_24980);
nor UO_2167 (O_2167,N_24931,N_24932);
xor UO_2168 (O_2168,N_24526,N_24876);
xor UO_2169 (O_2169,N_24734,N_24517);
or UO_2170 (O_2170,N_24719,N_24953);
and UO_2171 (O_2171,N_24837,N_24876);
and UO_2172 (O_2172,N_24713,N_24730);
nand UO_2173 (O_2173,N_24513,N_24699);
or UO_2174 (O_2174,N_24909,N_24887);
nor UO_2175 (O_2175,N_24912,N_24765);
or UO_2176 (O_2176,N_24659,N_24813);
nand UO_2177 (O_2177,N_24569,N_24824);
xnor UO_2178 (O_2178,N_24615,N_24797);
or UO_2179 (O_2179,N_24869,N_24559);
nor UO_2180 (O_2180,N_24921,N_24617);
or UO_2181 (O_2181,N_24653,N_24656);
or UO_2182 (O_2182,N_24694,N_24758);
and UO_2183 (O_2183,N_24933,N_24545);
and UO_2184 (O_2184,N_24642,N_24543);
and UO_2185 (O_2185,N_24629,N_24849);
xnor UO_2186 (O_2186,N_24502,N_24652);
xor UO_2187 (O_2187,N_24862,N_24538);
nor UO_2188 (O_2188,N_24869,N_24899);
nand UO_2189 (O_2189,N_24733,N_24738);
or UO_2190 (O_2190,N_24767,N_24661);
nand UO_2191 (O_2191,N_24900,N_24748);
xnor UO_2192 (O_2192,N_24552,N_24890);
and UO_2193 (O_2193,N_24901,N_24669);
or UO_2194 (O_2194,N_24586,N_24619);
and UO_2195 (O_2195,N_24613,N_24522);
and UO_2196 (O_2196,N_24630,N_24564);
nand UO_2197 (O_2197,N_24592,N_24735);
or UO_2198 (O_2198,N_24595,N_24931);
and UO_2199 (O_2199,N_24766,N_24602);
or UO_2200 (O_2200,N_24736,N_24697);
nand UO_2201 (O_2201,N_24805,N_24532);
nor UO_2202 (O_2202,N_24861,N_24702);
and UO_2203 (O_2203,N_24728,N_24960);
nor UO_2204 (O_2204,N_24847,N_24513);
xnor UO_2205 (O_2205,N_24941,N_24952);
nor UO_2206 (O_2206,N_24724,N_24901);
or UO_2207 (O_2207,N_24784,N_24868);
nor UO_2208 (O_2208,N_24630,N_24771);
nor UO_2209 (O_2209,N_24706,N_24930);
and UO_2210 (O_2210,N_24837,N_24887);
or UO_2211 (O_2211,N_24792,N_24727);
or UO_2212 (O_2212,N_24871,N_24917);
and UO_2213 (O_2213,N_24879,N_24862);
xor UO_2214 (O_2214,N_24938,N_24782);
nand UO_2215 (O_2215,N_24917,N_24815);
or UO_2216 (O_2216,N_24981,N_24932);
nor UO_2217 (O_2217,N_24593,N_24772);
nor UO_2218 (O_2218,N_24660,N_24906);
nor UO_2219 (O_2219,N_24544,N_24771);
xor UO_2220 (O_2220,N_24990,N_24931);
or UO_2221 (O_2221,N_24655,N_24529);
and UO_2222 (O_2222,N_24932,N_24873);
xnor UO_2223 (O_2223,N_24914,N_24678);
nor UO_2224 (O_2224,N_24512,N_24759);
nor UO_2225 (O_2225,N_24625,N_24687);
xnor UO_2226 (O_2226,N_24520,N_24839);
and UO_2227 (O_2227,N_24608,N_24654);
xor UO_2228 (O_2228,N_24871,N_24522);
nand UO_2229 (O_2229,N_24957,N_24672);
nor UO_2230 (O_2230,N_24601,N_24566);
nor UO_2231 (O_2231,N_24817,N_24521);
nor UO_2232 (O_2232,N_24977,N_24943);
nand UO_2233 (O_2233,N_24561,N_24598);
and UO_2234 (O_2234,N_24987,N_24709);
nor UO_2235 (O_2235,N_24866,N_24740);
and UO_2236 (O_2236,N_24946,N_24630);
nand UO_2237 (O_2237,N_24614,N_24546);
nand UO_2238 (O_2238,N_24953,N_24930);
or UO_2239 (O_2239,N_24549,N_24757);
nand UO_2240 (O_2240,N_24830,N_24949);
nor UO_2241 (O_2241,N_24725,N_24772);
and UO_2242 (O_2242,N_24798,N_24925);
xor UO_2243 (O_2243,N_24803,N_24572);
or UO_2244 (O_2244,N_24897,N_24975);
or UO_2245 (O_2245,N_24792,N_24582);
xor UO_2246 (O_2246,N_24537,N_24620);
nand UO_2247 (O_2247,N_24694,N_24844);
xnor UO_2248 (O_2248,N_24913,N_24565);
xor UO_2249 (O_2249,N_24967,N_24653);
and UO_2250 (O_2250,N_24735,N_24672);
xor UO_2251 (O_2251,N_24831,N_24791);
xor UO_2252 (O_2252,N_24600,N_24810);
or UO_2253 (O_2253,N_24733,N_24568);
xnor UO_2254 (O_2254,N_24700,N_24781);
nand UO_2255 (O_2255,N_24578,N_24992);
nand UO_2256 (O_2256,N_24517,N_24990);
or UO_2257 (O_2257,N_24989,N_24570);
nor UO_2258 (O_2258,N_24795,N_24670);
and UO_2259 (O_2259,N_24942,N_24594);
and UO_2260 (O_2260,N_24504,N_24942);
and UO_2261 (O_2261,N_24531,N_24816);
or UO_2262 (O_2262,N_24603,N_24539);
nor UO_2263 (O_2263,N_24840,N_24894);
nor UO_2264 (O_2264,N_24512,N_24579);
or UO_2265 (O_2265,N_24891,N_24881);
and UO_2266 (O_2266,N_24956,N_24842);
or UO_2267 (O_2267,N_24863,N_24887);
or UO_2268 (O_2268,N_24790,N_24858);
or UO_2269 (O_2269,N_24849,N_24566);
nand UO_2270 (O_2270,N_24813,N_24542);
or UO_2271 (O_2271,N_24984,N_24558);
nand UO_2272 (O_2272,N_24768,N_24892);
or UO_2273 (O_2273,N_24662,N_24943);
and UO_2274 (O_2274,N_24982,N_24680);
or UO_2275 (O_2275,N_24547,N_24857);
nor UO_2276 (O_2276,N_24598,N_24791);
nand UO_2277 (O_2277,N_24853,N_24855);
nand UO_2278 (O_2278,N_24797,N_24995);
and UO_2279 (O_2279,N_24533,N_24979);
or UO_2280 (O_2280,N_24715,N_24716);
or UO_2281 (O_2281,N_24709,N_24965);
nor UO_2282 (O_2282,N_24519,N_24901);
or UO_2283 (O_2283,N_24634,N_24757);
nand UO_2284 (O_2284,N_24992,N_24579);
nor UO_2285 (O_2285,N_24904,N_24567);
nand UO_2286 (O_2286,N_24866,N_24949);
xnor UO_2287 (O_2287,N_24552,N_24980);
or UO_2288 (O_2288,N_24506,N_24714);
xnor UO_2289 (O_2289,N_24774,N_24848);
xor UO_2290 (O_2290,N_24555,N_24508);
nor UO_2291 (O_2291,N_24894,N_24769);
or UO_2292 (O_2292,N_24611,N_24963);
xor UO_2293 (O_2293,N_24641,N_24847);
nand UO_2294 (O_2294,N_24587,N_24549);
and UO_2295 (O_2295,N_24665,N_24905);
and UO_2296 (O_2296,N_24772,N_24549);
nor UO_2297 (O_2297,N_24567,N_24805);
or UO_2298 (O_2298,N_24853,N_24863);
or UO_2299 (O_2299,N_24843,N_24780);
nor UO_2300 (O_2300,N_24650,N_24978);
xnor UO_2301 (O_2301,N_24717,N_24773);
xnor UO_2302 (O_2302,N_24501,N_24900);
and UO_2303 (O_2303,N_24661,N_24727);
and UO_2304 (O_2304,N_24949,N_24992);
and UO_2305 (O_2305,N_24905,N_24899);
nand UO_2306 (O_2306,N_24643,N_24624);
nor UO_2307 (O_2307,N_24575,N_24980);
xor UO_2308 (O_2308,N_24726,N_24529);
xor UO_2309 (O_2309,N_24948,N_24511);
nor UO_2310 (O_2310,N_24870,N_24584);
xor UO_2311 (O_2311,N_24637,N_24918);
nand UO_2312 (O_2312,N_24892,N_24555);
nand UO_2313 (O_2313,N_24672,N_24901);
nor UO_2314 (O_2314,N_24898,N_24871);
xor UO_2315 (O_2315,N_24714,N_24511);
nand UO_2316 (O_2316,N_24928,N_24551);
xnor UO_2317 (O_2317,N_24610,N_24818);
xor UO_2318 (O_2318,N_24962,N_24831);
or UO_2319 (O_2319,N_24656,N_24796);
xor UO_2320 (O_2320,N_24644,N_24542);
xor UO_2321 (O_2321,N_24773,N_24795);
nand UO_2322 (O_2322,N_24685,N_24536);
nand UO_2323 (O_2323,N_24962,N_24606);
and UO_2324 (O_2324,N_24562,N_24824);
and UO_2325 (O_2325,N_24678,N_24679);
or UO_2326 (O_2326,N_24840,N_24649);
and UO_2327 (O_2327,N_24566,N_24675);
nand UO_2328 (O_2328,N_24833,N_24967);
nand UO_2329 (O_2329,N_24550,N_24583);
nor UO_2330 (O_2330,N_24638,N_24774);
and UO_2331 (O_2331,N_24793,N_24736);
and UO_2332 (O_2332,N_24529,N_24764);
nor UO_2333 (O_2333,N_24986,N_24565);
nor UO_2334 (O_2334,N_24500,N_24947);
and UO_2335 (O_2335,N_24629,N_24926);
and UO_2336 (O_2336,N_24764,N_24788);
and UO_2337 (O_2337,N_24688,N_24503);
xor UO_2338 (O_2338,N_24686,N_24707);
xnor UO_2339 (O_2339,N_24916,N_24607);
xor UO_2340 (O_2340,N_24806,N_24962);
xnor UO_2341 (O_2341,N_24990,N_24967);
nor UO_2342 (O_2342,N_24827,N_24516);
and UO_2343 (O_2343,N_24774,N_24803);
nand UO_2344 (O_2344,N_24745,N_24851);
nor UO_2345 (O_2345,N_24659,N_24989);
nor UO_2346 (O_2346,N_24966,N_24869);
nor UO_2347 (O_2347,N_24539,N_24968);
nand UO_2348 (O_2348,N_24576,N_24579);
or UO_2349 (O_2349,N_24863,N_24536);
xor UO_2350 (O_2350,N_24642,N_24708);
nand UO_2351 (O_2351,N_24708,N_24615);
nor UO_2352 (O_2352,N_24747,N_24634);
and UO_2353 (O_2353,N_24853,N_24623);
xor UO_2354 (O_2354,N_24654,N_24749);
xor UO_2355 (O_2355,N_24832,N_24947);
nand UO_2356 (O_2356,N_24541,N_24972);
or UO_2357 (O_2357,N_24886,N_24970);
nor UO_2358 (O_2358,N_24926,N_24766);
and UO_2359 (O_2359,N_24984,N_24892);
nand UO_2360 (O_2360,N_24592,N_24955);
and UO_2361 (O_2361,N_24887,N_24566);
and UO_2362 (O_2362,N_24570,N_24626);
nand UO_2363 (O_2363,N_24619,N_24640);
nand UO_2364 (O_2364,N_24689,N_24562);
or UO_2365 (O_2365,N_24772,N_24633);
xnor UO_2366 (O_2366,N_24718,N_24612);
or UO_2367 (O_2367,N_24504,N_24945);
and UO_2368 (O_2368,N_24837,N_24632);
and UO_2369 (O_2369,N_24944,N_24871);
xnor UO_2370 (O_2370,N_24590,N_24913);
xnor UO_2371 (O_2371,N_24981,N_24607);
or UO_2372 (O_2372,N_24866,N_24979);
nand UO_2373 (O_2373,N_24888,N_24828);
nand UO_2374 (O_2374,N_24849,N_24621);
nand UO_2375 (O_2375,N_24786,N_24748);
and UO_2376 (O_2376,N_24960,N_24711);
or UO_2377 (O_2377,N_24764,N_24601);
nor UO_2378 (O_2378,N_24656,N_24821);
xnor UO_2379 (O_2379,N_24604,N_24603);
or UO_2380 (O_2380,N_24596,N_24628);
nor UO_2381 (O_2381,N_24630,N_24905);
nand UO_2382 (O_2382,N_24635,N_24617);
and UO_2383 (O_2383,N_24785,N_24911);
or UO_2384 (O_2384,N_24672,N_24613);
xor UO_2385 (O_2385,N_24710,N_24898);
or UO_2386 (O_2386,N_24919,N_24978);
nand UO_2387 (O_2387,N_24889,N_24578);
nand UO_2388 (O_2388,N_24704,N_24551);
nand UO_2389 (O_2389,N_24564,N_24889);
xnor UO_2390 (O_2390,N_24971,N_24844);
nor UO_2391 (O_2391,N_24682,N_24875);
xor UO_2392 (O_2392,N_24799,N_24672);
and UO_2393 (O_2393,N_24692,N_24950);
xor UO_2394 (O_2394,N_24545,N_24891);
and UO_2395 (O_2395,N_24521,N_24877);
or UO_2396 (O_2396,N_24818,N_24555);
nor UO_2397 (O_2397,N_24942,N_24759);
nand UO_2398 (O_2398,N_24917,N_24997);
and UO_2399 (O_2399,N_24823,N_24706);
nand UO_2400 (O_2400,N_24623,N_24851);
nor UO_2401 (O_2401,N_24959,N_24829);
nor UO_2402 (O_2402,N_24737,N_24884);
or UO_2403 (O_2403,N_24644,N_24582);
xnor UO_2404 (O_2404,N_24562,N_24668);
nand UO_2405 (O_2405,N_24843,N_24863);
nand UO_2406 (O_2406,N_24729,N_24648);
xnor UO_2407 (O_2407,N_24900,N_24794);
nand UO_2408 (O_2408,N_24860,N_24900);
and UO_2409 (O_2409,N_24932,N_24668);
nand UO_2410 (O_2410,N_24704,N_24723);
nor UO_2411 (O_2411,N_24852,N_24738);
and UO_2412 (O_2412,N_24695,N_24932);
and UO_2413 (O_2413,N_24825,N_24873);
nand UO_2414 (O_2414,N_24502,N_24672);
or UO_2415 (O_2415,N_24923,N_24790);
or UO_2416 (O_2416,N_24604,N_24715);
nor UO_2417 (O_2417,N_24634,N_24565);
nor UO_2418 (O_2418,N_24538,N_24670);
nor UO_2419 (O_2419,N_24781,N_24863);
xor UO_2420 (O_2420,N_24913,N_24657);
nor UO_2421 (O_2421,N_24912,N_24572);
nor UO_2422 (O_2422,N_24849,N_24735);
nor UO_2423 (O_2423,N_24987,N_24962);
nand UO_2424 (O_2424,N_24902,N_24575);
and UO_2425 (O_2425,N_24734,N_24698);
xnor UO_2426 (O_2426,N_24766,N_24695);
and UO_2427 (O_2427,N_24647,N_24742);
xor UO_2428 (O_2428,N_24508,N_24800);
xor UO_2429 (O_2429,N_24726,N_24583);
or UO_2430 (O_2430,N_24836,N_24813);
xor UO_2431 (O_2431,N_24782,N_24893);
xor UO_2432 (O_2432,N_24868,N_24763);
and UO_2433 (O_2433,N_24738,N_24776);
xor UO_2434 (O_2434,N_24620,N_24588);
nor UO_2435 (O_2435,N_24971,N_24940);
and UO_2436 (O_2436,N_24828,N_24914);
xnor UO_2437 (O_2437,N_24545,N_24860);
or UO_2438 (O_2438,N_24632,N_24737);
or UO_2439 (O_2439,N_24543,N_24788);
nor UO_2440 (O_2440,N_24865,N_24586);
xor UO_2441 (O_2441,N_24866,N_24737);
nor UO_2442 (O_2442,N_24611,N_24609);
and UO_2443 (O_2443,N_24556,N_24970);
and UO_2444 (O_2444,N_24677,N_24837);
and UO_2445 (O_2445,N_24783,N_24509);
nor UO_2446 (O_2446,N_24827,N_24649);
nand UO_2447 (O_2447,N_24927,N_24902);
or UO_2448 (O_2448,N_24981,N_24572);
or UO_2449 (O_2449,N_24820,N_24707);
xnor UO_2450 (O_2450,N_24751,N_24913);
and UO_2451 (O_2451,N_24518,N_24886);
nand UO_2452 (O_2452,N_24562,N_24643);
nand UO_2453 (O_2453,N_24911,N_24743);
nand UO_2454 (O_2454,N_24720,N_24807);
nand UO_2455 (O_2455,N_24555,N_24711);
or UO_2456 (O_2456,N_24986,N_24668);
or UO_2457 (O_2457,N_24715,N_24645);
nand UO_2458 (O_2458,N_24744,N_24634);
or UO_2459 (O_2459,N_24854,N_24500);
and UO_2460 (O_2460,N_24951,N_24602);
nand UO_2461 (O_2461,N_24701,N_24893);
or UO_2462 (O_2462,N_24788,N_24599);
xor UO_2463 (O_2463,N_24879,N_24628);
nor UO_2464 (O_2464,N_24660,N_24631);
xor UO_2465 (O_2465,N_24541,N_24747);
nor UO_2466 (O_2466,N_24684,N_24652);
xor UO_2467 (O_2467,N_24979,N_24543);
nand UO_2468 (O_2468,N_24729,N_24646);
nor UO_2469 (O_2469,N_24641,N_24501);
nand UO_2470 (O_2470,N_24966,N_24819);
or UO_2471 (O_2471,N_24627,N_24921);
and UO_2472 (O_2472,N_24557,N_24830);
nor UO_2473 (O_2473,N_24974,N_24805);
nand UO_2474 (O_2474,N_24577,N_24695);
xnor UO_2475 (O_2475,N_24977,N_24722);
and UO_2476 (O_2476,N_24733,N_24653);
and UO_2477 (O_2477,N_24843,N_24570);
or UO_2478 (O_2478,N_24537,N_24810);
or UO_2479 (O_2479,N_24585,N_24584);
nor UO_2480 (O_2480,N_24818,N_24596);
nor UO_2481 (O_2481,N_24831,N_24649);
nand UO_2482 (O_2482,N_24880,N_24982);
xnor UO_2483 (O_2483,N_24808,N_24944);
xor UO_2484 (O_2484,N_24922,N_24596);
xor UO_2485 (O_2485,N_24737,N_24546);
xnor UO_2486 (O_2486,N_24795,N_24804);
nand UO_2487 (O_2487,N_24736,N_24558);
nand UO_2488 (O_2488,N_24697,N_24754);
or UO_2489 (O_2489,N_24575,N_24797);
nor UO_2490 (O_2490,N_24745,N_24670);
xor UO_2491 (O_2491,N_24638,N_24757);
xor UO_2492 (O_2492,N_24951,N_24609);
and UO_2493 (O_2493,N_24870,N_24777);
and UO_2494 (O_2494,N_24957,N_24906);
or UO_2495 (O_2495,N_24568,N_24741);
nor UO_2496 (O_2496,N_24624,N_24507);
and UO_2497 (O_2497,N_24757,N_24642);
nand UO_2498 (O_2498,N_24676,N_24815);
nand UO_2499 (O_2499,N_24822,N_24842);
or UO_2500 (O_2500,N_24811,N_24898);
and UO_2501 (O_2501,N_24623,N_24785);
xnor UO_2502 (O_2502,N_24540,N_24505);
nor UO_2503 (O_2503,N_24512,N_24815);
xnor UO_2504 (O_2504,N_24989,N_24734);
and UO_2505 (O_2505,N_24623,N_24576);
and UO_2506 (O_2506,N_24875,N_24850);
and UO_2507 (O_2507,N_24961,N_24509);
or UO_2508 (O_2508,N_24692,N_24787);
nand UO_2509 (O_2509,N_24903,N_24852);
nor UO_2510 (O_2510,N_24961,N_24561);
xor UO_2511 (O_2511,N_24930,N_24747);
xor UO_2512 (O_2512,N_24722,N_24902);
or UO_2513 (O_2513,N_24915,N_24605);
nand UO_2514 (O_2514,N_24886,N_24784);
nand UO_2515 (O_2515,N_24666,N_24502);
or UO_2516 (O_2516,N_24969,N_24994);
nor UO_2517 (O_2517,N_24709,N_24819);
nand UO_2518 (O_2518,N_24594,N_24628);
nand UO_2519 (O_2519,N_24760,N_24860);
and UO_2520 (O_2520,N_24597,N_24980);
nand UO_2521 (O_2521,N_24969,N_24812);
or UO_2522 (O_2522,N_24806,N_24637);
nor UO_2523 (O_2523,N_24662,N_24836);
nor UO_2524 (O_2524,N_24616,N_24952);
nand UO_2525 (O_2525,N_24548,N_24669);
or UO_2526 (O_2526,N_24658,N_24734);
nand UO_2527 (O_2527,N_24816,N_24916);
nor UO_2528 (O_2528,N_24714,N_24602);
xnor UO_2529 (O_2529,N_24734,N_24628);
xnor UO_2530 (O_2530,N_24752,N_24664);
nor UO_2531 (O_2531,N_24996,N_24960);
and UO_2532 (O_2532,N_24639,N_24901);
nand UO_2533 (O_2533,N_24508,N_24905);
nor UO_2534 (O_2534,N_24545,N_24754);
and UO_2535 (O_2535,N_24870,N_24501);
xnor UO_2536 (O_2536,N_24850,N_24510);
xnor UO_2537 (O_2537,N_24852,N_24908);
xor UO_2538 (O_2538,N_24658,N_24850);
nor UO_2539 (O_2539,N_24537,N_24588);
nand UO_2540 (O_2540,N_24570,N_24861);
nand UO_2541 (O_2541,N_24659,N_24683);
nand UO_2542 (O_2542,N_24732,N_24855);
xnor UO_2543 (O_2543,N_24504,N_24846);
and UO_2544 (O_2544,N_24843,N_24835);
or UO_2545 (O_2545,N_24805,N_24972);
or UO_2546 (O_2546,N_24806,N_24582);
nor UO_2547 (O_2547,N_24733,N_24561);
nand UO_2548 (O_2548,N_24933,N_24775);
or UO_2549 (O_2549,N_24693,N_24543);
and UO_2550 (O_2550,N_24922,N_24547);
nand UO_2551 (O_2551,N_24526,N_24516);
nor UO_2552 (O_2552,N_24963,N_24518);
or UO_2553 (O_2553,N_24728,N_24551);
and UO_2554 (O_2554,N_24598,N_24651);
and UO_2555 (O_2555,N_24582,N_24672);
or UO_2556 (O_2556,N_24504,N_24783);
or UO_2557 (O_2557,N_24809,N_24613);
and UO_2558 (O_2558,N_24680,N_24990);
nand UO_2559 (O_2559,N_24618,N_24676);
nor UO_2560 (O_2560,N_24548,N_24791);
nor UO_2561 (O_2561,N_24955,N_24700);
or UO_2562 (O_2562,N_24784,N_24825);
xnor UO_2563 (O_2563,N_24912,N_24715);
or UO_2564 (O_2564,N_24940,N_24666);
and UO_2565 (O_2565,N_24824,N_24978);
xnor UO_2566 (O_2566,N_24854,N_24992);
and UO_2567 (O_2567,N_24973,N_24880);
xor UO_2568 (O_2568,N_24978,N_24782);
and UO_2569 (O_2569,N_24667,N_24617);
nor UO_2570 (O_2570,N_24847,N_24648);
nor UO_2571 (O_2571,N_24929,N_24621);
nand UO_2572 (O_2572,N_24843,N_24998);
nand UO_2573 (O_2573,N_24610,N_24900);
xor UO_2574 (O_2574,N_24919,N_24962);
xnor UO_2575 (O_2575,N_24758,N_24861);
xnor UO_2576 (O_2576,N_24939,N_24763);
nor UO_2577 (O_2577,N_24671,N_24946);
nor UO_2578 (O_2578,N_24521,N_24646);
or UO_2579 (O_2579,N_24703,N_24924);
and UO_2580 (O_2580,N_24566,N_24664);
or UO_2581 (O_2581,N_24675,N_24585);
nor UO_2582 (O_2582,N_24912,N_24582);
or UO_2583 (O_2583,N_24793,N_24650);
nor UO_2584 (O_2584,N_24659,N_24903);
nand UO_2585 (O_2585,N_24815,N_24942);
nand UO_2586 (O_2586,N_24899,N_24875);
and UO_2587 (O_2587,N_24894,N_24661);
nand UO_2588 (O_2588,N_24549,N_24852);
and UO_2589 (O_2589,N_24523,N_24922);
nor UO_2590 (O_2590,N_24855,N_24580);
nand UO_2591 (O_2591,N_24557,N_24630);
xor UO_2592 (O_2592,N_24662,N_24819);
or UO_2593 (O_2593,N_24646,N_24617);
and UO_2594 (O_2594,N_24998,N_24693);
and UO_2595 (O_2595,N_24919,N_24770);
xor UO_2596 (O_2596,N_24562,N_24590);
and UO_2597 (O_2597,N_24593,N_24820);
and UO_2598 (O_2598,N_24584,N_24963);
and UO_2599 (O_2599,N_24990,N_24866);
xnor UO_2600 (O_2600,N_24904,N_24959);
xor UO_2601 (O_2601,N_24622,N_24969);
or UO_2602 (O_2602,N_24846,N_24996);
nor UO_2603 (O_2603,N_24795,N_24550);
nor UO_2604 (O_2604,N_24714,N_24913);
xnor UO_2605 (O_2605,N_24981,N_24772);
or UO_2606 (O_2606,N_24976,N_24652);
nand UO_2607 (O_2607,N_24832,N_24637);
nor UO_2608 (O_2608,N_24956,N_24654);
or UO_2609 (O_2609,N_24568,N_24863);
and UO_2610 (O_2610,N_24849,N_24520);
and UO_2611 (O_2611,N_24840,N_24695);
nand UO_2612 (O_2612,N_24737,N_24878);
nor UO_2613 (O_2613,N_24681,N_24949);
xnor UO_2614 (O_2614,N_24807,N_24579);
or UO_2615 (O_2615,N_24864,N_24845);
xnor UO_2616 (O_2616,N_24977,N_24669);
nor UO_2617 (O_2617,N_24773,N_24720);
or UO_2618 (O_2618,N_24751,N_24513);
or UO_2619 (O_2619,N_24872,N_24780);
nor UO_2620 (O_2620,N_24553,N_24718);
nor UO_2621 (O_2621,N_24926,N_24795);
nor UO_2622 (O_2622,N_24554,N_24901);
xnor UO_2623 (O_2623,N_24665,N_24690);
nand UO_2624 (O_2624,N_24620,N_24632);
or UO_2625 (O_2625,N_24530,N_24653);
or UO_2626 (O_2626,N_24810,N_24987);
and UO_2627 (O_2627,N_24831,N_24621);
and UO_2628 (O_2628,N_24842,N_24714);
nor UO_2629 (O_2629,N_24926,N_24858);
nand UO_2630 (O_2630,N_24671,N_24955);
nor UO_2631 (O_2631,N_24568,N_24549);
xnor UO_2632 (O_2632,N_24612,N_24995);
xnor UO_2633 (O_2633,N_24930,N_24760);
nor UO_2634 (O_2634,N_24717,N_24949);
and UO_2635 (O_2635,N_24514,N_24934);
or UO_2636 (O_2636,N_24647,N_24659);
nand UO_2637 (O_2637,N_24723,N_24631);
xor UO_2638 (O_2638,N_24576,N_24910);
nor UO_2639 (O_2639,N_24954,N_24698);
nor UO_2640 (O_2640,N_24857,N_24732);
xnor UO_2641 (O_2641,N_24997,N_24838);
nor UO_2642 (O_2642,N_24867,N_24526);
nand UO_2643 (O_2643,N_24775,N_24618);
or UO_2644 (O_2644,N_24592,N_24715);
and UO_2645 (O_2645,N_24724,N_24617);
and UO_2646 (O_2646,N_24563,N_24727);
or UO_2647 (O_2647,N_24817,N_24955);
or UO_2648 (O_2648,N_24922,N_24962);
xnor UO_2649 (O_2649,N_24593,N_24881);
nand UO_2650 (O_2650,N_24608,N_24551);
nand UO_2651 (O_2651,N_24988,N_24902);
nand UO_2652 (O_2652,N_24666,N_24743);
and UO_2653 (O_2653,N_24890,N_24735);
and UO_2654 (O_2654,N_24576,N_24853);
nor UO_2655 (O_2655,N_24500,N_24540);
xnor UO_2656 (O_2656,N_24803,N_24619);
xnor UO_2657 (O_2657,N_24807,N_24860);
xor UO_2658 (O_2658,N_24781,N_24730);
nor UO_2659 (O_2659,N_24546,N_24599);
or UO_2660 (O_2660,N_24626,N_24721);
xor UO_2661 (O_2661,N_24758,N_24655);
xnor UO_2662 (O_2662,N_24717,N_24774);
or UO_2663 (O_2663,N_24661,N_24901);
xnor UO_2664 (O_2664,N_24983,N_24699);
nand UO_2665 (O_2665,N_24668,N_24520);
nand UO_2666 (O_2666,N_24528,N_24525);
and UO_2667 (O_2667,N_24739,N_24857);
nor UO_2668 (O_2668,N_24574,N_24746);
xor UO_2669 (O_2669,N_24854,N_24935);
xnor UO_2670 (O_2670,N_24657,N_24639);
nand UO_2671 (O_2671,N_24504,N_24708);
xor UO_2672 (O_2672,N_24735,N_24808);
and UO_2673 (O_2673,N_24568,N_24900);
or UO_2674 (O_2674,N_24907,N_24967);
nand UO_2675 (O_2675,N_24873,N_24720);
nand UO_2676 (O_2676,N_24765,N_24741);
nor UO_2677 (O_2677,N_24573,N_24513);
and UO_2678 (O_2678,N_24832,N_24597);
nand UO_2679 (O_2679,N_24620,N_24855);
nor UO_2680 (O_2680,N_24730,N_24508);
and UO_2681 (O_2681,N_24653,N_24845);
or UO_2682 (O_2682,N_24633,N_24926);
xnor UO_2683 (O_2683,N_24933,N_24704);
and UO_2684 (O_2684,N_24601,N_24683);
xnor UO_2685 (O_2685,N_24940,N_24848);
nor UO_2686 (O_2686,N_24829,N_24679);
nand UO_2687 (O_2687,N_24837,N_24590);
nor UO_2688 (O_2688,N_24728,N_24881);
xor UO_2689 (O_2689,N_24643,N_24638);
and UO_2690 (O_2690,N_24636,N_24632);
and UO_2691 (O_2691,N_24930,N_24609);
and UO_2692 (O_2692,N_24827,N_24605);
nor UO_2693 (O_2693,N_24546,N_24919);
or UO_2694 (O_2694,N_24571,N_24686);
nor UO_2695 (O_2695,N_24582,N_24771);
and UO_2696 (O_2696,N_24590,N_24765);
xor UO_2697 (O_2697,N_24692,N_24648);
nor UO_2698 (O_2698,N_24821,N_24953);
or UO_2699 (O_2699,N_24869,N_24557);
xor UO_2700 (O_2700,N_24644,N_24639);
xor UO_2701 (O_2701,N_24651,N_24889);
and UO_2702 (O_2702,N_24559,N_24713);
xor UO_2703 (O_2703,N_24735,N_24792);
or UO_2704 (O_2704,N_24876,N_24934);
nor UO_2705 (O_2705,N_24740,N_24842);
or UO_2706 (O_2706,N_24858,N_24675);
nand UO_2707 (O_2707,N_24522,N_24548);
or UO_2708 (O_2708,N_24599,N_24610);
and UO_2709 (O_2709,N_24590,N_24619);
nor UO_2710 (O_2710,N_24663,N_24503);
nor UO_2711 (O_2711,N_24966,N_24645);
nor UO_2712 (O_2712,N_24735,N_24859);
xnor UO_2713 (O_2713,N_24714,N_24856);
and UO_2714 (O_2714,N_24684,N_24507);
xor UO_2715 (O_2715,N_24841,N_24975);
xor UO_2716 (O_2716,N_24804,N_24811);
or UO_2717 (O_2717,N_24601,N_24949);
nand UO_2718 (O_2718,N_24888,N_24822);
nand UO_2719 (O_2719,N_24513,N_24709);
nand UO_2720 (O_2720,N_24842,N_24578);
xnor UO_2721 (O_2721,N_24761,N_24749);
nor UO_2722 (O_2722,N_24790,N_24663);
nand UO_2723 (O_2723,N_24590,N_24605);
nand UO_2724 (O_2724,N_24993,N_24936);
and UO_2725 (O_2725,N_24812,N_24637);
and UO_2726 (O_2726,N_24508,N_24995);
nor UO_2727 (O_2727,N_24786,N_24974);
nand UO_2728 (O_2728,N_24776,N_24611);
xor UO_2729 (O_2729,N_24903,N_24668);
xor UO_2730 (O_2730,N_24814,N_24536);
nand UO_2731 (O_2731,N_24921,N_24622);
nor UO_2732 (O_2732,N_24903,N_24970);
and UO_2733 (O_2733,N_24748,N_24574);
nand UO_2734 (O_2734,N_24731,N_24972);
xor UO_2735 (O_2735,N_24869,N_24674);
or UO_2736 (O_2736,N_24686,N_24857);
xor UO_2737 (O_2737,N_24931,N_24847);
nand UO_2738 (O_2738,N_24767,N_24561);
and UO_2739 (O_2739,N_24883,N_24715);
nand UO_2740 (O_2740,N_24809,N_24956);
or UO_2741 (O_2741,N_24543,N_24841);
nor UO_2742 (O_2742,N_24734,N_24866);
xor UO_2743 (O_2743,N_24525,N_24790);
nor UO_2744 (O_2744,N_24673,N_24815);
xor UO_2745 (O_2745,N_24591,N_24706);
or UO_2746 (O_2746,N_24955,N_24791);
nor UO_2747 (O_2747,N_24923,N_24920);
or UO_2748 (O_2748,N_24838,N_24890);
or UO_2749 (O_2749,N_24702,N_24687);
or UO_2750 (O_2750,N_24719,N_24641);
xor UO_2751 (O_2751,N_24507,N_24511);
nand UO_2752 (O_2752,N_24563,N_24769);
xnor UO_2753 (O_2753,N_24757,N_24652);
nand UO_2754 (O_2754,N_24621,N_24900);
nand UO_2755 (O_2755,N_24898,N_24784);
xnor UO_2756 (O_2756,N_24564,N_24572);
and UO_2757 (O_2757,N_24585,N_24517);
xor UO_2758 (O_2758,N_24971,N_24645);
or UO_2759 (O_2759,N_24888,N_24684);
xnor UO_2760 (O_2760,N_24692,N_24821);
or UO_2761 (O_2761,N_24965,N_24761);
and UO_2762 (O_2762,N_24518,N_24826);
nor UO_2763 (O_2763,N_24868,N_24730);
xnor UO_2764 (O_2764,N_24690,N_24866);
nand UO_2765 (O_2765,N_24527,N_24580);
nor UO_2766 (O_2766,N_24599,N_24574);
xnor UO_2767 (O_2767,N_24511,N_24889);
xor UO_2768 (O_2768,N_24630,N_24903);
xor UO_2769 (O_2769,N_24953,N_24608);
or UO_2770 (O_2770,N_24993,N_24550);
nor UO_2771 (O_2771,N_24627,N_24613);
nor UO_2772 (O_2772,N_24583,N_24723);
xnor UO_2773 (O_2773,N_24901,N_24907);
or UO_2774 (O_2774,N_24812,N_24625);
or UO_2775 (O_2775,N_24918,N_24644);
or UO_2776 (O_2776,N_24598,N_24973);
nand UO_2777 (O_2777,N_24502,N_24671);
and UO_2778 (O_2778,N_24523,N_24737);
xor UO_2779 (O_2779,N_24802,N_24839);
or UO_2780 (O_2780,N_24708,N_24986);
or UO_2781 (O_2781,N_24605,N_24898);
and UO_2782 (O_2782,N_24521,N_24637);
and UO_2783 (O_2783,N_24879,N_24952);
and UO_2784 (O_2784,N_24744,N_24705);
and UO_2785 (O_2785,N_24961,N_24744);
and UO_2786 (O_2786,N_24705,N_24809);
xnor UO_2787 (O_2787,N_24994,N_24749);
xnor UO_2788 (O_2788,N_24809,N_24605);
and UO_2789 (O_2789,N_24646,N_24912);
nand UO_2790 (O_2790,N_24509,N_24938);
xnor UO_2791 (O_2791,N_24705,N_24868);
nor UO_2792 (O_2792,N_24733,N_24564);
xnor UO_2793 (O_2793,N_24833,N_24933);
nor UO_2794 (O_2794,N_24607,N_24766);
and UO_2795 (O_2795,N_24769,N_24836);
and UO_2796 (O_2796,N_24963,N_24570);
and UO_2797 (O_2797,N_24730,N_24627);
nand UO_2798 (O_2798,N_24849,N_24853);
xnor UO_2799 (O_2799,N_24678,N_24670);
xor UO_2800 (O_2800,N_24762,N_24551);
xnor UO_2801 (O_2801,N_24560,N_24823);
xnor UO_2802 (O_2802,N_24754,N_24808);
and UO_2803 (O_2803,N_24570,N_24893);
and UO_2804 (O_2804,N_24672,N_24999);
or UO_2805 (O_2805,N_24520,N_24601);
and UO_2806 (O_2806,N_24865,N_24925);
or UO_2807 (O_2807,N_24705,N_24876);
xnor UO_2808 (O_2808,N_24957,N_24925);
xor UO_2809 (O_2809,N_24732,N_24734);
xnor UO_2810 (O_2810,N_24720,N_24840);
xor UO_2811 (O_2811,N_24966,N_24962);
or UO_2812 (O_2812,N_24744,N_24922);
nor UO_2813 (O_2813,N_24681,N_24917);
or UO_2814 (O_2814,N_24676,N_24934);
nor UO_2815 (O_2815,N_24554,N_24586);
nand UO_2816 (O_2816,N_24856,N_24508);
or UO_2817 (O_2817,N_24993,N_24738);
and UO_2818 (O_2818,N_24638,N_24543);
and UO_2819 (O_2819,N_24772,N_24770);
nor UO_2820 (O_2820,N_24758,N_24605);
nor UO_2821 (O_2821,N_24990,N_24935);
and UO_2822 (O_2822,N_24902,N_24925);
and UO_2823 (O_2823,N_24879,N_24898);
and UO_2824 (O_2824,N_24568,N_24798);
and UO_2825 (O_2825,N_24995,N_24506);
nand UO_2826 (O_2826,N_24930,N_24540);
xnor UO_2827 (O_2827,N_24692,N_24546);
and UO_2828 (O_2828,N_24943,N_24679);
xnor UO_2829 (O_2829,N_24673,N_24804);
nor UO_2830 (O_2830,N_24605,N_24962);
nand UO_2831 (O_2831,N_24564,N_24529);
nor UO_2832 (O_2832,N_24719,N_24573);
nand UO_2833 (O_2833,N_24566,N_24997);
or UO_2834 (O_2834,N_24647,N_24888);
xor UO_2835 (O_2835,N_24754,N_24841);
and UO_2836 (O_2836,N_24813,N_24633);
and UO_2837 (O_2837,N_24835,N_24957);
nor UO_2838 (O_2838,N_24845,N_24613);
nand UO_2839 (O_2839,N_24717,N_24837);
and UO_2840 (O_2840,N_24963,N_24600);
nand UO_2841 (O_2841,N_24963,N_24859);
xor UO_2842 (O_2842,N_24992,N_24710);
and UO_2843 (O_2843,N_24639,N_24525);
and UO_2844 (O_2844,N_24529,N_24630);
nor UO_2845 (O_2845,N_24619,N_24747);
nor UO_2846 (O_2846,N_24728,N_24864);
xor UO_2847 (O_2847,N_24945,N_24718);
nand UO_2848 (O_2848,N_24733,N_24997);
and UO_2849 (O_2849,N_24542,N_24828);
xnor UO_2850 (O_2850,N_24651,N_24781);
nand UO_2851 (O_2851,N_24579,N_24991);
nor UO_2852 (O_2852,N_24922,N_24718);
or UO_2853 (O_2853,N_24686,N_24856);
and UO_2854 (O_2854,N_24746,N_24783);
xnor UO_2855 (O_2855,N_24610,N_24623);
or UO_2856 (O_2856,N_24815,N_24930);
nand UO_2857 (O_2857,N_24661,N_24622);
nand UO_2858 (O_2858,N_24642,N_24960);
and UO_2859 (O_2859,N_24671,N_24544);
nor UO_2860 (O_2860,N_24680,N_24956);
xnor UO_2861 (O_2861,N_24969,N_24773);
and UO_2862 (O_2862,N_24842,N_24700);
or UO_2863 (O_2863,N_24778,N_24871);
and UO_2864 (O_2864,N_24620,N_24865);
nand UO_2865 (O_2865,N_24871,N_24851);
and UO_2866 (O_2866,N_24935,N_24730);
and UO_2867 (O_2867,N_24653,N_24776);
xor UO_2868 (O_2868,N_24928,N_24875);
or UO_2869 (O_2869,N_24609,N_24950);
or UO_2870 (O_2870,N_24674,N_24828);
xnor UO_2871 (O_2871,N_24747,N_24726);
or UO_2872 (O_2872,N_24841,N_24656);
and UO_2873 (O_2873,N_24842,N_24552);
xnor UO_2874 (O_2874,N_24941,N_24749);
xnor UO_2875 (O_2875,N_24513,N_24691);
xor UO_2876 (O_2876,N_24905,N_24994);
nand UO_2877 (O_2877,N_24706,N_24804);
xor UO_2878 (O_2878,N_24803,N_24742);
xor UO_2879 (O_2879,N_24635,N_24553);
nor UO_2880 (O_2880,N_24698,N_24953);
nand UO_2881 (O_2881,N_24642,N_24571);
nand UO_2882 (O_2882,N_24592,N_24694);
xor UO_2883 (O_2883,N_24646,N_24988);
nand UO_2884 (O_2884,N_24981,N_24588);
nand UO_2885 (O_2885,N_24980,N_24981);
and UO_2886 (O_2886,N_24700,N_24691);
and UO_2887 (O_2887,N_24960,N_24831);
xor UO_2888 (O_2888,N_24828,N_24985);
and UO_2889 (O_2889,N_24802,N_24912);
or UO_2890 (O_2890,N_24965,N_24738);
xor UO_2891 (O_2891,N_24588,N_24865);
nand UO_2892 (O_2892,N_24802,N_24862);
or UO_2893 (O_2893,N_24924,N_24548);
and UO_2894 (O_2894,N_24935,N_24503);
nor UO_2895 (O_2895,N_24528,N_24988);
nand UO_2896 (O_2896,N_24990,N_24583);
nand UO_2897 (O_2897,N_24698,N_24787);
and UO_2898 (O_2898,N_24868,N_24886);
nor UO_2899 (O_2899,N_24576,N_24924);
and UO_2900 (O_2900,N_24533,N_24798);
nor UO_2901 (O_2901,N_24679,N_24747);
or UO_2902 (O_2902,N_24793,N_24839);
nor UO_2903 (O_2903,N_24873,N_24619);
xnor UO_2904 (O_2904,N_24958,N_24927);
or UO_2905 (O_2905,N_24802,N_24885);
xnor UO_2906 (O_2906,N_24711,N_24968);
nor UO_2907 (O_2907,N_24881,N_24857);
or UO_2908 (O_2908,N_24837,N_24709);
nand UO_2909 (O_2909,N_24970,N_24601);
nand UO_2910 (O_2910,N_24604,N_24503);
nor UO_2911 (O_2911,N_24712,N_24999);
xor UO_2912 (O_2912,N_24970,N_24627);
nor UO_2913 (O_2913,N_24656,N_24920);
and UO_2914 (O_2914,N_24983,N_24767);
nand UO_2915 (O_2915,N_24693,N_24807);
xor UO_2916 (O_2916,N_24916,N_24862);
xor UO_2917 (O_2917,N_24959,N_24925);
or UO_2918 (O_2918,N_24568,N_24545);
nand UO_2919 (O_2919,N_24909,N_24849);
nor UO_2920 (O_2920,N_24543,N_24739);
or UO_2921 (O_2921,N_24966,N_24739);
xor UO_2922 (O_2922,N_24797,N_24860);
nand UO_2923 (O_2923,N_24544,N_24936);
or UO_2924 (O_2924,N_24688,N_24526);
and UO_2925 (O_2925,N_24916,N_24575);
xnor UO_2926 (O_2926,N_24570,N_24517);
nand UO_2927 (O_2927,N_24751,N_24791);
xnor UO_2928 (O_2928,N_24926,N_24648);
nand UO_2929 (O_2929,N_24908,N_24877);
or UO_2930 (O_2930,N_24697,N_24808);
xnor UO_2931 (O_2931,N_24964,N_24578);
xnor UO_2932 (O_2932,N_24932,N_24585);
nand UO_2933 (O_2933,N_24877,N_24819);
nand UO_2934 (O_2934,N_24504,N_24793);
nand UO_2935 (O_2935,N_24514,N_24720);
nand UO_2936 (O_2936,N_24540,N_24908);
nor UO_2937 (O_2937,N_24616,N_24573);
xnor UO_2938 (O_2938,N_24981,N_24878);
xor UO_2939 (O_2939,N_24960,N_24534);
and UO_2940 (O_2940,N_24916,N_24931);
xnor UO_2941 (O_2941,N_24938,N_24842);
xor UO_2942 (O_2942,N_24573,N_24733);
or UO_2943 (O_2943,N_24796,N_24983);
nor UO_2944 (O_2944,N_24887,N_24773);
or UO_2945 (O_2945,N_24731,N_24546);
or UO_2946 (O_2946,N_24614,N_24552);
xor UO_2947 (O_2947,N_24746,N_24675);
xor UO_2948 (O_2948,N_24534,N_24944);
and UO_2949 (O_2949,N_24923,N_24780);
and UO_2950 (O_2950,N_24857,N_24562);
nor UO_2951 (O_2951,N_24801,N_24863);
and UO_2952 (O_2952,N_24575,N_24884);
nor UO_2953 (O_2953,N_24831,N_24636);
nor UO_2954 (O_2954,N_24509,N_24569);
xnor UO_2955 (O_2955,N_24525,N_24811);
or UO_2956 (O_2956,N_24831,N_24508);
nor UO_2957 (O_2957,N_24604,N_24978);
nor UO_2958 (O_2958,N_24887,N_24876);
and UO_2959 (O_2959,N_24770,N_24795);
and UO_2960 (O_2960,N_24681,N_24903);
and UO_2961 (O_2961,N_24840,N_24813);
and UO_2962 (O_2962,N_24956,N_24921);
or UO_2963 (O_2963,N_24545,N_24851);
nand UO_2964 (O_2964,N_24762,N_24722);
nand UO_2965 (O_2965,N_24577,N_24559);
xor UO_2966 (O_2966,N_24665,N_24706);
nor UO_2967 (O_2967,N_24733,N_24933);
and UO_2968 (O_2968,N_24909,N_24765);
nand UO_2969 (O_2969,N_24556,N_24654);
or UO_2970 (O_2970,N_24897,N_24749);
or UO_2971 (O_2971,N_24817,N_24530);
nor UO_2972 (O_2972,N_24640,N_24967);
nand UO_2973 (O_2973,N_24661,N_24995);
and UO_2974 (O_2974,N_24904,N_24541);
nand UO_2975 (O_2975,N_24821,N_24893);
nand UO_2976 (O_2976,N_24748,N_24571);
xor UO_2977 (O_2977,N_24589,N_24564);
nand UO_2978 (O_2978,N_24500,N_24526);
nor UO_2979 (O_2979,N_24725,N_24917);
or UO_2980 (O_2980,N_24789,N_24814);
nand UO_2981 (O_2981,N_24660,N_24944);
nand UO_2982 (O_2982,N_24723,N_24681);
nor UO_2983 (O_2983,N_24941,N_24722);
nor UO_2984 (O_2984,N_24550,N_24802);
or UO_2985 (O_2985,N_24521,N_24685);
nor UO_2986 (O_2986,N_24694,N_24904);
nor UO_2987 (O_2987,N_24816,N_24957);
nand UO_2988 (O_2988,N_24952,N_24680);
nand UO_2989 (O_2989,N_24752,N_24656);
and UO_2990 (O_2990,N_24611,N_24686);
nor UO_2991 (O_2991,N_24524,N_24921);
and UO_2992 (O_2992,N_24635,N_24915);
or UO_2993 (O_2993,N_24669,N_24624);
xnor UO_2994 (O_2994,N_24539,N_24982);
and UO_2995 (O_2995,N_24722,N_24534);
nor UO_2996 (O_2996,N_24907,N_24855);
nand UO_2997 (O_2997,N_24932,N_24830);
xor UO_2998 (O_2998,N_24544,N_24837);
nand UO_2999 (O_2999,N_24527,N_24531);
endmodule