module basic_1500_15000_2000_15_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_807,In_1374);
or U1 (N_1,In_969,In_1400);
nand U2 (N_2,In_1023,In_246);
and U3 (N_3,In_1437,In_940);
nor U4 (N_4,In_487,In_881);
nand U5 (N_5,In_1480,In_1092);
nor U6 (N_6,In_1000,In_224);
nand U7 (N_7,In_1043,In_1141);
and U8 (N_8,In_417,In_308);
nor U9 (N_9,In_361,In_680);
and U10 (N_10,In_471,In_1354);
nand U11 (N_11,In_1415,In_952);
nor U12 (N_12,In_1129,In_1010);
nand U13 (N_13,In_1309,In_998);
nor U14 (N_14,In_551,In_967);
and U15 (N_15,In_1060,In_359);
nor U16 (N_16,In_547,In_597);
or U17 (N_17,In_94,In_221);
nor U18 (N_18,In_839,In_1422);
and U19 (N_19,In_1169,In_38);
xnor U20 (N_20,In_1139,In_61);
nand U21 (N_21,In_12,In_847);
nor U22 (N_22,In_32,In_600);
and U23 (N_23,In_1020,In_173);
and U24 (N_24,In_926,In_357);
and U25 (N_25,In_1119,In_1191);
nand U26 (N_26,In_791,In_13);
and U27 (N_27,In_852,In_6);
nor U28 (N_28,In_884,In_1409);
nor U29 (N_29,In_1499,In_548);
nor U30 (N_30,In_57,In_976);
nand U31 (N_31,In_1061,In_701);
nand U32 (N_32,In_718,In_725);
nor U33 (N_33,In_953,In_669);
nand U34 (N_34,In_981,In_327);
and U35 (N_35,In_764,In_894);
and U36 (N_36,In_1182,In_438);
or U37 (N_37,In_1161,In_1219);
nand U38 (N_38,In_75,In_305);
nand U39 (N_39,In_444,In_1026);
nor U40 (N_40,In_157,In_1240);
or U41 (N_41,In_275,In_1270);
or U42 (N_42,In_538,In_1394);
xnor U43 (N_43,In_1097,In_290);
xnor U44 (N_44,In_933,In_523);
or U45 (N_45,In_777,In_694);
nand U46 (N_46,In_567,In_161);
xnor U47 (N_47,In_106,In_436);
nand U48 (N_48,In_549,In_326);
or U49 (N_49,In_95,In_1176);
xor U50 (N_50,In_1086,In_1089);
nand U51 (N_51,In_963,In_1143);
nor U52 (N_52,In_1302,In_318);
nor U53 (N_53,In_2,In_146);
or U54 (N_54,In_1223,In_292);
and U55 (N_55,In_24,In_100);
nand U56 (N_56,In_1458,In_469);
and U57 (N_57,In_617,In_1450);
nand U58 (N_58,In_29,In_664);
and U59 (N_59,In_416,In_844);
or U60 (N_60,In_973,In_813);
nor U61 (N_61,In_1245,In_826);
and U62 (N_62,In_151,In_561);
or U63 (N_63,In_961,In_463);
and U64 (N_64,In_528,In_1416);
nor U65 (N_65,In_1208,In_584);
and U66 (N_66,In_451,In_332);
and U67 (N_67,In_810,In_1375);
nor U68 (N_68,In_811,In_165);
or U69 (N_69,In_572,In_1293);
and U70 (N_70,In_1483,In_608);
nor U71 (N_71,In_465,In_77);
and U72 (N_72,In_866,In_905);
and U73 (N_73,In_995,In_480);
nor U74 (N_74,In_162,In_1457);
or U75 (N_75,In_709,In_365);
or U76 (N_76,In_501,In_535);
and U77 (N_77,In_988,In_544);
nor U78 (N_78,In_1075,In_1484);
nand U79 (N_79,In_534,In_1482);
and U80 (N_80,In_1443,In_223);
xor U81 (N_81,In_303,In_354);
nand U82 (N_82,In_1327,In_1113);
and U83 (N_83,In_748,In_687);
and U84 (N_84,In_634,In_319);
and U85 (N_85,In_1142,In_248);
or U86 (N_86,In_496,In_758);
or U87 (N_87,In_155,In_181);
or U88 (N_88,In_1105,In_1073);
nor U89 (N_89,In_986,In_1071);
nand U90 (N_90,In_271,In_796);
and U91 (N_91,In_1085,In_73);
nand U92 (N_92,In_682,In_1306);
nand U93 (N_93,In_663,In_234);
xnor U94 (N_94,In_595,In_1417);
or U95 (N_95,In_1404,In_203);
and U96 (N_96,In_1288,In_1384);
or U97 (N_97,In_1467,In_1299);
or U98 (N_98,In_1432,In_490);
nand U99 (N_99,In_21,In_139);
or U100 (N_100,In_1214,In_814);
and U101 (N_101,In_662,In_1326);
nor U102 (N_102,In_524,In_999);
xnor U103 (N_103,In_312,In_222);
and U104 (N_104,In_765,In_779);
or U105 (N_105,In_838,In_968);
and U106 (N_106,In_1407,In_1249);
nand U107 (N_107,In_1455,In_606);
nor U108 (N_108,In_1285,In_179);
and U109 (N_109,In_674,In_775);
nand U110 (N_110,In_1423,In_792);
nand U111 (N_111,In_1030,In_1213);
xnor U112 (N_112,In_1007,In_1068);
and U113 (N_113,In_1134,In_786);
and U114 (N_114,In_486,In_1031);
nand U115 (N_115,In_209,In_768);
xor U116 (N_116,In_1470,In_1449);
nand U117 (N_117,In_728,In_336);
and U118 (N_118,In_520,In_377);
nand U119 (N_119,In_562,In_956);
nand U120 (N_120,In_717,In_1307);
or U121 (N_121,In_1392,In_304);
nand U122 (N_122,In_289,In_641);
and U123 (N_123,In_526,In_205);
xnor U124 (N_124,In_315,In_1198);
nand U125 (N_125,In_175,In_875);
nand U126 (N_126,In_590,In_1255);
nor U127 (N_127,In_262,In_1202);
nand U128 (N_128,In_59,In_1475);
nand U129 (N_129,In_873,In_1229);
nand U130 (N_130,In_172,In_242);
nor U131 (N_131,In_936,In_787);
or U132 (N_132,In_375,In_1103);
or U133 (N_133,In_610,In_340);
xnor U134 (N_134,In_228,In_631);
nand U135 (N_135,In_1230,In_372);
and U136 (N_136,In_1149,In_227);
or U137 (N_137,In_543,In_1199);
or U138 (N_138,In_1122,In_458);
nand U139 (N_139,In_169,In_346);
or U140 (N_140,In_1002,In_1076);
or U141 (N_141,In_1385,In_233);
nand U142 (N_142,In_1107,In_341);
and U143 (N_143,In_1368,In_1174);
and U144 (N_144,In_843,In_1402);
nor U145 (N_145,In_592,In_1059);
and U146 (N_146,In_892,In_1295);
nor U147 (N_147,In_239,In_96);
nor U148 (N_148,In_269,In_612);
nand U149 (N_149,In_696,In_620);
or U150 (N_150,In_1039,In_1300);
or U151 (N_151,In_994,In_1273);
and U152 (N_152,In_86,In_984);
nand U153 (N_153,In_34,In_427);
or U154 (N_154,In_187,In_293);
nand U155 (N_155,In_1410,In_1494);
or U156 (N_156,In_1284,In_1337);
nand U157 (N_157,In_726,In_916);
and U158 (N_158,In_756,In_1244);
or U159 (N_159,In_752,In_1253);
or U160 (N_160,In_982,In_83);
and U161 (N_161,In_1361,In_236);
nand U162 (N_162,In_499,In_1172);
nor U163 (N_163,In_938,In_174);
nor U164 (N_164,In_84,In_960);
nand U165 (N_165,In_314,In_951);
or U166 (N_166,In_371,In_502);
and U167 (N_167,In_589,In_1379);
nor U168 (N_168,In_655,In_350);
xor U169 (N_169,In_1011,In_795);
or U170 (N_170,In_863,In_1234);
nor U171 (N_171,In_1135,In_1232);
nand U172 (N_172,In_1491,In_216);
xnor U173 (N_173,In_835,In_26);
and U174 (N_174,In_644,In_676);
or U175 (N_175,In_909,In_1261);
nand U176 (N_176,In_586,In_492);
nand U177 (N_177,In_754,In_887);
or U178 (N_178,In_1221,In_351);
nand U179 (N_179,In_734,In_1012);
nand U180 (N_180,In_434,In_468);
or U181 (N_181,In_51,In_947);
nand U182 (N_182,In_335,In_1117);
or U183 (N_183,In_781,In_1388);
nand U184 (N_184,In_1123,In_53);
and U185 (N_185,In_398,In_237);
or U186 (N_186,In_99,In_230);
nand U187 (N_187,In_1325,In_334);
or U188 (N_188,In_623,In_603);
nand U189 (N_189,In_1497,In_553);
or U190 (N_190,In_702,In_1358);
xnor U191 (N_191,In_429,In_1469);
and U192 (N_192,In_516,In_352);
nor U193 (N_193,In_895,In_798);
and U194 (N_194,In_1398,In_1035);
or U195 (N_195,In_1005,In_900);
and U196 (N_196,In_1314,In_642);
and U197 (N_197,In_363,In_251);
xor U198 (N_198,In_911,In_706);
or U199 (N_199,In_670,In_632);
or U200 (N_200,In_1492,In_879);
and U201 (N_201,In_921,In_395);
and U202 (N_202,In_1356,In_1266);
and U203 (N_203,In_651,In_1339);
nor U204 (N_204,In_1095,In_131);
and U205 (N_205,In_198,In_972);
or U206 (N_206,In_250,In_74);
nor U207 (N_207,In_773,In_1046);
or U208 (N_208,In_240,In_679);
nand U209 (N_209,In_15,In_48);
or U210 (N_210,In_393,In_367);
or U211 (N_211,In_903,In_1347);
xnor U212 (N_212,In_724,In_806);
nand U213 (N_213,In_1247,In_1308);
xnor U214 (N_214,In_115,In_527);
nand U215 (N_215,In_1056,In_3);
and U216 (N_216,In_1003,In_270);
nor U217 (N_217,In_145,In_122);
nor U218 (N_218,In_1233,In_959);
and U219 (N_219,In_1393,In_1496);
xnor U220 (N_220,In_691,In_435);
nand U221 (N_221,In_1070,In_1424);
nor U222 (N_222,In_397,In_882);
nor U223 (N_223,In_78,In_915);
nor U224 (N_224,In_253,In_871);
and U225 (N_225,In_1114,In_753);
nor U226 (N_226,In_282,In_1252);
xnor U227 (N_227,In_168,In_1246);
nand U228 (N_228,In_355,In_574);
nor U229 (N_229,In_188,In_569);
or U230 (N_230,In_957,In_116);
xnor U231 (N_231,In_575,In_420);
and U232 (N_232,In_576,In_192);
xnor U233 (N_233,In_573,In_98);
or U234 (N_234,In_1460,In_1188);
and U235 (N_235,In_439,In_320);
and U236 (N_236,In_539,In_1439);
xor U237 (N_237,In_625,In_422);
nand U238 (N_238,In_736,In_594);
or U239 (N_239,In_788,In_404);
nand U240 (N_240,In_1321,In_751);
or U241 (N_241,In_828,In_1153);
or U242 (N_242,In_1436,In_133);
or U243 (N_243,In_159,In_735);
and U244 (N_244,In_285,In_178);
nand U245 (N_245,In_189,In_307);
and U246 (N_246,In_783,In_280);
nand U247 (N_247,In_441,In_703);
and U248 (N_248,In_517,In_598);
nor U249 (N_249,In_729,In_1196);
or U250 (N_250,In_910,In_426);
and U251 (N_251,In_1420,In_217);
xor U252 (N_252,In_1224,In_732);
and U253 (N_253,In_1048,In_914);
nand U254 (N_254,In_191,In_1231);
nor U255 (N_255,In_506,In_1133);
or U256 (N_256,In_123,In_347);
or U257 (N_257,In_409,In_297);
or U258 (N_258,In_1167,In_1360);
nor U259 (N_259,In_407,In_424);
or U260 (N_260,In_1180,In_503);
nand U261 (N_261,In_313,In_1069);
nor U262 (N_262,In_1151,In_804);
and U263 (N_263,In_349,In_697);
and U264 (N_264,In_68,In_1256);
or U265 (N_265,In_287,In_533);
nand U266 (N_266,In_370,In_128);
and U267 (N_267,In_849,In_103);
and U268 (N_268,In_495,In_1330);
nor U269 (N_269,In_1237,In_1222);
and U270 (N_270,In_445,In_288);
xor U271 (N_271,In_1215,In_1225);
nor U272 (N_272,In_1088,In_117);
nand U273 (N_273,In_842,In_1485);
nor U274 (N_274,In_30,In_816);
and U275 (N_275,In_944,In_1185);
xor U276 (N_276,In_60,In_430);
nor U277 (N_277,In_942,In_985);
xor U278 (N_278,In_1454,In_328);
or U279 (N_279,In_1238,In_1344);
or U280 (N_280,In_746,In_1236);
and U281 (N_281,In_1,In_802);
nor U282 (N_282,In_996,In_265);
xor U283 (N_283,In_1064,In_1444);
or U284 (N_284,In_599,In_1459);
nand U285 (N_285,In_653,In_244);
nor U286 (N_286,In_72,In_1132);
nand U287 (N_287,In_109,In_1399);
or U288 (N_288,In_376,In_552);
and U289 (N_289,In_79,In_1322);
xor U290 (N_290,In_353,In_379);
nand U291 (N_291,In_411,In_955);
nor U292 (N_292,In_1148,In_1016);
and U293 (N_293,In_1463,In_1258);
and U294 (N_294,In_107,In_245);
nor U295 (N_295,In_659,In_1465);
and U296 (N_296,In_325,In_711);
and U297 (N_297,In_1051,In_1468);
nand U298 (N_298,In_97,In_1029);
nand U299 (N_299,In_971,In_554);
and U300 (N_300,In_31,In_950);
xor U301 (N_301,In_120,In_477);
or U302 (N_302,In_587,In_629);
or U303 (N_303,In_789,In_323);
and U304 (N_304,In_470,In_943);
or U305 (N_305,In_284,In_154);
xnor U306 (N_306,In_830,In_46);
and U307 (N_307,In_1489,In_514);
nand U308 (N_308,In_200,In_782);
and U309 (N_309,In_418,In_33);
xnor U310 (N_310,In_90,In_5);
xnor U311 (N_311,In_212,In_428);
nand U312 (N_312,In_505,In_722);
nand U313 (N_313,In_827,In_152);
xnor U314 (N_314,In_977,In_475);
or U315 (N_315,In_868,In_615);
or U316 (N_316,In_1034,In_1033);
or U317 (N_317,In_1419,In_1216);
xnor U318 (N_318,In_119,In_721);
or U319 (N_319,In_808,In_1476);
nand U320 (N_320,In_738,In_1189);
nand U321 (N_321,In_47,In_111);
or U322 (N_322,In_1163,In_1257);
and U323 (N_323,In_1057,In_196);
and U324 (N_324,In_1197,In_688);
and U325 (N_325,In_531,In_767);
or U326 (N_326,In_616,In_472);
or U327 (N_327,In_1078,In_461);
nor U328 (N_328,In_309,In_563);
nand U329 (N_329,In_1279,In_613);
nor U330 (N_330,In_949,In_193);
nor U331 (N_331,In_784,In_1274);
or U332 (N_332,In_1292,In_383);
xor U333 (N_333,In_507,In_19);
xor U334 (N_334,In_932,In_519);
nand U335 (N_335,In_364,In_1106);
or U336 (N_336,In_1091,In_333);
and U337 (N_337,In_633,In_394);
or U338 (N_338,In_1352,In_1022);
nand U339 (N_339,In_730,In_919);
nor U340 (N_340,In_4,In_941);
and U341 (N_341,In_1116,In_1334);
xor U342 (N_342,In_668,In_382);
and U343 (N_343,In_772,In_449);
or U344 (N_344,In_356,In_760);
or U345 (N_345,In_67,In_1186);
or U346 (N_346,In_425,In_602);
and U347 (N_347,In_1235,In_521);
or U348 (N_348,In_42,In_1187);
nand U349 (N_349,In_997,In_1280);
nand U350 (N_350,In_298,In_1156);
xor U351 (N_351,In_1286,In_1104);
or U352 (N_352,In_1190,In_980);
nor U353 (N_353,In_665,In_140);
or U354 (N_354,In_1380,In_1019);
and U355 (N_355,In_1008,In_965);
nand U356 (N_356,In_1389,In_105);
xnor U357 (N_357,In_17,In_821);
and U358 (N_358,In_1150,In_1137);
or U359 (N_359,In_818,In_466);
nor U360 (N_360,In_1067,In_1453);
xnor U361 (N_361,In_1390,In_494);
nor U362 (N_362,In_443,In_624);
xor U363 (N_363,In_433,In_301);
nand U364 (N_364,In_295,In_928);
or U365 (N_365,In_1277,In_1146);
nand U366 (N_366,In_1272,In_693);
or U367 (N_367,In_785,In_1166);
or U368 (N_368,In_1498,In_137);
nand U369 (N_369,In_185,In_81);
or U370 (N_370,In_1428,In_1265);
or U371 (N_371,In_1298,In_1006);
and U372 (N_372,In_759,In_306);
and U373 (N_373,In_1473,In_1363);
nor U374 (N_374,In_860,In_18);
and U375 (N_375,In_1296,In_1477);
and U376 (N_376,In_92,In_102);
and U377 (N_377,In_1332,In_630);
nand U378 (N_378,In_565,In_368);
and U379 (N_379,In_453,In_831);
xnor U380 (N_380,In_862,In_1228);
and U381 (N_381,In_1461,In_927);
or U382 (N_382,In_931,In_247);
nand U383 (N_383,In_1184,In_1278);
nand U384 (N_384,In_226,In_646);
and U385 (N_385,In_337,In_626);
or U386 (N_386,In_690,In_747);
and U387 (N_387,In_1206,In_708);
or U388 (N_388,In_546,In_899);
nor U389 (N_389,In_1269,In_43);
and U390 (N_390,In_640,In_266);
nand U391 (N_391,In_614,In_672);
nand U392 (N_392,In_761,In_657);
and U393 (N_393,In_403,In_945);
xor U394 (N_394,In_618,In_848);
nor U395 (N_395,In_778,In_1304);
nand U396 (N_396,In_699,In_448);
nand U397 (N_397,In_126,In_1421);
nor U398 (N_398,In_948,In_129);
nand U399 (N_399,In_621,In_1411);
or U400 (N_400,In_497,In_583);
or U401 (N_401,In_199,In_322);
nor U402 (N_402,In_525,In_124);
nand U403 (N_403,In_385,In_1038);
or U404 (N_404,In_885,In_254);
or U405 (N_405,In_1001,In_800);
nor U406 (N_406,In_1096,In_857);
nand U407 (N_407,In_190,In_1047);
and U408 (N_408,In_374,In_628);
nor U409 (N_409,In_321,In_231);
nand U410 (N_410,In_66,In_1041);
or U411 (N_411,In_581,In_1124);
nand U412 (N_412,In_388,In_437);
or U413 (N_413,In_698,In_1353);
nor U414 (N_414,In_125,In_147);
and U415 (N_415,In_80,In_1145);
xor U416 (N_416,In_1397,In_1065);
xor U417 (N_417,In_978,In_1178);
nand U418 (N_418,In_316,In_541);
nand U419 (N_419,In_170,In_537);
nor U420 (N_420,In_714,In_744);
nor U421 (N_421,In_7,In_158);
nor U422 (N_422,In_845,In_854);
nand U423 (N_423,In_870,In_118);
and U424 (N_424,In_560,In_1173);
nor U425 (N_425,In_888,In_1200);
or U426 (N_426,In_134,In_1426);
nor U427 (N_427,In_1204,In_743);
or U428 (N_428,In_1217,In_1479);
nor U429 (N_429,In_637,In_63);
xnor U430 (N_430,In_1209,In_329);
or U431 (N_431,In_638,In_255);
xor U432 (N_432,In_1045,In_1319);
and U433 (N_433,In_467,In_966);
nand U434 (N_434,In_1136,In_1282);
nand U435 (N_435,In_647,In_858);
and U436 (N_436,In_1168,In_815);
or U437 (N_437,In_585,In_1170);
and U438 (N_438,In_1155,In_832);
xnor U439 (N_439,In_85,In_1021);
xnor U440 (N_440,In_294,In_10);
and U441 (N_441,In_1183,In_1372);
nor U442 (N_442,In_16,In_1101);
nor U443 (N_443,In_975,In_588);
and U444 (N_444,In_686,In_1218);
and U445 (N_445,In_419,In_908);
and U446 (N_446,In_0,In_917);
nand U447 (N_447,In_260,In_654);
nand U448 (N_448,In_311,In_1287);
nand U449 (N_449,In_201,In_1418);
or U450 (N_450,In_979,In_799);
or U451 (N_451,In_1084,In_1162);
nor U452 (N_452,In_542,In_1291);
or U453 (N_453,In_923,In_283);
nor U454 (N_454,In_897,In_1464);
nand U455 (N_455,In_296,In_493);
nor U456 (N_456,In_142,In_489);
or U457 (N_457,In_431,In_762);
and U458 (N_458,In_1248,In_177);
or U459 (N_459,In_731,In_872);
and U460 (N_460,In_512,In_144);
nor U461 (N_461,In_1239,In_906);
nor U462 (N_462,In_1451,In_925);
nor U463 (N_463,In_167,In_1366);
xnor U464 (N_464,In_661,In_1171);
or U465 (N_465,In_1301,In_1147);
xor U466 (N_466,In_564,In_101);
nand U467 (N_467,In_384,In_1452);
nor U468 (N_468,In_1433,In_396);
nor U469 (N_469,In_391,In_360);
and U470 (N_470,In_210,In_1125);
or U471 (N_471,In_330,In_1427);
xor U472 (N_472,In_958,In_1448);
xnor U473 (N_473,In_874,In_1130);
nor U474 (N_474,In_593,In_1495);
nor U475 (N_475,In_912,In_1446);
or U476 (N_476,In_893,In_1466);
and U477 (N_477,In_1343,In_902);
and U478 (N_478,In_1112,In_281);
nand U479 (N_479,In_267,In_1318);
nor U480 (N_480,In_1276,In_695);
and U481 (N_481,In_510,In_1430);
or U482 (N_482,In_770,In_1362);
nand U483 (N_483,In_700,In_1425);
nand U484 (N_484,In_206,In_607);
and U485 (N_485,In_163,In_596);
or U486 (N_486,In_91,In_257);
nor U487 (N_487,In_1227,In_650);
xor U488 (N_488,In_184,In_498);
xnor U489 (N_489,In_402,In_28);
xnor U490 (N_490,In_851,In_1317);
nor U491 (N_491,In_559,In_1431);
nand U492 (N_492,In_890,In_415);
and U493 (N_493,In_50,In_1111);
xnor U494 (N_494,In_1378,In_675);
or U495 (N_495,In_276,In_183);
and U496 (N_496,In_836,In_666);
nor U497 (N_497,In_913,In_529);
or U498 (N_498,In_1462,In_1471);
nand U499 (N_499,In_56,In_1315);
nor U500 (N_500,In_252,In_1371);
or U501 (N_501,In_1401,In_1128);
or U502 (N_502,In_62,In_723);
and U503 (N_503,In_716,In_1364);
or U504 (N_504,In_934,In_1211);
or U505 (N_505,In_324,In_518);
nand U506 (N_506,In_1267,In_1127);
nand U507 (N_507,In_1036,In_1062);
xor U508 (N_508,In_898,In_1412);
and U509 (N_509,In_571,In_1164);
nand U510 (N_510,In_278,In_677);
xnor U511 (N_511,In_1447,In_954);
and U512 (N_512,In_114,In_11);
and U513 (N_513,In_462,In_386);
nand U514 (N_514,In_719,In_1336);
or U515 (N_515,In_479,In_331);
or U516 (N_516,In_504,In_1083);
nand U517 (N_517,In_373,In_645);
or U518 (N_518,In_755,In_1100);
or U519 (N_519,In_478,In_622);
and U520 (N_520,In_577,In_924);
nand U521 (N_521,In_1396,In_482);
xor U522 (N_522,In_1338,In_1342);
and U523 (N_523,In_801,In_1383);
or U524 (N_524,In_1203,In_1121);
xnor U525 (N_525,In_202,In_148);
or U526 (N_526,In_1009,In_14);
or U527 (N_527,In_1259,In_962);
or U528 (N_528,In_40,In_1120);
xor U529 (N_529,In_604,In_635);
nor U530 (N_530,In_1207,In_1079);
xor U531 (N_531,In_121,In_1251);
nor U532 (N_532,In_970,In_69);
nor U533 (N_533,In_1310,In_286);
or U534 (N_534,In_648,In_1320);
nand U535 (N_535,In_1094,In_745);
xor U536 (N_536,In_180,In_45);
nand U537 (N_537,In_766,In_1212);
or U538 (N_538,In_89,In_591);
xnor U539 (N_539,In_508,In_1037);
xor U540 (N_540,In_156,In_1263);
nand U541 (N_541,In_1359,In_1478);
or U542 (N_542,In_809,In_1138);
and U543 (N_543,In_713,In_1395);
nor U544 (N_544,In_989,In_1063);
nor U545 (N_545,In_93,In_749);
or U546 (N_546,In_387,In_901);
and U547 (N_547,In_1115,In_1264);
or U548 (N_548,In_652,In_937);
nor U549 (N_549,In_1442,In_1289);
or U550 (N_550,In_1015,In_1024);
and U551 (N_551,In_1386,In_678);
or U552 (N_552,In_392,In_1414);
or U553 (N_553,In_344,In_611);
or U554 (N_554,In_545,In_39);
nor U555 (N_555,In_249,In_1241);
or U556 (N_556,In_757,In_649);
nor U557 (N_557,In_1365,In_164);
or U558 (N_558,In_1486,In_859);
nor U559 (N_559,In_195,In_609);
xnor U560 (N_560,In_401,In_1316);
nand U561 (N_561,In_1014,In_259);
nand U562 (N_562,In_141,In_110);
xnor U563 (N_563,In_473,In_20);
or U564 (N_564,In_1165,In_579);
xor U565 (N_565,In_1297,In_491);
xnor U566 (N_566,In_457,In_215);
nor U567 (N_567,In_219,In_214);
and U568 (N_568,In_446,In_841);
or U569 (N_569,In_840,In_408);
nor U570 (N_570,In_601,In_1367);
and U571 (N_571,In_299,In_88);
nand U572 (N_572,In_166,In_1355);
nand U573 (N_573,In_474,In_343);
and U574 (N_574,In_1262,In_317);
nor U575 (N_575,In_1025,In_389);
and U576 (N_576,In_1077,In_797);
or U577 (N_577,In_1093,In_930);
xnor U578 (N_578,In_780,In_338);
or U579 (N_579,In_1098,In_636);
nand U580 (N_580,In_1054,In_1004);
xnor U581 (N_581,In_1440,In_1429);
nand U582 (N_582,In_1403,In_1382);
and U583 (N_583,In_658,In_856);
nand U584 (N_584,In_27,In_264);
nand U585 (N_585,In_272,In_149);
or U586 (N_586,In_741,In_513);
or U587 (N_587,In_987,In_310);
nand U588 (N_588,In_1271,In_1487);
and U589 (N_589,In_812,In_65);
xor U590 (N_590,In_823,In_660);
xnor U591 (N_591,In_1072,In_208);
nand U592 (N_592,In_771,In_1108);
and U593 (N_593,In_667,In_71);
nand U594 (N_594,In_423,In_1329);
nand U595 (N_595,In_256,In_869);
nand U596 (N_596,In_639,In_64);
nor U597 (N_597,In_990,In_550);
nor U598 (N_598,In_220,In_861);
and U599 (N_599,In_263,In_1053);
and U600 (N_600,In_794,In_380);
nand U601 (N_601,In_1243,In_1376);
and U602 (N_602,In_1481,In_1159);
or U603 (N_603,In_44,In_727);
nor U604 (N_604,In_720,In_1377);
or U605 (N_605,In_578,In_399);
nand U606 (N_606,In_22,In_1042);
nand U607 (N_607,In_566,In_1242);
nor U608 (N_608,In_362,In_1028);
nor U609 (N_609,In_825,In_452);
nand U610 (N_610,In_243,In_488);
and U611 (N_611,In_820,In_1405);
nand U612 (N_612,In_182,In_378);
and U613 (N_613,In_127,In_1160);
nor U614 (N_614,In_833,In_710);
nor U615 (N_615,In_557,In_25);
nor U616 (N_616,In_1305,In_582);
nand U617 (N_617,In_1177,In_1192);
xnor U618 (N_618,In_817,In_345);
nand U619 (N_619,In_805,In_238);
xnor U620 (N_620,In_803,In_1250);
and U621 (N_621,In_211,In_113);
and U622 (N_622,In_1032,In_138);
or U623 (N_623,In_414,In_1406);
nand U624 (N_624,In_712,In_1040);
or U625 (N_625,In_150,In_865);
or U626 (N_626,In_9,In_160);
nand U627 (N_627,In_1472,In_733);
or U628 (N_628,In_1152,In_1348);
nand U629 (N_629,In_459,In_907);
nor U630 (N_630,In_186,In_400);
and U631 (N_631,In_213,In_405);
xnor U632 (N_632,In_1074,In_500);
or U633 (N_633,In_929,In_1313);
or U634 (N_634,In_450,In_300);
and U635 (N_635,In_1373,In_671);
nand U636 (N_636,In_1201,In_580);
nor U637 (N_637,In_837,In_1220);
and U638 (N_638,In_1294,In_1154);
and U639 (N_639,In_1018,In_277);
and U640 (N_640,In_704,In_763);
nor U641 (N_641,In_54,In_878);
xor U642 (N_642,In_130,In_568);
and U643 (N_643,In_522,In_58);
nor U644 (N_644,In_939,In_76);
and U645 (N_645,In_454,In_1281);
nor U646 (N_646,In_1087,In_685);
xnor U647 (N_647,In_1179,In_108);
or U648 (N_648,In_790,In_1175);
nor U649 (N_649,In_348,In_35);
nor U650 (N_650,In_824,In_1140);
or U651 (N_651,In_464,In_37);
nand U652 (N_652,In_1345,In_1050);
or U653 (N_653,In_8,In_421);
or U654 (N_654,In_536,In_737);
nand U655 (N_655,In_1194,In_1080);
nand U656 (N_656,In_681,In_1058);
or U657 (N_657,In_1210,In_456);
nand U658 (N_658,In_515,In_769);
xnor U659 (N_659,In_992,In_1226);
and U660 (N_660,In_1488,In_36);
nand U661 (N_661,In_683,In_1445);
and U662 (N_662,In_918,In_1254);
and U663 (N_663,In_619,In_964);
or U664 (N_664,In_867,In_1260);
nand U665 (N_665,In_705,In_136);
or U666 (N_666,In_509,In_232);
nand U667 (N_667,In_993,In_532);
or U668 (N_668,In_935,In_1102);
nor U669 (N_669,In_511,In_740);
nand U670 (N_670,In_715,In_1490);
and U671 (N_671,In_171,In_1351);
and U672 (N_672,In_1109,In_883);
and U673 (N_673,In_1118,In_1346);
nor U674 (N_674,In_104,In_793);
nand U675 (N_675,In_904,In_112);
xor U676 (N_676,In_229,In_643);
xor U677 (N_677,In_1441,In_55);
nand U678 (N_678,In_846,In_1311);
nand U679 (N_679,In_1090,In_1312);
nor U680 (N_680,In_1044,In_739);
or U681 (N_681,In_440,In_656);
nand U682 (N_682,In_1158,In_1110);
nand U683 (N_683,In_1349,In_886);
nand U684 (N_684,In_1456,In_274);
or U685 (N_685,In_1082,In_627);
nor U686 (N_686,In_750,In_1408);
and U687 (N_687,In_1324,In_880);
or U688 (N_688,In_197,In_742);
or U689 (N_689,In_1055,In_1381);
nand U690 (N_690,In_1328,In_52);
xor U691 (N_691,In_850,In_1413);
or U692 (N_692,In_455,In_366);
nand U693 (N_693,In_1493,In_82);
or U694 (N_694,In_891,In_1387);
nor U695 (N_695,In_1181,In_447);
and U696 (N_696,In_555,In_1333);
nor U697 (N_697,In_1357,In_1126);
nor U698 (N_698,In_1331,In_1066);
and U699 (N_699,In_1081,In_1268);
and U700 (N_700,In_261,In_829);
and U701 (N_701,In_864,In_1283);
or U702 (N_702,In_1391,In_241);
or U703 (N_703,In_258,In_87);
nand U704 (N_704,In_819,In_460);
and U705 (N_705,In_1438,In_268);
nand U706 (N_706,In_876,In_49);
and U707 (N_707,In_390,In_774);
or U708 (N_708,In_369,In_481);
or U709 (N_709,In_70,In_1017);
nand U710 (N_710,In_1027,In_556);
or U711 (N_711,In_822,In_889);
nor U712 (N_712,In_225,In_689);
and U713 (N_713,In_776,In_132);
xnor U714 (N_714,In_485,In_207);
or U715 (N_715,In_983,In_143);
nor U716 (N_716,In_558,In_1290);
or U717 (N_717,In_853,In_153);
nor U718 (N_718,In_381,In_1099);
nor U719 (N_719,In_432,In_218);
xor U720 (N_720,In_834,In_1157);
or U721 (N_721,In_540,In_1435);
and U722 (N_722,In_135,In_877);
and U723 (N_723,In_176,In_530);
and U724 (N_724,In_1369,In_279);
nor U725 (N_725,In_291,In_1144);
and U726 (N_726,In_1350,In_358);
or U727 (N_727,In_1335,In_406);
xnor U728 (N_728,In_1434,In_302);
or U729 (N_729,In_1303,In_605);
nor U730 (N_730,In_410,In_1205);
or U731 (N_731,In_1341,In_1275);
nand U732 (N_732,In_23,In_1323);
xor U733 (N_733,In_1131,In_920);
and U734 (N_734,In_442,In_204);
nor U735 (N_735,In_570,In_194);
nor U736 (N_736,In_896,In_1474);
and U737 (N_737,In_673,In_707);
and U738 (N_738,In_946,In_41);
xor U739 (N_739,In_1370,In_273);
nand U740 (N_740,In_342,In_922);
nand U741 (N_741,In_1340,In_476);
and U742 (N_742,In_974,In_484);
and U743 (N_743,In_339,In_1193);
nor U744 (N_744,In_412,In_1013);
xnor U745 (N_745,In_1195,In_235);
or U746 (N_746,In_991,In_692);
and U747 (N_747,In_1052,In_483);
nor U748 (N_748,In_684,In_855);
nand U749 (N_749,In_1049,In_413);
xnor U750 (N_750,In_850,In_1282);
or U751 (N_751,In_337,In_231);
nand U752 (N_752,In_1451,In_759);
or U753 (N_753,In_330,In_1185);
and U754 (N_754,In_165,In_823);
and U755 (N_755,In_830,In_1100);
or U756 (N_756,In_883,In_550);
or U757 (N_757,In_152,In_870);
nor U758 (N_758,In_838,In_830);
and U759 (N_759,In_1478,In_1441);
nor U760 (N_760,In_770,In_1290);
xnor U761 (N_761,In_1262,In_962);
nand U762 (N_762,In_1401,In_70);
or U763 (N_763,In_462,In_734);
and U764 (N_764,In_241,In_45);
and U765 (N_765,In_1467,In_1490);
or U766 (N_766,In_755,In_1144);
and U767 (N_767,In_1110,In_481);
nand U768 (N_768,In_1164,In_419);
and U769 (N_769,In_1213,In_918);
or U770 (N_770,In_964,In_729);
xor U771 (N_771,In_25,In_165);
nand U772 (N_772,In_1092,In_1245);
xnor U773 (N_773,In_911,In_942);
and U774 (N_774,In_278,In_451);
nor U775 (N_775,In_1214,In_565);
nor U776 (N_776,In_888,In_73);
and U777 (N_777,In_1331,In_200);
nor U778 (N_778,In_1209,In_611);
nor U779 (N_779,In_848,In_815);
or U780 (N_780,In_408,In_1328);
and U781 (N_781,In_1127,In_949);
or U782 (N_782,In_1338,In_129);
or U783 (N_783,In_1459,In_913);
nand U784 (N_784,In_136,In_1042);
nor U785 (N_785,In_1093,In_1296);
and U786 (N_786,In_350,In_50);
and U787 (N_787,In_1077,In_1108);
and U788 (N_788,In_1303,In_931);
nor U789 (N_789,In_629,In_1355);
or U790 (N_790,In_1457,In_36);
or U791 (N_791,In_1332,In_423);
or U792 (N_792,In_1184,In_473);
or U793 (N_793,In_978,In_290);
nand U794 (N_794,In_1052,In_88);
or U795 (N_795,In_234,In_1472);
nor U796 (N_796,In_1487,In_1199);
xnor U797 (N_797,In_733,In_227);
nor U798 (N_798,In_408,In_933);
or U799 (N_799,In_787,In_88);
or U800 (N_800,In_673,In_1268);
and U801 (N_801,In_325,In_1079);
and U802 (N_802,In_338,In_164);
nor U803 (N_803,In_169,In_792);
and U804 (N_804,In_184,In_992);
nor U805 (N_805,In_542,In_1189);
or U806 (N_806,In_999,In_1101);
or U807 (N_807,In_816,In_964);
nand U808 (N_808,In_356,In_387);
nor U809 (N_809,In_349,In_281);
nand U810 (N_810,In_936,In_1207);
or U811 (N_811,In_982,In_1223);
nor U812 (N_812,In_1082,In_1230);
or U813 (N_813,In_1403,In_325);
nand U814 (N_814,In_98,In_167);
nand U815 (N_815,In_1352,In_1462);
nor U816 (N_816,In_857,In_293);
nor U817 (N_817,In_1329,In_1360);
and U818 (N_818,In_361,In_240);
nand U819 (N_819,In_676,In_68);
xnor U820 (N_820,In_1007,In_70);
nor U821 (N_821,In_782,In_343);
or U822 (N_822,In_1172,In_349);
nor U823 (N_823,In_1318,In_1411);
and U824 (N_824,In_1467,In_264);
and U825 (N_825,In_190,In_749);
or U826 (N_826,In_986,In_646);
nor U827 (N_827,In_663,In_886);
nor U828 (N_828,In_264,In_1426);
and U829 (N_829,In_314,In_1202);
nor U830 (N_830,In_872,In_1305);
nor U831 (N_831,In_200,In_103);
nand U832 (N_832,In_906,In_1431);
nand U833 (N_833,In_1323,In_990);
or U834 (N_834,In_569,In_1051);
xnor U835 (N_835,In_822,In_579);
or U836 (N_836,In_836,In_791);
or U837 (N_837,In_1189,In_1269);
nor U838 (N_838,In_20,In_970);
xnor U839 (N_839,In_872,In_1343);
nand U840 (N_840,In_1123,In_1235);
nor U841 (N_841,In_148,In_1126);
nand U842 (N_842,In_774,In_1346);
and U843 (N_843,In_795,In_194);
nand U844 (N_844,In_1280,In_1269);
xnor U845 (N_845,In_1460,In_95);
nand U846 (N_846,In_775,In_56);
xor U847 (N_847,In_606,In_320);
and U848 (N_848,In_209,In_497);
nor U849 (N_849,In_1429,In_741);
nor U850 (N_850,In_1490,In_211);
and U851 (N_851,In_163,In_854);
and U852 (N_852,In_300,In_534);
or U853 (N_853,In_891,In_1417);
nor U854 (N_854,In_438,In_290);
and U855 (N_855,In_1461,In_625);
nand U856 (N_856,In_1044,In_636);
and U857 (N_857,In_1418,In_799);
and U858 (N_858,In_1119,In_31);
and U859 (N_859,In_525,In_867);
and U860 (N_860,In_17,In_499);
xor U861 (N_861,In_1360,In_205);
or U862 (N_862,In_1457,In_548);
nor U863 (N_863,In_1358,In_1133);
or U864 (N_864,In_519,In_1124);
nand U865 (N_865,In_1088,In_1148);
nor U866 (N_866,In_908,In_317);
nand U867 (N_867,In_1292,In_261);
and U868 (N_868,In_489,In_178);
or U869 (N_869,In_134,In_331);
and U870 (N_870,In_834,In_30);
and U871 (N_871,In_1307,In_529);
xor U872 (N_872,In_55,In_1113);
nand U873 (N_873,In_426,In_1343);
and U874 (N_874,In_1288,In_989);
nand U875 (N_875,In_1408,In_772);
nand U876 (N_876,In_482,In_53);
nor U877 (N_877,In_606,In_583);
and U878 (N_878,In_1057,In_45);
or U879 (N_879,In_976,In_713);
and U880 (N_880,In_40,In_1378);
or U881 (N_881,In_99,In_460);
nor U882 (N_882,In_871,In_368);
nand U883 (N_883,In_1407,In_1260);
xor U884 (N_884,In_30,In_1492);
xor U885 (N_885,In_318,In_1340);
or U886 (N_886,In_246,In_1460);
or U887 (N_887,In_1097,In_1458);
or U888 (N_888,In_689,In_1441);
nand U889 (N_889,In_227,In_766);
nor U890 (N_890,In_1049,In_1010);
nand U891 (N_891,In_619,In_1226);
nand U892 (N_892,In_1064,In_1107);
and U893 (N_893,In_1319,In_1011);
xor U894 (N_894,In_884,In_621);
nand U895 (N_895,In_911,In_371);
nor U896 (N_896,In_1080,In_610);
or U897 (N_897,In_161,In_511);
xnor U898 (N_898,In_983,In_1114);
nor U899 (N_899,In_1006,In_856);
nor U900 (N_900,In_1491,In_224);
nand U901 (N_901,In_1269,In_211);
nand U902 (N_902,In_1038,In_708);
or U903 (N_903,In_285,In_836);
and U904 (N_904,In_617,In_1021);
nand U905 (N_905,In_1157,In_18);
nor U906 (N_906,In_785,In_651);
and U907 (N_907,In_1251,In_503);
nor U908 (N_908,In_937,In_1339);
nand U909 (N_909,In_24,In_671);
xnor U910 (N_910,In_443,In_763);
nor U911 (N_911,In_468,In_1075);
nand U912 (N_912,In_1439,In_1355);
nand U913 (N_913,In_201,In_1141);
or U914 (N_914,In_1283,In_543);
xnor U915 (N_915,In_1171,In_1052);
nor U916 (N_916,In_481,In_1283);
and U917 (N_917,In_873,In_271);
nor U918 (N_918,In_1191,In_1103);
nand U919 (N_919,In_1271,In_1395);
nand U920 (N_920,In_1392,In_67);
or U921 (N_921,In_1161,In_1343);
nand U922 (N_922,In_432,In_582);
nand U923 (N_923,In_1342,In_448);
nor U924 (N_924,In_475,In_404);
or U925 (N_925,In_520,In_1428);
nor U926 (N_926,In_86,In_1371);
nor U927 (N_927,In_868,In_842);
and U928 (N_928,In_1240,In_395);
nor U929 (N_929,In_317,In_1020);
or U930 (N_930,In_292,In_196);
nand U931 (N_931,In_1385,In_1142);
nand U932 (N_932,In_681,In_1051);
xor U933 (N_933,In_380,In_873);
nor U934 (N_934,In_96,In_19);
nor U935 (N_935,In_564,In_1299);
or U936 (N_936,In_639,In_1346);
nor U937 (N_937,In_298,In_679);
nor U938 (N_938,In_893,In_437);
nand U939 (N_939,In_272,In_26);
or U940 (N_940,In_1481,In_352);
xnor U941 (N_941,In_1089,In_574);
and U942 (N_942,In_1427,In_635);
and U943 (N_943,In_1055,In_1208);
or U944 (N_944,In_641,In_1263);
or U945 (N_945,In_280,In_1169);
nor U946 (N_946,In_1204,In_1474);
and U947 (N_947,In_1193,In_410);
or U948 (N_948,In_181,In_300);
nand U949 (N_949,In_1447,In_808);
nor U950 (N_950,In_1289,In_1042);
nor U951 (N_951,In_88,In_274);
xor U952 (N_952,In_748,In_1056);
nand U953 (N_953,In_755,In_1163);
and U954 (N_954,In_1105,In_719);
or U955 (N_955,In_515,In_966);
nor U956 (N_956,In_478,In_1174);
and U957 (N_957,In_1331,In_875);
or U958 (N_958,In_678,In_1294);
nand U959 (N_959,In_207,In_714);
nor U960 (N_960,In_682,In_1245);
or U961 (N_961,In_1019,In_1195);
nor U962 (N_962,In_650,In_859);
nand U963 (N_963,In_977,In_592);
or U964 (N_964,In_15,In_318);
or U965 (N_965,In_315,In_1138);
nand U966 (N_966,In_506,In_584);
and U967 (N_967,In_304,In_809);
nor U968 (N_968,In_410,In_1456);
nand U969 (N_969,In_745,In_505);
and U970 (N_970,In_413,In_687);
and U971 (N_971,In_1484,In_310);
and U972 (N_972,In_1187,In_1184);
nor U973 (N_973,In_568,In_1358);
xor U974 (N_974,In_472,In_1331);
or U975 (N_975,In_1008,In_1397);
and U976 (N_976,In_91,In_1014);
nand U977 (N_977,In_310,In_446);
or U978 (N_978,In_1261,In_20);
nand U979 (N_979,In_610,In_96);
and U980 (N_980,In_551,In_266);
nor U981 (N_981,In_374,In_1393);
nand U982 (N_982,In_841,In_457);
and U983 (N_983,In_265,In_1306);
nand U984 (N_984,In_675,In_447);
and U985 (N_985,In_1194,In_1280);
and U986 (N_986,In_638,In_463);
nand U987 (N_987,In_834,In_1413);
nor U988 (N_988,In_1041,In_957);
and U989 (N_989,In_685,In_1224);
nor U990 (N_990,In_173,In_413);
xnor U991 (N_991,In_1354,In_78);
nand U992 (N_992,In_369,In_613);
and U993 (N_993,In_1401,In_679);
xnor U994 (N_994,In_1115,In_321);
nand U995 (N_995,In_1395,In_1213);
nor U996 (N_996,In_301,In_432);
nand U997 (N_997,In_103,In_123);
nand U998 (N_998,In_1387,In_1300);
or U999 (N_999,In_696,In_749);
nor U1000 (N_1000,N_618,N_286);
or U1001 (N_1001,N_127,N_399);
or U1002 (N_1002,N_590,N_948);
nor U1003 (N_1003,N_664,N_607);
and U1004 (N_1004,N_25,N_594);
and U1005 (N_1005,N_728,N_702);
xnor U1006 (N_1006,N_787,N_557);
and U1007 (N_1007,N_703,N_932);
nor U1008 (N_1008,N_410,N_54);
nor U1009 (N_1009,N_281,N_340);
nand U1010 (N_1010,N_640,N_271);
nand U1011 (N_1011,N_124,N_733);
nor U1012 (N_1012,N_236,N_168);
and U1013 (N_1013,N_441,N_626);
and U1014 (N_1014,N_167,N_817);
nand U1015 (N_1015,N_82,N_798);
and U1016 (N_1016,N_136,N_867);
or U1017 (N_1017,N_976,N_678);
nand U1018 (N_1018,N_114,N_674);
and U1019 (N_1019,N_103,N_216);
nor U1020 (N_1020,N_391,N_994);
nor U1021 (N_1021,N_879,N_934);
nor U1022 (N_1022,N_229,N_218);
or U1023 (N_1023,N_889,N_820);
and U1024 (N_1024,N_148,N_722);
xor U1025 (N_1025,N_108,N_790);
xor U1026 (N_1026,N_219,N_356);
nor U1027 (N_1027,N_427,N_40);
nor U1028 (N_1028,N_824,N_378);
or U1029 (N_1029,N_936,N_525);
and U1030 (N_1030,N_969,N_331);
or U1031 (N_1031,N_380,N_263);
nand U1032 (N_1032,N_895,N_428);
or U1033 (N_1033,N_848,N_488);
nor U1034 (N_1034,N_1,N_294);
nor U1035 (N_1035,N_291,N_395);
xnor U1036 (N_1036,N_914,N_650);
or U1037 (N_1037,N_111,N_169);
nor U1038 (N_1038,N_486,N_581);
nor U1039 (N_1039,N_516,N_966);
xor U1040 (N_1040,N_6,N_116);
and U1041 (N_1041,N_933,N_632);
nand U1042 (N_1042,N_579,N_426);
nand U1043 (N_1043,N_425,N_446);
xnor U1044 (N_1044,N_361,N_953);
nand U1045 (N_1045,N_155,N_66);
or U1046 (N_1046,N_792,N_503);
nand U1047 (N_1047,N_133,N_849);
nor U1048 (N_1048,N_520,N_444);
or U1049 (N_1049,N_173,N_959);
nor U1050 (N_1050,N_962,N_660);
nand U1051 (N_1051,N_203,N_107);
nor U1052 (N_1052,N_891,N_705);
nand U1053 (N_1053,N_862,N_911);
nand U1054 (N_1054,N_95,N_414);
nand U1055 (N_1055,N_839,N_987);
xnor U1056 (N_1056,N_611,N_42);
or U1057 (N_1057,N_559,N_573);
nor U1058 (N_1058,N_756,N_711);
or U1059 (N_1059,N_368,N_81);
nand U1060 (N_1060,N_970,N_975);
nand U1061 (N_1061,N_4,N_697);
nand U1062 (N_1062,N_188,N_997);
or U1063 (N_1063,N_985,N_898);
and U1064 (N_1064,N_699,N_471);
and U1065 (N_1065,N_350,N_35);
and U1066 (N_1066,N_869,N_726);
or U1067 (N_1067,N_7,N_893);
and U1068 (N_1068,N_298,N_299);
nand U1069 (N_1069,N_314,N_113);
nor U1070 (N_1070,N_125,N_715);
nand U1071 (N_1071,N_724,N_585);
xnor U1072 (N_1072,N_877,N_473);
xnor U1073 (N_1073,N_465,N_179);
or U1074 (N_1074,N_77,N_762);
xor U1075 (N_1075,N_161,N_913);
nand U1076 (N_1076,N_900,N_905);
and U1077 (N_1077,N_600,N_661);
xor U1078 (N_1078,N_138,N_199);
or U1079 (N_1079,N_55,N_770);
or U1080 (N_1080,N_121,N_625);
and U1081 (N_1081,N_595,N_819);
nor U1082 (N_1082,N_400,N_170);
or U1083 (N_1083,N_261,N_589);
nor U1084 (N_1084,N_177,N_463);
or U1085 (N_1085,N_289,N_739);
nor U1086 (N_1086,N_135,N_100);
nand U1087 (N_1087,N_137,N_126);
nor U1088 (N_1088,N_531,N_878);
and U1089 (N_1089,N_897,N_751);
or U1090 (N_1090,N_815,N_822);
xor U1091 (N_1091,N_194,N_417);
nor U1092 (N_1092,N_608,N_193);
or U1093 (N_1093,N_231,N_612);
xor U1094 (N_1094,N_651,N_556);
and U1095 (N_1095,N_569,N_880);
and U1096 (N_1096,N_840,N_220);
and U1097 (N_1097,N_307,N_498);
nand U1098 (N_1098,N_892,N_712);
nor U1099 (N_1099,N_282,N_580);
and U1100 (N_1100,N_48,N_799);
or U1101 (N_1101,N_980,N_338);
nor U1102 (N_1102,N_487,N_430);
and U1103 (N_1103,N_431,N_649);
nor U1104 (N_1104,N_535,N_260);
and U1105 (N_1105,N_637,N_662);
nand U1106 (N_1106,N_552,N_492);
nor U1107 (N_1107,N_311,N_690);
or U1108 (N_1108,N_795,N_484);
nor U1109 (N_1109,N_514,N_527);
and U1110 (N_1110,N_285,N_894);
xor U1111 (N_1111,N_719,N_935);
xnor U1112 (N_1112,N_205,N_293);
or U1113 (N_1113,N_224,N_388);
or U1114 (N_1114,N_825,N_49);
xnor U1115 (N_1115,N_477,N_554);
nor U1116 (N_1116,N_39,N_254);
xnor U1117 (N_1117,N_646,N_351);
nand U1118 (N_1118,N_13,N_19);
nor U1119 (N_1119,N_720,N_404);
xor U1120 (N_1120,N_478,N_258);
nor U1121 (N_1121,N_863,N_511);
nand U1122 (N_1122,N_567,N_575);
or U1123 (N_1123,N_782,N_506);
and U1124 (N_1124,N_382,N_807);
nor U1125 (N_1125,N_460,N_371);
nand U1126 (N_1126,N_445,N_960);
nor U1127 (N_1127,N_729,N_154);
nand U1128 (N_1128,N_922,N_616);
nor U1129 (N_1129,N_51,N_67);
or U1130 (N_1130,N_367,N_232);
nor U1131 (N_1131,N_234,N_887);
and U1132 (N_1132,N_313,N_735);
nand U1133 (N_1133,N_747,N_659);
xnor U1134 (N_1134,N_686,N_475);
and U1135 (N_1135,N_207,N_206);
nor U1136 (N_1136,N_504,N_539);
xnor U1137 (N_1137,N_283,N_944);
xnor U1138 (N_1138,N_160,N_680);
nor U1139 (N_1139,N_904,N_571);
or U1140 (N_1140,N_93,N_939);
or U1141 (N_1141,N_376,N_278);
nand U1142 (N_1142,N_406,N_90);
and U1143 (N_1143,N_749,N_890);
and U1144 (N_1144,N_10,N_33);
and U1145 (N_1145,N_85,N_467);
or U1146 (N_1146,N_109,N_639);
xor U1147 (N_1147,N_295,N_968);
or U1148 (N_1148,N_725,N_708);
or U1149 (N_1149,N_786,N_204);
nand U1150 (N_1150,N_946,N_472);
and U1151 (N_1151,N_112,N_192);
or U1152 (N_1152,N_494,N_65);
xnor U1153 (N_1153,N_978,N_779);
and U1154 (N_1154,N_238,N_8);
and U1155 (N_1155,N_622,N_437);
and U1156 (N_1156,N_620,N_252);
nor U1157 (N_1157,N_122,N_507);
nor U1158 (N_1158,N_627,N_588);
nor U1159 (N_1159,N_584,N_115);
and U1160 (N_1160,N_663,N_163);
or U1161 (N_1161,N_587,N_954);
nand U1162 (N_1162,N_518,N_866);
nand U1163 (N_1163,N_439,N_644);
xor U1164 (N_1164,N_26,N_306);
or U1165 (N_1165,N_619,N_777);
and U1166 (N_1166,N_718,N_865);
or U1167 (N_1167,N_459,N_316);
nand U1168 (N_1168,N_450,N_732);
nor U1169 (N_1169,N_772,N_609);
or U1170 (N_1170,N_642,N_783);
nor U1171 (N_1171,N_146,N_424);
nand U1172 (N_1172,N_211,N_265);
and U1173 (N_1173,N_208,N_268);
nor U1174 (N_1174,N_166,N_131);
or U1175 (N_1175,N_117,N_931);
and U1176 (N_1176,N_916,N_24);
nand U1177 (N_1177,N_906,N_244);
nor U1178 (N_1178,N_752,N_951);
nand U1179 (N_1179,N_123,N_270);
nor U1180 (N_1180,N_563,N_704);
xnor U1181 (N_1181,N_657,N_280);
or U1182 (N_1182,N_604,N_876);
and U1183 (N_1183,N_185,N_264);
nor U1184 (N_1184,N_16,N_334);
nor U1185 (N_1185,N_476,N_746);
nand U1186 (N_1186,N_755,N_390);
or U1187 (N_1187,N_730,N_920);
or U1188 (N_1188,N_566,N_249);
and U1189 (N_1189,N_748,N_707);
or U1190 (N_1190,N_360,N_583);
nand U1191 (N_1191,N_423,N_63);
nand U1192 (N_1192,N_700,N_50);
and U1193 (N_1193,N_734,N_741);
and U1194 (N_1194,N_78,N_383);
xor U1195 (N_1195,N_709,N_23);
and U1196 (N_1196,N_189,N_989);
and U1197 (N_1197,N_530,N_673);
nand U1198 (N_1198,N_451,N_5);
or U1199 (N_1199,N_793,N_176);
and U1200 (N_1200,N_499,N_836);
and U1201 (N_1201,N_621,N_140);
or U1202 (N_1202,N_455,N_648);
nor U1203 (N_1203,N_297,N_780);
xnor U1204 (N_1204,N_788,N_462);
and U1205 (N_1205,N_676,N_397);
xnor U1206 (N_1206,N_977,N_757);
or U1207 (N_1207,N_183,N_631);
or U1208 (N_1208,N_346,N_603);
nand U1209 (N_1209,N_32,N_101);
nand U1210 (N_1210,N_949,N_352);
nand U1211 (N_1211,N_191,N_829);
or U1212 (N_1212,N_420,N_613);
and U1213 (N_1213,N_28,N_277);
and U1214 (N_1214,N_534,N_551);
or U1215 (N_1215,N_689,N_309);
xor U1216 (N_1216,N_60,N_358);
or U1217 (N_1217,N_810,N_841);
nor U1218 (N_1218,N_667,N_828);
and U1219 (N_1219,N_21,N_458);
or U1220 (N_1220,N_129,N_921);
and U1221 (N_1221,N_992,N_64);
nand U1222 (N_1222,N_442,N_979);
nand U1223 (N_1223,N_778,N_528);
nor U1224 (N_1224,N_687,N_447);
nor U1225 (N_1225,N_89,N_186);
or U1226 (N_1226,N_636,N_88);
nor U1227 (N_1227,N_61,N_804);
nand U1228 (N_1228,N_405,N_41);
nor U1229 (N_1229,N_775,N_86);
nand U1230 (N_1230,N_469,N_957);
and U1231 (N_1231,N_149,N_940);
and U1232 (N_1232,N_403,N_481);
nor U1233 (N_1233,N_14,N_562);
or U1234 (N_1234,N_927,N_72);
or U1235 (N_1235,N_731,N_134);
or U1236 (N_1236,N_74,N_461);
nand U1237 (N_1237,N_243,N_744);
and U1238 (N_1238,N_982,N_990);
and U1239 (N_1239,N_118,N_312);
and U1240 (N_1240,N_529,N_102);
and U1241 (N_1241,N_105,N_402);
or U1242 (N_1242,N_303,N_235);
or U1243 (N_1243,N_345,N_513);
or U1244 (N_1244,N_760,N_858);
or U1245 (N_1245,N_596,N_578);
or U1246 (N_1246,N_130,N_643);
nor U1247 (N_1247,N_438,N_999);
or U1248 (N_1248,N_723,N_242);
nand U1249 (N_1249,N_485,N_468);
nand U1250 (N_1250,N_682,N_685);
nand U1251 (N_1251,N_267,N_961);
nand U1252 (N_1252,N_34,N_342);
nor U1253 (N_1253,N_698,N_986);
nor U1254 (N_1254,N_805,N_577);
or U1255 (N_1255,N_918,N_572);
and U1256 (N_1256,N_681,N_813);
and U1257 (N_1257,N_721,N_943);
or U1258 (N_1258,N_677,N_500);
nand U1259 (N_1259,N_991,N_753);
nor U1260 (N_1260,N_217,N_175);
and U1261 (N_1261,N_771,N_310);
nor U1262 (N_1262,N_493,N_292);
xor U1263 (N_1263,N_262,N_187);
nor U1264 (N_1264,N_198,N_683);
xor U1265 (N_1265,N_381,N_318);
xnor U1266 (N_1266,N_347,N_925);
and U1267 (N_1267,N_964,N_882);
nor U1268 (N_1268,N_370,N_190);
nor U1269 (N_1269,N_323,N_266);
and U1270 (N_1270,N_706,N_502);
or U1271 (N_1271,N_870,N_76);
nand U1272 (N_1272,N_963,N_328);
and U1273 (N_1273,N_791,N_623);
nor U1274 (N_1274,N_389,N_510);
or U1275 (N_1275,N_326,N_174);
or U1276 (N_1276,N_765,N_348);
nand U1277 (N_1277,N_945,N_561);
or U1278 (N_1278,N_830,N_213);
and U1279 (N_1279,N_246,N_509);
nand U1280 (N_1280,N_57,N_222);
nor U1281 (N_1281,N_816,N_809);
and U1282 (N_1282,N_157,N_550);
nor U1283 (N_1283,N_432,N_415);
xor U1284 (N_1284,N_330,N_320);
nand U1285 (N_1285,N_287,N_296);
or U1286 (N_1286,N_110,N_714);
or U1287 (N_1287,N_716,N_106);
or U1288 (N_1288,N_856,N_668);
xor U1289 (N_1289,N_495,N_408);
nor U1290 (N_1290,N_907,N_200);
nor U1291 (N_1291,N_272,N_541);
xor U1292 (N_1292,N_240,N_901);
and U1293 (N_1293,N_727,N_36);
and U1294 (N_1294,N_602,N_259);
nand U1295 (N_1295,N_653,N_926);
nand U1296 (N_1296,N_2,N_874);
nor U1297 (N_1297,N_119,N_253);
nand U1298 (N_1298,N_302,N_832);
xor U1299 (N_1299,N_924,N_542);
and U1300 (N_1300,N_322,N_821);
nor U1301 (N_1301,N_958,N_407);
nand U1302 (N_1302,N_75,N_0);
and U1303 (N_1303,N_20,N_864);
and U1304 (N_1304,N_372,N_142);
and U1305 (N_1305,N_339,N_656);
nor U1306 (N_1306,N_411,N_491);
and U1307 (N_1307,N_421,N_104);
xnor U1308 (N_1308,N_938,N_956);
nor U1309 (N_1309,N_181,N_274);
and U1310 (N_1310,N_9,N_457);
nand U1311 (N_1311,N_508,N_353);
nand U1312 (N_1312,N_851,N_479);
nor U1313 (N_1313,N_794,N_324);
and U1314 (N_1314,N_955,N_98);
xor U1315 (N_1315,N_92,N_496);
or U1316 (N_1316,N_433,N_670);
and U1317 (N_1317,N_152,N_517);
xor U1318 (N_1318,N_172,N_996);
or U1319 (N_1319,N_99,N_796);
nor U1320 (N_1320,N_256,N_385);
nand U1321 (N_1321,N_610,N_629);
or U1322 (N_1322,N_449,N_52);
nand U1323 (N_1323,N_327,N_827);
and U1324 (N_1324,N_436,N_941);
and U1325 (N_1325,N_141,N_568);
or U1326 (N_1326,N_315,N_929);
nand U1327 (N_1327,N_758,N_558);
or U1328 (N_1328,N_846,N_781);
or U1329 (N_1329,N_881,N_418);
or U1330 (N_1330,N_290,N_624);
xnor U1331 (N_1331,N_652,N_373);
and U1332 (N_1332,N_87,N_967);
nand U1333 (N_1333,N_548,N_132);
and U1334 (N_1334,N_91,N_31);
and U1335 (N_1335,N_392,N_344);
nand U1336 (N_1336,N_750,N_845);
or U1337 (N_1337,N_784,N_37);
xor U1338 (N_1338,N_482,N_973);
nor U1339 (N_1339,N_523,N_761);
or U1340 (N_1340,N_544,N_288);
and U1341 (N_1341,N_855,N_743);
xnor U1342 (N_1342,N_79,N_776);
nor U1343 (N_1343,N_713,N_165);
nor U1344 (N_1344,N_490,N_416);
or U1345 (N_1345,N_440,N_823);
nor U1346 (N_1346,N_972,N_615);
and U1347 (N_1347,N_574,N_226);
or U1348 (N_1348,N_645,N_362);
nand U1349 (N_1349,N_560,N_337);
xnor U1350 (N_1350,N_343,N_665);
and U1351 (N_1351,N_47,N_470);
and U1352 (N_1352,N_717,N_654);
xor U1353 (N_1353,N_852,N_909);
nand U1354 (N_1354,N_386,N_538);
or U1355 (N_1355,N_857,N_928);
or U1356 (N_1356,N_868,N_497);
or U1357 (N_1357,N_215,N_837);
or U1358 (N_1358,N_519,N_196);
and U1359 (N_1359,N_301,N_354);
or U1360 (N_1360,N_452,N_464);
and U1361 (N_1361,N_888,N_671);
or U1362 (N_1362,N_570,N_628);
nand U1363 (N_1363,N_885,N_145);
nor U1364 (N_1364,N_308,N_545);
and U1365 (N_1365,N_273,N_474);
nand U1366 (N_1366,N_71,N_30);
xnor U1367 (N_1367,N_802,N_147);
nand U1368 (N_1368,N_785,N_736);
nor U1369 (N_1369,N_582,N_228);
and U1370 (N_1370,N_696,N_917);
nand U1371 (N_1371,N_773,N_591);
and U1372 (N_1372,N_429,N_279);
or U1373 (N_1373,N_694,N_413);
or U1374 (N_1374,N_156,N_422);
nand U1375 (N_1375,N_97,N_740);
and U1376 (N_1376,N_526,N_319);
or U1377 (N_1377,N_801,N_11);
and U1378 (N_1378,N_764,N_164);
nand U1379 (N_1379,N_453,N_693);
xnor U1380 (N_1380,N_902,N_396);
nor U1381 (N_1381,N_701,N_903);
or U1382 (N_1382,N_230,N_988);
nor U1383 (N_1383,N_143,N_409);
or U1384 (N_1384,N_162,N_896);
and U1385 (N_1385,N_742,N_329);
or U1386 (N_1386,N_915,N_128);
nor U1387 (N_1387,N_871,N_349);
and U1388 (N_1388,N_592,N_838);
nand U1389 (N_1389,N_873,N_239);
or U1390 (N_1390,N_336,N_365);
or U1391 (N_1391,N_952,N_15);
nand U1392 (N_1392,N_835,N_923);
and U1393 (N_1393,N_672,N_767);
nor U1394 (N_1394,N_178,N_543);
xnor U1395 (N_1395,N_435,N_635);
xor U1396 (N_1396,N_3,N_214);
and U1397 (N_1397,N_44,N_180);
xor U1398 (N_1398,N_284,N_223);
nand U1399 (N_1399,N_384,N_355);
nor U1400 (N_1400,N_317,N_606);
nand U1401 (N_1401,N_335,N_853);
nor U1402 (N_1402,N_666,N_647);
or U1403 (N_1403,N_818,N_859);
xor U1404 (N_1404,N_547,N_251);
or U1405 (N_1405,N_159,N_375);
nand U1406 (N_1406,N_96,N_466);
or U1407 (N_1407,N_257,N_56);
nor U1408 (N_1408,N_212,N_598);
or U1409 (N_1409,N_221,N_658);
xor U1410 (N_1410,N_533,N_241);
and U1411 (N_1411,N_393,N_12);
and U1412 (N_1412,N_942,N_321);
or U1413 (N_1413,N_225,N_379);
nand U1414 (N_1414,N_505,N_374);
and U1415 (N_1415,N_971,N_59);
and U1416 (N_1416,N_248,N_861);
or U1417 (N_1417,N_811,N_831);
nand U1418 (N_1418,N_899,N_883);
and U1419 (N_1419,N_184,N_872);
and U1420 (N_1420,N_930,N_710);
and U1421 (N_1421,N_29,N_332);
and U1422 (N_1422,N_363,N_150);
or U1423 (N_1423,N_633,N_454);
or U1424 (N_1424,N_522,N_769);
nand U1425 (N_1425,N_369,N_549);
nor U1426 (N_1426,N_808,N_387);
and U1427 (N_1427,N_800,N_641);
nand U1428 (N_1428,N_675,N_669);
or U1429 (N_1429,N_919,N_443);
or U1430 (N_1430,N_974,N_182);
nand U1431 (N_1431,N_419,N_38);
nand U1432 (N_1432,N_201,N_908);
and U1433 (N_1433,N_69,N_512);
nand U1434 (N_1434,N_515,N_605);
and U1435 (N_1435,N_139,N_73);
and U1436 (N_1436,N_434,N_684);
or U1437 (N_1437,N_394,N_614);
and U1438 (N_1438,N_843,N_655);
nor U1439 (N_1439,N_333,N_195);
nand U1440 (N_1440,N_456,N_599);
and U1441 (N_1441,N_70,N_981);
and U1442 (N_1442,N_22,N_255);
or U1443 (N_1443,N_910,N_983);
or U1444 (N_1444,N_826,N_630);
or U1445 (N_1445,N_237,N_357);
and U1446 (N_1446,N_377,N_768);
xor U1447 (N_1447,N_850,N_58);
nand U1448 (N_1448,N_46,N_984);
or U1449 (N_1449,N_275,N_202);
nand U1450 (N_1450,N_833,N_83);
nand U1451 (N_1451,N_276,N_763);
nor U1452 (N_1452,N_300,N_84);
nor U1453 (N_1453,N_597,N_448);
nor U1454 (N_1454,N_68,N_227);
and U1455 (N_1455,N_27,N_171);
or U1456 (N_1456,N_521,N_158);
nor U1457 (N_1457,N_80,N_480);
and U1458 (N_1458,N_540,N_412);
nor U1459 (N_1459,N_738,N_45);
nor U1460 (N_1460,N_245,N_884);
nor U1461 (N_1461,N_17,N_993);
and U1462 (N_1462,N_501,N_737);
xnor U1463 (N_1463,N_886,N_53);
or U1464 (N_1464,N_912,N_269);
nor U1465 (N_1465,N_995,N_759);
and U1466 (N_1466,N_814,N_947);
nor U1467 (N_1467,N_564,N_553);
and U1468 (N_1468,N_489,N_197);
or U1469 (N_1469,N_601,N_847);
or U1470 (N_1470,N_18,N_62);
nand U1471 (N_1471,N_854,N_247);
nor U1472 (N_1472,N_695,N_233);
nand U1473 (N_1473,N_679,N_341);
xor U1474 (N_1474,N_860,N_565);
nor U1475 (N_1475,N_789,N_210);
nand U1476 (N_1476,N_555,N_812);
and U1477 (N_1477,N_634,N_844);
nand U1478 (N_1478,N_875,N_617);
nor U1479 (N_1479,N_305,N_524);
or U1480 (N_1480,N_304,N_797);
or U1481 (N_1481,N_842,N_691);
or U1482 (N_1482,N_754,N_745);
or U1483 (N_1483,N_638,N_546);
or U1484 (N_1484,N_43,N_937);
nor U1485 (N_1485,N_401,N_536);
nor U1486 (N_1486,N_688,N_532);
or U1487 (N_1487,N_965,N_120);
nor U1488 (N_1488,N_153,N_250);
and U1489 (N_1489,N_483,N_366);
nor U1490 (N_1490,N_803,N_593);
or U1491 (N_1491,N_325,N_692);
nor U1492 (N_1492,N_586,N_774);
and U1493 (N_1493,N_359,N_834);
xor U1494 (N_1494,N_144,N_998);
or U1495 (N_1495,N_806,N_151);
nand U1496 (N_1496,N_364,N_950);
and U1497 (N_1497,N_209,N_398);
nor U1498 (N_1498,N_766,N_576);
nand U1499 (N_1499,N_94,N_537);
nand U1500 (N_1500,N_371,N_139);
and U1501 (N_1501,N_974,N_418);
or U1502 (N_1502,N_800,N_724);
nand U1503 (N_1503,N_137,N_121);
or U1504 (N_1504,N_168,N_530);
or U1505 (N_1505,N_469,N_234);
xor U1506 (N_1506,N_866,N_379);
nand U1507 (N_1507,N_797,N_792);
or U1508 (N_1508,N_996,N_871);
xnor U1509 (N_1509,N_561,N_650);
xnor U1510 (N_1510,N_527,N_565);
or U1511 (N_1511,N_70,N_899);
nor U1512 (N_1512,N_787,N_746);
nor U1513 (N_1513,N_873,N_870);
nand U1514 (N_1514,N_85,N_18);
xnor U1515 (N_1515,N_507,N_678);
nand U1516 (N_1516,N_551,N_463);
xnor U1517 (N_1517,N_250,N_545);
nor U1518 (N_1518,N_117,N_432);
or U1519 (N_1519,N_542,N_15);
and U1520 (N_1520,N_399,N_93);
xnor U1521 (N_1521,N_409,N_961);
nor U1522 (N_1522,N_50,N_186);
nand U1523 (N_1523,N_776,N_787);
xnor U1524 (N_1524,N_302,N_892);
and U1525 (N_1525,N_905,N_971);
nand U1526 (N_1526,N_946,N_406);
or U1527 (N_1527,N_739,N_924);
nand U1528 (N_1528,N_463,N_710);
and U1529 (N_1529,N_925,N_577);
xnor U1530 (N_1530,N_430,N_81);
or U1531 (N_1531,N_185,N_588);
and U1532 (N_1532,N_213,N_425);
or U1533 (N_1533,N_276,N_436);
or U1534 (N_1534,N_612,N_168);
nand U1535 (N_1535,N_784,N_496);
xnor U1536 (N_1536,N_250,N_143);
and U1537 (N_1537,N_578,N_213);
nor U1538 (N_1538,N_867,N_206);
nand U1539 (N_1539,N_227,N_828);
xnor U1540 (N_1540,N_2,N_197);
nand U1541 (N_1541,N_735,N_319);
xnor U1542 (N_1542,N_565,N_928);
nand U1543 (N_1543,N_235,N_468);
nor U1544 (N_1544,N_789,N_477);
nor U1545 (N_1545,N_353,N_571);
and U1546 (N_1546,N_354,N_178);
nand U1547 (N_1547,N_873,N_950);
nand U1548 (N_1548,N_282,N_237);
nor U1549 (N_1549,N_71,N_917);
nand U1550 (N_1550,N_64,N_283);
and U1551 (N_1551,N_496,N_9);
nor U1552 (N_1552,N_208,N_613);
nand U1553 (N_1553,N_281,N_867);
or U1554 (N_1554,N_193,N_51);
or U1555 (N_1555,N_589,N_195);
and U1556 (N_1556,N_437,N_288);
nor U1557 (N_1557,N_792,N_282);
nor U1558 (N_1558,N_434,N_767);
nor U1559 (N_1559,N_883,N_876);
and U1560 (N_1560,N_145,N_204);
nor U1561 (N_1561,N_272,N_80);
or U1562 (N_1562,N_285,N_711);
nor U1563 (N_1563,N_31,N_279);
xnor U1564 (N_1564,N_247,N_301);
xnor U1565 (N_1565,N_229,N_630);
nor U1566 (N_1566,N_514,N_497);
or U1567 (N_1567,N_551,N_943);
nor U1568 (N_1568,N_196,N_944);
nor U1569 (N_1569,N_387,N_398);
nor U1570 (N_1570,N_178,N_199);
nand U1571 (N_1571,N_527,N_951);
nand U1572 (N_1572,N_569,N_415);
and U1573 (N_1573,N_200,N_742);
and U1574 (N_1574,N_938,N_369);
xor U1575 (N_1575,N_819,N_457);
xnor U1576 (N_1576,N_463,N_72);
or U1577 (N_1577,N_907,N_416);
xor U1578 (N_1578,N_994,N_626);
or U1579 (N_1579,N_105,N_289);
nor U1580 (N_1580,N_232,N_699);
nor U1581 (N_1581,N_566,N_442);
or U1582 (N_1582,N_193,N_44);
or U1583 (N_1583,N_278,N_864);
nand U1584 (N_1584,N_584,N_707);
and U1585 (N_1585,N_648,N_212);
or U1586 (N_1586,N_20,N_969);
nor U1587 (N_1587,N_988,N_164);
or U1588 (N_1588,N_752,N_42);
and U1589 (N_1589,N_550,N_905);
and U1590 (N_1590,N_35,N_805);
and U1591 (N_1591,N_955,N_625);
nor U1592 (N_1592,N_878,N_657);
or U1593 (N_1593,N_579,N_320);
nand U1594 (N_1594,N_688,N_682);
xnor U1595 (N_1595,N_666,N_225);
and U1596 (N_1596,N_895,N_810);
nand U1597 (N_1597,N_225,N_317);
xnor U1598 (N_1598,N_474,N_446);
xnor U1599 (N_1599,N_79,N_222);
nor U1600 (N_1600,N_12,N_594);
and U1601 (N_1601,N_257,N_937);
nor U1602 (N_1602,N_932,N_314);
or U1603 (N_1603,N_403,N_654);
xor U1604 (N_1604,N_433,N_651);
nand U1605 (N_1605,N_435,N_572);
nand U1606 (N_1606,N_423,N_968);
nand U1607 (N_1607,N_948,N_797);
nor U1608 (N_1608,N_565,N_26);
nor U1609 (N_1609,N_797,N_685);
nand U1610 (N_1610,N_459,N_735);
nand U1611 (N_1611,N_374,N_753);
nand U1612 (N_1612,N_370,N_469);
nand U1613 (N_1613,N_598,N_848);
or U1614 (N_1614,N_332,N_665);
and U1615 (N_1615,N_465,N_457);
xor U1616 (N_1616,N_378,N_700);
and U1617 (N_1617,N_884,N_133);
nor U1618 (N_1618,N_342,N_54);
xor U1619 (N_1619,N_378,N_197);
nor U1620 (N_1620,N_34,N_621);
nand U1621 (N_1621,N_603,N_524);
xnor U1622 (N_1622,N_321,N_596);
or U1623 (N_1623,N_856,N_690);
nor U1624 (N_1624,N_398,N_321);
nand U1625 (N_1625,N_618,N_461);
and U1626 (N_1626,N_650,N_520);
xor U1627 (N_1627,N_456,N_609);
nor U1628 (N_1628,N_295,N_249);
and U1629 (N_1629,N_270,N_819);
nand U1630 (N_1630,N_647,N_365);
or U1631 (N_1631,N_951,N_920);
and U1632 (N_1632,N_106,N_655);
nor U1633 (N_1633,N_391,N_304);
or U1634 (N_1634,N_327,N_4);
and U1635 (N_1635,N_671,N_585);
and U1636 (N_1636,N_873,N_929);
and U1637 (N_1637,N_368,N_338);
or U1638 (N_1638,N_2,N_326);
and U1639 (N_1639,N_395,N_719);
and U1640 (N_1640,N_229,N_659);
nor U1641 (N_1641,N_743,N_927);
and U1642 (N_1642,N_503,N_369);
or U1643 (N_1643,N_336,N_877);
or U1644 (N_1644,N_230,N_868);
or U1645 (N_1645,N_153,N_19);
and U1646 (N_1646,N_413,N_138);
or U1647 (N_1647,N_495,N_43);
nor U1648 (N_1648,N_148,N_855);
nor U1649 (N_1649,N_633,N_243);
and U1650 (N_1650,N_800,N_191);
nor U1651 (N_1651,N_541,N_709);
nand U1652 (N_1652,N_593,N_565);
nor U1653 (N_1653,N_731,N_620);
nor U1654 (N_1654,N_239,N_948);
or U1655 (N_1655,N_994,N_604);
and U1656 (N_1656,N_556,N_937);
or U1657 (N_1657,N_456,N_345);
and U1658 (N_1658,N_453,N_27);
or U1659 (N_1659,N_134,N_951);
xnor U1660 (N_1660,N_409,N_832);
nor U1661 (N_1661,N_120,N_333);
or U1662 (N_1662,N_551,N_896);
and U1663 (N_1663,N_453,N_829);
and U1664 (N_1664,N_536,N_391);
or U1665 (N_1665,N_894,N_94);
or U1666 (N_1666,N_537,N_41);
nand U1667 (N_1667,N_916,N_670);
nand U1668 (N_1668,N_137,N_532);
nor U1669 (N_1669,N_886,N_776);
xor U1670 (N_1670,N_465,N_641);
or U1671 (N_1671,N_715,N_71);
nor U1672 (N_1672,N_704,N_511);
nand U1673 (N_1673,N_536,N_967);
nor U1674 (N_1674,N_283,N_623);
and U1675 (N_1675,N_460,N_818);
xor U1676 (N_1676,N_893,N_803);
xnor U1677 (N_1677,N_427,N_128);
and U1678 (N_1678,N_454,N_956);
and U1679 (N_1679,N_169,N_316);
xnor U1680 (N_1680,N_851,N_463);
and U1681 (N_1681,N_706,N_774);
nor U1682 (N_1682,N_60,N_62);
nand U1683 (N_1683,N_91,N_965);
and U1684 (N_1684,N_174,N_483);
xnor U1685 (N_1685,N_113,N_348);
or U1686 (N_1686,N_441,N_328);
nor U1687 (N_1687,N_544,N_796);
nand U1688 (N_1688,N_336,N_715);
nand U1689 (N_1689,N_23,N_428);
or U1690 (N_1690,N_444,N_139);
and U1691 (N_1691,N_657,N_561);
nand U1692 (N_1692,N_655,N_43);
or U1693 (N_1693,N_927,N_840);
and U1694 (N_1694,N_140,N_799);
nand U1695 (N_1695,N_337,N_740);
xnor U1696 (N_1696,N_402,N_549);
nand U1697 (N_1697,N_906,N_875);
nor U1698 (N_1698,N_771,N_366);
nand U1699 (N_1699,N_723,N_502);
xnor U1700 (N_1700,N_383,N_936);
or U1701 (N_1701,N_5,N_21);
nor U1702 (N_1702,N_815,N_347);
and U1703 (N_1703,N_665,N_420);
xnor U1704 (N_1704,N_16,N_461);
nand U1705 (N_1705,N_183,N_583);
nor U1706 (N_1706,N_490,N_170);
and U1707 (N_1707,N_283,N_716);
and U1708 (N_1708,N_463,N_238);
nor U1709 (N_1709,N_334,N_145);
nand U1710 (N_1710,N_544,N_954);
xnor U1711 (N_1711,N_595,N_462);
xnor U1712 (N_1712,N_599,N_573);
nor U1713 (N_1713,N_237,N_796);
and U1714 (N_1714,N_189,N_537);
nor U1715 (N_1715,N_761,N_403);
or U1716 (N_1716,N_206,N_399);
or U1717 (N_1717,N_991,N_945);
or U1718 (N_1718,N_277,N_674);
nor U1719 (N_1719,N_612,N_448);
nor U1720 (N_1720,N_519,N_587);
nor U1721 (N_1721,N_28,N_959);
nand U1722 (N_1722,N_909,N_807);
nor U1723 (N_1723,N_18,N_489);
xnor U1724 (N_1724,N_54,N_753);
nor U1725 (N_1725,N_226,N_170);
and U1726 (N_1726,N_86,N_728);
nor U1727 (N_1727,N_624,N_881);
or U1728 (N_1728,N_227,N_171);
or U1729 (N_1729,N_102,N_522);
nor U1730 (N_1730,N_652,N_69);
and U1731 (N_1731,N_555,N_924);
or U1732 (N_1732,N_579,N_39);
and U1733 (N_1733,N_44,N_805);
nor U1734 (N_1734,N_770,N_83);
xor U1735 (N_1735,N_705,N_858);
and U1736 (N_1736,N_496,N_805);
nand U1737 (N_1737,N_275,N_124);
nor U1738 (N_1738,N_761,N_749);
xor U1739 (N_1739,N_28,N_753);
and U1740 (N_1740,N_656,N_692);
xor U1741 (N_1741,N_75,N_156);
xor U1742 (N_1742,N_674,N_406);
nor U1743 (N_1743,N_480,N_708);
and U1744 (N_1744,N_335,N_121);
or U1745 (N_1745,N_295,N_458);
and U1746 (N_1746,N_933,N_104);
nand U1747 (N_1747,N_375,N_503);
and U1748 (N_1748,N_889,N_286);
and U1749 (N_1749,N_563,N_646);
nor U1750 (N_1750,N_985,N_700);
nand U1751 (N_1751,N_67,N_367);
or U1752 (N_1752,N_800,N_526);
nor U1753 (N_1753,N_548,N_350);
nor U1754 (N_1754,N_836,N_682);
or U1755 (N_1755,N_992,N_135);
nor U1756 (N_1756,N_470,N_662);
and U1757 (N_1757,N_361,N_956);
and U1758 (N_1758,N_956,N_302);
nor U1759 (N_1759,N_444,N_741);
and U1760 (N_1760,N_104,N_999);
nor U1761 (N_1761,N_335,N_549);
xor U1762 (N_1762,N_948,N_125);
and U1763 (N_1763,N_138,N_680);
or U1764 (N_1764,N_948,N_456);
nor U1765 (N_1765,N_670,N_355);
and U1766 (N_1766,N_527,N_550);
or U1767 (N_1767,N_119,N_797);
or U1768 (N_1768,N_608,N_571);
or U1769 (N_1769,N_393,N_559);
and U1770 (N_1770,N_703,N_304);
nand U1771 (N_1771,N_604,N_957);
nand U1772 (N_1772,N_681,N_65);
nor U1773 (N_1773,N_690,N_68);
xnor U1774 (N_1774,N_917,N_666);
nand U1775 (N_1775,N_421,N_486);
nor U1776 (N_1776,N_752,N_48);
nand U1777 (N_1777,N_864,N_739);
nor U1778 (N_1778,N_933,N_916);
and U1779 (N_1779,N_107,N_7);
or U1780 (N_1780,N_929,N_69);
and U1781 (N_1781,N_249,N_314);
xor U1782 (N_1782,N_4,N_25);
or U1783 (N_1783,N_104,N_716);
or U1784 (N_1784,N_742,N_696);
nor U1785 (N_1785,N_831,N_792);
and U1786 (N_1786,N_599,N_150);
or U1787 (N_1787,N_615,N_481);
nand U1788 (N_1788,N_492,N_315);
or U1789 (N_1789,N_357,N_278);
or U1790 (N_1790,N_902,N_46);
nand U1791 (N_1791,N_849,N_393);
and U1792 (N_1792,N_956,N_924);
or U1793 (N_1793,N_414,N_897);
nor U1794 (N_1794,N_588,N_488);
or U1795 (N_1795,N_708,N_699);
nor U1796 (N_1796,N_974,N_173);
and U1797 (N_1797,N_846,N_271);
and U1798 (N_1798,N_367,N_602);
and U1799 (N_1799,N_923,N_598);
or U1800 (N_1800,N_79,N_493);
and U1801 (N_1801,N_817,N_197);
nand U1802 (N_1802,N_196,N_248);
and U1803 (N_1803,N_799,N_642);
xnor U1804 (N_1804,N_221,N_724);
nand U1805 (N_1805,N_273,N_986);
nand U1806 (N_1806,N_596,N_590);
nor U1807 (N_1807,N_897,N_772);
xor U1808 (N_1808,N_793,N_70);
and U1809 (N_1809,N_324,N_999);
nand U1810 (N_1810,N_964,N_397);
nor U1811 (N_1811,N_962,N_360);
nand U1812 (N_1812,N_982,N_646);
nor U1813 (N_1813,N_90,N_553);
and U1814 (N_1814,N_982,N_397);
xnor U1815 (N_1815,N_746,N_108);
nor U1816 (N_1816,N_929,N_374);
nand U1817 (N_1817,N_154,N_912);
nor U1818 (N_1818,N_485,N_3);
nor U1819 (N_1819,N_696,N_190);
nor U1820 (N_1820,N_497,N_572);
xor U1821 (N_1821,N_880,N_458);
nand U1822 (N_1822,N_193,N_329);
nand U1823 (N_1823,N_623,N_529);
or U1824 (N_1824,N_187,N_546);
and U1825 (N_1825,N_65,N_675);
nor U1826 (N_1826,N_981,N_485);
and U1827 (N_1827,N_203,N_291);
xnor U1828 (N_1828,N_839,N_233);
and U1829 (N_1829,N_725,N_31);
and U1830 (N_1830,N_206,N_787);
or U1831 (N_1831,N_917,N_771);
and U1832 (N_1832,N_55,N_350);
xnor U1833 (N_1833,N_632,N_883);
nor U1834 (N_1834,N_251,N_867);
nand U1835 (N_1835,N_165,N_808);
or U1836 (N_1836,N_21,N_885);
nor U1837 (N_1837,N_703,N_819);
or U1838 (N_1838,N_97,N_135);
nand U1839 (N_1839,N_787,N_696);
nor U1840 (N_1840,N_761,N_463);
nor U1841 (N_1841,N_242,N_670);
nor U1842 (N_1842,N_532,N_774);
nor U1843 (N_1843,N_774,N_732);
or U1844 (N_1844,N_99,N_852);
and U1845 (N_1845,N_921,N_424);
and U1846 (N_1846,N_988,N_436);
nand U1847 (N_1847,N_335,N_66);
nand U1848 (N_1848,N_2,N_553);
nand U1849 (N_1849,N_635,N_378);
nand U1850 (N_1850,N_980,N_254);
and U1851 (N_1851,N_828,N_780);
nor U1852 (N_1852,N_905,N_765);
xor U1853 (N_1853,N_924,N_497);
nor U1854 (N_1854,N_134,N_664);
xor U1855 (N_1855,N_98,N_759);
and U1856 (N_1856,N_958,N_38);
nor U1857 (N_1857,N_188,N_427);
and U1858 (N_1858,N_608,N_398);
nand U1859 (N_1859,N_612,N_992);
nor U1860 (N_1860,N_424,N_173);
and U1861 (N_1861,N_122,N_47);
and U1862 (N_1862,N_832,N_30);
nor U1863 (N_1863,N_675,N_876);
or U1864 (N_1864,N_969,N_46);
xor U1865 (N_1865,N_658,N_566);
or U1866 (N_1866,N_268,N_261);
xnor U1867 (N_1867,N_408,N_590);
or U1868 (N_1868,N_672,N_120);
and U1869 (N_1869,N_892,N_867);
xnor U1870 (N_1870,N_701,N_138);
xor U1871 (N_1871,N_76,N_122);
and U1872 (N_1872,N_600,N_671);
nor U1873 (N_1873,N_883,N_551);
xor U1874 (N_1874,N_531,N_113);
and U1875 (N_1875,N_327,N_270);
and U1876 (N_1876,N_588,N_77);
or U1877 (N_1877,N_199,N_429);
nand U1878 (N_1878,N_573,N_699);
and U1879 (N_1879,N_574,N_538);
or U1880 (N_1880,N_482,N_208);
or U1881 (N_1881,N_255,N_560);
xor U1882 (N_1882,N_902,N_743);
and U1883 (N_1883,N_446,N_976);
nor U1884 (N_1884,N_290,N_803);
xnor U1885 (N_1885,N_353,N_838);
nor U1886 (N_1886,N_201,N_140);
nor U1887 (N_1887,N_996,N_931);
or U1888 (N_1888,N_258,N_984);
and U1889 (N_1889,N_959,N_170);
nor U1890 (N_1890,N_466,N_551);
or U1891 (N_1891,N_540,N_927);
and U1892 (N_1892,N_550,N_399);
or U1893 (N_1893,N_212,N_634);
and U1894 (N_1894,N_264,N_965);
nor U1895 (N_1895,N_404,N_354);
nand U1896 (N_1896,N_835,N_904);
or U1897 (N_1897,N_376,N_632);
nand U1898 (N_1898,N_136,N_51);
nor U1899 (N_1899,N_943,N_101);
and U1900 (N_1900,N_773,N_462);
nor U1901 (N_1901,N_923,N_167);
and U1902 (N_1902,N_648,N_451);
and U1903 (N_1903,N_670,N_140);
or U1904 (N_1904,N_631,N_395);
nor U1905 (N_1905,N_117,N_97);
nand U1906 (N_1906,N_294,N_829);
and U1907 (N_1907,N_634,N_570);
and U1908 (N_1908,N_485,N_557);
nor U1909 (N_1909,N_816,N_421);
or U1910 (N_1910,N_445,N_628);
xnor U1911 (N_1911,N_265,N_281);
and U1912 (N_1912,N_611,N_78);
or U1913 (N_1913,N_761,N_178);
and U1914 (N_1914,N_106,N_756);
xnor U1915 (N_1915,N_681,N_84);
and U1916 (N_1916,N_161,N_784);
and U1917 (N_1917,N_720,N_128);
nor U1918 (N_1918,N_894,N_342);
and U1919 (N_1919,N_599,N_910);
nand U1920 (N_1920,N_640,N_480);
or U1921 (N_1921,N_608,N_910);
xnor U1922 (N_1922,N_611,N_658);
or U1923 (N_1923,N_580,N_418);
nand U1924 (N_1924,N_78,N_675);
and U1925 (N_1925,N_447,N_289);
nand U1926 (N_1926,N_851,N_123);
xor U1927 (N_1927,N_900,N_960);
nand U1928 (N_1928,N_731,N_535);
nor U1929 (N_1929,N_979,N_199);
and U1930 (N_1930,N_25,N_198);
nand U1931 (N_1931,N_922,N_702);
or U1932 (N_1932,N_740,N_982);
nor U1933 (N_1933,N_215,N_770);
xor U1934 (N_1934,N_24,N_870);
nor U1935 (N_1935,N_836,N_799);
or U1936 (N_1936,N_310,N_776);
nor U1937 (N_1937,N_277,N_609);
nand U1938 (N_1938,N_806,N_312);
nor U1939 (N_1939,N_25,N_63);
nor U1940 (N_1940,N_674,N_646);
xnor U1941 (N_1941,N_565,N_818);
nor U1942 (N_1942,N_47,N_326);
nand U1943 (N_1943,N_117,N_550);
xor U1944 (N_1944,N_855,N_323);
or U1945 (N_1945,N_327,N_217);
nand U1946 (N_1946,N_746,N_546);
and U1947 (N_1947,N_906,N_474);
nor U1948 (N_1948,N_400,N_143);
nand U1949 (N_1949,N_197,N_884);
and U1950 (N_1950,N_298,N_594);
nand U1951 (N_1951,N_489,N_906);
nor U1952 (N_1952,N_380,N_366);
xor U1953 (N_1953,N_975,N_541);
or U1954 (N_1954,N_626,N_38);
and U1955 (N_1955,N_772,N_738);
nand U1956 (N_1956,N_520,N_90);
nand U1957 (N_1957,N_406,N_267);
and U1958 (N_1958,N_714,N_277);
nor U1959 (N_1959,N_207,N_741);
nand U1960 (N_1960,N_277,N_193);
nor U1961 (N_1961,N_738,N_314);
or U1962 (N_1962,N_583,N_709);
xor U1963 (N_1963,N_173,N_63);
and U1964 (N_1964,N_89,N_46);
nor U1965 (N_1965,N_760,N_179);
nand U1966 (N_1966,N_483,N_571);
nand U1967 (N_1967,N_399,N_685);
and U1968 (N_1968,N_783,N_955);
nand U1969 (N_1969,N_179,N_320);
and U1970 (N_1970,N_283,N_525);
or U1971 (N_1971,N_480,N_51);
xnor U1972 (N_1972,N_533,N_950);
or U1973 (N_1973,N_298,N_421);
or U1974 (N_1974,N_978,N_639);
nand U1975 (N_1975,N_774,N_744);
xnor U1976 (N_1976,N_505,N_269);
nor U1977 (N_1977,N_636,N_538);
and U1978 (N_1978,N_156,N_90);
and U1979 (N_1979,N_499,N_846);
and U1980 (N_1980,N_606,N_750);
nand U1981 (N_1981,N_387,N_302);
nand U1982 (N_1982,N_726,N_699);
or U1983 (N_1983,N_956,N_8);
or U1984 (N_1984,N_926,N_265);
xor U1985 (N_1985,N_360,N_279);
or U1986 (N_1986,N_126,N_638);
nand U1987 (N_1987,N_480,N_575);
or U1988 (N_1988,N_266,N_30);
nor U1989 (N_1989,N_388,N_698);
or U1990 (N_1990,N_243,N_230);
nand U1991 (N_1991,N_429,N_65);
and U1992 (N_1992,N_908,N_861);
and U1993 (N_1993,N_512,N_415);
nor U1994 (N_1994,N_65,N_388);
nand U1995 (N_1995,N_909,N_16);
xor U1996 (N_1996,N_431,N_702);
and U1997 (N_1997,N_907,N_723);
nand U1998 (N_1998,N_390,N_254);
and U1999 (N_1999,N_649,N_635);
and U2000 (N_2000,N_1709,N_1602);
xnor U2001 (N_2001,N_1201,N_1881);
and U2002 (N_2002,N_1642,N_1540);
or U2003 (N_2003,N_1756,N_1838);
and U2004 (N_2004,N_1697,N_1781);
nor U2005 (N_2005,N_1200,N_1524);
xor U2006 (N_2006,N_1089,N_1630);
and U2007 (N_2007,N_1773,N_1960);
nand U2008 (N_2008,N_1387,N_1302);
or U2009 (N_2009,N_1030,N_1862);
nand U2010 (N_2010,N_1261,N_1520);
nor U2011 (N_2011,N_1803,N_1438);
or U2012 (N_2012,N_1156,N_1922);
nand U2013 (N_2013,N_1472,N_1945);
nor U2014 (N_2014,N_1561,N_1804);
and U2015 (N_2015,N_1651,N_1508);
and U2016 (N_2016,N_1372,N_1071);
xnor U2017 (N_2017,N_1955,N_1616);
xor U2018 (N_2018,N_1331,N_1677);
xnor U2019 (N_2019,N_1327,N_1815);
and U2020 (N_2020,N_1622,N_1356);
or U2021 (N_2021,N_1348,N_1659);
nand U2022 (N_2022,N_1653,N_1464);
nor U2023 (N_2023,N_1539,N_1150);
nand U2024 (N_2024,N_1696,N_1909);
nor U2025 (N_2025,N_1538,N_1517);
nor U2026 (N_2026,N_1559,N_1031);
nand U2027 (N_2027,N_1205,N_1418);
nor U2028 (N_2028,N_1995,N_1388);
or U2029 (N_2029,N_1063,N_1411);
and U2030 (N_2030,N_1637,N_1913);
nand U2031 (N_2031,N_1688,N_1161);
nand U2032 (N_2032,N_1082,N_1184);
or U2033 (N_2033,N_1260,N_1301);
and U2034 (N_2034,N_1239,N_1413);
nand U2035 (N_2035,N_1127,N_1450);
or U2036 (N_2036,N_1212,N_1046);
and U2037 (N_2037,N_1243,N_1820);
and U2038 (N_2038,N_1056,N_1436);
or U2039 (N_2039,N_1510,N_1810);
nand U2040 (N_2040,N_1178,N_1818);
and U2041 (N_2041,N_1976,N_1505);
or U2042 (N_2042,N_1021,N_1812);
nand U2043 (N_2043,N_1307,N_1858);
nor U2044 (N_2044,N_1042,N_1888);
nand U2045 (N_2045,N_1249,N_1589);
nor U2046 (N_2046,N_1774,N_1091);
and U2047 (N_2047,N_1816,N_1430);
and U2048 (N_2048,N_1577,N_1417);
nand U2049 (N_2049,N_1065,N_1710);
nand U2050 (N_2050,N_1720,N_1667);
and U2051 (N_2051,N_1138,N_1078);
nand U2052 (N_2052,N_1730,N_1608);
and U2053 (N_2053,N_1236,N_1408);
and U2054 (N_2054,N_1185,N_1219);
or U2055 (N_2055,N_1886,N_1823);
nand U2056 (N_2056,N_1546,N_1959);
nor U2057 (N_2057,N_1530,N_1344);
nand U2058 (N_2058,N_1754,N_1347);
and U2059 (N_2059,N_1639,N_1587);
or U2060 (N_2060,N_1900,N_1597);
and U2061 (N_2061,N_1176,N_1225);
or U2062 (N_2062,N_1140,N_1682);
or U2063 (N_2063,N_1401,N_1994);
nor U2064 (N_2064,N_1376,N_1547);
xor U2065 (N_2065,N_1453,N_1181);
nor U2066 (N_2066,N_1088,N_1163);
nand U2067 (N_2067,N_1332,N_1375);
nand U2068 (N_2068,N_1476,N_1005);
nor U2069 (N_2069,N_1317,N_1188);
nor U2070 (N_2070,N_1255,N_1654);
nand U2071 (N_2071,N_1809,N_1992);
nor U2072 (N_2072,N_1873,N_1040);
and U2073 (N_2073,N_1121,N_1641);
and U2074 (N_2074,N_1565,N_1813);
xnor U2075 (N_2075,N_1570,N_1165);
or U2076 (N_2076,N_1445,N_1320);
or U2077 (N_2077,N_1323,N_1226);
and U2078 (N_2078,N_1549,N_1170);
or U2079 (N_2079,N_1883,N_1407);
or U2080 (N_2080,N_1433,N_1652);
and U2081 (N_2081,N_1805,N_1284);
or U2082 (N_2082,N_1930,N_1942);
nor U2083 (N_2083,N_1488,N_1670);
nor U2084 (N_2084,N_1234,N_1341);
nor U2085 (N_2085,N_1786,N_1834);
nand U2086 (N_2086,N_1275,N_1590);
or U2087 (N_2087,N_1131,N_1772);
xnor U2088 (N_2088,N_1802,N_1534);
nor U2089 (N_2089,N_1403,N_1033);
and U2090 (N_2090,N_1048,N_1601);
nand U2091 (N_2091,N_1175,N_1265);
nand U2092 (N_2092,N_1563,N_1721);
xor U2093 (N_2093,N_1429,N_1342);
nand U2094 (N_2094,N_1791,N_1489);
and U2095 (N_2095,N_1471,N_1735);
nor U2096 (N_2096,N_1680,N_1704);
nor U2097 (N_2097,N_1075,N_1258);
nor U2098 (N_2098,N_1951,N_1545);
nand U2099 (N_2099,N_1984,N_1643);
nand U2100 (N_2100,N_1358,N_1001);
xor U2101 (N_2101,N_1998,N_1645);
nor U2102 (N_2102,N_1070,N_1668);
or U2103 (N_2103,N_1167,N_1211);
and U2104 (N_2104,N_1953,N_1828);
or U2105 (N_2105,N_1830,N_1058);
and U2106 (N_2106,N_1292,N_1421);
or U2107 (N_2107,N_1354,N_1442);
xor U2108 (N_2108,N_1890,N_1957);
or U2109 (N_2109,N_1855,N_1365);
nor U2110 (N_2110,N_1829,N_1297);
nor U2111 (N_2111,N_1064,N_1541);
or U2112 (N_2112,N_1963,N_1085);
nand U2113 (N_2113,N_1194,N_1183);
nand U2114 (N_2114,N_1568,N_1468);
nor U2115 (N_2115,N_1198,N_1775);
nor U2116 (N_2116,N_1555,N_1002);
xor U2117 (N_2117,N_1398,N_1853);
or U2118 (N_2118,N_1092,N_1726);
or U2119 (N_2119,N_1947,N_1764);
nor U2120 (N_2120,N_1594,N_1192);
nor U2121 (N_2121,N_1766,N_1700);
nor U2122 (N_2122,N_1961,N_1072);
nor U2123 (N_2123,N_1705,N_1123);
nand U2124 (N_2124,N_1459,N_1842);
nand U2125 (N_2125,N_1940,N_1245);
nor U2126 (N_2126,N_1363,N_1920);
and U2127 (N_2127,N_1385,N_1152);
or U2128 (N_2128,N_1511,N_1314);
and U2129 (N_2129,N_1738,N_1397);
or U2130 (N_2130,N_1485,N_1729);
nor U2131 (N_2131,N_1043,N_1330);
or U2132 (N_2132,N_1887,N_1015);
nand U2133 (N_2133,N_1558,N_1349);
nor U2134 (N_2134,N_1507,N_1045);
nand U2135 (N_2135,N_1980,N_1733);
and U2136 (N_2136,N_1270,N_1311);
nor U2137 (N_2137,N_1598,N_1025);
or U2138 (N_2138,N_1262,N_1898);
and U2139 (N_2139,N_1708,N_1061);
nor U2140 (N_2140,N_1609,N_1119);
nand U2141 (N_2141,N_1083,N_1811);
xor U2142 (N_2142,N_1990,N_1964);
nand U2143 (N_2143,N_1400,N_1991);
nand U2144 (N_2144,N_1744,N_1932);
nor U2145 (N_2145,N_1346,N_1849);
nor U2146 (N_2146,N_1190,N_1142);
or U2147 (N_2147,N_1007,N_1195);
nor U2148 (N_2148,N_1610,N_1108);
or U2149 (N_2149,N_1415,N_1474);
nor U2150 (N_2150,N_1217,N_1747);
and U2151 (N_2151,N_1079,N_1921);
nor U2152 (N_2152,N_1215,N_1516);
nor U2153 (N_2153,N_1066,N_1615);
xnor U2154 (N_2154,N_1867,N_1454);
nand U2155 (N_2155,N_1084,N_1286);
nand U2156 (N_2156,N_1595,N_1420);
or U2157 (N_2157,N_1869,N_1483);
nor U2158 (N_2158,N_1655,N_1985);
nand U2159 (N_2159,N_1305,N_1714);
nor U2160 (N_2160,N_1288,N_1294);
xnor U2161 (N_2161,N_1521,N_1322);
and U2162 (N_2162,N_1694,N_1216);
and U2163 (N_2163,N_1634,N_1593);
or U2164 (N_2164,N_1209,N_1392);
and U2165 (N_2165,N_1529,N_1582);
or U2166 (N_2166,N_1177,N_1795);
nor U2167 (N_2167,N_1599,N_1160);
and U2168 (N_2168,N_1479,N_1782);
nand U2169 (N_2169,N_1281,N_1456);
nand U2170 (N_2170,N_1298,N_1711);
nor U2171 (N_2171,N_1220,N_1164);
xnor U2172 (N_2172,N_1067,N_1449);
and U2173 (N_2173,N_1780,N_1278);
or U2174 (N_2174,N_1441,N_1443);
or U2175 (N_2175,N_1807,N_1856);
and U2176 (N_2176,N_1826,N_1621);
and U2177 (N_2177,N_1154,N_1968);
xnor U2178 (N_2178,N_1444,N_1470);
and U2179 (N_2179,N_1204,N_1303);
nor U2180 (N_2180,N_1076,N_1857);
xor U2181 (N_2181,N_1939,N_1394);
nand U2182 (N_2182,N_1293,N_1871);
xor U2183 (N_2183,N_1918,N_1573);
nand U2184 (N_2184,N_1843,N_1877);
xor U2185 (N_2185,N_1618,N_1875);
nor U2186 (N_2186,N_1971,N_1414);
nand U2187 (N_2187,N_1748,N_1325);
nor U2188 (N_2188,N_1081,N_1876);
xor U2189 (N_2189,N_1916,N_1784);
or U2190 (N_2190,N_1997,N_1724);
nor U2191 (N_2191,N_1681,N_1351);
nor U2192 (N_2192,N_1901,N_1907);
or U2193 (N_2193,N_1227,N_1073);
xor U2194 (N_2194,N_1647,N_1231);
and U2195 (N_2195,N_1552,N_1528);
xnor U2196 (N_2196,N_1941,N_1895);
nand U2197 (N_2197,N_1580,N_1241);
nor U2198 (N_2198,N_1310,N_1989);
and U2199 (N_2199,N_1824,N_1448);
and U2200 (N_2200,N_1787,N_1999);
nor U2201 (N_2201,N_1113,N_1461);
nand U2202 (N_2202,N_1676,N_1844);
nand U2203 (N_2203,N_1504,N_1519);
and U2204 (N_2204,N_1244,N_1228);
and U2205 (N_2205,N_1465,N_1208);
nor U2206 (N_2206,N_1586,N_1410);
nor U2207 (N_2207,N_1831,N_1972);
or U2208 (N_2208,N_1290,N_1369);
or U2209 (N_2209,N_1583,N_1371);
nand U2210 (N_2210,N_1825,N_1133);
nand U2211 (N_2211,N_1703,N_1050);
or U2212 (N_2212,N_1143,N_1657);
and U2213 (N_2213,N_1962,N_1207);
nor U2214 (N_2214,N_1362,N_1739);
nor U2215 (N_2215,N_1350,N_1671);
nand U2216 (N_2216,N_1817,N_1731);
or U2217 (N_2217,N_1762,N_1835);
nand U2218 (N_2218,N_1276,N_1891);
nand U2219 (N_2219,N_1462,N_1906);
nor U2220 (N_2220,N_1296,N_1093);
nor U2221 (N_2221,N_1291,N_1402);
nor U2222 (N_2222,N_1147,N_1256);
or U2223 (N_2223,N_1306,N_1144);
nor U2224 (N_2224,N_1861,N_1359);
nor U2225 (N_2225,N_1117,N_1024);
or U2226 (N_2226,N_1148,N_1525);
nand U2227 (N_2227,N_1832,N_1193);
nor U2228 (N_2228,N_1683,N_1800);
xnor U2229 (N_2229,N_1702,N_1218);
nand U2230 (N_2230,N_1578,N_1460);
and U2231 (N_2231,N_1591,N_1224);
or U2232 (N_2232,N_1478,N_1658);
xnor U2233 (N_2233,N_1770,N_1435);
nor U2234 (N_2234,N_1467,N_1821);
xor U2235 (N_2235,N_1051,N_1706);
nor U2236 (N_2236,N_1788,N_1419);
and U2237 (N_2237,N_1522,N_1814);
nor U2238 (N_2238,N_1202,N_1316);
nand U2239 (N_2239,N_1159,N_1172);
nor U2240 (N_2240,N_1189,N_1874);
and U2241 (N_2241,N_1503,N_1870);
or U2242 (N_2242,N_1425,N_1656);
and U2243 (N_2243,N_1675,N_1125);
nand U2244 (N_2244,N_1099,N_1743);
nand U2245 (N_2245,N_1685,N_1789);
and U2246 (N_2246,N_1380,N_1267);
or U2247 (N_2247,N_1017,N_1364);
nor U2248 (N_2248,N_1299,N_1513);
and U2249 (N_2249,N_1384,N_1182);
xnor U2250 (N_2250,N_1315,N_1692);
nor U2251 (N_2251,N_1734,N_1259);
xnor U2252 (N_2252,N_1978,N_1531);
or U2253 (N_2253,N_1560,N_1396);
nand U2254 (N_2254,N_1864,N_1406);
or U2255 (N_2255,N_1661,N_1649);
nor U2256 (N_2256,N_1247,N_1034);
or U2257 (N_2257,N_1571,N_1389);
nor U2258 (N_2258,N_1378,N_1339);
nand U2259 (N_2259,N_1946,N_1012);
or U2260 (N_2260,N_1624,N_1248);
nor U2261 (N_2261,N_1983,N_1210);
nor U2262 (N_2262,N_1492,N_1695);
nand U2263 (N_2263,N_1626,N_1785);
nand U2264 (N_2264,N_1028,N_1037);
nand U2265 (N_2265,N_1309,N_1105);
nor U2266 (N_2266,N_1986,N_1699);
nor U2267 (N_2267,N_1579,N_1722);
xnor U2268 (N_2268,N_1086,N_1679);
or U2269 (N_2269,N_1010,N_1761);
nor U2270 (N_2270,N_1822,N_1221);
or U2271 (N_2271,N_1892,N_1979);
nand U2272 (N_2272,N_1155,N_1575);
and U2273 (N_2273,N_1011,N_1282);
nor U2274 (N_2274,N_1678,N_1557);
and U2275 (N_2275,N_1130,N_1952);
nand U2276 (N_2276,N_1057,N_1324);
nor U2277 (N_2277,N_1493,N_1405);
nor U2278 (N_2278,N_1638,N_1126);
or U2279 (N_2279,N_1426,N_1059);
nor U2280 (N_2280,N_1274,N_1080);
and U2281 (N_2281,N_1340,N_1242);
nand U2282 (N_2282,N_1736,N_1118);
nor U2283 (N_2283,N_1484,N_1854);
nor U2284 (N_2284,N_1318,N_1285);
or U2285 (N_2285,N_1924,N_1923);
or U2286 (N_2286,N_1689,N_1171);
or U2287 (N_2287,N_1687,N_1473);
or U2288 (N_2288,N_1926,N_1797);
nor U2289 (N_2289,N_1796,N_1166);
xnor U2290 (N_2290,N_1783,N_1567);
xnor U2291 (N_2291,N_1455,N_1588);
nand U2292 (N_2292,N_1847,N_1232);
nor U2293 (N_2293,N_1878,N_1701);
nand U2294 (N_2294,N_1122,N_1840);
or U2295 (N_2295,N_1937,N_1269);
nor U2296 (N_2296,N_1973,N_1191);
and U2297 (N_2297,N_1745,N_1771);
or U2298 (N_2298,N_1872,N_1600);
nand U2299 (N_2299,N_1728,N_1049);
nand U2300 (N_2300,N_1345,N_1304);
and U2301 (N_2301,N_1422,N_1068);
nand U2302 (N_2302,N_1753,N_1819);
nand U2303 (N_2303,N_1103,N_1612);
and U2304 (N_2304,N_1112,N_1313);
xnor U2305 (N_2305,N_1446,N_1663);
and U2306 (N_2306,N_1662,N_1929);
nand U2307 (N_2307,N_1954,N_1798);
nand U2308 (N_2308,N_1903,N_1533);
xnor U2309 (N_2309,N_1319,N_1115);
and U2310 (N_2310,N_1135,N_1712);
or U2311 (N_2311,N_1919,N_1749);
or U2312 (N_2312,N_1253,N_1790);
xnor U2313 (N_2313,N_1069,N_1273);
nand U2314 (N_2314,N_1370,N_1335);
nand U2315 (N_2315,N_1605,N_1146);
or U2316 (N_2316,N_1447,N_1416);
and U2317 (N_2317,N_1312,N_1087);
or U2318 (N_2318,N_1882,N_1969);
or U2319 (N_2319,N_1614,N_1725);
nor U2320 (N_2320,N_1910,N_1022);
xnor U2321 (N_2321,N_1427,N_1128);
nand U2322 (N_2322,N_1633,N_1434);
nor U2323 (N_2323,N_1627,N_1606);
or U2324 (N_2324,N_1684,N_1965);
and U2325 (N_2325,N_1038,N_1514);
nand U2326 (N_2326,N_1632,N_1987);
and U2327 (N_2327,N_1287,N_1026);
nand U2328 (N_2328,N_1020,N_1196);
or U2329 (N_2329,N_1382,N_1719);
or U2330 (N_2330,N_1768,N_1333);
nor U2331 (N_2331,N_1077,N_1613);
and U2332 (N_2332,N_1263,N_1357);
nor U2333 (N_2333,N_1611,N_1343);
nand U2334 (N_2334,N_1399,N_1004);
xor U2335 (N_2335,N_1238,N_1686);
nor U2336 (N_2336,N_1794,N_1581);
and U2337 (N_2337,N_1707,N_1257);
nand U2338 (N_2338,N_1691,N_1767);
nand U2339 (N_2339,N_1868,N_1074);
or U2340 (N_2340,N_1102,N_1596);
and U2341 (N_2341,N_1062,N_1793);
nor U2342 (N_2342,N_1029,N_1635);
and U2343 (N_2343,N_1090,N_1237);
or U2344 (N_2344,N_1837,N_1741);
nor U2345 (N_2345,N_1569,N_1377);
nor U2346 (N_2346,N_1035,N_1660);
nor U2347 (N_2347,N_1114,N_1168);
or U2348 (N_2348,N_1373,N_1173);
nor U2349 (N_2349,N_1566,N_1254);
xor U2350 (N_2350,N_1203,N_1629);
and U2351 (N_2351,N_1698,N_1604);
nand U2352 (N_2352,N_1329,N_1475);
nor U2353 (N_2353,N_1151,N_1268);
and U2354 (N_2354,N_1763,N_1617);
nor U2355 (N_2355,N_1851,N_1506);
nor U2356 (N_2356,N_1355,N_1027);
nor U2357 (N_2357,N_1925,N_1423);
xor U2358 (N_2358,N_1585,N_1230);
nor U2359 (N_2359,N_1915,N_1880);
and U2360 (N_2360,N_1912,N_1153);
nand U2361 (N_2361,N_1672,N_1481);
nor U2362 (N_2362,N_1496,N_1993);
nor U2363 (N_2363,N_1098,N_1482);
and U2364 (N_2364,N_1897,N_1554);
nand U2365 (N_2365,N_1097,N_1272);
or U2366 (N_2366,N_1179,N_1096);
nor U2367 (N_2367,N_1866,N_1246);
nor U2368 (N_2368,N_1381,N_1233);
nor U2369 (N_2369,N_1466,N_1336);
nand U2370 (N_2370,N_1116,N_1859);
or U2371 (N_2371,N_1542,N_1640);
nand U2372 (N_2372,N_1041,N_1948);
nand U2373 (N_2373,N_1905,N_1337);
xnor U2374 (N_2374,N_1666,N_1379);
nand U2375 (N_2375,N_1499,N_1956);
nor U2376 (N_2376,N_1222,N_1206);
nor U2377 (N_2377,N_1603,N_1141);
or U2378 (N_2378,N_1509,N_1740);
nor U2379 (N_2379,N_1512,N_1145);
and U2380 (N_2380,N_1526,N_1223);
or U2381 (N_2381,N_1395,N_1548);
xor U2382 (N_2382,N_1412,N_1523);
or U2383 (N_2383,N_1949,N_1032);
and U2384 (N_2384,N_1494,N_1852);
or U2385 (N_2385,N_1039,N_1009);
nor U2386 (N_2386,N_1631,N_1564);
nand U2387 (N_2387,N_1052,N_1180);
nand U2388 (N_2388,N_1518,N_1006);
or U2389 (N_2389,N_1760,N_1982);
nor U2390 (N_2390,N_1537,N_1690);
nand U2391 (N_2391,N_1746,N_1352);
or U2392 (N_2392,N_1132,N_1742);
or U2393 (N_2393,N_1250,N_1644);
nor U2394 (N_2394,N_1139,N_1836);
or U2395 (N_2395,N_1428,N_1996);
or U2396 (N_2396,N_1648,N_1646);
xor U2397 (N_2397,N_1879,N_1197);
nor U2398 (N_2398,N_1752,N_1487);
and U2399 (N_2399,N_1409,N_1715);
nand U2400 (N_2400,N_1008,N_1016);
nor U2401 (N_2401,N_1899,N_1556);
nand U2402 (N_2402,N_1502,N_1765);
and U2403 (N_2403,N_1491,N_1755);
nor U2404 (N_2404,N_1252,N_1893);
nor U2405 (N_2405,N_1884,N_1391);
or U2406 (N_2406,N_1914,N_1107);
nor U2407 (N_2407,N_1584,N_1535);
nor U2408 (N_2408,N_1498,N_1936);
nor U2409 (N_2409,N_1833,N_1623);
xor U2410 (N_2410,N_1500,N_1917);
and U2411 (N_2411,N_1367,N_1023);
and U2412 (N_2412,N_1366,N_1863);
nor U2413 (N_2413,N_1944,N_1393);
nand U2414 (N_2414,N_1106,N_1055);
or U2415 (N_2415,N_1328,N_1865);
or U2416 (N_2416,N_1778,N_1360);
or U2417 (N_2417,N_1266,N_1149);
and U2418 (N_2418,N_1095,N_1186);
nor U2419 (N_2419,N_1137,N_1124);
and U2420 (N_2420,N_1003,N_1777);
and U2421 (N_2421,N_1750,N_1636);
or U2422 (N_2422,N_1437,N_1845);
xnor U2423 (N_2423,N_1120,N_1967);
nor U2424 (N_2424,N_1162,N_1334);
and U2425 (N_2425,N_1495,N_1271);
or U2426 (N_2426,N_1943,N_1440);
nor U2427 (N_2427,N_1673,N_1723);
nand U2428 (N_2428,N_1850,N_1693);
nand U2429 (N_2429,N_1279,N_1169);
or U2430 (N_2430,N_1501,N_1966);
or U2431 (N_2431,N_1839,N_1716);
or U2432 (N_2432,N_1187,N_1806);
and U2433 (N_2433,N_1758,N_1572);
and U2434 (N_2434,N_1550,N_1368);
and U2435 (N_2435,N_1574,N_1497);
xor U2436 (N_2436,N_1737,N_1933);
and U2437 (N_2437,N_1620,N_1353);
or U2438 (N_2438,N_1213,N_1515);
nand U2439 (N_2439,N_1439,N_1158);
nor U2440 (N_2440,N_1235,N_1477);
and U2441 (N_2441,N_1251,N_1060);
nor U2442 (N_2442,N_1326,N_1894);
xnor U2443 (N_2443,N_1101,N_1283);
and U2444 (N_2444,N_1136,N_1717);
and U2445 (N_2445,N_1988,N_1665);
nand U2446 (N_2446,N_1543,N_1669);
nor U2447 (N_2447,N_1551,N_1848);
and U2448 (N_2448,N_1532,N_1129);
and U2449 (N_2449,N_1214,N_1769);
and U2450 (N_2450,N_1846,N_1607);
nand U2451 (N_2451,N_1361,N_1240);
nor U2452 (N_2452,N_1970,N_1280);
nand U2453 (N_2453,N_1732,N_1902);
nand U2454 (N_2454,N_1451,N_1432);
or U2455 (N_2455,N_1779,N_1490);
and U2456 (N_2456,N_1792,N_1553);
or U2457 (N_2457,N_1801,N_1458);
nand U2458 (N_2458,N_1431,N_1808);
nor U2459 (N_2459,N_1592,N_1759);
or U2460 (N_2460,N_1981,N_1860);
nand U2461 (N_2461,N_1338,N_1841);
nand U2462 (N_2462,N_1727,N_1457);
xnor U2463 (N_2463,N_1958,N_1134);
and U2464 (N_2464,N_1014,N_1664);
and U2465 (N_2465,N_1308,N_1019);
and U2466 (N_2466,N_1718,N_1013);
nand U2467 (N_2467,N_1018,N_1576);
and U2468 (N_2468,N_1928,N_1713);
nor U2469 (N_2469,N_1480,N_1452);
and U2470 (N_2470,N_1469,N_1628);
or U2471 (N_2471,N_1264,N_1625);
nor U2472 (N_2472,N_1751,N_1295);
or U2473 (N_2473,N_1289,N_1927);
nor U2474 (N_2474,N_1404,N_1300);
and U2475 (N_2475,N_1321,N_1827);
and U2476 (N_2476,N_1109,N_1911);
and U2477 (N_2477,N_1938,N_1094);
nor U2478 (N_2478,N_1463,N_1757);
and U2479 (N_2479,N_1053,N_1904);
and U2480 (N_2480,N_1044,N_1889);
xor U2481 (N_2481,N_1386,N_1054);
nor U2482 (N_2482,N_1157,N_1527);
nand U2483 (N_2483,N_1374,N_1934);
nand U2484 (N_2484,N_1619,N_1674);
and U2485 (N_2485,N_1383,N_1174);
nor U2486 (N_2486,N_1000,N_1199);
nand U2487 (N_2487,N_1424,N_1536);
and U2488 (N_2488,N_1885,N_1100);
nor U2489 (N_2489,N_1776,N_1935);
nand U2490 (N_2490,N_1110,N_1229);
nand U2491 (N_2491,N_1977,N_1799);
and U2492 (N_2492,N_1277,N_1896);
nor U2493 (N_2493,N_1908,N_1974);
and U2494 (N_2494,N_1650,N_1486);
and U2495 (N_2495,N_1036,N_1931);
xnor U2496 (N_2496,N_1111,N_1975);
xor U2497 (N_2497,N_1544,N_1104);
nor U2498 (N_2498,N_1950,N_1047);
and U2499 (N_2499,N_1562,N_1390);
nand U2500 (N_2500,N_1581,N_1503);
nor U2501 (N_2501,N_1317,N_1601);
or U2502 (N_2502,N_1384,N_1410);
or U2503 (N_2503,N_1670,N_1900);
nand U2504 (N_2504,N_1406,N_1018);
nor U2505 (N_2505,N_1537,N_1891);
and U2506 (N_2506,N_1358,N_1536);
nor U2507 (N_2507,N_1739,N_1724);
nor U2508 (N_2508,N_1006,N_1054);
and U2509 (N_2509,N_1478,N_1227);
nand U2510 (N_2510,N_1449,N_1789);
or U2511 (N_2511,N_1352,N_1065);
or U2512 (N_2512,N_1422,N_1187);
nand U2513 (N_2513,N_1679,N_1507);
or U2514 (N_2514,N_1857,N_1363);
nand U2515 (N_2515,N_1612,N_1016);
nand U2516 (N_2516,N_1018,N_1205);
nor U2517 (N_2517,N_1359,N_1833);
nand U2518 (N_2518,N_1771,N_1165);
nand U2519 (N_2519,N_1781,N_1326);
nand U2520 (N_2520,N_1383,N_1741);
and U2521 (N_2521,N_1060,N_1353);
nand U2522 (N_2522,N_1086,N_1091);
xnor U2523 (N_2523,N_1109,N_1576);
and U2524 (N_2524,N_1641,N_1337);
nand U2525 (N_2525,N_1689,N_1373);
nand U2526 (N_2526,N_1094,N_1536);
nor U2527 (N_2527,N_1965,N_1358);
or U2528 (N_2528,N_1256,N_1776);
and U2529 (N_2529,N_1660,N_1367);
nor U2530 (N_2530,N_1218,N_1642);
and U2531 (N_2531,N_1301,N_1691);
and U2532 (N_2532,N_1822,N_1485);
and U2533 (N_2533,N_1085,N_1486);
nor U2534 (N_2534,N_1800,N_1838);
or U2535 (N_2535,N_1630,N_1433);
nor U2536 (N_2536,N_1014,N_1096);
xor U2537 (N_2537,N_1055,N_1379);
xor U2538 (N_2538,N_1271,N_1022);
xnor U2539 (N_2539,N_1710,N_1412);
nand U2540 (N_2540,N_1106,N_1874);
nand U2541 (N_2541,N_1365,N_1084);
nor U2542 (N_2542,N_1826,N_1210);
nor U2543 (N_2543,N_1031,N_1014);
nor U2544 (N_2544,N_1831,N_1856);
and U2545 (N_2545,N_1869,N_1400);
or U2546 (N_2546,N_1312,N_1364);
and U2547 (N_2547,N_1914,N_1962);
or U2548 (N_2548,N_1929,N_1315);
nand U2549 (N_2549,N_1786,N_1636);
and U2550 (N_2550,N_1686,N_1048);
and U2551 (N_2551,N_1176,N_1320);
nand U2552 (N_2552,N_1990,N_1781);
or U2553 (N_2553,N_1031,N_1896);
or U2554 (N_2554,N_1640,N_1399);
and U2555 (N_2555,N_1523,N_1920);
or U2556 (N_2556,N_1469,N_1168);
and U2557 (N_2557,N_1020,N_1823);
nand U2558 (N_2558,N_1505,N_1763);
nand U2559 (N_2559,N_1646,N_1600);
nand U2560 (N_2560,N_1753,N_1951);
nor U2561 (N_2561,N_1832,N_1944);
nand U2562 (N_2562,N_1272,N_1072);
xnor U2563 (N_2563,N_1141,N_1242);
and U2564 (N_2564,N_1048,N_1813);
xnor U2565 (N_2565,N_1956,N_1172);
nand U2566 (N_2566,N_1856,N_1405);
nor U2567 (N_2567,N_1517,N_1970);
or U2568 (N_2568,N_1631,N_1497);
and U2569 (N_2569,N_1611,N_1843);
and U2570 (N_2570,N_1040,N_1091);
or U2571 (N_2571,N_1852,N_1931);
and U2572 (N_2572,N_1468,N_1251);
nand U2573 (N_2573,N_1506,N_1086);
or U2574 (N_2574,N_1525,N_1612);
and U2575 (N_2575,N_1147,N_1819);
nand U2576 (N_2576,N_1024,N_1387);
and U2577 (N_2577,N_1360,N_1720);
xnor U2578 (N_2578,N_1817,N_1269);
xor U2579 (N_2579,N_1552,N_1495);
and U2580 (N_2580,N_1974,N_1936);
and U2581 (N_2581,N_1977,N_1789);
and U2582 (N_2582,N_1390,N_1581);
nor U2583 (N_2583,N_1743,N_1594);
or U2584 (N_2584,N_1605,N_1362);
and U2585 (N_2585,N_1792,N_1747);
nor U2586 (N_2586,N_1204,N_1758);
and U2587 (N_2587,N_1126,N_1234);
nand U2588 (N_2588,N_1683,N_1184);
or U2589 (N_2589,N_1011,N_1934);
and U2590 (N_2590,N_1369,N_1372);
and U2591 (N_2591,N_1275,N_1070);
or U2592 (N_2592,N_1135,N_1531);
xnor U2593 (N_2593,N_1095,N_1098);
nand U2594 (N_2594,N_1257,N_1664);
nand U2595 (N_2595,N_1669,N_1131);
nand U2596 (N_2596,N_1373,N_1569);
xor U2597 (N_2597,N_1027,N_1889);
and U2598 (N_2598,N_1179,N_1243);
nor U2599 (N_2599,N_1229,N_1038);
and U2600 (N_2600,N_1347,N_1594);
or U2601 (N_2601,N_1509,N_1823);
and U2602 (N_2602,N_1034,N_1099);
nand U2603 (N_2603,N_1064,N_1900);
xnor U2604 (N_2604,N_1498,N_1295);
nand U2605 (N_2605,N_1070,N_1170);
nor U2606 (N_2606,N_1985,N_1690);
nand U2607 (N_2607,N_1793,N_1950);
nand U2608 (N_2608,N_1557,N_1146);
xor U2609 (N_2609,N_1660,N_1610);
or U2610 (N_2610,N_1897,N_1491);
nand U2611 (N_2611,N_1191,N_1368);
nand U2612 (N_2612,N_1608,N_1361);
or U2613 (N_2613,N_1264,N_1803);
nor U2614 (N_2614,N_1912,N_1815);
nor U2615 (N_2615,N_1755,N_1686);
and U2616 (N_2616,N_1737,N_1393);
nor U2617 (N_2617,N_1058,N_1418);
nor U2618 (N_2618,N_1506,N_1491);
nand U2619 (N_2619,N_1264,N_1727);
nand U2620 (N_2620,N_1969,N_1954);
or U2621 (N_2621,N_1916,N_1141);
and U2622 (N_2622,N_1980,N_1299);
nand U2623 (N_2623,N_1494,N_1027);
and U2624 (N_2624,N_1807,N_1157);
xor U2625 (N_2625,N_1416,N_1953);
or U2626 (N_2626,N_1620,N_1983);
xor U2627 (N_2627,N_1030,N_1829);
and U2628 (N_2628,N_1786,N_1957);
xnor U2629 (N_2629,N_1224,N_1057);
nand U2630 (N_2630,N_1655,N_1331);
nor U2631 (N_2631,N_1512,N_1558);
xnor U2632 (N_2632,N_1704,N_1993);
nand U2633 (N_2633,N_1185,N_1695);
or U2634 (N_2634,N_1768,N_1661);
or U2635 (N_2635,N_1959,N_1095);
or U2636 (N_2636,N_1697,N_1883);
and U2637 (N_2637,N_1110,N_1825);
nand U2638 (N_2638,N_1929,N_1097);
nor U2639 (N_2639,N_1371,N_1671);
and U2640 (N_2640,N_1590,N_1983);
and U2641 (N_2641,N_1297,N_1637);
and U2642 (N_2642,N_1997,N_1440);
and U2643 (N_2643,N_1902,N_1296);
xnor U2644 (N_2644,N_1052,N_1403);
and U2645 (N_2645,N_1282,N_1627);
or U2646 (N_2646,N_1638,N_1144);
nand U2647 (N_2647,N_1094,N_1479);
or U2648 (N_2648,N_1467,N_1518);
and U2649 (N_2649,N_1520,N_1558);
xnor U2650 (N_2650,N_1396,N_1685);
and U2651 (N_2651,N_1172,N_1495);
nand U2652 (N_2652,N_1497,N_1173);
or U2653 (N_2653,N_1840,N_1973);
xor U2654 (N_2654,N_1390,N_1858);
nand U2655 (N_2655,N_1905,N_1351);
or U2656 (N_2656,N_1389,N_1601);
xnor U2657 (N_2657,N_1894,N_1058);
or U2658 (N_2658,N_1359,N_1559);
nor U2659 (N_2659,N_1475,N_1336);
nand U2660 (N_2660,N_1525,N_1702);
or U2661 (N_2661,N_1066,N_1459);
nand U2662 (N_2662,N_1878,N_1177);
nand U2663 (N_2663,N_1134,N_1199);
nand U2664 (N_2664,N_1114,N_1375);
nor U2665 (N_2665,N_1856,N_1814);
and U2666 (N_2666,N_1255,N_1991);
nor U2667 (N_2667,N_1812,N_1963);
nor U2668 (N_2668,N_1925,N_1143);
and U2669 (N_2669,N_1296,N_1818);
nor U2670 (N_2670,N_1010,N_1227);
or U2671 (N_2671,N_1322,N_1299);
nor U2672 (N_2672,N_1793,N_1156);
or U2673 (N_2673,N_1164,N_1163);
nor U2674 (N_2674,N_1642,N_1016);
and U2675 (N_2675,N_1300,N_1390);
xor U2676 (N_2676,N_1167,N_1674);
xor U2677 (N_2677,N_1066,N_1242);
or U2678 (N_2678,N_1268,N_1392);
nand U2679 (N_2679,N_1029,N_1078);
and U2680 (N_2680,N_1224,N_1041);
or U2681 (N_2681,N_1184,N_1132);
nor U2682 (N_2682,N_1191,N_1728);
nand U2683 (N_2683,N_1374,N_1599);
xor U2684 (N_2684,N_1780,N_1052);
nand U2685 (N_2685,N_1466,N_1923);
and U2686 (N_2686,N_1178,N_1500);
and U2687 (N_2687,N_1136,N_1164);
nand U2688 (N_2688,N_1770,N_1354);
and U2689 (N_2689,N_1742,N_1464);
and U2690 (N_2690,N_1110,N_1776);
or U2691 (N_2691,N_1912,N_1574);
nand U2692 (N_2692,N_1918,N_1405);
nand U2693 (N_2693,N_1847,N_1164);
and U2694 (N_2694,N_1158,N_1354);
nand U2695 (N_2695,N_1133,N_1707);
nand U2696 (N_2696,N_1724,N_1067);
nor U2697 (N_2697,N_1681,N_1285);
and U2698 (N_2698,N_1313,N_1653);
or U2699 (N_2699,N_1548,N_1116);
or U2700 (N_2700,N_1896,N_1085);
nor U2701 (N_2701,N_1975,N_1639);
nor U2702 (N_2702,N_1275,N_1581);
and U2703 (N_2703,N_1052,N_1111);
or U2704 (N_2704,N_1080,N_1038);
nor U2705 (N_2705,N_1159,N_1347);
nand U2706 (N_2706,N_1245,N_1115);
nand U2707 (N_2707,N_1414,N_1713);
xnor U2708 (N_2708,N_1122,N_1957);
or U2709 (N_2709,N_1436,N_1511);
nor U2710 (N_2710,N_1802,N_1418);
and U2711 (N_2711,N_1522,N_1793);
or U2712 (N_2712,N_1976,N_1904);
nand U2713 (N_2713,N_1049,N_1277);
or U2714 (N_2714,N_1926,N_1189);
nand U2715 (N_2715,N_1124,N_1959);
nand U2716 (N_2716,N_1350,N_1147);
nor U2717 (N_2717,N_1296,N_1479);
or U2718 (N_2718,N_1522,N_1820);
nand U2719 (N_2719,N_1875,N_1805);
or U2720 (N_2720,N_1033,N_1828);
nor U2721 (N_2721,N_1009,N_1562);
and U2722 (N_2722,N_1131,N_1039);
xor U2723 (N_2723,N_1064,N_1002);
or U2724 (N_2724,N_1374,N_1026);
nor U2725 (N_2725,N_1442,N_1771);
or U2726 (N_2726,N_1878,N_1601);
or U2727 (N_2727,N_1055,N_1844);
and U2728 (N_2728,N_1570,N_1244);
nor U2729 (N_2729,N_1276,N_1824);
and U2730 (N_2730,N_1695,N_1590);
nand U2731 (N_2731,N_1952,N_1509);
or U2732 (N_2732,N_1075,N_1132);
xor U2733 (N_2733,N_1137,N_1170);
and U2734 (N_2734,N_1282,N_1738);
and U2735 (N_2735,N_1953,N_1675);
or U2736 (N_2736,N_1017,N_1985);
nand U2737 (N_2737,N_1199,N_1303);
xor U2738 (N_2738,N_1855,N_1750);
and U2739 (N_2739,N_1051,N_1058);
or U2740 (N_2740,N_1675,N_1500);
or U2741 (N_2741,N_1748,N_1305);
or U2742 (N_2742,N_1852,N_1938);
or U2743 (N_2743,N_1044,N_1807);
or U2744 (N_2744,N_1704,N_1835);
or U2745 (N_2745,N_1617,N_1050);
and U2746 (N_2746,N_1657,N_1885);
nor U2747 (N_2747,N_1926,N_1476);
nand U2748 (N_2748,N_1484,N_1980);
xnor U2749 (N_2749,N_1027,N_1160);
nor U2750 (N_2750,N_1012,N_1692);
and U2751 (N_2751,N_1447,N_1538);
nand U2752 (N_2752,N_1231,N_1746);
and U2753 (N_2753,N_1770,N_1531);
or U2754 (N_2754,N_1928,N_1006);
or U2755 (N_2755,N_1165,N_1314);
and U2756 (N_2756,N_1247,N_1640);
or U2757 (N_2757,N_1384,N_1355);
and U2758 (N_2758,N_1024,N_1274);
or U2759 (N_2759,N_1744,N_1237);
nor U2760 (N_2760,N_1894,N_1142);
and U2761 (N_2761,N_1325,N_1730);
or U2762 (N_2762,N_1494,N_1909);
xnor U2763 (N_2763,N_1084,N_1199);
and U2764 (N_2764,N_1442,N_1163);
nand U2765 (N_2765,N_1888,N_1994);
or U2766 (N_2766,N_1707,N_1385);
nor U2767 (N_2767,N_1432,N_1043);
and U2768 (N_2768,N_1933,N_1464);
nand U2769 (N_2769,N_1054,N_1830);
xnor U2770 (N_2770,N_1989,N_1421);
and U2771 (N_2771,N_1040,N_1274);
nor U2772 (N_2772,N_1317,N_1491);
nand U2773 (N_2773,N_1949,N_1906);
or U2774 (N_2774,N_1128,N_1047);
nor U2775 (N_2775,N_1326,N_1818);
or U2776 (N_2776,N_1519,N_1497);
nor U2777 (N_2777,N_1255,N_1095);
nand U2778 (N_2778,N_1529,N_1192);
nand U2779 (N_2779,N_1229,N_1014);
xor U2780 (N_2780,N_1641,N_1640);
nor U2781 (N_2781,N_1795,N_1282);
and U2782 (N_2782,N_1323,N_1429);
or U2783 (N_2783,N_1546,N_1487);
and U2784 (N_2784,N_1326,N_1976);
nand U2785 (N_2785,N_1017,N_1916);
nand U2786 (N_2786,N_1452,N_1790);
nand U2787 (N_2787,N_1186,N_1112);
xor U2788 (N_2788,N_1640,N_1158);
xor U2789 (N_2789,N_1280,N_1871);
nor U2790 (N_2790,N_1167,N_1999);
or U2791 (N_2791,N_1347,N_1582);
nand U2792 (N_2792,N_1514,N_1998);
and U2793 (N_2793,N_1004,N_1060);
and U2794 (N_2794,N_1161,N_1963);
nand U2795 (N_2795,N_1751,N_1023);
or U2796 (N_2796,N_1237,N_1188);
nor U2797 (N_2797,N_1415,N_1014);
nand U2798 (N_2798,N_1215,N_1776);
nand U2799 (N_2799,N_1455,N_1096);
and U2800 (N_2800,N_1628,N_1263);
nor U2801 (N_2801,N_1018,N_1440);
and U2802 (N_2802,N_1393,N_1421);
xnor U2803 (N_2803,N_1474,N_1721);
xnor U2804 (N_2804,N_1704,N_1591);
or U2805 (N_2805,N_1209,N_1815);
nand U2806 (N_2806,N_1788,N_1768);
or U2807 (N_2807,N_1418,N_1600);
nor U2808 (N_2808,N_1333,N_1947);
nor U2809 (N_2809,N_1470,N_1564);
or U2810 (N_2810,N_1042,N_1572);
xor U2811 (N_2811,N_1127,N_1029);
nand U2812 (N_2812,N_1381,N_1185);
and U2813 (N_2813,N_1634,N_1254);
nand U2814 (N_2814,N_1691,N_1113);
nand U2815 (N_2815,N_1449,N_1675);
and U2816 (N_2816,N_1416,N_1204);
nor U2817 (N_2817,N_1550,N_1319);
nand U2818 (N_2818,N_1011,N_1671);
nor U2819 (N_2819,N_1660,N_1083);
or U2820 (N_2820,N_1323,N_1152);
xnor U2821 (N_2821,N_1234,N_1653);
and U2822 (N_2822,N_1154,N_1232);
nor U2823 (N_2823,N_1011,N_1336);
nor U2824 (N_2824,N_1624,N_1648);
xnor U2825 (N_2825,N_1201,N_1150);
and U2826 (N_2826,N_1884,N_1190);
and U2827 (N_2827,N_1520,N_1655);
or U2828 (N_2828,N_1995,N_1499);
xor U2829 (N_2829,N_1537,N_1832);
and U2830 (N_2830,N_1743,N_1242);
nor U2831 (N_2831,N_1467,N_1678);
or U2832 (N_2832,N_1135,N_1326);
nand U2833 (N_2833,N_1127,N_1268);
xnor U2834 (N_2834,N_1494,N_1953);
nor U2835 (N_2835,N_1088,N_1286);
nand U2836 (N_2836,N_1088,N_1707);
or U2837 (N_2837,N_1822,N_1562);
and U2838 (N_2838,N_1030,N_1050);
nor U2839 (N_2839,N_1816,N_1604);
xor U2840 (N_2840,N_1050,N_1405);
and U2841 (N_2841,N_1888,N_1169);
and U2842 (N_2842,N_1253,N_1819);
or U2843 (N_2843,N_1392,N_1798);
nand U2844 (N_2844,N_1155,N_1806);
nor U2845 (N_2845,N_1788,N_1461);
and U2846 (N_2846,N_1855,N_1761);
nor U2847 (N_2847,N_1475,N_1862);
and U2848 (N_2848,N_1271,N_1525);
xnor U2849 (N_2849,N_1984,N_1624);
or U2850 (N_2850,N_1632,N_1433);
and U2851 (N_2851,N_1388,N_1189);
or U2852 (N_2852,N_1619,N_1109);
nor U2853 (N_2853,N_1827,N_1715);
nand U2854 (N_2854,N_1142,N_1172);
nor U2855 (N_2855,N_1648,N_1898);
nor U2856 (N_2856,N_1986,N_1063);
and U2857 (N_2857,N_1111,N_1612);
and U2858 (N_2858,N_1360,N_1028);
nor U2859 (N_2859,N_1731,N_1552);
and U2860 (N_2860,N_1789,N_1627);
nor U2861 (N_2861,N_1451,N_1212);
or U2862 (N_2862,N_1983,N_1260);
nand U2863 (N_2863,N_1598,N_1286);
and U2864 (N_2864,N_1855,N_1655);
nor U2865 (N_2865,N_1447,N_1226);
nand U2866 (N_2866,N_1411,N_1326);
and U2867 (N_2867,N_1347,N_1607);
and U2868 (N_2868,N_1796,N_1553);
nor U2869 (N_2869,N_1603,N_1053);
nor U2870 (N_2870,N_1866,N_1398);
and U2871 (N_2871,N_1419,N_1225);
nand U2872 (N_2872,N_1188,N_1372);
or U2873 (N_2873,N_1492,N_1116);
and U2874 (N_2874,N_1054,N_1290);
or U2875 (N_2875,N_1183,N_1105);
xor U2876 (N_2876,N_1586,N_1541);
nor U2877 (N_2877,N_1039,N_1025);
xnor U2878 (N_2878,N_1188,N_1600);
and U2879 (N_2879,N_1528,N_1940);
and U2880 (N_2880,N_1412,N_1210);
and U2881 (N_2881,N_1334,N_1836);
xnor U2882 (N_2882,N_1177,N_1253);
nor U2883 (N_2883,N_1438,N_1644);
nor U2884 (N_2884,N_1828,N_1266);
and U2885 (N_2885,N_1008,N_1221);
or U2886 (N_2886,N_1253,N_1112);
and U2887 (N_2887,N_1596,N_1473);
nand U2888 (N_2888,N_1938,N_1360);
nor U2889 (N_2889,N_1109,N_1644);
and U2890 (N_2890,N_1147,N_1823);
or U2891 (N_2891,N_1774,N_1062);
xnor U2892 (N_2892,N_1399,N_1700);
nand U2893 (N_2893,N_1563,N_1088);
nand U2894 (N_2894,N_1153,N_1855);
or U2895 (N_2895,N_1624,N_1849);
nand U2896 (N_2896,N_1503,N_1981);
xnor U2897 (N_2897,N_1689,N_1484);
nor U2898 (N_2898,N_1051,N_1578);
xnor U2899 (N_2899,N_1733,N_1638);
xnor U2900 (N_2900,N_1393,N_1298);
nor U2901 (N_2901,N_1089,N_1550);
or U2902 (N_2902,N_1685,N_1720);
nand U2903 (N_2903,N_1129,N_1704);
nor U2904 (N_2904,N_1865,N_1700);
nor U2905 (N_2905,N_1132,N_1916);
or U2906 (N_2906,N_1586,N_1493);
nor U2907 (N_2907,N_1862,N_1746);
nor U2908 (N_2908,N_1110,N_1902);
or U2909 (N_2909,N_1649,N_1768);
or U2910 (N_2910,N_1113,N_1720);
nand U2911 (N_2911,N_1045,N_1436);
nand U2912 (N_2912,N_1748,N_1765);
and U2913 (N_2913,N_1436,N_1142);
nor U2914 (N_2914,N_1262,N_1890);
and U2915 (N_2915,N_1776,N_1426);
nor U2916 (N_2916,N_1657,N_1625);
nand U2917 (N_2917,N_1819,N_1756);
or U2918 (N_2918,N_1506,N_1463);
and U2919 (N_2919,N_1624,N_1841);
nor U2920 (N_2920,N_1468,N_1032);
nor U2921 (N_2921,N_1718,N_1039);
nand U2922 (N_2922,N_1568,N_1730);
nor U2923 (N_2923,N_1061,N_1387);
and U2924 (N_2924,N_1745,N_1959);
nor U2925 (N_2925,N_1672,N_1175);
and U2926 (N_2926,N_1040,N_1375);
and U2927 (N_2927,N_1310,N_1176);
nor U2928 (N_2928,N_1425,N_1177);
nor U2929 (N_2929,N_1650,N_1439);
and U2930 (N_2930,N_1535,N_1274);
xor U2931 (N_2931,N_1309,N_1604);
and U2932 (N_2932,N_1720,N_1647);
and U2933 (N_2933,N_1721,N_1276);
nor U2934 (N_2934,N_1947,N_1755);
nand U2935 (N_2935,N_1518,N_1023);
xnor U2936 (N_2936,N_1445,N_1667);
nor U2937 (N_2937,N_1359,N_1471);
nor U2938 (N_2938,N_1603,N_1451);
nand U2939 (N_2939,N_1263,N_1018);
and U2940 (N_2940,N_1863,N_1114);
xnor U2941 (N_2941,N_1914,N_1412);
and U2942 (N_2942,N_1114,N_1322);
nand U2943 (N_2943,N_1919,N_1836);
and U2944 (N_2944,N_1298,N_1844);
or U2945 (N_2945,N_1837,N_1984);
nand U2946 (N_2946,N_1026,N_1476);
xor U2947 (N_2947,N_1576,N_1441);
nand U2948 (N_2948,N_1759,N_1691);
nand U2949 (N_2949,N_1006,N_1865);
and U2950 (N_2950,N_1301,N_1708);
xor U2951 (N_2951,N_1147,N_1660);
and U2952 (N_2952,N_1871,N_1676);
nand U2953 (N_2953,N_1424,N_1317);
nand U2954 (N_2954,N_1832,N_1419);
nand U2955 (N_2955,N_1133,N_1865);
or U2956 (N_2956,N_1139,N_1634);
or U2957 (N_2957,N_1149,N_1405);
and U2958 (N_2958,N_1943,N_1710);
nand U2959 (N_2959,N_1556,N_1879);
xnor U2960 (N_2960,N_1786,N_1561);
xor U2961 (N_2961,N_1528,N_1676);
and U2962 (N_2962,N_1299,N_1512);
nand U2963 (N_2963,N_1825,N_1770);
nand U2964 (N_2964,N_1996,N_1604);
or U2965 (N_2965,N_1840,N_1098);
nor U2966 (N_2966,N_1747,N_1806);
nand U2967 (N_2967,N_1835,N_1755);
xor U2968 (N_2968,N_1380,N_1147);
nand U2969 (N_2969,N_1445,N_1165);
or U2970 (N_2970,N_1917,N_1858);
nor U2971 (N_2971,N_1414,N_1068);
nand U2972 (N_2972,N_1059,N_1574);
and U2973 (N_2973,N_1660,N_1429);
nand U2974 (N_2974,N_1819,N_1883);
and U2975 (N_2975,N_1784,N_1356);
nand U2976 (N_2976,N_1685,N_1142);
nor U2977 (N_2977,N_1168,N_1132);
and U2978 (N_2978,N_1549,N_1145);
nor U2979 (N_2979,N_1852,N_1941);
and U2980 (N_2980,N_1032,N_1988);
nor U2981 (N_2981,N_1807,N_1530);
and U2982 (N_2982,N_1893,N_1934);
and U2983 (N_2983,N_1620,N_1945);
nor U2984 (N_2984,N_1639,N_1957);
nand U2985 (N_2985,N_1125,N_1684);
xnor U2986 (N_2986,N_1483,N_1595);
xor U2987 (N_2987,N_1853,N_1887);
xor U2988 (N_2988,N_1371,N_1095);
nand U2989 (N_2989,N_1471,N_1135);
and U2990 (N_2990,N_1349,N_1140);
or U2991 (N_2991,N_1783,N_1105);
or U2992 (N_2992,N_1585,N_1561);
and U2993 (N_2993,N_1931,N_1387);
and U2994 (N_2994,N_1230,N_1435);
nand U2995 (N_2995,N_1359,N_1383);
and U2996 (N_2996,N_1258,N_1307);
nor U2997 (N_2997,N_1913,N_1547);
or U2998 (N_2998,N_1019,N_1842);
and U2999 (N_2999,N_1929,N_1154);
nand U3000 (N_3000,N_2076,N_2294);
nor U3001 (N_3001,N_2298,N_2747);
or U3002 (N_3002,N_2996,N_2173);
nand U3003 (N_3003,N_2965,N_2149);
nand U3004 (N_3004,N_2953,N_2084);
and U3005 (N_3005,N_2528,N_2887);
or U3006 (N_3006,N_2377,N_2192);
or U3007 (N_3007,N_2867,N_2566);
xnor U3008 (N_3008,N_2968,N_2337);
nand U3009 (N_3009,N_2099,N_2633);
and U3010 (N_3010,N_2007,N_2058);
nand U3011 (N_3011,N_2320,N_2104);
nor U3012 (N_3012,N_2804,N_2479);
or U3013 (N_3013,N_2782,N_2625);
xnor U3014 (N_3014,N_2982,N_2473);
nor U3015 (N_3015,N_2940,N_2460);
nor U3016 (N_3016,N_2878,N_2122);
and U3017 (N_3017,N_2132,N_2111);
and U3018 (N_3018,N_2009,N_2114);
nor U3019 (N_3019,N_2862,N_2484);
nand U3020 (N_3020,N_2253,N_2730);
or U3021 (N_3021,N_2427,N_2379);
or U3022 (N_3022,N_2643,N_2963);
nor U3023 (N_3023,N_2664,N_2561);
or U3024 (N_3024,N_2966,N_2644);
nor U3025 (N_3025,N_2502,N_2592);
or U3026 (N_3026,N_2131,N_2951);
or U3027 (N_3027,N_2938,N_2726);
nand U3028 (N_3028,N_2448,N_2639);
nand U3029 (N_3029,N_2001,N_2374);
and U3030 (N_3030,N_2929,N_2046);
or U3031 (N_3031,N_2093,N_2266);
xor U3032 (N_3032,N_2278,N_2039);
nor U3033 (N_3033,N_2956,N_2600);
nor U3034 (N_3034,N_2821,N_2063);
nor U3035 (N_3035,N_2736,N_2150);
and U3036 (N_3036,N_2013,N_2373);
xor U3037 (N_3037,N_2764,N_2026);
or U3038 (N_3038,N_2771,N_2977);
or U3039 (N_3039,N_2920,N_2067);
or U3040 (N_3040,N_2435,N_2092);
or U3041 (N_3041,N_2438,N_2523);
or U3042 (N_3042,N_2455,N_2692);
or U3043 (N_3043,N_2547,N_2156);
and U3044 (N_3044,N_2694,N_2748);
or U3045 (N_3045,N_2973,N_2816);
xor U3046 (N_3046,N_2714,N_2293);
and U3047 (N_3047,N_2638,N_2043);
and U3048 (N_3048,N_2230,N_2364);
nor U3049 (N_3049,N_2369,N_2321);
xnor U3050 (N_3050,N_2525,N_2786);
nand U3051 (N_3051,N_2045,N_2500);
and U3052 (N_3052,N_2077,N_2072);
nand U3053 (N_3053,N_2050,N_2174);
and U3054 (N_3054,N_2545,N_2283);
nor U3055 (N_3055,N_2272,N_2943);
nor U3056 (N_3056,N_2961,N_2734);
or U3057 (N_3057,N_2885,N_2555);
nor U3058 (N_3058,N_2517,N_2868);
or U3059 (N_3059,N_2739,N_2875);
or U3060 (N_3060,N_2971,N_2755);
and U3061 (N_3061,N_2387,N_2306);
or U3062 (N_3062,N_2095,N_2785);
and U3063 (N_3063,N_2129,N_2746);
nand U3064 (N_3064,N_2359,N_2705);
or U3065 (N_3065,N_2967,N_2216);
or U3066 (N_3066,N_2469,N_2146);
xor U3067 (N_3067,N_2014,N_2159);
or U3068 (N_3068,N_2891,N_2312);
nand U3069 (N_3069,N_2944,N_2499);
nor U3070 (N_3070,N_2004,N_2810);
nor U3071 (N_3071,N_2184,N_2932);
nand U3072 (N_3072,N_2605,N_2620);
nor U3073 (N_3073,N_2933,N_2419);
or U3074 (N_3074,N_2357,N_2258);
nor U3075 (N_3075,N_2686,N_2098);
or U3076 (N_3076,N_2934,N_2897);
and U3077 (N_3077,N_2650,N_2773);
nand U3078 (N_3078,N_2446,N_2840);
and U3079 (N_3079,N_2580,N_2511);
nand U3080 (N_3080,N_2022,N_2912);
and U3081 (N_3081,N_2531,N_2255);
nor U3082 (N_3082,N_2440,N_2708);
or U3083 (N_3083,N_2316,N_2861);
nor U3084 (N_3084,N_2880,N_2375);
or U3085 (N_3085,N_2397,N_2762);
nand U3086 (N_3086,N_2504,N_2205);
nand U3087 (N_3087,N_2035,N_2616);
and U3088 (N_3088,N_2823,N_2843);
and U3089 (N_3089,N_2097,N_2252);
and U3090 (N_3090,N_2952,N_2994);
or U3091 (N_3091,N_2116,N_2822);
nand U3092 (N_3092,N_2801,N_2703);
nor U3093 (N_3093,N_2695,N_2018);
or U3094 (N_3094,N_2593,N_2130);
or U3095 (N_3095,N_2323,N_2855);
or U3096 (N_3096,N_2220,N_2881);
or U3097 (N_3097,N_2573,N_2218);
nor U3098 (N_3098,N_2197,N_2453);
and U3099 (N_3099,N_2661,N_2059);
and U3100 (N_3100,N_2594,N_2815);
nor U3101 (N_3101,N_2548,N_2370);
nand U3102 (N_3102,N_2649,N_2800);
nor U3103 (N_3103,N_2466,N_2222);
xnor U3104 (N_3104,N_2556,N_2475);
and U3105 (N_3105,N_2494,N_2613);
nor U3106 (N_3106,N_2400,N_2617);
and U3107 (N_3107,N_2310,N_2346);
and U3108 (N_3108,N_2472,N_2535);
nor U3109 (N_3109,N_2154,N_2865);
or U3110 (N_3110,N_2203,N_2870);
nand U3111 (N_3111,N_2434,N_2731);
nand U3112 (N_3112,N_2962,N_2893);
and U3113 (N_3113,N_2352,N_2519);
nand U3114 (N_3114,N_2186,N_2894);
nand U3115 (N_3115,N_2949,N_2915);
or U3116 (N_3116,N_2096,N_2061);
or U3117 (N_3117,N_2081,N_2284);
xnor U3118 (N_3118,N_2117,N_2751);
and U3119 (N_3119,N_2838,N_2621);
or U3120 (N_3120,N_2091,N_2612);
nor U3121 (N_3121,N_2818,N_2927);
or U3122 (N_3122,N_2391,N_2136);
and U3123 (N_3123,N_2034,N_2313);
or U3124 (N_3124,N_2463,N_2596);
and U3125 (N_3125,N_2442,N_2615);
or U3126 (N_3126,N_2318,N_2238);
nand U3127 (N_3127,N_2299,N_2376);
and U3128 (N_3128,N_2470,N_2892);
nor U3129 (N_3129,N_2226,N_2425);
nor U3130 (N_3130,N_2082,N_2848);
or U3131 (N_3131,N_2295,N_2904);
or U3132 (N_3132,N_2948,N_2195);
or U3133 (N_3133,N_2683,N_2775);
and U3134 (N_3134,N_2054,N_2118);
nand U3135 (N_3135,N_2668,N_2214);
nor U3136 (N_3136,N_2171,N_2699);
and U3137 (N_3137,N_2085,N_2172);
or U3138 (N_3138,N_2654,N_2257);
and U3139 (N_3139,N_2324,N_2721);
or U3140 (N_3140,N_2231,N_2930);
or U3141 (N_3141,N_2431,N_2685);
nor U3142 (N_3142,N_2286,N_2152);
and U3143 (N_3143,N_2209,N_2767);
nor U3144 (N_3144,N_2339,N_2309);
nor U3145 (N_3145,N_2344,N_2492);
and U3146 (N_3146,N_2642,N_2872);
nand U3147 (N_3147,N_2048,N_2987);
xor U3148 (N_3148,N_2386,N_2353);
nor U3149 (N_3149,N_2845,N_2182);
xor U3150 (N_3150,N_2863,N_2655);
and U3151 (N_3151,N_2125,N_2498);
and U3152 (N_3152,N_2583,N_2859);
nand U3153 (N_3153,N_2327,N_2529);
and U3154 (N_3154,N_2662,N_2844);
nand U3155 (N_3155,N_2563,N_2889);
or U3156 (N_3156,N_2916,N_2345);
nand U3157 (N_3157,N_2491,N_2482);
nor U3158 (N_3158,N_2486,N_2441);
and U3159 (N_3159,N_2322,N_2354);
nor U3160 (N_3160,N_2011,N_2969);
and U3161 (N_3161,N_2540,N_2980);
and U3162 (N_3162,N_2200,N_2985);
nand U3163 (N_3163,N_2756,N_2138);
nor U3164 (N_3164,N_2213,N_2836);
nand U3165 (N_3165,N_2921,N_2032);
and U3166 (N_3166,N_2413,N_2825);
and U3167 (N_3167,N_2123,N_2340);
xor U3168 (N_3168,N_2185,N_2770);
and U3169 (N_3169,N_2070,N_2693);
and U3170 (N_3170,N_2995,N_2296);
or U3171 (N_3171,N_2317,N_2236);
nand U3172 (N_3172,N_2362,N_2056);
or U3173 (N_3173,N_2763,N_2459);
nor U3174 (N_3174,N_2575,N_2372);
or U3175 (N_3175,N_2304,N_2622);
nor U3176 (N_3176,N_2645,N_2414);
or U3177 (N_3177,N_2208,N_2135);
nor U3178 (N_3178,N_2140,N_2409);
or U3179 (N_3179,N_2017,N_2990);
or U3180 (N_3180,N_2811,N_2847);
nand U3181 (N_3181,N_2449,N_2590);
xor U3182 (N_3182,N_2623,N_2019);
and U3183 (N_3183,N_2513,N_2198);
nor U3184 (N_3184,N_2788,N_2603);
xnor U3185 (N_3185,N_2632,N_2006);
nand U3186 (N_3186,N_2935,N_2906);
or U3187 (N_3187,N_2351,N_2518);
or U3188 (N_3188,N_2290,N_2522);
nor U3189 (N_3189,N_2922,N_2853);
nand U3190 (N_3190,N_2740,N_2737);
nand U3191 (N_3191,N_2673,N_2779);
and U3192 (N_3192,N_2858,N_2270);
nor U3193 (N_3193,N_2170,N_2166);
or U3194 (N_3194,N_2311,N_2089);
or U3195 (N_3195,N_2071,N_2464);
nor U3196 (N_3196,N_2716,N_2724);
or U3197 (N_3197,N_2041,N_2772);
nand U3198 (N_3198,N_2688,N_2269);
nor U3199 (N_3199,N_2647,N_2147);
xor U3200 (N_3200,N_2974,N_2188);
or U3201 (N_3201,N_2565,N_2260);
nor U3202 (N_3202,N_2248,N_2646);
and U3203 (N_3203,N_2350,N_2275);
xnor U3204 (N_3204,N_2570,N_2991);
nand U3205 (N_3205,N_2201,N_2574);
nand U3206 (N_3206,N_2177,N_2520);
and U3207 (N_3207,N_2902,N_2834);
nand U3208 (N_3208,N_2793,N_2749);
nand U3209 (N_3209,N_2338,N_2835);
nor U3210 (N_3210,N_2381,N_2168);
nor U3211 (N_3211,N_2292,N_2088);
nand U3212 (N_3212,N_2718,N_2924);
nand U3213 (N_3213,N_2051,N_2681);
nor U3214 (N_3214,N_2189,N_2207);
or U3215 (N_3215,N_2280,N_2332);
nor U3216 (N_3216,N_2271,N_2584);
and U3217 (N_3217,N_2890,N_2802);
or U3218 (N_3218,N_2404,N_2595);
nor U3219 (N_3219,N_2175,N_2126);
nand U3220 (N_3220,N_2809,N_2947);
xnor U3221 (N_3221,N_2942,N_2732);
nand U3222 (N_3222,N_2497,N_2360);
or U3223 (N_3223,N_2833,N_2115);
and U3224 (N_3224,N_2079,N_2846);
and U3225 (N_3225,N_2153,N_2796);
nand U3226 (N_3226,N_2444,N_2120);
nor U3227 (N_3227,N_2342,N_2606);
and U3228 (N_3228,N_2042,N_2799);
nor U3229 (N_3229,N_2505,N_2759);
xor U3230 (N_3230,N_2109,N_2483);
and U3231 (N_3231,N_2585,N_2542);
or U3232 (N_3232,N_2060,N_2036);
or U3233 (N_3233,N_2326,N_2829);
nor U3234 (N_3234,N_2390,N_2443);
and U3235 (N_3235,N_2509,N_2065);
nor U3236 (N_3236,N_2554,N_2027);
nand U3237 (N_3237,N_2543,N_2588);
nand U3238 (N_3238,N_2553,N_2325);
nand U3239 (N_3239,N_2757,N_2589);
or U3240 (N_3240,N_2333,N_2276);
nor U3241 (N_3241,N_2101,N_2950);
nor U3242 (N_3242,N_2086,N_2564);
or U3243 (N_3243,N_2457,N_2134);
nand U3244 (N_3244,N_2908,N_2183);
nand U3245 (N_3245,N_2780,N_2480);
nand U3246 (N_3246,N_2485,N_2477);
or U3247 (N_3247,N_2331,N_2817);
nor U3248 (N_3248,N_2488,N_2378);
nor U3249 (N_3249,N_2000,N_2659);
xor U3250 (N_3250,N_2814,N_2384);
nor U3251 (N_3251,N_2674,N_2675);
nor U3252 (N_3252,N_2745,N_2478);
nor U3253 (N_3253,N_2083,N_2249);
and U3254 (N_3254,N_2682,N_2837);
nand U3255 (N_3255,N_2742,N_2784);
nand U3256 (N_3256,N_2402,N_2539);
xor U3257 (N_3257,N_2202,N_2960);
xor U3258 (N_3258,N_2066,N_2839);
and U3259 (N_3259,N_2075,N_2917);
nor U3260 (N_3260,N_2193,N_2094);
xnor U3261 (N_3261,N_2866,N_2926);
and U3262 (N_3262,N_2807,N_2989);
and U3263 (N_3263,N_2366,N_2429);
nor U3264 (N_3264,N_2781,N_2945);
nor U3265 (N_3265,N_2078,N_2450);
nor U3266 (N_3266,N_2828,N_2028);
and U3267 (N_3267,N_2671,N_2562);
nand U3268 (N_3268,N_2988,N_2383);
nor U3269 (N_3269,N_2999,N_2240);
and U3270 (N_3270,N_2667,N_2813);
nor U3271 (N_3271,N_2476,N_2744);
nor U3272 (N_3272,N_2160,N_2637);
nor U3273 (N_3273,N_2062,N_2964);
nand U3274 (N_3274,N_2805,N_2514);
nor U3275 (N_3275,N_2420,N_2510);
xor U3276 (N_3276,N_2627,N_2911);
nand U3277 (N_3277,N_2003,N_2481);
nor U3278 (N_3278,N_2761,N_2396);
nand U3279 (N_3279,N_2774,N_2158);
nand U3280 (N_3280,N_2191,N_2416);
nand U3281 (N_3281,N_2358,N_2163);
nor U3282 (N_3282,N_2678,N_2795);
or U3283 (N_3283,N_2112,N_2722);
nand U3284 (N_3284,N_2303,N_2907);
nor U3285 (N_3285,N_2288,N_2527);
or U3286 (N_3286,N_2819,N_2239);
or U3287 (N_3287,N_2841,N_2297);
or U3288 (N_3288,N_2005,N_2301);
nor U3289 (N_3289,N_2361,N_2720);
and U3290 (N_3290,N_2335,N_2194);
or U3291 (N_3291,N_2157,N_2106);
or U3292 (N_3292,N_2127,N_2913);
nor U3293 (N_3293,N_2367,N_2955);
nand U3294 (N_3294,N_2635,N_2055);
nand U3295 (N_3295,N_2010,N_2179);
xor U3296 (N_3296,N_2426,N_2347);
or U3297 (N_3297,N_2790,N_2133);
nand U3298 (N_3298,N_2957,N_2766);
or U3299 (N_3299,N_2029,N_2753);
and U3300 (N_3300,N_2723,N_2604);
or U3301 (N_3301,N_2851,N_2827);
nand U3302 (N_3302,N_2569,N_2735);
and U3303 (N_3303,N_2849,N_2824);
and U3304 (N_3304,N_2319,N_2521);
and U3305 (N_3305,N_2599,N_2701);
and U3306 (N_3306,N_2343,N_2456);
and U3307 (N_3307,N_2053,N_2710);
or U3308 (N_3308,N_2305,N_2430);
nand U3309 (N_3309,N_2958,N_2609);
xnor U3310 (N_3310,N_2246,N_2571);
nand U3311 (N_3311,N_2002,N_2368);
xor U3312 (N_3312,N_2141,N_2250);
or U3313 (N_3313,N_2047,N_2946);
or U3314 (N_3314,N_2919,N_2242);
nand U3315 (N_3315,N_2895,N_2355);
or U3316 (N_3316,N_2235,N_2244);
or U3317 (N_3317,N_2914,N_2672);
xnor U3318 (N_3318,N_2023,N_2899);
nand U3319 (N_3319,N_2648,N_2886);
nand U3320 (N_3320,N_2489,N_2388);
and U3321 (N_3321,N_2447,N_2607);
nor U3322 (N_3322,N_2237,N_2506);
nand U3323 (N_3323,N_2155,N_2787);
xnor U3324 (N_3324,N_2884,N_2107);
nor U3325 (N_3325,N_2532,N_2541);
or U3326 (N_3326,N_2546,N_2630);
nor U3327 (N_3327,N_2883,N_2660);
and U3328 (N_3328,N_2725,N_2549);
nor U3329 (N_3329,N_2128,N_2777);
nor U3330 (N_3330,N_2329,N_2572);
and U3331 (N_3331,N_2422,N_2210);
nor U3332 (N_3332,N_2262,N_2557);
nor U3333 (N_3333,N_2656,N_2382);
nand U3334 (N_3334,N_2826,N_2978);
and U3335 (N_3335,N_2080,N_2212);
xor U3336 (N_3336,N_2877,N_2064);
and U3337 (N_3337,N_2452,N_2040);
or U3338 (N_3338,N_2579,N_2052);
or U3339 (N_3339,N_2436,N_2233);
nor U3340 (N_3340,N_2167,N_2291);
xor U3341 (N_3341,N_2729,N_2265);
and U3342 (N_3342,N_2474,N_2769);
nand U3343 (N_3343,N_2385,N_2798);
nor U3344 (N_3344,N_2704,N_2432);
nand U3345 (N_3345,N_2015,N_2445);
and U3346 (N_3346,N_2407,N_2598);
or U3347 (N_3347,N_2487,N_2418);
nand U3348 (N_3348,N_2423,N_2854);
or U3349 (N_3349,N_2727,N_2229);
nand U3350 (N_3350,N_2970,N_2776);
and U3351 (N_3351,N_2119,N_2074);
or U3352 (N_3352,N_2879,N_2653);
xnor U3353 (N_3353,N_2954,N_2451);
xnor U3354 (N_3354,N_2399,N_2411);
nor U3355 (N_3355,N_2652,N_2640);
nor U3356 (N_3356,N_2698,N_2857);
nor U3357 (N_3357,N_2712,N_2669);
nor U3358 (N_3358,N_2241,N_2274);
or U3359 (N_3359,N_2108,N_2856);
or U3360 (N_3360,N_2069,N_2439);
and U3361 (N_3361,N_2679,N_2852);
xnor U3362 (N_3362,N_2273,N_2901);
nand U3363 (N_3363,N_2997,N_2808);
or U3364 (N_3364,N_2020,N_2334);
or U3365 (N_3365,N_2628,N_2690);
or U3366 (N_3366,N_2330,N_2228);
and U3367 (N_3367,N_2806,N_2433);
xnor U3368 (N_3368,N_2534,N_2882);
or U3369 (N_3369,N_2850,N_2289);
nor U3370 (N_3370,N_2582,N_2670);
nand U3371 (N_3371,N_2842,N_2719);
and U3372 (N_3372,N_2610,N_2760);
nor U3373 (N_3373,N_2939,N_2512);
and U3374 (N_3374,N_2490,N_2406);
and U3375 (N_3375,N_2389,N_2831);
or U3376 (N_3376,N_2794,N_2282);
nand U3377 (N_3377,N_2618,N_2164);
and U3378 (N_3378,N_2008,N_2392);
or U3379 (N_3379,N_2461,N_2873);
and U3380 (N_3380,N_2405,N_2715);
or U3381 (N_3381,N_2176,N_2812);
nor U3382 (N_3382,N_2137,N_2626);
nor U3383 (N_3383,N_2550,N_2636);
and U3384 (N_3384,N_2684,N_2256);
nand U3385 (N_3385,N_2918,N_2631);
or U3386 (N_3386,N_2738,N_2869);
or U3387 (N_3387,N_2984,N_2905);
and U3388 (N_3388,N_2619,N_2597);
nor U3389 (N_3389,N_2501,N_2601);
nand U3390 (N_3390,N_2371,N_2876);
nand U3391 (N_3391,N_2689,N_2178);
and U3392 (N_3392,N_2401,N_2666);
nand U3393 (N_3393,N_2768,N_2608);
nand U3394 (N_3394,N_2462,N_2049);
nor U3395 (N_3395,N_2243,N_2219);
nand U3396 (N_3396,N_2507,N_2765);
or U3397 (N_3397,N_2162,N_2789);
xor U3398 (N_3398,N_2874,N_2832);
nor U3399 (N_3399,N_2754,N_2700);
nor U3400 (N_3400,N_2936,N_2860);
xor U3401 (N_3401,N_2778,N_2910);
and U3402 (N_3402,N_2424,N_2687);
nand U3403 (N_3403,N_2830,N_2896);
nor U3404 (N_3404,N_2139,N_2224);
nor U3405 (N_3405,N_2021,N_2268);
nor U3406 (N_3406,N_2285,N_2415);
and U3407 (N_3407,N_2680,N_2454);
or U3408 (N_3408,N_2221,N_2783);
and U3409 (N_3409,N_2651,N_2791);
nor U3410 (N_3410,N_2713,N_2676);
nor U3411 (N_3411,N_2428,N_2394);
xor U3412 (N_3412,N_2044,N_2972);
nand U3413 (N_3413,N_2349,N_2533);
or U3414 (N_3414,N_2204,N_2803);
nor U3415 (N_3415,N_2979,N_2307);
and U3416 (N_3416,N_2417,N_2206);
nand U3417 (N_3417,N_2143,N_2033);
or U3418 (N_3418,N_2544,N_2663);
and U3419 (N_3419,N_2530,N_2380);
or U3420 (N_3420,N_2797,N_2611);
nor U3421 (N_3421,N_2254,N_2925);
and U3422 (N_3422,N_2888,N_2658);
nand U3423 (N_3423,N_2287,N_2551);
nor U3424 (N_3424,N_2277,N_2012);
and U3425 (N_3425,N_2581,N_2717);
nand U3426 (N_3426,N_2264,N_2728);
nand U3427 (N_3427,N_2261,N_2587);
and U3428 (N_3428,N_2758,N_2691);
or U3429 (N_3429,N_2871,N_2508);
xnor U3430 (N_3430,N_2165,N_2398);
nand U3431 (N_3431,N_2181,N_2196);
and U3432 (N_3432,N_2300,N_2976);
xor U3433 (N_3433,N_2403,N_2903);
or U3434 (N_3434,N_2931,N_2037);
nor U3435 (N_3435,N_2395,N_2538);
nor U3436 (N_3436,N_2308,N_2180);
and U3437 (N_3437,N_2234,N_2102);
and U3438 (N_3438,N_2232,N_2552);
nand U3439 (N_3439,N_2624,N_2493);
and U3440 (N_3440,N_2187,N_2030);
or U3441 (N_3441,N_2215,N_2524);
nand U3442 (N_3442,N_2665,N_2998);
and U3443 (N_3443,N_2024,N_2105);
and U3444 (N_3444,N_2567,N_2928);
or U3445 (N_3445,N_2314,N_2151);
xor U3446 (N_3446,N_2408,N_2302);
or U3447 (N_3447,N_2245,N_2161);
and U3448 (N_3448,N_2578,N_2016);
nand U3449 (N_3449,N_2752,N_2733);
nand U3450 (N_3450,N_2121,N_2471);
or U3451 (N_3451,N_2983,N_2941);
and U3452 (N_3452,N_2657,N_2923);
nand U3453 (N_3453,N_2199,N_2251);
and U3454 (N_3454,N_2909,N_2560);
nand U3455 (N_3455,N_2558,N_2315);
nor U3456 (N_3456,N_2864,N_2467);
xor U3457 (N_3457,N_2568,N_2336);
xnor U3458 (N_3458,N_2263,N_2743);
or U3459 (N_3459,N_2992,N_2468);
nor U3460 (N_3460,N_2937,N_2281);
or U3461 (N_3461,N_2090,N_2586);
and U3462 (N_3462,N_2792,N_2110);
or U3463 (N_3463,N_2217,N_2898);
or U3464 (N_3464,N_2421,N_2515);
or U3465 (N_3465,N_2073,N_2697);
and U3466 (N_3466,N_2100,N_2820);
or U3467 (N_3467,N_2741,N_2526);
and U3468 (N_3468,N_2458,N_2437);
or U3469 (N_3469,N_2328,N_2602);
or U3470 (N_3470,N_2169,N_2087);
or U3471 (N_3471,N_2031,N_2124);
and U3472 (N_3472,N_2363,N_2103);
xnor U3473 (N_3473,N_2144,N_2696);
xnor U3474 (N_3474,N_2227,N_2536);
nor U3475 (N_3475,N_2975,N_2711);
and U3476 (N_3476,N_2225,N_2993);
and U3477 (N_3477,N_2707,N_2677);
or U3478 (N_3478,N_2410,N_2614);
or U3479 (N_3479,N_2057,N_2267);
or U3480 (N_3480,N_2634,N_2341);
xnor U3481 (N_3481,N_2190,N_2113);
nor U3482 (N_3482,N_2503,N_2279);
and U3483 (N_3483,N_2356,N_2348);
or U3484 (N_3484,N_2576,N_2641);
nor U3485 (N_3485,N_2148,N_2706);
xnor U3486 (N_3486,N_2750,N_2516);
or U3487 (N_3487,N_2981,N_2702);
or U3488 (N_3488,N_2412,N_2709);
and U3489 (N_3489,N_2496,N_2465);
or U3490 (N_3490,N_2247,N_2211);
or U3491 (N_3491,N_2577,N_2495);
nand U3492 (N_3492,N_2537,N_2365);
nand U3493 (N_3493,N_2986,N_2591);
xnor U3494 (N_3494,N_2393,N_2959);
nand U3495 (N_3495,N_2142,N_2900);
nor U3496 (N_3496,N_2145,N_2559);
nor U3497 (N_3497,N_2223,N_2629);
nand U3498 (N_3498,N_2025,N_2259);
and U3499 (N_3499,N_2068,N_2038);
or U3500 (N_3500,N_2142,N_2916);
nor U3501 (N_3501,N_2010,N_2799);
nand U3502 (N_3502,N_2587,N_2274);
or U3503 (N_3503,N_2127,N_2255);
nor U3504 (N_3504,N_2310,N_2711);
nor U3505 (N_3505,N_2548,N_2303);
nand U3506 (N_3506,N_2929,N_2906);
and U3507 (N_3507,N_2716,N_2045);
or U3508 (N_3508,N_2774,N_2486);
nand U3509 (N_3509,N_2572,N_2641);
nor U3510 (N_3510,N_2467,N_2883);
or U3511 (N_3511,N_2861,N_2461);
or U3512 (N_3512,N_2762,N_2242);
and U3513 (N_3513,N_2027,N_2779);
or U3514 (N_3514,N_2398,N_2305);
and U3515 (N_3515,N_2816,N_2174);
or U3516 (N_3516,N_2316,N_2644);
nand U3517 (N_3517,N_2012,N_2177);
and U3518 (N_3518,N_2338,N_2089);
nand U3519 (N_3519,N_2924,N_2327);
nand U3520 (N_3520,N_2217,N_2443);
nor U3521 (N_3521,N_2776,N_2192);
and U3522 (N_3522,N_2738,N_2256);
or U3523 (N_3523,N_2073,N_2269);
and U3524 (N_3524,N_2353,N_2675);
nand U3525 (N_3525,N_2351,N_2272);
or U3526 (N_3526,N_2839,N_2514);
and U3527 (N_3527,N_2231,N_2786);
or U3528 (N_3528,N_2211,N_2274);
nor U3529 (N_3529,N_2195,N_2917);
nor U3530 (N_3530,N_2642,N_2008);
or U3531 (N_3531,N_2128,N_2208);
nor U3532 (N_3532,N_2292,N_2208);
and U3533 (N_3533,N_2186,N_2630);
and U3534 (N_3534,N_2293,N_2973);
nand U3535 (N_3535,N_2487,N_2230);
xnor U3536 (N_3536,N_2326,N_2890);
or U3537 (N_3537,N_2592,N_2101);
nor U3538 (N_3538,N_2452,N_2977);
and U3539 (N_3539,N_2909,N_2954);
or U3540 (N_3540,N_2102,N_2255);
and U3541 (N_3541,N_2051,N_2091);
and U3542 (N_3542,N_2214,N_2622);
nor U3543 (N_3543,N_2827,N_2848);
nor U3544 (N_3544,N_2980,N_2432);
nand U3545 (N_3545,N_2421,N_2713);
and U3546 (N_3546,N_2507,N_2693);
nor U3547 (N_3547,N_2726,N_2946);
and U3548 (N_3548,N_2790,N_2965);
nand U3549 (N_3549,N_2225,N_2685);
and U3550 (N_3550,N_2457,N_2763);
nand U3551 (N_3551,N_2446,N_2797);
or U3552 (N_3552,N_2277,N_2699);
nand U3553 (N_3553,N_2514,N_2744);
or U3554 (N_3554,N_2726,N_2845);
or U3555 (N_3555,N_2754,N_2235);
nand U3556 (N_3556,N_2434,N_2521);
xor U3557 (N_3557,N_2333,N_2115);
or U3558 (N_3558,N_2406,N_2062);
and U3559 (N_3559,N_2959,N_2909);
nand U3560 (N_3560,N_2672,N_2178);
nand U3561 (N_3561,N_2871,N_2603);
nand U3562 (N_3562,N_2867,N_2520);
or U3563 (N_3563,N_2916,N_2206);
nor U3564 (N_3564,N_2206,N_2941);
xor U3565 (N_3565,N_2378,N_2309);
xnor U3566 (N_3566,N_2412,N_2292);
nor U3567 (N_3567,N_2689,N_2441);
and U3568 (N_3568,N_2802,N_2589);
nand U3569 (N_3569,N_2880,N_2571);
nand U3570 (N_3570,N_2421,N_2615);
and U3571 (N_3571,N_2835,N_2857);
and U3572 (N_3572,N_2393,N_2878);
nand U3573 (N_3573,N_2601,N_2983);
nor U3574 (N_3574,N_2892,N_2122);
and U3575 (N_3575,N_2447,N_2198);
nor U3576 (N_3576,N_2132,N_2800);
xor U3577 (N_3577,N_2119,N_2184);
and U3578 (N_3578,N_2352,N_2873);
and U3579 (N_3579,N_2411,N_2319);
nand U3580 (N_3580,N_2280,N_2645);
nand U3581 (N_3581,N_2879,N_2795);
nor U3582 (N_3582,N_2114,N_2541);
and U3583 (N_3583,N_2647,N_2786);
and U3584 (N_3584,N_2085,N_2894);
xor U3585 (N_3585,N_2767,N_2976);
nand U3586 (N_3586,N_2950,N_2063);
and U3587 (N_3587,N_2418,N_2299);
or U3588 (N_3588,N_2515,N_2825);
or U3589 (N_3589,N_2376,N_2008);
and U3590 (N_3590,N_2796,N_2061);
and U3591 (N_3591,N_2771,N_2547);
xnor U3592 (N_3592,N_2247,N_2079);
nor U3593 (N_3593,N_2785,N_2671);
or U3594 (N_3594,N_2361,N_2541);
and U3595 (N_3595,N_2470,N_2131);
and U3596 (N_3596,N_2464,N_2443);
nand U3597 (N_3597,N_2129,N_2595);
and U3598 (N_3598,N_2428,N_2176);
or U3599 (N_3599,N_2861,N_2775);
nand U3600 (N_3600,N_2956,N_2627);
and U3601 (N_3601,N_2886,N_2219);
or U3602 (N_3602,N_2147,N_2475);
and U3603 (N_3603,N_2709,N_2184);
xnor U3604 (N_3604,N_2076,N_2862);
or U3605 (N_3605,N_2539,N_2098);
or U3606 (N_3606,N_2141,N_2112);
nand U3607 (N_3607,N_2484,N_2870);
nand U3608 (N_3608,N_2985,N_2123);
xnor U3609 (N_3609,N_2505,N_2791);
nand U3610 (N_3610,N_2787,N_2195);
and U3611 (N_3611,N_2298,N_2872);
nor U3612 (N_3612,N_2411,N_2074);
or U3613 (N_3613,N_2987,N_2194);
nand U3614 (N_3614,N_2496,N_2405);
and U3615 (N_3615,N_2704,N_2851);
and U3616 (N_3616,N_2757,N_2531);
nor U3617 (N_3617,N_2418,N_2283);
or U3618 (N_3618,N_2197,N_2304);
nand U3619 (N_3619,N_2458,N_2439);
xnor U3620 (N_3620,N_2445,N_2791);
nand U3621 (N_3621,N_2815,N_2589);
nand U3622 (N_3622,N_2108,N_2644);
xnor U3623 (N_3623,N_2004,N_2877);
nand U3624 (N_3624,N_2420,N_2045);
nor U3625 (N_3625,N_2253,N_2237);
nand U3626 (N_3626,N_2737,N_2764);
or U3627 (N_3627,N_2257,N_2391);
nand U3628 (N_3628,N_2463,N_2938);
nor U3629 (N_3629,N_2613,N_2063);
nand U3630 (N_3630,N_2209,N_2941);
nand U3631 (N_3631,N_2012,N_2548);
nand U3632 (N_3632,N_2109,N_2946);
or U3633 (N_3633,N_2202,N_2831);
and U3634 (N_3634,N_2102,N_2448);
nand U3635 (N_3635,N_2918,N_2638);
or U3636 (N_3636,N_2654,N_2811);
nand U3637 (N_3637,N_2333,N_2036);
nor U3638 (N_3638,N_2454,N_2035);
or U3639 (N_3639,N_2446,N_2220);
or U3640 (N_3640,N_2290,N_2712);
or U3641 (N_3641,N_2893,N_2116);
nand U3642 (N_3642,N_2324,N_2489);
or U3643 (N_3643,N_2352,N_2626);
and U3644 (N_3644,N_2407,N_2439);
and U3645 (N_3645,N_2913,N_2068);
or U3646 (N_3646,N_2903,N_2869);
and U3647 (N_3647,N_2456,N_2013);
and U3648 (N_3648,N_2353,N_2600);
or U3649 (N_3649,N_2418,N_2267);
nor U3650 (N_3650,N_2312,N_2587);
and U3651 (N_3651,N_2529,N_2804);
nand U3652 (N_3652,N_2155,N_2711);
or U3653 (N_3653,N_2686,N_2419);
or U3654 (N_3654,N_2120,N_2934);
and U3655 (N_3655,N_2972,N_2287);
nor U3656 (N_3656,N_2897,N_2615);
nor U3657 (N_3657,N_2727,N_2023);
nor U3658 (N_3658,N_2984,N_2912);
nor U3659 (N_3659,N_2720,N_2710);
and U3660 (N_3660,N_2549,N_2576);
or U3661 (N_3661,N_2260,N_2758);
nor U3662 (N_3662,N_2495,N_2012);
or U3663 (N_3663,N_2545,N_2247);
or U3664 (N_3664,N_2991,N_2538);
and U3665 (N_3665,N_2748,N_2239);
and U3666 (N_3666,N_2545,N_2661);
or U3667 (N_3667,N_2326,N_2185);
or U3668 (N_3668,N_2298,N_2385);
and U3669 (N_3669,N_2769,N_2027);
or U3670 (N_3670,N_2676,N_2735);
nor U3671 (N_3671,N_2067,N_2474);
and U3672 (N_3672,N_2078,N_2580);
or U3673 (N_3673,N_2665,N_2305);
nor U3674 (N_3674,N_2605,N_2333);
or U3675 (N_3675,N_2928,N_2059);
or U3676 (N_3676,N_2837,N_2912);
or U3677 (N_3677,N_2071,N_2565);
or U3678 (N_3678,N_2463,N_2274);
and U3679 (N_3679,N_2030,N_2459);
nand U3680 (N_3680,N_2942,N_2038);
or U3681 (N_3681,N_2135,N_2994);
nand U3682 (N_3682,N_2120,N_2604);
nor U3683 (N_3683,N_2992,N_2697);
or U3684 (N_3684,N_2932,N_2011);
and U3685 (N_3685,N_2287,N_2100);
and U3686 (N_3686,N_2653,N_2667);
nor U3687 (N_3687,N_2342,N_2803);
nor U3688 (N_3688,N_2846,N_2299);
xnor U3689 (N_3689,N_2726,N_2923);
and U3690 (N_3690,N_2654,N_2620);
nor U3691 (N_3691,N_2877,N_2346);
and U3692 (N_3692,N_2036,N_2779);
and U3693 (N_3693,N_2147,N_2455);
and U3694 (N_3694,N_2720,N_2594);
xnor U3695 (N_3695,N_2442,N_2669);
or U3696 (N_3696,N_2081,N_2429);
and U3697 (N_3697,N_2520,N_2192);
nor U3698 (N_3698,N_2997,N_2783);
nor U3699 (N_3699,N_2958,N_2963);
and U3700 (N_3700,N_2522,N_2486);
nand U3701 (N_3701,N_2988,N_2752);
and U3702 (N_3702,N_2647,N_2797);
and U3703 (N_3703,N_2771,N_2576);
or U3704 (N_3704,N_2774,N_2842);
and U3705 (N_3705,N_2073,N_2706);
or U3706 (N_3706,N_2886,N_2526);
and U3707 (N_3707,N_2591,N_2573);
nor U3708 (N_3708,N_2934,N_2807);
or U3709 (N_3709,N_2498,N_2098);
and U3710 (N_3710,N_2120,N_2555);
nor U3711 (N_3711,N_2763,N_2632);
or U3712 (N_3712,N_2791,N_2421);
nand U3713 (N_3713,N_2590,N_2405);
and U3714 (N_3714,N_2527,N_2298);
nor U3715 (N_3715,N_2383,N_2072);
and U3716 (N_3716,N_2943,N_2695);
or U3717 (N_3717,N_2901,N_2430);
nor U3718 (N_3718,N_2859,N_2757);
nor U3719 (N_3719,N_2195,N_2512);
nor U3720 (N_3720,N_2486,N_2271);
and U3721 (N_3721,N_2023,N_2189);
and U3722 (N_3722,N_2813,N_2208);
and U3723 (N_3723,N_2674,N_2168);
and U3724 (N_3724,N_2810,N_2869);
or U3725 (N_3725,N_2126,N_2599);
and U3726 (N_3726,N_2585,N_2399);
and U3727 (N_3727,N_2256,N_2842);
nor U3728 (N_3728,N_2518,N_2209);
and U3729 (N_3729,N_2396,N_2730);
or U3730 (N_3730,N_2513,N_2226);
and U3731 (N_3731,N_2703,N_2925);
and U3732 (N_3732,N_2983,N_2516);
nand U3733 (N_3733,N_2669,N_2004);
and U3734 (N_3734,N_2497,N_2644);
nand U3735 (N_3735,N_2129,N_2670);
nor U3736 (N_3736,N_2228,N_2130);
and U3737 (N_3737,N_2868,N_2750);
and U3738 (N_3738,N_2752,N_2368);
nand U3739 (N_3739,N_2179,N_2582);
nor U3740 (N_3740,N_2673,N_2111);
xnor U3741 (N_3741,N_2732,N_2169);
and U3742 (N_3742,N_2676,N_2795);
nor U3743 (N_3743,N_2827,N_2252);
xnor U3744 (N_3744,N_2048,N_2744);
or U3745 (N_3745,N_2925,N_2023);
and U3746 (N_3746,N_2058,N_2542);
or U3747 (N_3747,N_2631,N_2360);
nor U3748 (N_3748,N_2037,N_2731);
or U3749 (N_3749,N_2138,N_2314);
and U3750 (N_3750,N_2531,N_2665);
or U3751 (N_3751,N_2606,N_2321);
nand U3752 (N_3752,N_2570,N_2620);
xnor U3753 (N_3753,N_2641,N_2474);
nor U3754 (N_3754,N_2986,N_2253);
or U3755 (N_3755,N_2705,N_2976);
nand U3756 (N_3756,N_2375,N_2827);
and U3757 (N_3757,N_2062,N_2097);
and U3758 (N_3758,N_2956,N_2454);
xnor U3759 (N_3759,N_2070,N_2720);
xnor U3760 (N_3760,N_2143,N_2676);
nand U3761 (N_3761,N_2310,N_2799);
or U3762 (N_3762,N_2845,N_2882);
nand U3763 (N_3763,N_2254,N_2252);
nand U3764 (N_3764,N_2855,N_2151);
and U3765 (N_3765,N_2267,N_2311);
xor U3766 (N_3766,N_2300,N_2496);
nand U3767 (N_3767,N_2266,N_2469);
or U3768 (N_3768,N_2660,N_2268);
or U3769 (N_3769,N_2907,N_2740);
xor U3770 (N_3770,N_2688,N_2542);
or U3771 (N_3771,N_2009,N_2887);
xor U3772 (N_3772,N_2197,N_2940);
nor U3773 (N_3773,N_2277,N_2365);
and U3774 (N_3774,N_2746,N_2910);
and U3775 (N_3775,N_2664,N_2706);
and U3776 (N_3776,N_2646,N_2701);
and U3777 (N_3777,N_2110,N_2905);
or U3778 (N_3778,N_2863,N_2333);
nor U3779 (N_3779,N_2734,N_2916);
and U3780 (N_3780,N_2728,N_2792);
nor U3781 (N_3781,N_2684,N_2873);
and U3782 (N_3782,N_2552,N_2053);
nor U3783 (N_3783,N_2214,N_2697);
nor U3784 (N_3784,N_2214,N_2638);
nand U3785 (N_3785,N_2367,N_2158);
or U3786 (N_3786,N_2316,N_2231);
nand U3787 (N_3787,N_2700,N_2835);
nand U3788 (N_3788,N_2682,N_2960);
nand U3789 (N_3789,N_2093,N_2331);
nor U3790 (N_3790,N_2641,N_2432);
and U3791 (N_3791,N_2715,N_2074);
and U3792 (N_3792,N_2880,N_2767);
and U3793 (N_3793,N_2856,N_2424);
nor U3794 (N_3794,N_2013,N_2738);
nand U3795 (N_3795,N_2371,N_2341);
nor U3796 (N_3796,N_2185,N_2583);
nand U3797 (N_3797,N_2075,N_2367);
and U3798 (N_3798,N_2328,N_2074);
or U3799 (N_3799,N_2192,N_2857);
and U3800 (N_3800,N_2849,N_2898);
or U3801 (N_3801,N_2847,N_2572);
nor U3802 (N_3802,N_2635,N_2013);
nand U3803 (N_3803,N_2809,N_2147);
or U3804 (N_3804,N_2670,N_2057);
nor U3805 (N_3805,N_2796,N_2882);
or U3806 (N_3806,N_2633,N_2830);
nor U3807 (N_3807,N_2273,N_2362);
or U3808 (N_3808,N_2460,N_2624);
nor U3809 (N_3809,N_2942,N_2463);
nor U3810 (N_3810,N_2333,N_2049);
or U3811 (N_3811,N_2044,N_2196);
nand U3812 (N_3812,N_2343,N_2690);
nand U3813 (N_3813,N_2233,N_2547);
or U3814 (N_3814,N_2628,N_2301);
nor U3815 (N_3815,N_2454,N_2951);
and U3816 (N_3816,N_2823,N_2375);
nor U3817 (N_3817,N_2307,N_2737);
nand U3818 (N_3818,N_2531,N_2512);
or U3819 (N_3819,N_2765,N_2552);
nand U3820 (N_3820,N_2495,N_2547);
nor U3821 (N_3821,N_2689,N_2948);
nor U3822 (N_3822,N_2383,N_2976);
and U3823 (N_3823,N_2957,N_2634);
xor U3824 (N_3824,N_2866,N_2126);
and U3825 (N_3825,N_2816,N_2995);
nor U3826 (N_3826,N_2400,N_2263);
xor U3827 (N_3827,N_2730,N_2969);
or U3828 (N_3828,N_2346,N_2640);
or U3829 (N_3829,N_2596,N_2898);
or U3830 (N_3830,N_2245,N_2568);
nor U3831 (N_3831,N_2401,N_2682);
or U3832 (N_3832,N_2430,N_2203);
and U3833 (N_3833,N_2738,N_2317);
nor U3834 (N_3834,N_2779,N_2522);
nor U3835 (N_3835,N_2438,N_2769);
nor U3836 (N_3836,N_2644,N_2441);
or U3837 (N_3837,N_2023,N_2108);
nand U3838 (N_3838,N_2900,N_2562);
nor U3839 (N_3839,N_2212,N_2637);
nor U3840 (N_3840,N_2127,N_2766);
or U3841 (N_3841,N_2010,N_2175);
nand U3842 (N_3842,N_2056,N_2804);
or U3843 (N_3843,N_2756,N_2129);
xnor U3844 (N_3844,N_2556,N_2842);
and U3845 (N_3845,N_2270,N_2743);
or U3846 (N_3846,N_2486,N_2631);
or U3847 (N_3847,N_2140,N_2463);
nor U3848 (N_3848,N_2054,N_2932);
nand U3849 (N_3849,N_2867,N_2527);
and U3850 (N_3850,N_2263,N_2216);
nor U3851 (N_3851,N_2340,N_2984);
xnor U3852 (N_3852,N_2135,N_2262);
nor U3853 (N_3853,N_2833,N_2880);
nand U3854 (N_3854,N_2967,N_2485);
nor U3855 (N_3855,N_2244,N_2374);
nor U3856 (N_3856,N_2016,N_2402);
nor U3857 (N_3857,N_2739,N_2082);
xor U3858 (N_3858,N_2199,N_2183);
nand U3859 (N_3859,N_2340,N_2049);
or U3860 (N_3860,N_2350,N_2530);
nand U3861 (N_3861,N_2796,N_2905);
nand U3862 (N_3862,N_2589,N_2690);
nor U3863 (N_3863,N_2305,N_2233);
and U3864 (N_3864,N_2651,N_2988);
nand U3865 (N_3865,N_2790,N_2453);
nand U3866 (N_3866,N_2820,N_2657);
and U3867 (N_3867,N_2082,N_2703);
nor U3868 (N_3868,N_2184,N_2312);
and U3869 (N_3869,N_2877,N_2440);
xor U3870 (N_3870,N_2259,N_2236);
or U3871 (N_3871,N_2985,N_2734);
nand U3872 (N_3872,N_2236,N_2894);
and U3873 (N_3873,N_2908,N_2511);
nor U3874 (N_3874,N_2331,N_2924);
and U3875 (N_3875,N_2287,N_2025);
nand U3876 (N_3876,N_2499,N_2254);
or U3877 (N_3877,N_2416,N_2109);
or U3878 (N_3878,N_2928,N_2638);
nor U3879 (N_3879,N_2968,N_2746);
and U3880 (N_3880,N_2298,N_2751);
nand U3881 (N_3881,N_2522,N_2504);
nand U3882 (N_3882,N_2287,N_2638);
nor U3883 (N_3883,N_2767,N_2208);
or U3884 (N_3884,N_2761,N_2755);
xnor U3885 (N_3885,N_2635,N_2852);
and U3886 (N_3886,N_2149,N_2923);
nor U3887 (N_3887,N_2881,N_2702);
and U3888 (N_3888,N_2846,N_2187);
nor U3889 (N_3889,N_2211,N_2373);
and U3890 (N_3890,N_2115,N_2211);
and U3891 (N_3891,N_2117,N_2518);
nor U3892 (N_3892,N_2063,N_2131);
nand U3893 (N_3893,N_2426,N_2039);
xnor U3894 (N_3894,N_2392,N_2581);
and U3895 (N_3895,N_2266,N_2704);
and U3896 (N_3896,N_2272,N_2864);
nand U3897 (N_3897,N_2794,N_2153);
nor U3898 (N_3898,N_2458,N_2833);
or U3899 (N_3899,N_2161,N_2751);
xnor U3900 (N_3900,N_2666,N_2531);
xnor U3901 (N_3901,N_2774,N_2199);
and U3902 (N_3902,N_2998,N_2231);
and U3903 (N_3903,N_2729,N_2319);
or U3904 (N_3904,N_2506,N_2365);
nand U3905 (N_3905,N_2306,N_2653);
nand U3906 (N_3906,N_2763,N_2007);
nand U3907 (N_3907,N_2431,N_2531);
or U3908 (N_3908,N_2833,N_2966);
or U3909 (N_3909,N_2830,N_2933);
or U3910 (N_3910,N_2018,N_2243);
and U3911 (N_3911,N_2421,N_2622);
and U3912 (N_3912,N_2366,N_2986);
or U3913 (N_3913,N_2225,N_2181);
or U3914 (N_3914,N_2123,N_2179);
or U3915 (N_3915,N_2376,N_2394);
and U3916 (N_3916,N_2945,N_2344);
or U3917 (N_3917,N_2923,N_2421);
nand U3918 (N_3918,N_2851,N_2502);
nor U3919 (N_3919,N_2221,N_2127);
or U3920 (N_3920,N_2607,N_2975);
or U3921 (N_3921,N_2026,N_2524);
nor U3922 (N_3922,N_2285,N_2438);
nand U3923 (N_3923,N_2128,N_2754);
xor U3924 (N_3924,N_2245,N_2469);
nor U3925 (N_3925,N_2782,N_2046);
nand U3926 (N_3926,N_2858,N_2385);
or U3927 (N_3927,N_2222,N_2125);
nor U3928 (N_3928,N_2494,N_2823);
and U3929 (N_3929,N_2443,N_2843);
nor U3930 (N_3930,N_2798,N_2969);
xor U3931 (N_3931,N_2450,N_2930);
xor U3932 (N_3932,N_2225,N_2898);
nor U3933 (N_3933,N_2686,N_2930);
nor U3934 (N_3934,N_2824,N_2449);
nor U3935 (N_3935,N_2038,N_2499);
and U3936 (N_3936,N_2605,N_2188);
nand U3937 (N_3937,N_2715,N_2584);
nor U3938 (N_3938,N_2516,N_2165);
and U3939 (N_3939,N_2052,N_2978);
nand U3940 (N_3940,N_2297,N_2499);
and U3941 (N_3941,N_2036,N_2188);
xor U3942 (N_3942,N_2442,N_2278);
and U3943 (N_3943,N_2731,N_2019);
nor U3944 (N_3944,N_2975,N_2013);
and U3945 (N_3945,N_2923,N_2228);
nor U3946 (N_3946,N_2622,N_2498);
nor U3947 (N_3947,N_2993,N_2449);
or U3948 (N_3948,N_2320,N_2235);
nand U3949 (N_3949,N_2446,N_2386);
nand U3950 (N_3950,N_2560,N_2005);
xor U3951 (N_3951,N_2493,N_2495);
nand U3952 (N_3952,N_2752,N_2462);
and U3953 (N_3953,N_2910,N_2000);
and U3954 (N_3954,N_2066,N_2065);
and U3955 (N_3955,N_2243,N_2123);
nor U3956 (N_3956,N_2098,N_2903);
xnor U3957 (N_3957,N_2014,N_2559);
nor U3958 (N_3958,N_2553,N_2411);
xnor U3959 (N_3959,N_2844,N_2935);
and U3960 (N_3960,N_2141,N_2579);
nand U3961 (N_3961,N_2681,N_2107);
nand U3962 (N_3962,N_2974,N_2756);
nand U3963 (N_3963,N_2046,N_2080);
xnor U3964 (N_3964,N_2885,N_2280);
or U3965 (N_3965,N_2051,N_2323);
nor U3966 (N_3966,N_2644,N_2058);
nand U3967 (N_3967,N_2570,N_2320);
nand U3968 (N_3968,N_2868,N_2736);
nand U3969 (N_3969,N_2083,N_2084);
xnor U3970 (N_3970,N_2837,N_2688);
nor U3971 (N_3971,N_2387,N_2717);
or U3972 (N_3972,N_2103,N_2917);
nand U3973 (N_3973,N_2318,N_2827);
or U3974 (N_3974,N_2090,N_2105);
or U3975 (N_3975,N_2034,N_2498);
xnor U3976 (N_3976,N_2575,N_2654);
nor U3977 (N_3977,N_2612,N_2843);
nor U3978 (N_3978,N_2903,N_2452);
and U3979 (N_3979,N_2919,N_2848);
or U3980 (N_3980,N_2418,N_2178);
or U3981 (N_3981,N_2580,N_2975);
or U3982 (N_3982,N_2793,N_2005);
nor U3983 (N_3983,N_2388,N_2966);
nor U3984 (N_3984,N_2611,N_2867);
and U3985 (N_3985,N_2542,N_2383);
and U3986 (N_3986,N_2891,N_2208);
nand U3987 (N_3987,N_2433,N_2458);
xnor U3988 (N_3988,N_2351,N_2930);
and U3989 (N_3989,N_2458,N_2191);
or U3990 (N_3990,N_2048,N_2658);
xor U3991 (N_3991,N_2165,N_2823);
or U3992 (N_3992,N_2570,N_2215);
nor U3993 (N_3993,N_2562,N_2178);
nor U3994 (N_3994,N_2966,N_2728);
nor U3995 (N_3995,N_2720,N_2578);
and U3996 (N_3996,N_2792,N_2468);
or U3997 (N_3997,N_2365,N_2318);
or U3998 (N_3998,N_2858,N_2445);
or U3999 (N_3999,N_2224,N_2530);
nand U4000 (N_4000,N_3387,N_3686);
nand U4001 (N_4001,N_3421,N_3887);
nand U4002 (N_4002,N_3598,N_3735);
and U4003 (N_4003,N_3396,N_3720);
nor U4004 (N_4004,N_3769,N_3167);
and U4005 (N_4005,N_3064,N_3609);
and U4006 (N_4006,N_3631,N_3370);
or U4007 (N_4007,N_3157,N_3818);
xnor U4008 (N_4008,N_3416,N_3966);
or U4009 (N_4009,N_3853,N_3908);
nor U4010 (N_4010,N_3572,N_3653);
nand U4011 (N_4011,N_3923,N_3106);
nor U4012 (N_4012,N_3814,N_3329);
or U4013 (N_4013,N_3273,N_3304);
or U4014 (N_4014,N_3099,N_3988);
xnor U4015 (N_4015,N_3406,N_3776);
xnor U4016 (N_4016,N_3778,N_3932);
or U4017 (N_4017,N_3333,N_3436);
and U4018 (N_4018,N_3910,N_3994);
nor U4019 (N_4019,N_3664,N_3838);
and U4020 (N_4020,N_3420,N_3285);
nor U4021 (N_4021,N_3641,N_3309);
or U4022 (N_4022,N_3475,N_3193);
nor U4023 (N_4023,N_3467,N_3009);
and U4024 (N_4024,N_3753,N_3871);
or U4025 (N_4025,N_3086,N_3444);
xnor U4026 (N_4026,N_3974,N_3854);
and U4027 (N_4027,N_3177,N_3352);
or U4028 (N_4028,N_3052,N_3704);
and U4029 (N_4029,N_3105,N_3144);
or U4030 (N_4030,N_3522,N_3293);
nor U4031 (N_4031,N_3297,N_3063);
nor U4032 (N_4032,N_3365,N_3800);
and U4033 (N_4033,N_3441,N_3541);
and U4034 (N_4034,N_3795,N_3348);
nand U4035 (N_4035,N_3582,N_3514);
nor U4036 (N_4036,N_3862,N_3575);
xor U4037 (N_4037,N_3397,N_3104);
nand U4038 (N_4038,N_3740,N_3811);
nor U4039 (N_4039,N_3981,N_3788);
and U4040 (N_4040,N_3858,N_3823);
and U4041 (N_4041,N_3799,N_3107);
and U4042 (N_4042,N_3813,N_3069);
or U4043 (N_4043,N_3591,N_3801);
nand U4044 (N_4044,N_3497,N_3689);
or U4045 (N_4045,N_3516,N_3935);
xor U4046 (N_4046,N_3392,N_3618);
xor U4047 (N_4047,N_3526,N_3240);
nor U4048 (N_4048,N_3098,N_3471);
xnor U4049 (N_4049,N_3601,N_3235);
xnor U4050 (N_4050,N_3532,N_3041);
nand U4051 (N_4051,N_3132,N_3511);
and U4052 (N_4052,N_3611,N_3652);
or U4053 (N_4053,N_3496,N_3362);
and U4054 (N_4054,N_3973,N_3825);
or U4055 (N_4055,N_3787,N_3758);
or U4056 (N_4056,N_3116,N_3386);
nand U4057 (N_4057,N_3045,N_3894);
nor U4058 (N_4058,N_3832,N_3023);
nand U4059 (N_4059,N_3081,N_3487);
and U4060 (N_4060,N_3693,N_3508);
nor U4061 (N_4061,N_3223,N_3003);
and U4062 (N_4062,N_3166,N_3163);
and U4063 (N_4063,N_3569,N_3791);
nand U4064 (N_4064,N_3879,N_3488);
and U4065 (N_4065,N_3991,N_3890);
and U4066 (N_4066,N_3377,N_3793);
or U4067 (N_4067,N_3939,N_3750);
xnor U4068 (N_4068,N_3615,N_3250);
nand U4069 (N_4069,N_3903,N_3095);
nor U4070 (N_4070,N_3115,N_3028);
nor U4071 (N_4071,N_3480,N_3438);
and U4072 (N_4072,N_3427,N_3938);
xnor U4073 (N_4073,N_3660,N_3713);
xor U4074 (N_4074,N_3647,N_3902);
and U4075 (N_4075,N_3227,N_3243);
or U4076 (N_4076,N_3470,N_3145);
and U4077 (N_4077,N_3930,N_3958);
and U4078 (N_4078,N_3180,N_3186);
nor U4079 (N_4079,N_3752,N_3946);
nor U4080 (N_4080,N_3936,N_3563);
nand U4081 (N_4081,N_3049,N_3607);
and U4082 (N_4082,N_3411,N_3617);
nor U4083 (N_4083,N_3260,N_3739);
or U4084 (N_4084,N_3692,N_3307);
nor U4085 (N_4085,N_3619,N_3507);
nor U4086 (N_4086,N_3733,N_3032);
xnor U4087 (N_4087,N_3663,N_3108);
or U4088 (N_4088,N_3831,N_3812);
and U4089 (N_4089,N_3707,N_3662);
xnor U4090 (N_4090,N_3161,N_3816);
nor U4091 (N_4091,N_3817,N_3059);
or U4092 (N_4092,N_3082,N_3262);
or U4093 (N_4093,N_3238,N_3136);
nand U4094 (N_4094,N_3667,N_3738);
and U4095 (N_4095,N_3642,N_3583);
and U4096 (N_4096,N_3525,N_3863);
nand U4097 (N_4097,N_3356,N_3494);
and U4098 (N_4098,N_3548,N_3382);
or U4099 (N_4099,N_3864,N_3965);
and U4100 (N_4100,N_3056,N_3431);
nor U4101 (N_4101,N_3898,N_3876);
nor U4102 (N_4102,N_3141,N_3391);
nand U4103 (N_4103,N_3623,N_3715);
and U4104 (N_4104,N_3024,N_3389);
and U4105 (N_4105,N_3054,N_3709);
or U4106 (N_4106,N_3867,N_3101);
and U4107 (N_4107,N_3603,N_3326);
xor U4108 (N_4108,N_3531,N_3697);
and U4109 (N_4109,N_3192,N_3027);
xor U4110 (N_4110,N_3806,N_3628);
or U4111 (N_4111,N_3393,N_3530);
nand U4112 (N_4112,N_3513,N_3367);
or U4113 (N_4113,N_3668,N_3320);
nand U4114 (N_4114,N_3085,N_3636);
and U4115 (N_4115,N_3482,N_3445);
nor U4116 (N_4116,N_3498,N_3918);
and U4117 (N_4117,N_3160,N_3060);
xor U4118 (N_4118,N_3779,N_3906);
nand U4119 (N_4119,N_3589,N_3757);
or U4120 (N_4120,N_3544,N_3874);
and U4121 (N_4121,N_3378,N_3953);
nor U4122 (N_4122,N_3866,N_3634);
nor U4123 (N_4123,N_3162,N_3413);
nand U4124 (N_4124,N_3763,N_3998);
and U4125 (N_4125,N_3633,N_3435);
xor U4126 (N_4126,N_3784,N_3459);
and U4127 (N_4127,N_3460,N_3201);
nand U4128 (N_4128,N_3606,N_3143);
nand U4129 (N_4129,N_3643,N_3952);
nor U4130 (N_4130,N_3249,N_3982);
or U4131 (N_4131,N_3700,N_3680);
or U4132 (N_4132,N_3550,N_3635);
and U4133 (N_4133,N_3520,N_3417);
nor U4134 (N_4134,N_3368,N_3860);
nor U4135 (N_4135,N_3913,N_3675);
xnor U4136 (N_4136,N_3595,N_3156);
and U4137 (N_4137,N_3213,N_3454);
nor U4138 (N_4138,N_3334,N_3845);
xnor U4139 (N_4139,N_3179,N_3554);
nor U4140 (N_4140,N_3006,N_3729);
and U4141 (N_4141,N_3340,N_3899);
nand U4142 (N_4142,N_3029,N_3424);
or U4143 (N_4143,N_3640,N_3332);
nand U4144 (N_4144,N_3964,N_3978);
xnor U4145 (N_4145,N_3171,N_3540);
nand U4146 (N_4146,N_3351,N_3117);
or U4147 (N_4147,N_3884,N_3308);
or U4148 (N_4148,N_3244,N_3407);
nand U4149 (N_4149,N_3465,N_3093);
and U4150 (N_4150,N_3950,N_3521);
or U4151 (N_4151,N_3767,N_3280);
nor U4152 (N_4152,N_3001,N_3915);
nor U4153 (N_4153,N_3896,N_3716);
nor U4154 (N_4154,N_3967,N_3649);
and U4155 (N_4155,N_3736,N_3390);
and U4156 (N_4156,N_3528,N_3247);
or U4157 (N_4157,N_3466,N_3358);
or U4158 (N_4158,N_3418,N_3889);
nor U4159 (N_4159,N_3073,N_3610);
nand U4160 (N_4160,N_3168,N_3072);
or U4161 (N_4161,N_3252,N_3809);
nor U4162 (N_4162,N_3905,N_3159);
or U4163 (N_4163,N_3478,N_3518);
nand U4164 (N_4164,N_3783,N_3404);
nor U4165 (N_4165,N_3077,N_3463);
or U4166 (N_4166,N_3545,N_3139);
nor U4167 (N_4167,N_3847,N_3963);
or U4168 (N_4168,N_3364,N_3287);
xor U4169 (N_4169,N_3206,N_3555);
and U4170 (N_4170,N_3083,N_3158);
nor U4171 (N_4171,N_3302,N_3269);
nor U4172 (N_4172,N_3210,N_3588);
xor U4173 (N_4173,N_3926,N_3306);
and U4174 (N_4174,N_3219,N_3336);
or U4175 (N_4175,N_3870,N_3170);
or U4176 (N_4176,N_3030,N_3499);
nor U4177 (N_4177,N_3676,N_3533);
nand U4178 (N_4178,N_3587,N_3559);
nand U4179 (N_4179,N_3266,N_3992);
nor U4180 (N_4180,N_3682,N_3957);
and U4181 (N_4181,N_3872,N_3325);
and U4182 (N_4182,N_3921,N_3226);
and U4183 (N_4183,N_3922,N_3164);
nand U4184 (N_4184,N_3551,N_3688);
xor U4185 (N_4185,N_3313,N_3810);
nor U4186 (N_4186,N_3684,N_3924);
nor U4187 (N_4187,N_3415,N_3042);
or U4188 (N_4188,N_3855,N_3355);
and U4189 (N_4189,N_3673,N_3002);
or U4190 (N_4190,N_3299,N_3803);
nand U4191 (N_4191,N_3217,N_3360);
nor U4192 (N_4192,N_3840,N_3912);
nand U4193 (N_4193,N_3844,N_3706);
and U4194 (N_4194,N_3881,N_3792);
or U4195 (N_4195,N_3586,N_3962);
nor U4196 (N_4196,N_3549,N_3147);
or U4197 (N_4197,N_3639,N_3232);
nor U4198 (N_4198,N_3196,N_3919);
nand U4199 (N_4199,N_3119,N_3506);
xnor U4200 (N_4200,N_3129,N_3562);
and U4201 (N_4201,N_3696,N_3078);
or U4202 (N_4202,N_3625,N_3781);
nor U4203 (N_4203,N_3524,N_3019);
or U4204 (N_4204,N_3468,N_3985);
and U4205 (N_4205,N_3897,N_3376);
xor U4206 (N_4206,N_3578,N_3861);
nand U4207 (N_4207,N_3092,N_3353);
nor U4208 (N_4208,N_3339,N_3361);
nand U4209 (N_4209,N_3893,N_3597);
nor U4210 (N_4210,N_3112,N_3165);
nand U4211 (N_4211,N_3841,N_3359);
or U4212 (N_4212,N_3087,N_3409);
xor U4213 (N_4213,N_3058,N_3604);
nand U4214 (N_4214,N_3865,N_3181);
or U4215 (N_4215,N_3403,N_3286);
nand U4216 (N_4216,N_3314,N_3212);
and U4217 (N_4217,N_3802,N_3013);
or U4218 (N_4218,N_3830,N_3473);
nor U4219 (N_4219,N_3878,N_3677);
nand U4220 (N_4220,N_3674,N_3047);
nand U4221 (N_4221,N_3341,N_3651);
and U4222 (N_4222,N_3542,N_3798);
xor U4223 (N_4223,N_3630,N_3338);
xor U4224 (N_4224,N_3990,N_3256);
or U4225 (N_4225,N_3917,N_3395);
xor U4226 (N_4226,N_3311,N_3184);
nor U4227 (N_4227,N_3410,N_3268);
and U4228 (N_4228,N_3228,N_3661);
nand U4229 (N_4229,N_3654,N_3185);
nor U4230 (N_4230,N_3150,N_3986);
and U4231 (N_4231,N_3947,N_3678);
or U4232 (N_4232,N_3021,N_3146);
or U4233 (N_4233,N_3043,N_3679);
and U4234 (N_4234,N_3261,N_3379);
or U4235 (N_4235,N_3557,N_3851);
and U4236 (N_4236,N_3452,N_3349);
or U4237 (N_4237,N_3984,N_3836);
nor U4238 (N_4238,N_3949,N_3843);
nand U4239 (N_4239,N_3505,N_3567);
or U4240 (N_4240,N_3564,N_3330);
and U4241 (N_4241,N_3241,N_3584);
nor U4242 (N_4242,N_3613,N_3481);
nand U4243 (N_4243,N_3327,N_3580);
or U4244 (N_4244,N_3538,N_3321);
or U4245 (N_4245,N_3756,N_3242);
nor U4246 (N_4246,N_3423,N_3434);
xnor U4247 (N_4247,N_3515,N_3014);
nor U4248 (N_4248,N_3535,N_3565);
nor U4249 (N_4249,N_3945,N_3694);
and U4250 (N_4250,N_3195,N_3796);
xor U4251 (N_4251,N_3880,N_3182);
or U4252 (N_4252,N_3265,N_3127);
nand U4253 (N_4253,N_3560,N_3842);
nand U4254 (N_4254,N_3176,N_3931);
xnor U4255 (N_4255,N_3263,N_3373);
nor U4256 (N_4256,N_3122,N_3191);
nor U4257 (N_4257,N_3495,N_3071);
nor U4258 (N_4258,N_3296,N_3402);
and U4259 (N_4259,N_3608,N_3911);
and U4260 (N_4260,N_3558,N_3469);
or U4261 (N_4261,N_3999,N_3807);
xnor U4262 (N_4262,N_3222,N_3271);
and U4263 (N_4263,N_3303,N_3594);
or U4264 (N_4264,N_3067,N_3174);
nand U4265 (N_4265,N_3960,N_3972);
or U4266 (N_4266,N_3342,N_3476);
nand U4267 (N_4267,N_3500,N_3849);
and U4268 (N_4268,N_3820,N_3153);
nand U4269 (N_4269,N_3895,N_3732);
and U4270 (N_4270,N_3509,N_3717);
xnor U4271 (N_4271,N_3380,N_3489);
and U4272 (N_4272,N_3190,N_3237);
and U4273 (N_4273,N_3008,N_3149);
and U4274 (N_4274,N_3576,N_3432);
or U4275 (N_4275,N_3794,N_3512);
nor U4276 (N_4276,N_3666,N_3593);
or U4277 (N_4277,N_3909,N_3011);
and U4278 (N_4278,N_3109,N_3644);
or U4279 (N_4279,N_3833,N_3719);
nand U4280 (N_4280,N_3491,N_3221);
and U4281 (N_4281,N_3442,N_3780);
or U4282 (N_4282,N_3670,N_3264);
and U4283 (N_4283,N_3477,N_3394);
nand U4284 (N_4284,N_3133,N_3088);
and U4285 (N_4285,N_3343,N_3786);
xor U4286 (N_4286,N_3075,N_3169);
or U4287 (N_4287,N_3620,N_3076);
nor U4288 (N_4288,N_3037,N_3570);
xor U4289 (N_4289,N_3033,N_3455);
nor U4290 (N_4290,N_3187,N_3207);
nand U4291 (N_4291,N_3426,N_3474);
or U4292 (N_4292,N_3449,N_3288);
xor U4293 (N_4293,N_3944,N_3859);
and U4294 (N_4294,N_3900,N_3097);
or U4295 (N_4295,N_3768,N_3566);
or U4296 (N_4296,N_3022,N_3450);
nand U4297 (N_4297,N_3173,N_3821);
nand U4298 (N_4298,N_3026,N_3428);
nor U4299 (N_4299,N_3983,N_3130);
or U4300 (N_4300,N_3046,N_3592);
nor U4301 (N_4301,N_3989,N_3398);
xor U4302 (N_4302,N_3869,N_3258);
and U4303 (N_4303,N_3484,N_3742);
xnor U4304 (N_4304,N_3493,N_3062);
nor U4305 (N_4305,N_3537,N_3650);
nor U4306 (N_4306,N_3885,N_3301);
nor U4307 (N_4307,N_3070,N_3683);
and U4308 (N_4308,N_3699,N_3728);
or U4309 (N_4309,N_3724,N_3568);
or U4310 (N_4310,N_3178,N_3656);
or U4311 (N_4311,N_3773,N_3646);
xnor U4312 (N_4312,N_3084,N_3969);
and U4313 (N_4313,N_3315,N_3194);
xnor U4314 (N_4314,N_3048,N_3501);
nor U4315 (N_4315,N_3553,N_3142);
nor U4316 (N_4316,N_3961,N_3552);
nand U4317 (N_4317,N_3102,N_3230);
and U4318 (N_4318,N_3519,N_3637);
nor U4319 (N_4319,N_3039,N_3388);
nor U4320 (N_4320,N_3089,N_3034);
xnor U4321 (N_4321,N_3188,N_3727);
nand U4322 (N_4322,N_3711,N_3687);
and U4323 (N_4323,N_3135,N_3412);
nand U4324 (N_4324,N_3328,N_3714);
nand U4325 (N_4325,N_3708,N_3215);
nand U4326 (N_4326,N_3766,N_3722);
or U4327 (N_4327,N_3443,N_3581);
and U4328 (N_4328,N_3734,N_3725);
nor U4329 (N_4329,N_3492,N_3883);
nor U4330 (N_4330,N_3020,N_3038);
or U4331 (N_4331,N_3103,N_3824);
or U4332 (N_4332,N_3080,N_3829);
and U4333 (N_4333,N_3579,N_3134);
nor U4334 (N_4334,N_3638,N_3128);
xnor U4335 (N_4335,N_3970,N_3131);
nand U4336 (N_4336,N_3209,N_3543);
nor U4337 (N_4337,N_3626,N_3254);
nand U4338 (N_4338,N_3316,N_3272);
nand U4339 (N_4339,N_3120,N_3140);
nor U4340 (N_4340,N_3868,N_3721);
and U4341 (N_4341,N_3375,N_3053);
xnor U4342 (N_4342,N_3485,N_3121);
and U4343 (N_4343,N_3996,N_3202);
xnor U4344 (N_4344,N_3979,N_3453);
nor U4345 (N_4345,N_3018,N_3777);
xnor U4346 (N_4346,N_3705,N_3977);
nand U4347 (N_4347,N_3987,N_3624);
xnor U4348 (N_4348,N_3283,N_3502);
nor U4349 (N_4349,N_3956,N_3762);
or U4350 (N_4350,N_3017,N_3980);
nand U4351 (N_4351,N_3331,N_3886);
and U4352 (N_4352,N_3172,N_3312);
and U4353 (N_4353,N_3937,N_3834);
nand U4354 (N_4354,N_3672,N_3385);
or U4355 (N_4355,N_3951,N_3114);
or U4356 (N_4356,N_3224,N_3344);
nor U4357 (N_4357,N_3483,N_3590);
nor U4358 (N_4358,N_3203,N_3527);
nand U4359 (N_4359,N_3573,N_3968);
nand U4360 (N_4360,N_3826,N_3004);
and U4361 (N_4361,N_3621,N_3425);
nand U4362 (N_4362,N_3995,N_3510);
or U4363 (N_4363,N_3523,N_3245);
nor U4364 (N_4364,N_3384,N_3347);
nor U4365 (N_4365,N_3277,N_3730);
nor U4366 (N_4366,N_3929,N_3723);
and U4367 (N_4367,N_3371,N_3345);
or U4368 (N_4368,N_3955,N_3200);
nand U4369 (N_4369,N_3113,N_3892);
nor U4370 (N_4370,N_3671,N_3665);
or U4371 (N_4371,N_3175,N_3997);
nand U4372 (N_4372,N_3057,N_3298);
or U4373 (N_4373,N_3718,N_3400);
or U4374 (N_4374,N_3138,N_3925);
nor U4375 (N_4375,N_3292,N_3685);
nand U4376 (N_4376,N_3789,N_3975);
or U4377 (N_4377,N_3920,N_3771);
and U4378 (N_4378,N_3561,N_3529);
xnor U4379 (N_4379,N_3971,N_3472);
and U4380 (N_4380,N_3948,N_3440);
nand U4381 (N_4381,N_3458,N_3976);
nand U4382 (N_4382,N_3632,N_3775);
or U4383 (N_4383,N_3888,N_3448);
nor U4384 (N_4384,N_3805,N_3040);
and U4385 (N_4385,N_3600,N_3857);
nand U4386 (N_4386,N_3785,N_3819);
and U4387 (N_4387,N_3804,N_3051);
or U4388 (N_4388,N_3322,N_3659);
nor U4389 (N_4389,N_3765,N_3517);
and U4390 (N_4390,N_3839,N_3066);
and U4391 (N_4391,N_3695,N_3197);
and U4392 (N_4392,N_3790,N_3055);
nor U4393 (N_4393,N_3464,N_3236);
nand U4394 (N_4394,N_3914,N_3837);
nor U4395 (N_4395,N_3907,N_3614);
nor U4396 (N_4396,N_3933,N_3645);
nand U4397 (N_4397,N_3295,N_3747);
xnor U4398 (N_4398,N_3282,N_3943);
nor U4399 (N_4399,N_3381,N_3622);
and U4400 (N_4400,N_3737,N_3774);
nor U4401 (N_4401,N_3408,N_3031);
and U4402 (N_4402,N_3205,N_3616);
or U4403 (N_4403,N_3993,N_3754);
nor U4404 (N_4404,N_3074,N_3110);
xor U4405 (N_4405,N_3726,N_3025);
or U4406 (N_4406,N_3267,N_3731);
or U4407 (N_4407,N_3208,N_3148);
nand U4408 (N_4408,N_3751,N_3000);
nand U4409 (N_4409,N_3546,N_3366);
and U4410 (N_4410,N_3755,N_3204);
and U4411 (N_4411,N_3399,N_3189);
nor U4412 (N_4412,N_3852,N_3374);
nand U4413 (N_4413,N_3815,N_3005);
and U4414 (N_4414,N_3214,N_3012);
nand U4415 (N_4415,N_3255,N_3539);
and U4416 (N_4416,N_3536,N_3124);
nand U4417 (N_4417,N_3846,N_3571);
and U4418 (N_4418,N_3091,N_3710);
nand U4419 (N_4419,N_3916,N_3504);
nor U4420 (N_4420,N_3702,N_3904);
nand U4421 (N_4421,N_3300,N_3231);
nor U4422 (N_4422,N_3433,N_3940);
or U4423 (N_4423,N_3574,N_3761);
nand U4424 (N_4424,N_3954,N_3456);
nand U4425 (N_4425,N_3856,N_3848);
xnor U4426 (N_4426,N_3749,N_3959);
nand U4427 (N_4427,N_3486,N_3461);
nor U4428 (N_4428,N_3782,N_3891);
and U4429 (N_4429,N_3294,N_3764);
xnor U4430 (N_4430,N_3035,N_3629);
nor U4431 (N_4431,N_3934,N_3090);
nand U4432 (N_4432,N_3284,N_3490);
nor U4433 (N_4433,N_3743,N_3712);
nand U4434 (N_4434,N_3274,N_3827);
or U4435 (N_4435,N_3534,N_3828);
nand U4436 (N_4436,N_3151,N_3152);
nand U4437 (N_4437,N_3369,N_3218);
and U4438 (N_4438,N_3770,N_3276);
or U4439 (N_4439,N_3835,N_3257);
and U4440 (N_4440,N_3602,N_3248);
and U4441 (N_4441,N_3556,N_3291);
xor U4442 (N_4442,N_3346,N_3275);
and U4443 (N_4443,N_3419,N_3703);
and U4444 (N_4444,N_3808,N_3577);
nor U4445 (N_4445,N_3701,N_3759);
nor U4446 (N_4446,N_3401,N_3744);
nor U4447 (N_4447,N_3447,N_3289);
or U4448 (N_4448,N_3118,N_3941);
nand U4449 (N_4449,N_3137,N_3036);
nand U4450 (N_4450,N_3319,N_3669);
and U4451 (N_4451,N_3446,N_3942);
or U4452 (N_4452,N_3065,N_3015);
nand U4453 (N_4453,N_3503,N_3211);
or U4454 (N_4454,N_3324,N_3691);
nand U4455 (N_4455,N_3125,N_3229);
nand U4456 (N_4456,N_3126,N_3068);
and U4457 (N_4457,N_3317,N_3605);
and U4458 (N_4458,N_3698,N_3337);
nand U4459 (N_4459,N_3746,N_3061);
or U4460 (N_4460,N_3547,N_3016);
nor U4461 (N_4461,N_3901,N_3100);
nand U4462 (N_4462,N_3797,N_3183);
nand U4463 (N_4463,N_3429,N_3155);
and U4464 (N_4464,N_3310,N_3198);
and U4465 (N_4465,N_3430,N_3760);
nand U4466 (N_4466,N_3741,N_3681);
or U4467 (N_4467,N_3745,N_3437);
xnor U4468 (N_4468,N_3612,N_3259);
nor U4469 (N_4469,N_3010,N_3233);
and U4470 (N_4470,N_3596,N_3877);
nor U4471 (N_4471,N_3246,N_3875);
or U4472 (N_4472,N_3251,N_3479);
nand U4473 (N_4473,N_3225,N_3405);
nor U4474 (N_4474,N_3290,N_3648);
nor U4475 (N_4475,N_3279,N_3270);
nand U4476 (N_4476,N_3278,N_3822);
and U4477 (N_4477,N_3457,N_3323);
or U4478 (N_4478,N_3199,N_3585);
nand U4479 (N_4479,N_3350,N_3044);
xor U4480 (N_4480,N_3354,N_3094);
or U4481 (N_4481,N_3748,N_3627);
and U4482 (N_4482,N_3462,N_3414);
xor U4483 (N_4483,N_3927,N_3234);
nor U4484 (N_4484,N_3422,N_3882);
nor U4485 (N_4485,N_3451,N_3305);
or U4486 (N_4486,N_3658,N_3220);
and U4487 (N_4487,N_3216,N_3096);
nor U4488 (N_4488,N_3599,N_3873);
xor U4489 (N_4489,N_3335,N_3154);
nand U4490 (N_4490,N_3357,N_3363);
nand U4491 (N_4491,N_3050,N_3281);
and U4492 (N_4492,N_3655,N_3383);
xnor U4493 (N_4493,N_3253,N_3372);
nand U4494 (N_4494,N_3123,N_3928);
xor U4495 (N_4495,N_3079,N_3007);
and U4496 (N_4496,N_3772,N_3111);
or U4497 (N_4497,N_3439,N_3657);
nor U4498 (N_4498,N_3318,N_3239);
nand U4499 (N_4499,N_3850,N_3690);
nor U4500 (N_4500,N_3492,N_3904);
or U4501 (N_4501,N_3547,N_3665);
and U4502 (N_4502,N_3133,N_3551);
and U4503 (N_4503,N_3919,N_3472);
nand U4504 (N_4504,N_3335,N_3291);
nor U4505 (N_4505,N_3225,N_3843);
or U4506 (N_4506,N_3799,N_3980);
nand U4507 (N_4507,N_3750,N_3269);
nor U4508 (N_4508,N_3935,N_3350);
and U4509 (N_4509,N_3766,N_3683);
nor U4510 (N_4510,N_3713,N_3083);
nor U4511 (N_4511,N_3793,N_3227);
or U4512 (N_4512,N_3772,N_3938);
xnor U4513 (N_4513,N_3557,N_3193);
nand U4514 (N_4514,N_3956,N_3408);
nand U4515 (N_4515,N_3062,N_3489);
nand U4516 (N_4516,N_3889,N_3096);
nand U4517 (N_4517,N_3489,N_3054);
or U4518 (N_4518,N_3171,N_3139);
nand U4519 (N_4519,N_3990,N_3837);
or U4520 (N_4520,N_3972,N_3684);
or U4521 (N_4521,N_3908,N_3467);
nand U4522 (N_4522,N_3453,N_3531);
nor U4523 (N_4523,N_3403,N_3765);
nand U4524 (N_4524,N_3037,N_3930);
nand U4525 (N_4525,N_3581,N_3441);
or U4526 (N_4526,N_3327,N_3823);
and U4527 (N_4527,N_3447,N_3784);
nand U4528 (N_4528,N_3688,N_3187);
or U4529 (N_4529,N_3233,N_3324);
xnor U4530 (N_4530,N_3872,N_3303);
nor U4531 (N_4531,N_3896,N_3035);
nand U4532 (N_4532,N_3562,N_3344);
or U4533 (N_4533,N_3920,N_3877);
nor U4534 (N_4534,N_3106,N_3431);
nand U4535 (N_4535,N_3020,N_3611);
nor U4536 (N_4536,N_3815,N_3110);
and U4537 (N_4537,N_3284,N_3229);
nor U4538 (N_4538,N_3393,N_3191);
nand U4539 (N_4539,N_3795,N_3738);
and U4540 (N_4540,N_3768,N_3567);
and U4541 (N_4541,N_3369,N_3164);
nand U4542 (N_4542,N_3249,N_3076);
and U4543 (N_4543,N_3394,N_3768);
nor U4544 (N_4544,N_3753,N_3773);
and U4545 (N_4545,N_3330,N_3338);
and U4546 (N_4546,N_3530,N_3920);
nand U4547 (N_4547,N_3236,N_3072);
nand U4548 (N_4548,N_3550,N_3210);
and U4549 (N_4549,N_3650,N_3011);
or U4550 (N_4550,N_3418,N_3564);
nand U4551 (N_4551,N_3971,N_3461);
and U4552 (N_4552,N_3923,N_3887);
nand U4553 (N_4553,N_3906,N_3671);
nor U4554 (N_4554,N_3857,N_3559);
and U4555 (N_4555,N_3095,N_3778);
nor U4556 (N_4556,N_3826,N_3122);
or U4557 (N_4557,N_3283,N_3650);
or U4558 (N_4558,N_3171,N_3367);
nand U4559 (N_4559,N_3082,N_3823);
nand U4560 (N_4560,N_3946,N_3334);
nor U4561 (N_4561,N_3493,N_3043);
nor U4562 (N_4562,N_3026,N_3214);
or U4563 (N_4563,N_3416,N_3181);
or U4564 (N_4564,N_3111,N_3180);
or U4565 (N_4565,N_3962,N_3169);
or U4566 (N_4566,N_3019,N_3356);
nor U4567 (N_4567,N_3568,N_3092);
or U4568 (N_4568,N_3858,N_3874);
or U4569 (N_4569,N_3659,N_3835);
nand U4570 (N_4570,N_3438,N_3637);
nor U4571 (N_4571,N_3969,N_3942);
and U4572 (N_4572,N_3569,N_3127);
nand U4573 (N_4573,N_3495,N_3196);
nor U4574 (N_4574,N_3987,N_3784);
or U4575 (N_4575,N_3197,N_3730);
nor U4576 (N_4576,N_3480,N_3246);
nor U4577 (N_4577,N_3910,N_3340);
nand U4578 (N_4578,N_3346,N_3248);
xnor U4579 (N_4579,N_3180,N_3612);
nor U4580 (N_4580,N_3458,N_3267);
nor U4581 (N_4581,N_3734,N_3513);
nor U4582 (N_4582,N_3684,N_3418);
nor U4583 (N_4583,N_3764,N_3077);
nand U4584 (N_4584,N_3686,N_3893);
nor U4585 (N_4585,N_3215,N_3529);
or U4586 (N_4586,N_3790,N_3040);
nand U4587 (N_4587,N_3889,N_3481);
or U4588 (N_4588,N_3560,N_3109);
and U4589 (N_4589,N_3486,N_3293);
nand U4590 (N_4590,N_3086,N_3202);
nand U4591 (N_4591,N_3848,N_3576);
nor U4592 (N_4592,N_3460,N_3374);
and U4593 (N_4593,N_3778,N_3871);
nand U4594 (N_4594,N_3000,N_3014);
nand U4595 (N_4595,N_3633,N_3844);
nor U4596 (N_4596,N_3324,N_3903);
and U4597 (N_4597,N_3326,N_3913);
or U4598 (N_4598,N_3039,N_3713);
xnor U4599 (N_4599,N_3336,N_3230);
or U4600 (N_4600,N_3330,N_3204);
and U4601 (N_4601,N_3848,N_3389);
or U4602 (N_4602,N_3080,N_3769);
or U4603 (N_4603,N_3251,N_3515);
nand U4604 (N_4604,N_3840,N_3105);
nor U4605 (N_4605,N_3374,N_3501);
nand U4606 (N_4606,N_3721,N_3337);
and U4607 (N_4607,N_3441,N_3655);
nand U4608 (N_4608,N_3193,N_3292);
nor U4609 (N_4609,N_3830,N_3865);
and U4610 (N_4610,N_3187,N_3282);
and U4611 (N_4611,N_3000,N_3330);
nand U4612 (N_4612,N_3125,N_3790);
and U4613 (N_4613,N_3444,N_3644);
nand U4614 (N_4614,N_3826,N_3757);
nand U4615 (N_4615,N_3520,N_3809);
xor U4616 (N_4616,N_3476,N_3579);
xor U4617 (N_4617,N_3938,N_3740);
nand U4618 (N_4618,N_3795,N_3649);
or U4619 (N_4619,N_3070,N_3610);
xor U4620 (N_4620,N_3654,N_3014);
and U4621 (N_4621,N_3113,N_3131);
or U4622 (N_4622,N_3350,N_3190);
xor U4623 (N_4623,N_3620,N_3227);
and U4624 (N_4624,N_3712,N_3504);
or U4625 (N_4625,N_3141,N_3642);
or U4626 (N_4626,N_3984,N_3746);
nand U4627 (N_4627,N_3565,N_3477);
or U4628 (N_4628,N_3919,N_3547);
nor U4629 (N_4629,N_3041,N_3040);
nand U4630 (N_4630,N_3969,N_3135);
nand U4631 (N_4631,N_3156,N_3245);
or U4632 (N_4632,N_3723,N_3903);
or U4633 (N_4633,N_3997,N_3690);
and U4634 (N_4634,N_3534,N_3865);
xor U4635 (N_4635,N_3654,N_3504);
nor U4636 (N_4636,N_3156,N_3298);
nor U4637 (N_4637,N_3677,N_3720);
or U4638 (N_4638,N_3773,N_3190);
and U4639 (N_4639,N_3151,N_3450);
nand U4640 (N_4640,N_3657,N_3424);
or U4641 (N_4641,N_3029,N_3427);
or U4642 (N_4642,N_3904,N_3791);
or U4643 (N_4643,N_3764,N_3433);
or U4644 (N_4644,N_3764,N_3184);
nor U4645 (N_4645,N_3830,N_3775);
nor U4646 (N_4646,N_3516,N_3630);
xnor U4647 (N_4647,N_3045,N_3204);
nand U4648 (N_4648,N_3217,N_3203);
and U4649 (N_4649,N_3592,N_3767);
or U4650 (N_4650,N_3848,N_3528);
nand U4651 (N_4651,N_3885,N_3515);
nor U4652 (N_4652,N_3473,N_3517);
and U4653 (N_4653,N_3260,N_3209);
and U4654 (N_4654,N_3445,N_3304);
nor U4655 (N_4655,N_3248,N_3153);
nand U4656 (N_4656,N_3107,N_3115);
or U4657 (N_4657,N_3051,N_3716);
nor U4658 (N_4658,N_3813,N_3289);
or U4659 (N_4659,N_3894,N_3853);
nor U4660 (N_4660,N_3083,N_3719);
or U4661 (N_4661,N_3148,N_3949);
or U4662 (N_4662,N_3924,N_3211);
or U4663 (N_4663,N_3858,N_3149);
nand U4664 (N_4664,N_3648,N_3192);
or U4665 (N_4665,N_3274,N_3411);
or U4666 (N_4666,N_3257,N_3363);
nand U4667 (N_4667,N_3814,N_3749);
nand U4668 (N_4668,N_3351,N_3956);
nor U4669 (N_4669,N_3052,N_3761);
nor U4670 (N_4670,N_3486,N_3887);
nand U4671 (N_4671,N_3815,N_3503);
or U4672 (N_4672,N_3801,N_3844);
and U4673 (N_4673,N_3971,N_3919);
and U4674 (N_4674,N_3711,N_3983);
nor U4675 (N_4675,N_3596,N_3224);
xnor U4676 (N_4676,N_3682,N_3933);
and U4677 (N_4677,N_3510,N_3069);
and U4678 (N_4678,N_3167,N_3926);
and U4679 (N_4679,N_3711,N_3266);
or U4680 (N_4680,N_3259,N_3413);
nand U4681 (N_4681,N_3982,N_3456);
nor U4682 (N_4682,N_3963,N_3773);
and U4683 (N_4683,N_3888,N_3113);
nor U4684 (N_4684,N_3119,N_3163);
nand U4685 (N_4685,N_3919,N_3811);
or U4686 (N_4686,N_3277,N_3692);
or U4687 (N_4687,N_3410,N_3930);
or U4688 (N_4688,N_3095,N_3624);
nand U4689 (N_4689,N_3524,N_3698);
and U4690 (N_4690,N_3638,N_3963);
and U4691 (N_4691,N_3627,N_3746);
xor U4692 (N_4692,N_3533,N_3539);
nand U4693 (N_4693,N_3504,N_3438);
or U4694 (N_4694,N_3243,N_3394);
and U4695 (N_4695,N_3152,N_3627);
nor U4696 (N_4696,N_3513,N_3767);
nand U4697 (N_4697,N_3502,N_3508);
xor U4698 (N_4698,N_3506,N_3605);
nand U4699 (N_4699,N_3048,N_3341);
xor U4700 (N_4700,N_3581,N_3007);
or U4701 (N_4701,N_3370,N_3675);
nand U4702 (N_4702,N_3677,N_3705);
nor U4703 (N_4703,N_3656,N_3699);
nor U4704 (N_4704,N_3746,N_3469);
nand U4705 (N_4705,N_3529,N_3949);
or U4706 (N_4706,N_3291,N_3660);
or U4707 (N_4707,N_3339,N_3789);
nand U4708 (N_4708,N_3075,N_3919);
nor U4709 (N_4709,N_3032,N_3030);
nand U4710 (N_4710,N_3297,N_3893);
nor U4711 (N_4711,N_3358,N_3706);
xor U4712 (N_4712,N_3606,N_3706);
nand U4713 (N_4713,N_3519,N_3069);
nor U4714 (N_4714,N_3159,N_3493);
nor U4715 (N_4715,N_3336,N_3649);
or U4716 (N_4716,N_3103,N_3222);
or U4717 (N_4717,N_3993,N_3125);
nand U4718 (N_4718,N_3648,N_3391);
nand U4719 (N_4719,N_3586,N_3329);
and U4720 (N_4720,N_3304,N_3055);
or U4721 (N_4721,N_3004,N_3698);
nand U4722 (N_4722,N_3878,N_3300);
nor U4723 (N_4723,N_3486,N_3621);
nor U4724 (N_4724,N_3624,N_3018);
and U4725 (N_4725,N_3436,N_3690);
nor U4726 (N_4726,N_3729,N_3278);
or U4727 (N_4727,N_3411,N_3726);
and U4728 (N_4728,N_3508,N_3890);
xnor U4729 (N_4729,N_3188,N_3119);
nand U4730 (N_4730,N_3794,N_3809);
and U4731 (N_4731,N_3434,N_3240);
nand U4732 (N_4732,N_3317,N_3485);
nor U4733 (N_4733,N_3054,N_3358);
or U4734 (N_4734,N_3267,N_3356);
and U4735 (N_4735,N_3551,N_3484);
or U4736 (N_4736,N_3028,N_3905);
nor U4737 (N_4737,N_3066,N_3581);
nand U4738 (N_4738,N_3581,N_3220);
or U4739 (N_4739,N_3509,N_3336);
nand U4740 (N_4740,N_3871,N_3333);
nand U4741 (N_4741,N_3312,N_3150);
or U4742 (N_4742,N_3345,N_3176);
and U4743 (N_4743,N_3983,N_3987);
nor U4744 (N_4744,N_3320,N_3174);
and U4745 (N_4745,N_3218,N_3650);
and U4746 (N_4746,N_3011,N_3870);
nor U4747 (N_4747,N_3599,N_3923);
nand U4748 (N_4748,N_3550,N_3942);
or U4749 (N_4749,N_3288,N_3930);
nor U4750 (N_4750,N_3717,N_3690);
or U4751 (N_4751,N_3087,N_3462);
nand U4752 (N_4752,N_3871,N_3477);
nand U4753 (N_4753,N_3586,N_3706);
nor U4754 (N_4754,N_3127,N_3643);
nand U4755 (N_4755,N_3512,N_3722);
or U4756 (N_4756,N_3130,N_3773);
and U4757 (N_4757,N_3271,N_3923);
nor U4758 (N_4758,N_3130,N_3970);
nor U4759 (N_4759,N_3303,N_3630);
nand U4760 (N_4760,N_3903,N_3215);
or U4761 (N_4761,N_3440,N_3644);
nor U4762 (N_4762,N_3134,N_3892);
nor U4763 (N_4763,N_3806,N_3122);
and U4764 (N_4764,N_3400,N_3335);
and U4765 (N_4765,N_3938,N_3137);
nand U4766 (N_4766,N_3598,N_3984);
nor U4767 (N_4767,N_3580,N_3236);
or U4768 (N_4768,N_3145,N_3746);
xor U4769 (N_4769,N_3123,N_3984);
nor U4770 (N_4770,N_3086,N_3084);
nor U4771 (N_4771,N_3127,N_3720);
xor U4772 (N_4772,N_3270,N_3528);
nor U4773 (N_4773,N_3880,N_3332);
or U4774 (N_4774,N_3627,N_3234);
nor U4775 (N_4775,N_3648,N_3460);
or U4776 (N_4776,N_3308,N_3389);
nor U4777 (N_4777,N_3578,N_3432);
nor U4778 (N_4778,N_3428,N_3226);
or U4779 (N_4779,N_3174,N_3560);
nand U4780 (N_4780,N_3776,N_3969);
xor U4781 (N_4781,N_3954,N_3202);
nor U4782 (N_4782,N_3167,N_3345);
or U4783 (N_4783,N_3198,N_3937);
nor U4784 (N_4784,N_3908,N_3977);
nand U4785 (N_4785,N_3033,N_3287);
nand U4786 (N_4786,N_3155,N_3789);
or U4787 (N_4787,N_3181,N_3616);
or U4788 (N_4788,N_3083,N_3576);
or U4789 (N_4789,N_3070,N_3034);
or U4790 (N_4790,N_3485,N_3246);
and U4791 (N_4791,N_3262,N_3843);
nor U4792 (N_4792,N_3951,N_3093);
nand U4793 (N_4793,N_3189,N_3060);
and U4794 (N_4794,N_3871,N_3759);
and U4795 (N_4795,N_3463,N_3598);
or U4796 (N_4796,N_3802,N_3943);
nor U4797 (N_4797,N_3758,N_3803);
and U4798 (N_4798,N_3459,N_3291);
nand U4799 (N_4799,N_3181,N_3732);
nor U4800 (N_4800,N_3807,N_3648);
nand U4801 (N_4801,N_3333,N_3265);
nand U4802 (N_4802,N_3453,N_3223);
nor U4803 (N_4803,N_3109,N_3807);
nand U4804 (N_4804,N_3407,N_3736);
and U4805 (N_4805,N_3949,N_3181);
nand U4806 (N_4806,N_3609,N_3107);
nor U4807 (N_4807,N_3933,N_3167);
nand U4808 (N_4808,N_3242,N_3902);
nor U4809 (N_4809,N_3961,N_3815);
nand U4810 (N_4810,N_3090,N_3329);
or U4811 (N_4811,N_3361,N_3038);
or U4812 (N_4812,N_3950,N_3569);
nor U4813 (N_4813,N_3842,N_3877);
nor U4814 (N_4814,N_3053,N_3010);
or U4815 (N_4815,N_3940,N_3088);
or U4816 (N_4816,N_3090,N_3840);
nor U4817 (N_4817,N_3225,N_3524);
nor U4818 (N_4818,N_3681,N_3379);
nor U4819 (N_4819,N_3823,N_3084);
and U4820 (N_4820,N_3440,N_3270);
and U4821 (N_4821,N_3363,N_3810);
nor U4822 (N_4822,N_3527,N_3189);
and U4823 (N_4823,N_3809,N_3940);
and U4824 (N_4824,N_3473,N_3619);
or U4825 (N_4825,N_3904,N_3325);
and U4826 (N_4826,N_3172,N_3253);
nand U4827 (N_4827,N_3413,N_3303);
or U4828 (N_4828,N_3480,N_3089);
nand U4829 (N_4829,N_3986,N_3280);
and U4830 (N_4830,N_3089,N_3589);
or U4831 (N_4831,N_3304,N_3957);
nor U4832 (N_4832,N_3329,N_3650);
or U4833 (N_4833,N_3238,N_3694);
nor U4834 (N_4834,N_3758,N_3184);
or U4835 (N_4835,N_3892,N_3041);
and U4836 (N_4836,N_3883,N_3686);
and U4837 (N_4837,N_3476,N_3726);
nand U4838 (N_4838,N_3976,N_3776);
or U4839 (N_4839,N_3430,N_3677);
and U4840 (N_4840,N_3039,N_3226);
and U4841 (N_4841,N_3543,N_3829);
and U4842 (N_4842,N_3391,N_3981);
xor U4843 (N_4843,N_3680,N_3586);
and U4844 (N_4844,N_3661,N_3286);
nand U4845 (N_4845,N_3655,N_3303);
or U4846 (N_4846,N_3356,N_3499);
and U4847 (N_4847,N_3385,N_3120);
nor U4848 (N_4848,N_3469,N_3040);
nand U4849 (N_4849,N_3593,N_3139);
nor U4850 (N_4850,N_3631,N_3072);
nor U4851 (N_4851,N_3513,N_3341);
and U4852 (N_4852,N_3062,N_3377);
xnor U4853 (N_4853,N_3570,N_3973);
xnor U4854 (N_4854,N_3205,N_3189);
nor U4855 (N_4855,N_3937,N_3075);
xnor U4856 (N_4856,N_3259,N_3329);
nand U4857 (N_4857,N_3033,N_3837);
and U4858 (N_4858,N_3538,N_3584);
nand U4859 (N_4859,N_3016,N_3044);
xor U4860 (N_4860,N_3315,N_3947);
or U4861 (N_4861,N_3460,N_3369);
or U4862 (N_4862,N_3317,N_3899);
xor U4863 (N_4863,N_3390,N_3913);
xor U4864 (N_4864,N_3892,N_3434);
or U4865 (N_4865,N_3087,N_3147);
and U4866 (N_4866,N_3164,N_3962);
nor U4867 (N_4867,N_3210,N_3067);
or U4868 (N_4868,N_3792,N_3045);
or U4869 (N_4869,N_3337,N_3003);
and U4870 (N_4870,N_3812,N_3008);
nand U4871 (N_4871,N_3350,N_3086);
or U4872 (N_4872,N_3958,N_3060);
nor U4873 (N_4873,N_3874,N_3038);
nor U4874 (N_4874,N_3952,N_3723);
nor U4875 (N_4875,N_3787,N_3440);
nand U4876 (N_4876,N_3167,N_3692);
nand U4877 (N_4877,N_3028,N_3751);
or U4878 (N_4878,N_3646,N_3829);
xnor U4879 (N_4879,N_3500,N_3316);
xnor U4880 (N_4880,N_3034,N_3253);
or U4881 (N_4881,N_3086,N_3354);
nor U4882 (N_4882,N_3630,N_3646);
or U4883 (N_4883,N_3192,N_3037);
and U4884 (N_4884,N_3986,N_3316);
nor U4885 (N_4885,N_3875,N_3754);
or U4886 (N_4886,N_3255,N_3182);
or U4887 (N_4887,N_3490,N_3868);
nand U4888 (N_4888,N_3423,N_3522);
and U4889 (N_4889,N_3532,N_3981);
and U4890 (N_4890,N_3976,N_3983);
nor U4891 (N_4891,N_3113,N_3812);
xnor U4892 (N_4892,N_3466,N_3857);
nor U4893 (N_4893,N_3107,N_3070);
or U4894 (N_4894,N_3543,N_3289);
and U4895 (N_4895,N_3100,N_3938);
and U4896 (N_4896,N_3837,N_3189);
or U4897 (N_4897,N_3084,N_3475);
xor U4898 (N_4898,N_3280,N_3624);
or U4899 (N_4899,N_3292,N_3391);
xor U4900 (N_4900,N_3851,N_3392);
nor U4901 (N_4901,N_3108,N_3071);
or U4902 (N_4902,N_3239,N_3202);
nand U4903 (N_4903,N_3271,N_3209);
nand U4904 (N_4904,N_3040,N_3372);
xor U4905 (N_4905,N_3857,N_3026);
or U4906 (N_4906,N_3555,N_3078);
and U4907 (N_4907,N_3554,N_3021);
nand U4908 (N_4908,N_3032,N_3136);
xnor U4909 (N_4909,N_3311,N_3116);
or U4910 (N_4910,N_3431,N_3623);
or U4911 (N_4911,N_3212,N_3698);
and U4912 (N_4912,N_3682,N_3747);
and U4913 (N_4913,N_3235,N_3012);
nand U4914 (N_4914,N_3715,N_3912);
nor U4915 (N_4915,N_3868,N_3982);
or U4916 (N_4916,N_3355,N_3723);
nor U4917 (N_4917,N_3867,N_3148);
and U4918 (N_4918,N_3644,N_3573);
nand U4919 (N_4919,N_3657,N_3972);
or U4920 (N_4920,N_3824,N_3517);
or U4921 (N_4921,N_3039,N_3294);
nand U4922 (N_4922,N_3317,N_3377);
xnor U4923 (N_4923,N_3295,N_3342);
nor U4924 (N_4924,N_3170,N_3337);
nand U4925 (N_4925,N_3847,N_3018);
nor U4926 (N_4926,N_3689,N_3588);
nor U4927 (N_4927,N_3731,N_3473);
nor U4928 (N_4928,N_3211,N_3343);
or U4929 (N_4929,N_3384,N_3894);
nand U4930 (N_4930,N_3025,N_3071);
xor U4931 (N_4931,N_3330,N_3337);
or U4932 (N_4932,N_3644,N_3511);
and U4933 (N_4933,N_3463,N_3635);
nor U4934 (N_4934,N_3153,N_3977);
or U4935 (N_4935,N_3106,N_3830);
nand U4936 (N_4936,N_3230,N_3890);
and U4937 (N_4937,N_3919,N_3371);
nand U4938 (N_4938,N_3711,N_3246);
nand U4939 (N_4939,N_3918,N_3229);
nand U4940 (N_4940,N_3140,N_3801);
xor U4941 (N_4941,N_3398,N_3383);
and U4942 (N_4942,N_3025,N_3178);
or U4943 (N_4943,N_3203,N_3939);
nor U4944 (N_4944,N_3225,N_3738);
and U4945 (N_4945,N_3933,N_3803);
nand U4946 (N_4946,N_3191,N_3915);
nand U4947 (N_4947,N_3750,N_3963);
xnor U4948 (N_4948,N_3781,N_3795);
nand U4949 (N_4949,N_3233,N_3744);
and U4950 (N_4950,N_3765,N_3397);
nand U4951 (N_4951,N_3834,N_3617);
and U4952 (N_4952,N_3976,N_3825);
nor U4953 (N_4953,N_3816,N_3566);
or U4954 (N_4954,N_3578,N_3670);
or U4955 (N_4955,N_3055,N_3993);
nand U4956 (N_4956,N_3205,N_3971);
or U4957 (N_4957,N_3575,N_3427);
nand U4958 (N_4958,N_3823,N_3856);
nor U4959 (N_4959,N_3874,N_3661);
or U4960 (N_4960,N_3147,N_3951);
nor U4961 (N_4961,N_3991,N_3092);
or U4962 (N_4962,N_3749,N_3756);
nand U4963 (N_4963,N_3133,N_3359);
nand U4964 (N_4964,N_3460,N_3217);
and U4965 (N_4965,N_3009,N_3811);
and U4966 (N_4966,N_3445,N_3337);
xnor U4967 (N_4967,N_3072,N_3942);
nor U4968 (N_4968,N_3638,N_3677);
nand U4969 (N_4969,N_3650,N_3692);
or U4970 (N_4970,N_3489,N_3193);
or U4971 (N_4971,N_3718,N_3966);
nor U4972 (N_4972,N_3326,N_3690);
nand U4973 (N_4973,N_3578,N_3827);
nand U4974 (N_4974,N_3525,N_3349);
nor U4975 (N_4975,N_3821,N_3768);
and U4976 (N_4976,N_3600,N_3537);
nor U4977 (N_4977,N_3942,N_3715);
nor U4978 (N_4978,N_3913,N_3032);
nor U4979 (N_4979,N_3145,N_3042);
nor U4980 (N_4980,N_3907,N_3590);
xor U4981 (N_4981,N_3178,N_3193);
and U4982 (N_4982,N_3214,N_3614);
and U4983 (N_4983,N_3453,N_3029);
and U4984 (N_4984,N_3580,N_3631);
xnor U4985 (N_4985,N_3906,N_3170);
and U4986 (N_4986,N_3519,N_3638);
nor U4987 (N_4987,N_3455,N_3440);
nand U4988 (N_4988,N_3506,N_3059);
or U4989 (N_4989,N_3378,N_3561);
or U4990 (N_4990,N_3113,N_3402);
and U4991 (N_4991,N_3973,N_3870);
nor U4992 (N_4992,N_3858,N_3269);
nand U4993 (N_4993,N_3467,N_3155);
xor U4994 (N_4994,N_3076,N_3753);
nand U4995 (N_4995,N_3482,N_3424);
xor U4996 (N_4996,N_3382,N_3124);
xor U4997 (N_4997,N_3550,N_3077);
nor U4998 (N_4998,N_3174,N_3422);
nand U4999 (N_4999,N_3803,N_3439);
nor U5000 (N_5000,N_4326,N_4897);
nor U5001 (N_5001,N_4359,N_4608);
xnor U5002 (N_5002,N_4157,N_4284);
or U5003 (N_5003,N_4319,N_4810);
or U5004 (N_5004,N_4481,N_4297);
xnor U5005 (N_5005,N_4715,N_4040);
and U5006 (N_5006,N_4530,N_4698);
nand U5007 (N_5007,N_4364,N_4046);
and U5008 (N_5008,N_4438,N_4999);
or U5009 (N_5009,N_4491,N_4189);
or U5010 (N_5010,N_4376,N_4926);
nor U5011 (N_5011,N_4403,N_4766);
nor U5012 (N_5012,N_4785,N_4451);
xor U5013 (N_5013,N_4758,N_4298);
or U5014 (N_5014,N_4557,N_4240);
xnor U5015 (N_5015,N_4987,N_4583);
xnor U5016 (N_5016,N_4294,N_4652);
or U5017 (N_5017,N_4241,N_4814);
nand U5018 (N_5018,N_4008,N_4427);
and U5019 (N_5019,N_4514,N_4517);
nand U5020 (N_5020,N_4358,N_4220);
nand U5021 (N_5021,N_4551,N_4146);
and U5022 (N_5022,N_4378,N_4587);
or U5023 (N_5023,N_4743,N_4891);
nand U5024 (N_5024,N_4216,N_4187);
xor U5025 (N_5025,N_4420,N_4853);
nor U5026 (N_5026,N_4818,N_4574);
or U5027 (N_5027,N_4354,N_4951);
or U5028 (N_5028,N_4184,N_4556);
xnor U5029 (N_5029,N_4235,N_4841);
and U5030 (N_5030,N_4932,N_4499);
nand U5031 (N_5031,N_4836,N_4582);
nor U5032 (N_5032,N_4381,N_4212);
nand U5033 (N_5033,N_4397,N_4705);
nor U5034 (N_5034,N_4311,N_4479);
or U5035 (N_5035,N_4816,N_4067);
nor U5036 (N_5036,N_4324,N_4386);
nor U5037 (N_5037,N_4078,N_4800);
and U5038 (N_5038,N_4299,N_4533);
nand U5039 (N_5039,N_4928,N_4155);
and U5040 (N_5040,N_4461,N_4100);
nand U5041 (N_5041,N_4175,N_4309);
nand U5042 (N_5042,N_4173,N_4110);
nand U5043 (N_5043,N_4082,N_4779);
nor U5044 (N_5044,N_4988,N_4323);
or U5045 (N_5045,N_4858,N_4782);
nor U5046 (N_5046,N_4329,N_4979);
nor U5047 (N_5047,N_4660,N_4613);
nor U5048 (N_5048,N_4834,N_4925);
or U5049 (N_5049,N_4823,N_4000);
nor U5050 (N_5050,N_4279,N_4873);
or U5051 (N_5051,N_4150,N_4079);
nor U5052 (N_5052,N_4911,N_4941);
nand U5053 (N_5053,N_4111,N_4282);
and U5054 (N_5054,N_4103,N_4737);
nand U5055 (N_5055,N_4874,N_4751);
nor U5056 (N_5056,N_4048,N_4851);
nand U5057 (N_5057,N_4640,N_4736);
nand U5058 (N_5058,N_4576,N_4202);
xnor U5059 (N_5059,N_4559,N_4963);
xnor U5060 (N_5060,N_4983,N_4701);
nand U5061 (N_5061,N_4042,N_4607);
nor U5062 (N_5062,N_4729,N_4821);
or U5063 (N_5063,N_4986,N_4464);
nor U5064 (N_5064,N_4784,N_4207);
nand U5065 (N_5065,N_4585,N_4457);
or U5066 (N_5066,N_4492,N_4399);
nor U5067 (N_5067,N_4373,N_4203);
nand U5068 (N_5068,N_4690,N_4859);
and U5069 (N_5069,N_4706,N_4562);
nor U5070 (N_5070,N_4412,N_4208);
and U5071 (N_5071,N_4369,N_4915);
nand U5072 (N_5072,N_4436,N_4456);
or U5073 (N_5073,N_4218,N_4763);
nor U5074 (N_5074,N_4236,N_4962);
or U5075 (N_5075,N_4684,N_4720);
nand U5076 (N_5076,N_4422,N_4321);
and U5077 (N_5077,N_4382,N_4020);
nor U5078 (N_5078,N_4621,N_4136);
nor U5079 (N_5079,N_4888,N_4322);
nand U5080 (N_5080,N_4996,N_4027);
nor U5081 (N_5081,N_4016,N_4352);
and U5082 (N_5082,N_4808,N_4332);
nand U5083 (N_5083,N_4176,N_4346);
nor U5084 (N_5084,N_4072,N_4069);
and U5085 (N_5085,N_4351,N_4565);
or U5086 (N_5086,N_4964,N_4776);
and U5087 (N_5087,N_4980,N_4315);
or U5088 (N_5088,N_4474,N_4182);
nor U5089 (N_5089,N_4522,N_4091);
nor U5090 (N_5090,N_4878,N_4518);
nand U5091 (N_5091,N_4696,N_4722);
or U5092 (N_5092,N_4003,N_4919);
and U5093 (N_5093,N_4431,N_4270);
nand U5094 (N_5094,N_4250,N_4711);
or U5095 (N_5095,N_4374,N_4407);
and U5096 (N_5096,N_4985,N_4683);
xor U5097 (N_5097,N_4560,N_4300);
nand U5098 (N_5098,N_4174,N_4654);
and U5099 (N_5099,N_4248,N_4280);
nand U5100 (N_5100,N_4306,N_4658);
nand U5101 (N_5101,N_4880,N_4312);
and U5102 (N_5102,N_4114,N_4760);
nor U5103 (N_5103,N_4257,N_4748);
or U5104 (N_5104,N_4191,N_4030);
or U5105 (N_5105,N_4877,N_4510);
nand U5106 (N_5106,N_4338,N_4854);
nor U5107 (N_5107,N_4842,N_4876);
nor U5108 (N_5108,N_4889,N_4905);
and U5109 (N_5109,N_4239,N_4959);
nor U5110 (N_5110,N_4680,N_4883);
nand U5111 (N_5111,N_4575,N_4890);
or U5112 (N_5112,N_4966,N_4430);
and U5113 (N_5113,N_4090,N_4767);
and U5114 (N_5114,N_4224,N_4206);
nand U5115 (N_5115,N_4902,N_4945);
and U5116 (N_5116,N_4085,N_4256);
nor U5117 (N_5117,N_4290,N_4822);
nand U5118 (N_5118,N_4254,N_4154);
and U5119 (N_5119,N_4609,N_4862);
nand U5120 (N_5120,N_4170,N_4857);
xnor U5121 (N_5121,N_4672,N_4243);
nor U5122 (N_5122,N_4635,N_4264);
nor U5123 (N_5123,N_4958,N_4847);
or U5124 (N_5124,N_4846,N_4076);
and U5125 (N_5125,N_4527,N_4747);
xor U5126 (N_5126,N_4414,N_4591);
nor U5127 (N_5127,N_4277,N_4084);
or U5128 (N_5128,N_4707,N_4670);
xnor U5129 (N_5129,N_4327,N_4566);
or U5130 (N_5130,N_4147,N_4952);
nand U5131 (N_5131,N_4002,N_4981);
or U5132 (N_5132,N_4041,N_4601);
nor U5133 (N_5133,N_4716,N_4178);
nand U5134 (N_5134,N_4731,N_4960);
nor U5135 (N_5135,N_4480,N_4377);
nand U5136 (N_5136,N_4703,N_4893);
nand U5137 (N_5137,N_4795,N_4901);
and U5138 (N_5138,N_4093,N_4702);
nor U5139 (N_5139,N_4895,N_4555);
nand U5140 (N_5140,N_4483,N_4909);
and U5141 (N_5141,N_4128,N_4572);
xnor U5142 (N_5142,N_4471,N_4137);
nand U5143 (N_5143,N_4600,N_4472);
nor U5144 (N_5144,N_4389,N_4149);
nor U5145 (N_5145,N_4788,N_4970);
nor U5146 (N_5146,N_4022,N_4245);
and U5147 (N_5147,N_4063,N_4383);
or U5148 (N_5148,N_4615,N_4037);
nand U5149 (N_5149,N_4791,N_4444);
and U5150 (N_5150,N_4686,N_4167);
or U5151 (N_5151,N_4039,N_4501);
and U5152 (N_5152,N_4939,N_4695);
nor U5153 (N_5153,N_4283,N_4631);
nor U5154 (N_5154,N_4544,N_4169);
nand U5155 (N_5155,N_4789,N_4772);
nand U5156 (N_5156,N_4301,N_4797);
or U5157 (N_5157,N_4118,N_4950);
or U5158 (N_5158,N_4476,N_4594);
xnor U5159 (N_5159,N_4269,N_4317);
nand U5160 (N_5160,N_4503,N_4927);
nand U5161 (N_5161,N_4639,N_4343);
nor U5162 (N_5162,N_4535,N_4185);
nand U5163 (N_5163,N_4803,N_4825);
or U5164 (N_5164,N_4012,N_4098);
nor U5165 (N_5165,N_4028,N_4350);
and U5166 (N_5166,N_4164,N_4586);
nand U5167 (N_5167,N_4144,N_4253);
nor U5168 (N_5168,N_4805,N_4995);
or U5169 (N_5169,N_4429,N_4215);
and U5170 (N_5170,N_4832,N_4138);
nor U5171 (N_5171,N_4223,N_4620);
xor U5172 (N_5172,N_4467,N_4325);
nand U5173 (N_5173,N_4287,N_4840);
or U5174 (N_5174,N_4954,N_4071);
and U5175 (N_5175,N_4687,N_4596);
or U5176 (N_5176,N_4200,N_4777);
and U5177 (N_5177,N_4844,N_4630);
nor U5178 (N_5178,N_4913,N_4773);
nand U5179 (N_5179,N_4543,N_4538);
nor U5180 (N_5180,N_4267,N_4830);
nor U5181 (N_5181,N_4727,N_4525);
or U5182 (N_5182,N_4401,N_4227);
nor U5183 (N_5183,N_4056,N_4627);
nor U5184 (N_5184,N_4101,N_4644);
xor U5185 (N_5185,N_4034,N_4863);
or U5186 (N_5186,N_4095,N_4944);
or U5187 (N_5187,N_4771,N_4837);
or U5188 (N_5188,N_4550,N_4367);
or U5189 (N_5189,N_4334,N_4387);
or U5190 (N_5190,N_4192,N_4682);
xnor U5191 (N_5191,N_4740,N_4997);
and U5192 (N_5192,N_4829,N_4026);
or U5193 (N_5193,N_4708,N_4335);
nand U5194 (N_5194,N_4807,N_4469);
xnor U5195 (N_5195,N_4511,N_4819);
or U5196 (N_5196,N_4709,N_4247);
nor U5197 (N_5197,N_4508,N_4141);
nor U5198 (N_5198,N_4379,N_4083);
nor U5199 (N_5199,N_4734,N_4599);
nand U5200 (N_5200,N_4903,N_4460);
or U5201 (N_5201,N_4139,N_4904);
or U5202 (N_5202,N_4233,N_4130);
nor U5203 (N_5203,N_4602,N_4140);
nor U5204 (N_5204,N_4418,N_4077);
or U5205 (N_5205,N_4875,N_4342);
or U5206 (N_5206,N_4907,N_4674);
nand U5207 (N_5207,N_4755,N_4122);
nand U5208 (N_5208,N_4009,N_4453);
nor U5209 (N_5209,N_4942,N_4619);
and U5210 (N_5210,N_4442,N_4211);
or U5211 (N_5211,N_4852,N_4628);
and U5212 (N_5212,N_4019,N_4432);
nand U5213 (N_5213,N_4624,N_4029);
xnor U5214 (N_5214,N_4380,N_4368);
nand U5215 (N_5215,N_4662,N_4573);
or U5216 (N_5216,N_4281,N_4523);
and U5217 (N_5217,N_4035,N_4423);
or U5218 (N_5218,N_4894,N_4498);
and U5219 (N_5219,N_4470,N_4293);
nand U5220 (N_5220,N_4465,N_4567);
nor U5221 (N_5221,N_4676,N_4831);
nand U5222 (N_5222,N_4428,N_4363);
nor U5223 (N_5223,N_4713,N_4879);
nand U5224 (N_5224,N_4590,N_4679);
nor U5225 (N_5225,N_4552,N_4536);
nand U5226 (N_5226,N_4145,N_4838);
nand U5227 (N_5227,N_4217,N_4296);
and U5228 (N_5228,N_4260,N_4104);
xnor U5229 (N_5229,N_4811,N_4441);
xnor U5230 (N_5230,N_4244,N_4232);
or U5231 (N_5231,N_4865,N_4790);
xnor U5232 (N_5232,N_4168,N_4947);
nand U5233 (N_5233,N_4833,N_4765);
nor U5234 (N_5234,N_4246,N_4869);
nand U5235 (N_5235,N_4070,N_4806);
xor U5236 (N_5236,N_4937,N_4540);
and U5237 (N_5237,N_4728,N_4933);
nand U5238 (N_5238,N_4308,N_4017);
or U5239 (N_5239,N_4448,N_4675);
and U5240 (N_5240,N_4058,N_4489);
nand U5241 (N_5241,N_4957,N_4802);
nor U5242 (N_5242,N_4305,N_4882);
xor U5243 (N_5243,N_4746,N_4977);
or U5244 (N_5244,N_4867,N_4195);
and U5245 (N_5245,N_4120,N_4661);
or U5246 (N_5246,N_4316,N_4158);
nor U5247 (N_5247,N_4390,N_4064);
and U5248 (N_5248,N_4384,N_4724);
nand U5249 (N_5249,N_4458,N_4099);
nand U5250 (N_5250,N_4792,N_4234);
xnor U5251 (N_5251,N_4799,N_4375);
or U5252 (N_5252,N_4775,N_4370);
and U5253 (N_5253,N_4025,N_4922);
or U5254 (N_5254,N_4578,N_4497);
xor U5255 (N_5255,N_4450,N_4010);
nor U5256 (N_5256,N_4165,N_4973);
or U5257 (N_5257,N_4314,N_4513);
nand U5258 (N_5258,N_4692,N_4953);
nor U5259 (N_5259,N_4463,N_4249);
nand U5260 (N_5260,N_4618,N_4752);
nor U5261 (N_5261,N_4998,N_4569);
nor U5262 (N_5262,N_4188,N_4754);
and U5263 (N_5263,N_4406,N_4581);
nor U5264 (N_5264,N_4900,N_4437);
and U5265 (N_5265,N_4417,N_4295);
and U5266 (N_5266,N_4113,N_4946);
nor U5267 (N_5267,N_4395,N_4744);
nand U5268 (N_5268,N_4699,N_4860);
nand U5269 (N_5269,N_4204,N_4198);
or U5270 (N_5270,N_4357,N_4749);
xor U5271 (N_5271,N_4402,N_4826);
or U5272 (N_5272,N_4331,N_4303);
or U5273 (N_5273,N_4057,N_4221);
and U5274 (N_5274,N_4940,N_4991);
nor U5275 (N_5275,N_4595,N_4087);
or U5276 (N_5276,N_4712,N_4887);
and U5277 (N_5277,N_4049,N_4770);
nor U5278 (N_5278,N_4313,N_4885);
nand U5279 (N_5279,N_4718,N_4774);
nand U5280 (N_5280,N_4112,N_4126);
nand U5281 (N_5281,N_4493,N_4183);
and U5282 (N_5282,N_4759,N_4421);
xnor U5283 (N_5283,N_4360,N_4982);
nor U5284 (N_5284,N_4571,N_4968);
nor U5285 (N_5285,N_4866,N_4180);
nand U5286 (N_5286,N_4646,N_4892);
nor U5287 (N_5287,N_4864,N_4605);
and U5288 (N_5288,N_4735,N_4186);
xnor U5289 (N_5289,N_4115,N_4589);
nor U5290 (N_5290,N_4433,N_4507);
xor U5291 (N_5291,N_4961,N_4156);
or U5292 (N_5292,N_4129,N_4745);
and U5293 (N_5293,N_4488,N_4532);
or U5294 (N_5294,N_4161,N_4673);
and U5295 (N_5295,N_4127,N_4768);
or U5296 (N_5296,N_4967,N_4333);
xnor U5297 (N_5297,N_4344,N_4546);
and U5298 (N_5298,N_4632,N_4160);
nor U5299 (N_5299,N_4622,N_4278);
nor U5300 (N_5300,N_4539,N_4753);
xor U5301 (N_5301,N_4693,N_4005);
and U5302 (N_5302,N_4534,N_4142);
nand U5303 (N_5303,N_4181,N_4445);
or U5304 (N_5304,N_4623,N_4584);
or U5305 (N_5305,N_4362,N_4588);
or U5306 (N_5306,N_4975,N_4124);
and U5307 (N_5307,N_4993,N_4201);
nand U5308 (N_5308,N_4353,N_4153);
and U5309 (N_5309,N_4400,N_4657);
xor U5310 (N_5310,N_4738,N_4526);
nor U5311 (N_5311,N_4171,N_4725);
nor U5312 (N_5312,N_4835,N_4055);
nand U5313 (N_5313,N_4219,N_4916);
nor U5314 (N_5314,N_4047,N_4691);
nor U5315 (N_5315,N_4271,N_4398);
or U5316 (N_5316,N_4252,N_4531);
and U5317 (N_5317,N_4405,N_4131);
nand U5318 (N_5318,N_4506,N_4750);
xor U5319 (N_5319,N_4310,N_4872);
nor U5320 (N_5320,N_4769,N_4021);
nand U5321 (N_5321,N_4366,N_4132);
nand U5322 (N_5322,N_4638,N_4861);
or U5323 (N_5323,N_4340,N_4656);
nand U5324 (N_5324,N_4462,N_4106);
nand U5325 (N_5325,N_4719,N_4614);
and U5326 (N_5326,N_4669,N_4984);
and U5327 (N_5327,N_4651,N_4910);
nor U5328 (N_5328,N_4649,N_4561);
and U5329 (N_5329,N_4440,N_4936);
and U5330 (N_5330,N_4410,N_4579);
or U5331 (N_5331,N_4547,N_4906);
nor U5332 (N_5332,N_4004,N_4655);
and U5333 (N_5333,N_4163,N_4681);
or U5334 (N_5334,N_4116,N_4949);
or U5335 (N_5335,N_4337,N_4152);
nand U5336 (N_5336,N_4473,N_4468);
nor U5337 (N_5337,N_4018,N_4794);
and U5338 (N_5338,N_4650,N_4545);
nand U5339 (N_5339,N_4285,N_4194);
xnor U5340 (N_5340,N_4036,N_4653);
xor U5341 (N_5341,N_4917,N_4558);
and U5342 (N_5342,N_4274,N_4385);
or U5343 (N_5343,N_4272,N_4006);
and U5344 (N_5344,N_4918,N_4213);
nor U5345 (N_5345,N_4809,N_4061);
and U5346 (N_5346,N_4528,N_4974);
and U5347 (N_5347,N_4148,N_4336);
nor U5348 (N_5348,N_4914,N_4320);
or U5349 (N_5349,N_4225,N_4265);
nand U5350 (N_5350,N_4598,N_4081);
and U5351 (N_5351,N_4812,N_4289);
nor U5352 (N_5352,N_4286,N_4956);
or U5353 (N_5353,N_4971,N_4663);
or U5354 (N_5354,N_4097,N_4409);
and U5355 (N_5355,N_4109,N_4330);
or U5356 (N_5356,N_4339,N_4276);
nand U5357 (N_5357,N_4226,N_4238);
and U5358 (N_5358,N_4732,N_4086);
nor U5359 (N_5359,N_4664,N_4426);
nor U5360 (N_5360,N_4815,N_4080);
and U5361 (N_5361,N_4392,N_4935);
nor U5362 (N_5362,N_4443,N_4636);
nor U5363 (N_5363,N_4839,N_4075);
nor U5364 (N_5364,N_4262,N_4490);
nor U5365 (N_5365,N_4920,N_4850);
nor U5366 (N_5366,N_4447,N_4486);
nand U5367 (N_5367,N_4466,N_4721);
and U5368 (N_5368,N_4452,N_4261);
nor U5369 (N_5369,N_4482,N_4487);
nor U5370 (N_5370,N_4856,N_4637);
and U5371 (N_5371,N_4787,N_4827);
or U5372 (N_5372,N_4045,N_4820);
nor U5373 (N_5373,N_4347,N_4989);
nor U5374 (N_5374,N_4500,N_4242);
nand U5375 (N_5375,N_4912,N_4934);
xnor U5376 (N_5376,N_4610,N_4355);
or U5377 (N_5377,N_4259,N_4001);
and U5378 (N_5378,N_4439,N_4563);
nand U5379 (N_5379,N_4641,N_4520);
nand U5380 (N_5380,N_4258,N_4849);
nor U5381 (N_5381,N_4549,N_4938);
and U5382 (N_5382,N_4778,N_4229);
xor U5383 (N_5383,N_4793,N_4396);
nor U5384 (N_5384,N_4726,N_4929);
nand U5385 (N_5385,N_4475,N_4921);
and U5386 (N_5386,N_4930,N_4307);
nor U5387 (N_5387,N_4123,N_4043);
nor U5388 (N_5388,N_4704,N_4554);
or U5389 (N_5389,N_4255,N_4739);
or U5390 (N_5390,N_4089,N_4742);
nand U5391 (N_5391,N_4496,N_4023);
nand U5392 (N_5392,N_4197,N_4015);
and U5393 (N_5393,N_4616,N_4896);
nor U5394 (N_5394,N_4214,N_4612);
nand U5395 (N_5395,N_4054,N_4884);
or U5396 (N_5396,N_4521,N_4349);
and U5397 (N_5397,N_4923,N_4592);
nand U5398 (N_5398,N_4516,N_4074);
nand U5399 (N_5399,N_4062,N_4757);
nand U5400 (N_5400,N_4484,N_4446);
nor U5401 (N_5401,N_4976,N_4193);
and U5402 (N_5402,N_4568,N_4786);
nor U5403 (N_5403,N_4263,N_4570);
xor U5404 (N_5404,N_4541,N_4341);
nand U5405 (N_5405,N_4119,N_4564);
nand U5406 (N_5406,N_4345,N_4014);
or U5407 (N_5407,N_4828,N_4647);
or U5408 (N_5408,N_4972,N_4371);
and U5409 (N_5409,N_4404,N_4205);
nand U5410 (N_5410,N_4714,N_4965);
nor U5411 (N_5411,N_4485,N_4053);
or U5412 (N_5412,N_4391,N_4143);
nand U5413 (N_5413,N_4494,N_4007);
and U5414 (N_5414,N_4764,N_4667);
or U5415 (N_5415,N_4275,N_4228);
and U5416 (N_5416,N_4088,N_4813);
nand U5417 (N_5417,N_4762,N_4288);
or U5418 (N_5418,N_4166,N_4065);
xnor U5419 (N_5419,N_4730,N_4666);
nand U5420 (N_5420,N_4529,N_4723);
nand U5421 (N_5421,N_4700,N_4013);
nand U5422 (N_5422,N_4665,N_4924);
or U5423 (N_5423,N_4931,N_4495);
nor U5424 (N_5424,N_4394,N_4780);
or U5425 (N_5425,N_4733,N_4978);
nand U5426 (N_5426,N_4689,N_4577);
xnor U5427 (N_5427,N_4617,N_4134);
nor U5428 (N_5428,N_4121,N_4668);
nand U5429 (N_5429,N_4291,N_4304);
or U5430 (N_5430,N_4626,N_4824);
or U5431 (N_5431,N_4419,N_4994);
and U5432 (N_5432,N_4172,N_4886);
nor U5433 (N_5433,N_4230,N_4044);
nand U5434 (N_5434,N_4125,N_4210);
and U5435 (N_5435,N_4449,N_4604);
nor U5436 (N_5436,N_4302,N_4505);
nor U5437 (N_5437,N_4455,N_4943);
and U5438 (N_5438,N_4108,N_4868);
and U5439 (N_5439,N_4969,N_4190);
nor U5440 (N_5440,N_4454,N_4266);
nand U5441 (N_5441,N_4059,N_4955);
or U5442 (N_5442,N_4783,N_4524);
nor U5443 (N_5443,N_4372,N_4361);
nor U5444 (N_5444,N_4151,N_4990);
nand U5445 (N_5445,N_4024,N_4292);
or U5446 (N_5446,N_4717,N_4504);
nor U5447 (N_5447,N_4502,N_4781);
xor U5448 (N_5448,N_4710,N_4629);
xnor U5449 (N_5449,N_4094,N_4694);
nor U5450 (N_5450,N_4633,N_4411);
and U5451 (N_5451,N_4642,N_4611);
and U5452 (N_5452,N_4060,N_4553);
or U5453 (N_5453,N_4542,N_4424);
nor U5454 (N_5454,N_4870,N_4548);
or U5455 (N_5455,N_4133,N_4671);
xnor U5456 (N_5456,N_4603,N_4318);
nor U5457 (N_5457,N_4512,N_4107);
or U5458 (N_5458,N_4509,N_4537);
nand U5459 (N_5459,N_4268,N_4096);
and U5460 (N_5460,N_4625,N_4231);
nor U5461 (N_5461,N_4908,N_4117);
or U5462 (N_5462,N_4992,N_4222);
and U5463 (N_5463,N_4804,N_4871);
and U5464 (N_5464,N_4685,N_4051);
and U5465 (N_5465,N_4199,N_4688);
nand U5466 (N_5466,N_4697,N_4580);
and U5467 (N_5467,N_4434,N_4066);
and U5468 (N_5468,N_4179,N_4593);
nand U5469 (N_5469,N_4848,N_4032);
nor U5470 (N_5470,N_4659,N_4817);
nand U5471 (N_5471,N_4388,N_4678);
nor U5472 (N_5472,N_4092,N_4801);
xor U5473 (N_5473,N_4519,N_4477);
nand U5474 (N_5474,N_4761,N_4251);
nand U5475 (N_5475,N_4606,N_4237);
and U5476 (N_5476,N_4209,N_4031);
nor U5477 (N_5477,N_4416,N_4898);
xor U5478 (N_5478,N_4515,N_4597);
nor U5479 (N_5479,N_4478,N_4328);
nor U5480 (N_5480,N_4393,N_4011);
and U5481 (N_5481,N_4899,N_4677);
nor U5482 (N_5482,N_4459,N_4634);
or U5483 (N_5483,N_4348,N_4756);
or U5484 (N_5484,N_4798,N_4408);
nor U5485 (N_5485,N_4273,N_4356);
xor U5486 (N_5486,N_4162,N_4645);
nor U5487 (N_5487,N_4435,N_4177);
or U5488 (N_5488,N_4135,N_4033);
or U5489 (N_5489,N_4415,N_4068);
and U5490 (N_5490,N_4796,N_4643);
or U5491 (N_5491,N_4881,N_4196);
and U5492 (N_5492,N_4102,N_4073);
nor U5493 (N_5493,N_4948,N_4038);
xnor U5494 (N_5494,N_4413,N_4843);
nand U5495 (N_5495,N_4855,N_4648);
and U5496 (N_5496,N_4050,N_4845);
nor U5497 (N_5497,N_4741,N_4159);
nand U5498 (N_5498,N_4365,N_4052);
and U5499 (N_5499,N_4425,N_4105);
xor U5500 (N_5500,N_4788,N_4070);
and U5501 (N_5501,N_4403,N_4364);
or U5502 (N_5502,N_4617,N_4360);
nand U5503 (N_5503,N_4137,N_4855);
nor U5504 (N_5504,N_4551,N_4212);
xnor U5505 (N_5505,N_4272,N_4890);
and U5506 (N_5506,N_4481,N_4131);
or U5507 (N_5507,N_4493,N_4572);
and U5508 (N_5508,N_4310,N_4964);
xnor U5509 (N_5509,N_4213,N_4104);
nor U5510 (N_5510,N_4617,N_4098);
nand U5511 (N_5511,N_4393,N_4786);
xnor U5512 (N_5512,N_4601,N_4763);
and U5513 (N_5513,N_4613,N_4025);
nor U5514 (N_5514,N_4290,N_4183);
and U5515 (N_5515,N_4399,N_4682);
or U5516 (N_5516,N_4259,N_4438);
xor U5517 (N_5517,N_4824,N_4996);
nor U5518 (N_5518,N_4803,N_4719);
nor U5519 (N_5519,N_4916,N_4942);
nand U5520 (N_5520,N_4633,N_4486);
and U5521 (N_5521,N_4520,N_4327);
nor U5522 (N_5522,N_4615,N_4758);
nand U5523 (N_5523,N_4302,N_4878);
or U5524 (N_5524,N_4009,N_4335);
xnor U5525 (N_5525,N_4778,N_4342);
nand U5526 (N_5526,N_4367,N_4947);
nor U5527 (N_5527,N_4174,N_4874);
nand U5528 (N_5528,N_4041,N_4479);
or U5529 (N_5529,N_4547,N_4176);
or U5530 (N_5530,N_4662,N_4289);
nor U5531 (N_5531,N_4139,N_4270);
xnor U5532 (N_5532,N_4342,N_4590);
nor U5533 (N_5533,N_4344,N_4094);
xnor U5534 (N_5534,N_4636,N_4204);
and U5535 (N_5535,N_4043,N_4984);
xnor U5536 (N_5536,N_4636,N_4460);
and U5537 (N_5537,N_4173,N_4795);
and U5538 (N_5538,N_4416,N_4366);
or U5539 (N_5539,N_4846,N_4601);
or U5540 (N_5540,N_4713,N_4069);
or U5541 (N_5541,N_4408,N_4760);
xor U5542 (N_5542,N_4080,N_4670);
nand U5543 (N_5543,N_4565,N_4864);
nor U5544 (N_5544,N_4027,N_4091);
nand U5545 (N_5545,N_4919,N_4741);
nor U5546 (N_5546,N_4970,N_4882);
and U5547 (N_5547,N_4337,N_4623);
nor U5548 (N_5548,N_4520,N_4730);
nand U5549 (N_5549,N_4165,N_4462);
or U5550 (N_5550,N_4086,N_4017);
and U5551 (N_5551,N_4576,N_4651);
or U5552 (N_5552,N_4576,N_4488);
xor U5553 (N_5553,N_4315,N_4331);
or U5554 (N_5554,N_4066,N_4908);
xnor U5555 (N_5555,N_4425,N_4947);
nand U5556 (N_5556,N_4745,N_4741);
xnor U5557 (N_5557,N_4118,N_4986);
and U5558 (N_5558,N_4059,N_4954);
nand U5559 (N_5559,N_4770,N_4399);
and U5560 (N_5560,N_4587,N_4305);
or U5561 (N_5561,N_4182,N_4966);
nor U5562 (N_5562,N_4773,N_4386);
nor U5563 (N_5563,N_4247,N_4423);
nand U5564 (N_5564,N_4274,N_4982);
or U5565 (N_5565,N_4721,N_4835);
xor U5566 (N_5566,N_4190,N_4757);
and U5567 (N_5567,N_4932,N_4802);
xnor U5568 (N_5568,N_4374,N_4878);
or U5569 (N_5569,N_4369,N_4227);
or U5570 (N_5570,N_4579,N_4528);
nand U5571 (N_5571,N_4652,N_4824);
nor U5572 (N_5572,N_4159,N_4612);
nand U5573 (N_5573,N_4420,N_4650);
nand U5574 (N_5574,N_4467,N_4617);
or U5575 (N_5575,N_4172,N_4047);
xor U5576 (N_5576,N_4144,N_4167);
or U5577 (N_5577,N_4516,N_4284);
or U5578 (N_5578,N_4488,N_4670);
and U5579 (N_5579,N_4157,N_4388);
nand U5580 (N_5580,N_4862,N_4953);
xnor U5581 (N_5581,N_4071,N_4516);
nand U5582 (N_5582,N_4230,N_4323);
nor U5583 (N_5583,N_4721,N_4981);
and U5584 (N_5584,N_4867,N_4148);
nor U5585 (N_5585,N_4590,N_4568);
xor U5586 (N_5586,N_4052,N_4906);
or U5587 (N_5587,N_4517,N_4248);
and U5588 (N_5588,N_4018,N_4037);
or U5589 (N_5589,N_4912,N_4054);
and U5590 (N_5590,N_4458,N_4000);
and U5591 (N_5591,N_4284,N_4491);
nor U5592 (N_5592,N_4710,N_4034);
or U5593 (N_5593,N_4044,N_4278);
nand U5594 (N_5594,N_4431,N_4542);
nor U5595 (N_5595,N_4781,N_4219);
and U5596 (N_5596,N_4289,N_4496);
xor U5597 (N_5597,N_4976,N_4404);
and U5598 (N_5598,N_4487,N_4747);
or U5599 (N_5599,N_4402,N_4815);
and U5600 (N_5600,N_4774,N_4895);
nor U5601 (N_5601,N_4066,N_4425);
and U5602 (N_5602,N_4321,N_4868);
or U5603 (N_5603,N_4031,N_4659);
and U5604 (N_5604,N_4828,N_4105);
and U5605 (N_5605,N_4532,N_4949);
xnor U5606 (N_5606,N_4369,N_4091);
xnor U5607 (N_5607,N_4316,N_4792);
nand U5608 (N_5608,N_4706,N_4377);
or U5609 (N_5609,N_4189,N_4328);
nand U5610 (N_5610,N_4157,N_4929);
and U5611 (N_5611,N_4723,N_4784);
and U5612 (N_5612,N_4894,N_4610);
and U5613 (N_5613,N_4540,N_4034);
xor U5614 (N_5614,N_4506,N_4624);
nand U5615 (N_5615,N_4315,N_4946);
nand U5616 (N_5616,N_4804,N_4824);
nand U5617 (N_5617,N_4089,N_4064);
or U5618 (N_5618,N_4066,N_4144);
and U5619 (N_5619,N_4141,N_4146);
nand U5620 (N_5620,N_4777,N_4758);
and U5621 (N_5621,N_4482,N_4391);
nor U5622 (N_5622,N_4889,N_4517);
nand U5623 (N_5623,N_4686,N_4570);
nor U5624 (N_5624,N_4052,N_4583);
nand U5625 (N_5625,N_4389,N_4471);
or U5626 (N_5626,N_4957,N_4885);
xnor U5627 (N_5627,N_4331,N_4623);
xor U5628 (N_5628,N_4538,N_4966);
and U5629 (N_5629,N_4617,N_4558);
nand U5630 (N_5630,N_4580,N_4620);
nand U5631 (N_5631,N_4701,N_4295);
xor U5632 (N_5632,N_4821,N_4255);
or U5633 (N_5633,N_4582,N_4837);
or U5634 (N_5634,N_4859,N_4352);
nor U5635 (N_5635,N_4896,N_4068);
and U5636 (N_5636,N_4327,N_4419);
nor U5637 (N_5637,N_4096,N_4078);
or U5638 (N_5638,N_4110,N_4872);
and U5639 (N_5639,N_4277,N_4151);
xor U5640 (N_5640,N_4177,N_4989);
or U5641 (N_5641,N_4912,N_4832);
xor U5642 (N_5642,N_4622,N_4015);
or U5643 (N_5643,N_4391,N_4234);
nand U5644 (N_5644,N_4023,N_4032);
nor U5645 (N_5645,N_4714,N_4928);
nor U5646 (N_5646,N_4896,N_4333);
or U5647 (N_5647,N_4421,N_4681);
nor U5648 (N_5648,N_4932,N_4797);
or U5649 (N_5649,N_4006,N_4967);
nand U5650 (N_5650,N_4627,N_4655);
and U5651 (N_5651,N_4586,N_4731);
and U5652 (N_5652,N_4296,N_4483);
nor U5653 (N_5653,N_4623,N_4325);
and U5654 (N_5654,N_4480,N_4922);
nor U5655 (N_5655,N_4229,N_4513);
nor U5656 (N_5656,N_4050,N_4211);
nand U5657 (N_5657,N_4039,N_4262);
nand U5658 (N_5658,N_4012,N_4796);
nand U5659 (N_5659,N_4699,N_4513);
and U5660 (N_5660,N_4297,N_4271);
nor U5661 (N_5661,N_4228,N_4464);
nor U5662 (N_5662,N_4449,N_4862);
xnor U5663 (N_5663,N_4823,N_4599);
or U5664 (N_5664,N_4082,N_4540);
or U5665 (N_5665,N_4854,N_4362);
xnor U5666 (N_5666,N_4264,N_4145);
and U5667 (N_5667,N_4850,N_4368);
xnor U5668 (N_5668,N_4028,N_4886);
nand U5669 (N_5669,N_4405,N_4177);
nor U5670 (N_5670,N_4803,N_4118);
or U5671 (N_5671,N_4996,N_4592);
xnor U5672 (N_5672,N_4798,N_4239);
xnor U5673 (N_5673,N_4986,N_4122);
or U5674 (N_5674,N_4794,N_4645);
nor U5675 (N_5675,N_4649,N_4104);
nand U5676 (N_5676,N_4631,N_4086);
nor U5677 (N_5677,N_4389,N_4007);
nand U5678 (N_5678,N_4062,N_4477);
and U5679 (N_5679,N_4372,N_4171);
xnor U5680 (N_5680,N_4524,N_4267);
nand U5681 (N_5681,N_4291,N_4109);
nor U5682 (N_5682,N_4690,N_4251);
xor U5683 (N_5683,N_4127,N_4584);
nor U5684 (N_5684,N_4048,N_4328);
and U5685 (N_5685,N_4888,N_4327);
nand U5686 (N_5686,N_4377,N_4957);
nor U5687 (N_5687,N_4860,N_4748);
or U5688 (N_5688,N_4027,N_4973);
or U5689 (N_5689,N_4319,N_4521);
and U5690 (N_5690,N_4407,N_4124);
and U5691 (N_5691,N_4433,N_4413);
and U5692 (N_5692,N_4665,N_4271);
or U5693 (N_5693,N_4580,N_4531);
nand U5694 (N_5694,N_4745,N_4699);
xnor U5695 (N_5695,N_4990,N_4397);
nand U5696 (N_5696,N_4810,N_4890);
nand U5697 (N_5697,N_4194,N_4447);
xnor U5698 (N_5698,N_4893,N_4427);
nand U5699 (N_5699,N_4450,N_4108);
and U5700 (N_5700,N_4850,N_4337);
nand U5701 (N_5701,N_4244,N_4147);
nor U5702 (N_5702,N_4176,N_4123);
and U5703 (N_5703,N_4509,N_4047);
and U5704 (N_5704,N_4423,N_4078);
nor U5705 (N_5705,N_4354,N_4624);
nand U5706 (N_5706,N_4025,N_4469);
nand U5707 (N_5707,N_4434,N_4959);
nor U5708 (N_5708,N_4249,N_4623);
or U5709 (N_5709,N_4936,N_4221);
and U5710 (N_5710,N_4458,N_4467);
or U5711 (N_5711,N_4358,N_4974);
or U5712 (N_5712,N_4834,N_4717);
or U5713 (N_5713,N_4383,N_4648);
nor U5714 (N_5714,N_4040,N_4648);
nand U5715 (N_5715,N_4852,N_4158);
or U5716 (N_5716,N_4803,N_4706);
nor U5717 (N_5717,N_4469,N_4302);
or U5718 (N_5718,N_4073,N_4394);
and U5719 (N_5719,N_4021,N_4014);
and U5720 (N_5720,N_4592,N_4467);
or U5721 (N_5721,N_4170,N_4907);
nor U5722 (N_5722,N_4529,N_4731);
nand U5723 (N_5723,N_4945,N_4564);
nor U5724 (N_5724,N_4170,N_4333);
nor U5725 (N_5725,N_4694,N_4052);
and U5726 (N_5726,N_4061,N_4645);
xnor U5727 (N_5727,N_4210,N_4478);
nor U5728 (N_5728,N_4954,N_4383);
nand U5729 (N_5729,N_4078,N_4900);
xor U5730 (N_5730,N_4168,N_4839);
nor U5731 (N_5731,N_4659,N_4463);
and U5732 (N_5732,N_4778,N_4121);
or U5733 (N_5733,N_4803,N_4013);
and U5734 (N_5734,N_4618,N_4419);
nor U5735 (N_5735,N_4025,N_4169);
or U5736 (N_5736,N_4985,N_4756);
nand U5737 (N_5737,N_4476,N_4536);
and U5738 (N_5738,N_4516,N_4680);
or U5739 (N_5739,N_4870,N_4126);
nand U5740 (N_5740,N_4200,N_4327);
nand U5741 (N_5741,N_4619,N_4993);
or U5742 (N_5742,N_4720,N_4790);
nand U5743 (N_5743,N_4371,N_4432);
and U5744 (N_5744,N_4152,N_4891);
nand U5745 (N_5745,N_4822,N_4908);
and U5746 (N_5746,N_4461,N_4603);
or U5747 (N_5747,N_4237,N_4981);
nand U5748 (N_5748,N_4606,N_4282);
nand U5749 (N_5749,N_4573,N_4048);
or U5750 (N_5750,N_4019,N_4642);
and U5751 (N_5751,N_4358,N_4700);
nand U5752 (N_5752,N_4745,N_4651);
nor U5753 (N_5753,N_4788,N_4554);
and U5754 (N_5754,N_4916,N_4448);
nand U5755 (N_5755,N_4697,N_4280);
nand U5756 (N_5756,N_4912,N_4383);
nand U5757 (N_5757,N_4282,N_4967);
or U5758 (N_5758,N_4376,N_4824);
xor U5759 (N_5759,N_4195,N_4792);
nor U5760 (N_5760,N_4341,N_4221);
xnor U5761 (N_5761,N_4273,N_4607);
and U5762 (N_5762,N_4274,N_4600);
nand U5763 (N_5763,N_4980,N_4337);
or U5764 (N_5764,N_4647,N_4975);
nor U5765 (N_5765,N_4865,N_4875);
and U5766 (N_5766,N_4654,N_4305);
or U5767 (N_5767,N_4931,N_4189);
xor U5768 (N_5768,N_4339,N_4590);
nor U5769 (N_5769,N_4319,N_4190);
and U5770 (N_5770,N_4629,N_4972);
nand U5771 (N_5771,N_4827,N_4406);
nor U5772 (N_5772,N_4728,N_4614);
or U5773 (N_5773,N_4471,N_4781);
nand U5774 (N_5774,N_4277,N_4858);
and U5775 (N_5775,N_4218,N_4122);
or U5776 (N_5776,N_4885,N_4119);
or U5777 (N_5777,N_4187,N_4242);
xnor U5778 (N_5778,N_4089,N_4017);
nand U5779 (N_5779,N_4402,N_4733);
or U5780 (N_5780,N_4755,N_4413);
xnor U5781 (N_5781,N_4704,N_4339);
nand U5782 (N_5782,N_4726,N_4827);
nand U5783 (N_5783,N_4560,N_4228);
and U5784 (N_5784,N_4441,N_4272);
xnor U5785 (N_5785,N_4655,N_4371);
or U5786 (N_5786,N_4038,N_4494);
xnor U5787 (N_5787,N_4742,N_4074);
nand U5788 (N_5788,N_4515,N_4190);
nor U5789 (N_5789,N_4582,N_4984);
nand U5790 (N_5790,N_4124,N_4478);
nor U5791 (N_5791,N_4854,N_4113);
or U5792 (N_5792,N_4407,N_4806);
and U5793 (N_5793,N_4431,N_4386);
or U5794 (N_5794,N_4874,N_4161);
or U5795 (N_5795,N_4049,N_4361);
nand U5796 (N_5796,N_4402,N_4322);
nor U5797 (N_5797,N_4058,N_4865);
or U5798 (N_5798,N_4784,N_4566);
nor U5799 (N_5799,N_4178,N_4912);
and U5800 (N_5800,N_4069,N_4179);
nor U5801 (N_5801,N_4971,N_4823);
nor U5802 (N_5802,N_4795,N_4522);
or U5803 (N_5803,N_4467,N_4665);
or U5804 (N_5804,N_4617,N_4048);
xor U5805 (N_5805,N_4551,N_4561);
and U5806 (N_5806,N_4011,N_4376);
or U5807 (N_5807,N_4899,N_4747);
or U5808 (N_5808,N_4923,N_4682);
nand U5809 (N_5809,N_4046,N_4210);
or U5810 (N_5810,N_4600,N_4007);
nand U5811 (N_5811,N_4601,N_4398);
and U5812 (N_5812,N_4428,N_4722);
and U5813 (N_5813,N_4348,N_4969);
or U5814 (N_5814,N_4471,N_4095);
and U5815 (N_5815,N_4170,N_4338);
or U5816 (N_5816,N_4332,N_4130);
and U5817 (N_5817,N_4308,N_4856);
nor U5818 (N_5818,N_4865,N_4361);
and U5819 (N_5819,N_4062,N_4137);
or U5820 (N_5820,N_4688,N_4270);
xor U5821 (N_5821,N_4051,N_4617);
nand U5822 (N_5822,N_4906,N_4874);
and U5823 (N_5823,N_4675,N_4918);
nor U5824 (N_5824,N_4050,N_4064);
nor U5825 (N_5825,N_4237,N_4449);
or U5826 (N_5826,N_4444,N_4985);
nor U5827 (N_5827,N_4266,N_4840);
xnor U5828 (N_5828,N_4666,N_4718);
nor U5829 (N_5829,N_4016,N_4601);
and U5830 (N_5830,N_4161,N_4708);
or U5831 (N_5831,N_4968,N_4838);
nor U5832 (N_5832,N_4694,N_4682);
nand U5833 (N_5833,N_4220,N_4564);
nand U5834 (N_5834,N_4834,N_4046);
nand U5835 (N_5835,N_4398,N_4623);
or U5836 (N_5836,N_4155,N_4486);
or U5837 (N_5837,N_4148,N_4714);
and U5838 (N_5838,N_4151,N_4705);
or U5839 (N_5839,N_4648,N_4512);
nor U5840 (N_5840,N_4365,N_4346);
nand U5841 (N_5841,N_4646,N_4373);
nor U5842 (N_5842,N_4126,N_4443);
nand U5843 (N_5843,N_4995,N_4086);
xor U5844 (N_5844,N_4435,N_4728);
or U5845 (N_5845,N_4369,N_4202);
or U5846 (N_5846,N_4145,N_4532);
nor U5847 (N_5847,N_4829,N_4401);
nand U5848 (N_5848,N_4390,N_4089);
nor U5849 (N_5849,N_4084,N_4786);
and U5850 (N_5850,N_4225,N_4982);
nor U5851 (N_5851,N_4896,N_4889);
nor U5852 (N_5852,N_4721,N_4400);
nor U5853 (N_5853,N_4189,N_4200);
xnor U5854 (N_5854,N_4523,N_4940);
or U5855 (N_5855,N_4075,N_4031);
or U5856 (N_5856,N_4539,N_4800);
nand U5857 (N_5857,N_4512,N_4328);
nand U5858 (N_5858,N_4281,N_4584);
nor U5859 (N_5859,N_4567,N_4746);
and U5860 (N_5860,N_4789,N_4817);
or U5861 (N_5861,N_4348,N_4060);
xor U5862 (N_5862,N_4145,N_4682);
and U5863 (N_5863,N_4388,N_4796);
or U5864 (N_5864,N_4744,N_4812);
or U5865 (N_5865,N_4121,N_4028);
and U5866 (N_5866,N_4855,N_4397);
nand U5867 (N_5867,N_4451,N_4149);
nand U5868 (N_5868,N_4314,N_4322);
nor U5869 (N_5869,N_4642,N_4739);
nand U5870 (N_5870,N_4061,N_4767);
and U5871 (N_5871,N_4291,N_4590);
nor U5872 (N_5872,N_4351,N_4525);
or U5873 (N_5873,N_4534,N_4095);
and U5874 (N_5874,N_4481,N_4550);
and U5875 (N_5875,N_4614,N_4302);
nand U5876 (N_5876,N_4076,N_4062);
nor U5877 (N_5877,N_4119,N_4741);
and U5878 (N_5878,N_4706,N_4997);
nor U5879 (N_5879,N_4960,N_4766);
and U5880 (N_5880,N_4618,N_4978);
xnor U5881 (N_5881,N_4279,N_4995);
xnor U5882 (N_5882,N_4835,N_4145);
nand U5883 (N_5883,N_4137,N_4407);
nor U5884 (N_5884,N_4323,N_4446);
nand U5885 (N_5885,N_4509,N_4905);
nor U5886 (N_5886,N_4437,N_4578);
nand U5887 (N_5887,N_4563,N_4551);
and U5888 (N_5888,N_4961,N_4024);
nand U5889 (N_5889,N_4809,N_4814);
nor U5890 (N_5890,N_4850,N_4633);
nand U5891 (N_5891,N_4122,N_4483);
nor U5892 (N_5892,N_4882,N_4545);
nand U5893 (N_5893,N_4742,N_4300);
or U5894 (N_5894,N_4593,N_4241);
nand U5895 (N_5895,N_4127,N_4433);
and U5896 (N_5896,N_4394,N_4669);
xnor U5897 (N_5897,N_4226,N_4417);
and U5898 (N_5898,N_4512,N_4919);
and U5899 (N_5899,N_4779,N_4179);
xnor U5900 (N_5900,N_4527,N_4916);
nand U5901 (N_5901,N_4236,N_4213);
nor U5902 (N_5902,N_4740,N_4658);
nand U5903 (N_5903,N_4491,N_4648);
or U5904 (N_5904,N_4666,N_4468);
and U5905 (N_5905,N_4842,N_4659);
or U5906 (N_5906,N_4182,N_4159);
nand U5907 (N_5907,N_4105,N_4637);
xnor U5908 (N_5908,N_4823,N_4154);
nor U5909 (N_5909,N_4325,N_4798);
nor U5910 (N_5910,N_4451,N_4932);
nand U5911 (N_5911,N_4201,N_4318);
xor U5912 (N_5912,N_4345,N_4110);
and U5913 (N_5913,N_4906,N_4145);
and U5914 (N_5914,N_4257,N_4595);
and U5915 (N_5915,N_4068,N_4192);
nor U5916 (N_5916,N_4572,N_4539);
nor U5917 (N_5917,N_4750,N_4118);
or U5918 (N_5918,N_4038,N_4650);
and U5919 (N_5919,N_4771,N_4052);
nand U5920 (N_5920,N_4219,N_4037);
nor U5921 (N_5921,N_4315,N_4430);
nor U5922 (N_5922,N_4354,N_4117);
nor U5923 (N_5923,N_4071,N_4667);
nor U5924 (N_5924,N_4127,N_4785);
nor U5925 (N_5925,N_4898,N_4473);
nand U5926 (N_5926,N_4831,N_4006);
xor U5927 (N_5927,N_4185,N_4033);
xnor U5928 (N_5928,N_4698,N_4816);
nand U5929 (N_5929,N_4370,N_4867);
or U5930 (N_5930,N_4557,N_4215);
nand U5931 (N_5931,N_4456,N_4235);
nor U5932 (N_5932,N_4429,N_4200);
and U5933 (N_5933,N_4034,N_4188);
nor U5934 (N_5934,N_4038,N_4029);
or U5935 (N_5935,N_4645,N_4859);
xor U5936 (N_5936,N_4388,N_4265);
or U5937 (N_5937,N_4306,N_4069);
xor U5938 (N_5938,N_4541,N_4621);
nand U5939 (N_5939,N_4220,N_4461);
and U5940 (N_5940,N_4061,N_4094);
nand U5941 (N_5941,N_4372,N_4824);
and U5942 (N_5942,N_4727,N_4106);
nor U5943 (N_5943,N_4789,N_4678);
nand U5944 (N_5944,N_4336,N_4491);
nor U5945 (N_5945,N_4784,N_4146);
nand U5946 (N_5946,N_4559,N_4166);
nand U5947 (N_5947,N_4188,N_4298);
nor U5948 (N_5948,N_4353,N_4974);
nand U5949 (N_5949,N_4794,N_4623);
or U5950 (N_5950,N_4563,N_4150);
and U5951 (N_5951,N_4089,N_4671);
and U5952 (N_5952,N_4581,N_4875);
or U5953 (N_5953,N_4874,N_4060);
xor U5954 (N_5954,N_4609,N_4549);
and U5955 (N_5955,N_4656,N_4347);
and U5956 (N_5956,N_4632,N_4324);
nor U5957 (N_5957,N_4151,N_4443);
xor U5958 (N_5958,N_4495,N_4829);
nand U5959 (N_5959,N_4228,N_4060);
and U5960 (N_5960,N_4897,N_4622);
nand U5961 (N_5961,N_4508,N_4359);
nor U5962 (N_5962,N_4683,N_4414);
and U5963 (N_5963,N_4848,N_4150);
or U5964 (N_5964,N_4706,N_4769);
and U5965 (N_5965,N_4340,N_4502);
xor U5966 (N_5966,N_4822,N_4475);
xor U5967 (N_5967,N_4744,N_4444);
nor U5968 (N_5968,N_4554,N_4209);
or U5969 (N_5969,N_4743,N_4734);
or U5970 (N_5970,N_4771,N_4673);
nor U5971 (N_5971,N_4373,N_4991);
or U5972 (N_5972,N_4616,N_4998);
or U5973 (N_5973,N_4299,N_4325);
nor U5974 (N_5974,N_4815,N_4678);
nor U5975 (N_5975,N_4316,N_4219);
or U5976 (N_5976,N_4687,N_4560);
xor U5977 (N_5977,N_4620,N_4308);
and U5978 (N_5978,N_4372,N_4901);
or U5979 (N_5979,N_4472,N_4585);
xnor U5980 (N_5980,N_4177,N_4747);
nand U5981 (N_5981,N_4880,N_4111);
xnor U5982 (N_5982,N_4131,N_4355);
and U5983 (N_5983,N_4609,N_4696);
or U5984 (N_5984,N_4022,N_4757);
or U5985 (N_5985,N_4243,N_4287);
or U5986 (N_5986,N_4371,N_4940);
nor U5987 (N_5987,N_4848,N_4134);
nor U5988 (N_5988,N_4876,N_4439);
and U5989 (N_5989,N_4188,N_4343);
nor U5990 (N_5990,N_4948,N_4416);
xnor U5991 (N_5991,N_4429,N_4678);
xor U5992 (N_5992,N_4796,N_4520);
and U5993 (N_5993,N_4608,N_4544);
or U5994 (N_5994,N_4229,N_4288);
nand U5995 (N_5995,N_4353,N_4272);
or U5996 (N_5996,N_4260,N_4490);
nor U5997 (N_5997,N_4713,N_4006);
nor U5998 (N_5998,N_4498,N_4082);
nand U5999 (N_5999,N_4758,N_4305);
nand U6000 (N_6000,N_5591,N_5103);
and U6001 (N_6001,N_5886,N_5534);
and U6002 (N_6002,N_5795,N_5529);
nor U6003 (N_6003,N_5739,N_5492);
xnor U6004 (N_6004,N_5349,N_5320);
nor U6005 (N_6005,N_5404,N_5427);
nand U6006 (N_6006,N_5242,N_5636);
and U6007 (N_6007,N_5957,N_5179);
and U6008 (N_6008,N_5050,N_5025);
nand U6009 (N_6009,N_5020,N_5912);
nand U6010 (N_6010,N_5840,N_5006);
nand U6011 (N_6011,N_5546,N_5657);
or U6012 (N_6012,N_5641,N_5462);
or U6013 (N_6013,N_5222,N_5350);
nand U6014 (N_6014,N_5868,N_5112);
nor U6015 (N_6015,N_5152,N_5576);
and U6016 (N_6016,N_5519,N_5361);
and U6017 (N_6017,N_5642,N_5022);
and U6018 (N_6018,N_5769,N_5544);
nor U6019 (N_6019,N_5786,N_5168);
xnor U6020 (N_6020,N_5843,N_5167);
or U6021 (N_6021,N_5805,N_5719);
nand U6022 (N_6022,N_5144,N_5091);
nand U6023 (N_6023,N_5881,N_5558);
or U6024 (N_6024,N_5491,N_5667);
and U6025 (N_6025,N_5720,N_5663);
and U6026 (N_6026,N_5696,N_5594);
or U6027 (N_6027,N_5999,N_5151);
and U6028 (N_6028,N_5851,N_5804);
and U6029 (N_6029,N_5631,N_5753);
nand U6030 (N_6030,N_5467,N_5056);
nand U6031 (N_6031,N_5426,N_5824);
xnor U6032 (N_6032,N_5399,N_5400);
and U6033 (N_6033,N_5441,N_5428);
and U6034 (N_6034,N_5549,N_5319);
and U6035 (N_6035,N_5405,N_5950);
or U6036 (N_6036,N_5872,N_5810);
nor U6037 (N_6037,N_5601,N_5045);
nor U6038 (N_6038,N_5928,N_5030);
and U6039 (N_6039,N_5272,N_5058);
or U6040 (N_6040,N_5187,N_5785);
or U6041 (N_6041,N_5311,N_5789);
and U6042 (N_6042,N_5722,N_5488);
and U6043 (N_6043,N_5165,N_5575);
nor U6044 (N_6044,N_5634,N_5163);
nand U6045 (N_6045,N_5962,N_5891);
or U6046 (N_6046,N_5147,N_5260);
nor U6047 (N_6047,N_5371,N_5816);
and U6048 (N_6048,N_5509,N_5172);
nor U6049 (N_6049,N_5264,N_5117);
nor U6050 (N_6050,N_5366,N_5827);
and U6051 (N_6051,N_5628,N_5666);
xor U6052 (N_6052,N_5969,N_5880);
nand U6053 (N_6053,N_5624,N_5815);
or U6054 (N_6054,N_5162,N_5286);
nor U6055 (N_6055,N_5934,N_5439);
and U6056 (N_6056,N_5487,N_5894);
nand U6057 (N_6057,N_5126,N_5166);
or U6058 (N_6058,N_5976,N_5330);
nor U6059 (N_6059,N_5185,N_5751);
xor U6060 (N_6060,N_5215,N_5563);
and U6061 (N_6061,N_5143,N_5502);
nor U6062 (N_6062,N_5196,N_5859);
nand U6063 (N_6063,N_5714,N_5858);
or U6064 (N_6064,N_5532,N_5271);
nor U6065 (N_6065,N_5246,N_5370);
or U6066 (N_6066,N_5908,N_5567);
nand U6067 (N_6067,N_5228,N_5718);
nor U6068 (N_6068,N_5302,N_5472);
or U6069 (N_6069,N_5064,N_5335);
and U6070 (N_6070,N_5105,N_5750);
nor U6071 (N_6071,N_5277,N_5419);
nor U6072 (N_6072,N_5903,N_5229);
and U6073 (N_6073,N_5063,N_5687);
and U6074 (N_6074,N_5692,N_5807);
nor U6075 (N_6075,N_5744,N_5884);
nor U6076 (N_6076,N_5792,N_5516);
or U6077 (N_6077,N_5447,N_5520);
xnor U6078 (N_6078,N_5240,N_5153);
nor U6079 (N_6079,N_5609,N_5398);
xor U6080 (N_6080,N_5086,N_5579);
nand U6081 (N_6081,N_5885,N_5620);
nor U6082 (N_6082,N_5643,N_5759);
nand U6083 (N_6083,N_5026,N_5413);
and U6084 (N_6084,N_5363,N_5263);
nor U6085 (N_6085,N_5616,N_5721);
and U6086 (N_6086,N_5497,N_5300);
nor U6087 (N_6087,N_5498,N_5604);
nor U6088 (N_6088,N_5675,N_5446);
nor U6089 (N_6089,N_5774,N_5844);
nor U6090 (N_6090,N_5464,N_5727);
or U6091 (N_6091,N_5775,N_5932);
and U6092 (N_6092,N_5474,N_5925);
xor U6093 (N_6093,N_5809,N_5205);
nor U6094 (N_6094,N_5640,N_5996);
or U6095 (N_6095,N_5638,N_5612);
xor U6096 (N_6096,N_5997,N_5541);
nor U6097 (N_6097,N_5777,N_5623);
and U6098 (N_6098,N_5084,N_5926);
nand U6099 (N_6099,N_5128,N_5494);
nor U6100 (N_6100,N_5918,N_5290);
or U6101 (N_6101,N_5647,N_5160);
nor U6102 (N_6102,N_5417,N_5983);
and U6103 (N_6103,N_5731,N_5995);
nor U6104 (N_6104,N_5883,N_5676);
and U6105 (N_6105,N_5923,N_5099);
nand U6106 (N_6106,N_5372,N_5632);
and U6107 (N_6107,N_5454,N_5104);
nor U6108 (N_6108,N_5629,N_5814);
and U6109 (N_6109,N_5208,N_5289);
nand U6110 (N_6110,N_5484,N_5113);
xor U6111 (N_6111,N_5946,N_5724);
or U6112 (N_6112,N_5501,N_5080);
nand U6113 (N_6113,N_5390,N_5040);
nor U6114 (N_6114,N_5414,N_5314);
and U6115 (N_6115,N_5012,N_5075);
or U6116 (N_6116,N_5793,N_5929);
nand U6117 (N_6117,N_5955,N_5452);
xor U6118 (N_6118,N_5115,N_5834);
nand U6119 (N_6119,N_5017,N_5737);
and U6120 (N_6120,N_5486,N_5967);
nor U6121 (N_6121,N_5280,N_5244);
and U6122 (N_6122,N_5085,N_5703);
nor U6123 (N_6123,N_5865,N_5161);
or U6124 (N_6124,N_5791,N_5965);
nor U6125 (N_6125,N_5735,N_5583);
nor U6126 (N_6126,N_5867,N_5566);
and U6127 (N_6127,N_5038,N_5057);
and U6128 (N_6128,N_5909,N_5922);
nand U6129 (N_6129,N_5433,N_5819);
and U6130 (N_6130,N_5788,N_5557);
xnor U6131 (N_6131,N_5705,N_5312);
nor U6132 (N_6132,N_5811,N_5990);
or U6133 (N_6133,N_5619,N_5939);
nand U6134 (N_6134,N_5911,N_5268);
and U6135 (N_6135,N_5212,N_5145);
or U6136 (N_6136,N_5453,N_5537);
or U6137 (N_6137,N_5729,N_5987);
or U6138 (N_6138,N_5421,N_5364);
nor U6139 (N_6139,N_5917,N_5668);
or U6140 (N_6140,N_5087,N_5456);
or U6141 (N_6141,N_5373,N_5924);
and U6142 (N_6142,N_5307,N_5547);
nand U6143 (N_6143,N_5670,N_5748);
nand U6144 (N_6144,N_5961,N_5175);
nor U6145 (N_6145,N_5689,N_5321);
or U6146 (N_6146,N_5470,N_5071);
and U6147 (N_6147,N_5396,N_5561);
nand U6148 (N_6148,N_5651,N_5202);
nor U6149 (N_6149,N_5970,N_5968);
nand U6150 (N_6150,N_5513,N_5463);
nand U6151 (N_6151,N_5257,N_5344);
or U6152 (N_6152,N_5174,N_5232);
and U6153 (N_6153,N_5386,N_5897);
or U6154 (N_6154,N_5284,N_5008);
xor U6155 (N_6155,N_5083,N_5746);
nor U6156 (N_6156,N_5713,N_5424);
nor U6157 (N_6157,N_5481,N_5605);
xnor U6158 (N_6158,N_5322,N_5047);
or U6159 (N_6159,N_5381,N_5276);
nor U6160 (N_6160,N_5125,N_5102);
xnor U6161 (N_6161,N_5131,N_5402);
nand U6162 (N_6162,N_5921,N_5798);
nand U6163 (N_6163,N_5599,N_5028);
nand U6164 (N_6164,N_5830,N_5904);
or U6165 (N_6165,N_5051,N_5432);
and U6166 (N_6166,N_5587,N_5665);
nand U6167 (N_6167,N_5570,N_5796);
nand U6168 (N_6168,N_5833,N_5374);
xnor U6169 (N_6169,N_5565,N_5251);
xor U6170 (N_6170,N_5706,N_5096);
or U6171 (N_6171,N_5407,N_5613);
nor U6172 (N_6172,N_5140,N_5614);
and U6173 (N_6173,N_5707,N_5274);
xor U6174 (N_6174,N_5054,N_5150);
nand U6175 (N_6175,N_5820,N_5683);
and U6176 (N_6176,N_5773,N_5298);
and U6177 (N_6177,N_5496,N_5316);
nor U6178 (N_6178,N_5238,N_5979);
nor U6179 (N_6179,N_5233,N_5269);
nand U6180 (N_6180,N_5283,N_5677);
nor U6181 (N_6181,N_5226,N_5101);
or U6182 (N_6182,N_5986,N_5552);
nor U6183 (N_6183,N_5114,N_5449);
nand U6184 (N_6184,N_5896,N_5664);
nand U6185 (N_6185,N_5533,N_5031);
or U6186 (N_6186,N_5034,N_5392);
xor U6187 (N_6187,N_5653,N_5806);
and U6188 (N_6188,N_5313,N_5015);
and U6189 (N_6189,N_5383,N_5403);
nor U6190 (N_6190,N_5410,N_5148);
nor U6191 (N_6191,N_5935,N_5648);
and U6192 (N_6192,N_5985,N_5236);
or U6193 (N_6193,N_5483,N_5297);
nor U6194 (N_6194,N_5443,N_5507);
nor U6195 (N_6195,N_5137,N_5695);
xnor U6196 (N_6196,N_5401,N_5035);
nand U6197 (N_6197,N_5699,N_5182);
nand U6198 (N_6198,N_5243,N_5776);
or U6199 (N_6199,N_5517,N_5149);
and U6200 (N_6200,N_5645,N_5072);
nand U6201 (N_6201,N_5255,N_5018);
nand U6202 (N_6202,N_5480,N_5615);
nand U6203 (N_6203,N_5241,N_5756);
nor U6204 (N_6204,N_5237,N_5625);
or U6205 (N_6205,N_5523,N_5210);
xor U6206 (N_6206,N_5375,N_5134);
xor U6207 (N_6207,N_5438,N_5039);
or U6208 (N_6208,N_5138,N_5301);
nor U6209 (N_6209,N_5994,N_5078);
xor U6210 (N_6210,N_5581,N_5841);
or U6211 (N_6211,N_5948,N_5317);
nand U6212 (N_6212,N_5279,N_5697);
and U6213 (N_6213,N_5434,N_5879);
or U6214 (N_6214,N_5021,N_5393);
or U6215 (N_6215,N_5573,N_5649);
nor U6216 (N_6216,N_5036,N_5089);
or U6217 (N_6217,N_5338,N_5919);
or U6218 (N_6218,N_5678,N_5493);
xnor U6219 (N_6219,N_5914,N_5800);
or U6220 (N_6220,N_5329,N_5861);
and U6221 (N_6221,N_5192,N_5870);
xor U6222 (N_6222,N_5554,N_5963);
nor U6223 (N_6223,N_5808,N_5977);
xor U6224 (N_6224,N_5539,N_5589);
nand U6225 (N_6225,N_5133,N_5755);
nor U6226 (N_6226,N_5941,N_5551);
or U6227 (N_6227,N_5639,N_5460);
or U6228 (N_6228,N_5216,N_5906);
or U6229 (N_6229,N_5423,N_5180);
and U6230 (N_6230,N_5288,N_5770);
nand U6231 (N_6231,N_5817,N_5445);
nor U6232 (N_6232,N_5002,N_5309);
and U6233 (N_6233,N_5526,N_5760);
nor U6234 (N_6234,N_5450,N_5866);
nor U6235 (N_6235,N_5094,N_5875);
nor U6236 (N_6236,N_5082,N_5701);
nor U6237 (N_6237,N_5333,N_5754);
and U6238 (N_6238,N_5540,N_5876);
or U6239 (N_6239,N_5869,N_5448);
nand U6240 (N_6240,N_5409,N_5933);
nor U6241 (N_6241,N_5231,N_5521);
nor U6242 (N_6242,N_5690,N_5218);
nor U6243 (N_6243,N_5019,N_5042);
and U6244 (N_6244,N_5530,N_5440);
xnor U6245 (N_6245,N_5959,N_5013);
nand U6246 (N_6246,N_5170,N_5254);
nor U6247 (N_6247,N_5303,N_5674);
and U6248 (N_6248,N_5607,N_5525);
or U6249 (N_6249,N_5359,N_5097);
or U6250 (N_6250,N_5761,N_5331);
nand U6251 (N_6251,N_5499,N_5204);
or U6252 (N_6252,N_5074,N_5848);
and U6253 (N_6253,N_5458,N_5181);
or U6254 (N_6254,N_5693,N_5949);
nand U6255 (N_6255,N_5273,N_5387);
xnor U6256 (N_6256,N_5069,N_5700);
nor U6257 (N_6257,N_5295,N_5945);
and U6258 (N_6258,N_5466,N_5037);
or U6259 (N_6259,N_5459,N_5734);
and U6260 (N_6260,N_5076,N_5442);
and U6261 (N_6261,N_5016,N_5984);
or U6262 (N_6262,N_5790,N_5758);
nand U6263 (N_6263,N_5802,N_5553);
or U6264 (N_6264,N_5960,N_5650);
nand U6265 (N_6265,N_5477,N_5764);
xor U6266 (N_6266,N_5646,N_5818);
nand U6267 (N_6267,N_5262,N_5951);
or U6268 (N_6268,N_5577,N_5055);
nand U6269 (N_6269,N_5813,N_5473);
and U6270 (N_6270,N_5435,N_5412);
xnor U6271 (N_6271,N_5337,N_5489);
nor U6272 (N_6272,N_5200,N_5849);
or U6273 (N_6273,N_5888,N_5797);
nand U6274 (N_6274,N_5942,N_5654);
nor U6275 (N_6275,N_5588,N_5235);
or U6276 (N_6276,N_5053,N_5355);
nand U6277 (N_6277,N_5081,N_5169);
nand U6278 (N_6278,N_5468,N_5230);
nor U6279 (N_6279,N_5092,N_5415);
xnor U6280 (N_6280,N_5506,N_5562);
nor U6281 (N_6281,N_5304,N_5847);
nor U6282 (N_6282,N_5839,N_5377);
or U6283 (N_6283,N_5586,N_5061);
or U6284 (N_6284,N_5600,N_5451);
or U6285 (N_6285,N_5176,N_5457);
nor U6286 (N_6286,N_5902,N_5900);
nor U6287 (N_6287,N_5001,N_5173);
nor U6288 (N_6288,N_5004,N_5033);
nand U6289 (N_6289,N_5079,N_5568);
or U6290 (N_6290,N_5673,N_5384);
nand U6291 (N_6291,N_5211,N_5065);
and U6292 (N_6292,N_5278,N_5275);
or U6293 (N_6293,N_5005,N_5679);
and U6294 (N_6294,N_5669,N_5027);
nand U6295 (N_6295,N_5772,N_5191);
nor U6296 (N_6296,N_5156,N_5158);
nor U6297 (N_6297,N_5346,N_5937);
xnor U6298 (N_6298,N_5266,N_5771);
or U6299 (N_6299,N_5757,N_5093);
and U6300 (N_6300,N_5123,N_5512);
nand U6301 (N_6301,N_5365,N_5476);
or U6302 (N_6302,N_5854,N_5927);
xor U6303 (N_6303,N_5686,N_5340);
nand U6304 (N_6304,N_5555,N_5662);
and U6305 (N_6305,N_5048,N_5608);
xor U6306 (N_6306,N_5478,N_5837);
nand U6307 (N_6307,N_5610,N_5406);
nor U6308 (N_6308,N_5711,N_5318);
and U6309 (N_6309,N_5510,N_5622);
nor U6310 (N_6310,N_5991,N_5659);
and U6311 (N_6311,N_5936,N_5437);
nand U6312 (N_6312,N_5702,N_5907);
nand U6313 (N_6313,N_5611,N_5343);
nor U6314 (N_6314,N_5070,N_5766);
nand U6315 (N_6315,N_5245,N_5014);
and U6316 (N_6316,N_5627,N_5877);
and U6317 (N_6317,N_5598,N_5431);
or U6318 (N_6318,N_5716,N_5095);
nand U6319 (N_6319,N_5527,N_5603);
nor U6320 (N_6320,N_5305,N_5626);
and U6321 (N_6321,N_5342,N_5652);
nand U6322 (N_6322,N_5916,N_5726);
and U6323 (N_6323,N_5252,N_5195);
or U6324 (N_6324,N_5569,N_5832);
or U6325 (N_6325,N_5890,N_5709);
or U6326 (N_6326,N_5325,N_5154);
and U6327 (N_6327,N_5835,N_5436);
nand U6328 (N_6328,N_5857,N_5485);
and U6329 (N_6329,N_5124,N_5385);
nand U6330 (N_6330,N_5281,N_5127);
and U6331 (N_6331,N_5360,N_5339);
nand U6332 (N_6332,N_5024,N_5710);
or U6333 (N_6333,N_5862,N_5073);
or U6334 (N_6334,N_5972,N_5299);
or U6335 (N_6335,N_5362,N_5352);
and U6336 (N_6336,N_5119,N_5060);
or U6337 (N_6337,N_5068,N_5584);
nand U6338 (N_6338,N_5201,N_5511);
nor U6339 (N_6339,N_5618,N_5090);
and U6340 (N_6340,N_5253,N_5111);
and U6341 (N_6341,N_5762,N_5495);
nand U6342 (N_6342,N_5712,N_5787);
and U6343 (N_6343,N_5524,N_5188);
and U6344 (N_6344,N_5121,N_5285);
or U6345 (N_6345,N_5465,N_5256);
nor U6346 (N_6346,N_5429,N_5602);
and U6347 (N_6347,N_5422,N_5784);
or U6348 (N_6348,N_5100,N_5671);
nor U6349 (N_6349,N_5694,N_5077);
and U6350 (N_6350,N_5416,N_5590);
or U6351 (N_6351,N_5633,N_5873);
and U6352 (N_6352,N_5225,N_5864);
nand U6353 (N_6353,N_5556,N_5536);
nor U6354 (N_6354,N_5444,N_5655);
and U6355 (N_6355,N_5294,N_5292);
nand U6356 (N_6356,N_5110,N_5159);
and U6357 (N_6357,N_5838,N_5249);
nand U6358 (N_6358,N_5106,N_5691);
nor U6359 (N_6359,N_5369,N_5178);
nor U6360 (N_6360,N_5358,N_5003);
nand U6361 (N_6361,N_5247,N_5136);
nor U6362 (N_6362,N_5736,N_5098);
nor U6363 (N_6363,N_5571,N_5905);
or U6364 (N_6364,N_5522,N_5198);
nor U6365 (N_6365,N_5310,N_5973);
or U6366 (N_6366,N_5913,N_5560);
or U6367 (N_6367,N_5688,N_5822);
or U6368 (N_6368,N_5010,N_5860);
or U6369 (N_6369,N_5550,N_5964);
or U6370 (N_6370,N_5129,N_5479);
or U6371 (N_6371,N_5206,N_5471);
nand U6372 (N_6372,N_5621,N_5812);
nand U6373 (N_6373,N_5681,N_5515);
and U6374 (N_6374,N_5596,N_5542);
and U6375 (N_6375,N_5482,N_5425);
and U6376 (N_6376,N_5826,N_5966);
and U6377 (N_6377,N_5000,N_5234);
or U6378 (N_6378,N_5209,N_5043);
or U6379 (N_6379,N_5852,N_5146);
or U6380 (N_6380,N_5763,N_5177);
nor U6381 (N_6381,N_5430,N_5794);
or U6382 (N_6382,N_5742,N_5958);
nor U6383 (N_6383,N_5856,N_5863);
or U6384 (N_6384,N_5380,N_5368);
nand U6385 (N_6385,N_5258,N_5717);
and U6386 (N_6386,N_5730,N_5504);
nand U6387 (N_6387,N_5052,N_5203);
nand U6388 (N_6388,N_5142,N_5782);
nor U6389 (N_6389,N_5637,N_5778);
nand U6390 (N_6390,N_5846,N_5518);
nor U6391 (N_6391,N_5293,N_5455);
and U6392 (N_6392,N_5988,N_5326);
and U6393 (N_6393,N_5221,N_5656);
nor U6394 (N_6394,N_5943,N_5324);
nor U6395 (N_6395,N_5411,N_5120);
nor U6396 (N_6396,N_5500,N_5901);
nand U6397 (N_6397,N_5975,N_5853);
nor U6398 (N_6398,N_5270,N_5155);
nand U6399 (N_6399,N_5508,N_5213);
xor U6400 (N_6400,N_5336,N_5395);
and U6401 (N_6401,N_5382,N_5118);
nand U6402 (N_6402,N_5184,N_5892);
xnor U6403 (N_6403,N_5041,N_5780);
or U6404 (N_6404,N_5559,N_5193);
and U6405 (N_6405,N_5171,N_5930);
and U6406 (N_6406,N_5978,N_5680);
nand U6407 (N_6407,N_5954,N_5938);
or U6408 (N_6408,N_5475,N_5332);
or U6409 (N_6409,N_5842,N_5397);
and U6410 (N_6410,N_5408,N_5836);
or U6411 (N_6411,N_5825,N_5592);
nor U6412 (N_6412,N_5059,N_5250);
nor U6413 (N_6413,N_5564,N_5893);
xnor U6414 (N_6414,N_5606,N_5183);
nor U6415 (N_6415,N_5108,N_5528);
nor U6416 (N_6416,N_5032,N_5956);
xor U6417 (N_6417,N_5217,N_5389);
nor U6418 (N_6418,N_5328,N_5351);
nor U6419 (N_6419,N_5347,N_5469);
nand U6420 (N_6420,N_5503,N_5265);
nor U6421 (N_6421,N_5135,N_5871);
nor U6422 (N_6422,N_5378,N_5803);
or U6423 (N_6423,N_5779,N_5698);
nor U6424 (N_6424,N_5660,N_5418);
and U6425 (N_6425,N_5765,N_5593);
and U6426 (N_6426,N_5882,N_5940);
nand U6427 (N_6427,N_5207,N_5672);
or U6428 (N_6428,N_5821,N_5974);
nand U6429 (N_6429,N_5219,N_5315);
xnor U6430 (N_6430,N_5732,N_5572);
nor U6431 (N_6431,N_5296,N_5376);
nand U6432 (N_6432,N_5831,N_5224);
nor U6433 (N_6433,N_5580,N_5189);
nor U6434 (N_6434,N_5878,N_5781);
xnor U6435 (N_6435,N_5029,N_5980);
nor U6436 (N_6436,N_5823,N_5752);
nand U6437 (N_6437,N_5538,N_5595);
or U6438 (N_6438,N_5248,N_5199);
and U6439 (N_6439,N_5661,N_5740);
and U6440 (N_6440,N_5543,N_5682);
and U6441 (N_6441,N_5490,N_5505);
nand U6442 (N_6442,N_5239,N_5139);
nand U6443 (N_6443,N_5971,N_5630);
nand U6444 (N_6444,N_5011,N_5214);
nand U6445 (N_6445,N_5749,N_5617);
or U6446 (N_6446,N_5887,N_5067);
and U6447 (N_6447,N_5341,N_5130);
xnor U6448 (N_6448,N_5874,N_5845);
nand U6449 (N_6449,N_5088,N_5910);
and U6450 (N_6450,N_5574,N_5828);
xor U6451 (N_6451,N_5783,N_5981);
or U6452 (N_6452,N_5379,N_5334);
nor U6453 (N_6453,N_5291,N_5194);
and U6454 (N_6454,N_5723,N_5715);
or U6455 (N_6455,N_5947,N_5220);
or U6456 (N_6456,N_5741,N_5282);
or U6457 (N_6457,N_5998,N_5684);
or U6458 (N_6458,N_5461,N_5357);
or U6459 (N_6459,N_5747,N_5308);
or U6460 (N_6460,N_5704,N_5708);
and U6461 (N_6461,N_5186,N_5931);
and U6462 (N_6462,N_5354,N_5141);
and U6463 (N_6463,N_5046,N_5306);
or U6464 (N_6464,N_5267,N_5953);
nand U6465 (N_6465,N_5323,N_5733);
nor U6466 (N_6466,N_5007,N_5197);
and U6467 (N_6467,N_5545,N_5116);
nand U6468 (N_6468,N_5348,N_5367);
and U6469 (N_6469,N_5685,N_5259);
or U6470 (N_6470,N_5190,N_5768);
nand U6471 (N_6471,N_5582,N_5915);
nand U6472 (N_6472,N_5585,N_5394);
or U6473 (N_6473,N_5899,N_5122);
and U6474 (N_6474,N_5049,N_5044);
nand U6475 (N_6475,N_5801,N_5944);
and U6476 (N_6476,N_5388,N_5895);
nand U6477 (N_6477,N_5982,N_5745);
nor U6478 (N_6478,N_5855,N_5531);
or U6479 (N_6479,N_5952,N_5658);
or U6480 (N_6480,N_5535,N_5992);
nor U6481 (N_6481,N_5728,N_5920);
or U6482 (N_6482,N_5066,N_5635);
or U6483 (N_6483,N_5514,N_5850);
and U6484 (N_6484,N_5023,N_5644);
or U6485 (N_6485,N_5132,N_5578);
and U6486 (N_6486,N_5889,N_5009);
nand U6487 (N_6487,N_5223,N_5107);
nand U6488 (N_6488,N_5164,N_5353);
nand U6489 (N_6489,N_5327,N_5993);
nor U6490 (N_6490,N_5227,N_5420);
or U6491 (N_6491,N_5738,N_5356);
and U6492 (N_6492,N_5062,N_5109);
and U6493 (N_6493,N_5597,N_5261);
and U6494 (N_6494,N_5287,N_5157);
nand U6495 (N_6495,N_5548,N_5743);
nand U6496 (N_6496,N_5767,N_5829);
and U6497 (N_6497,N_5799,N_5391);
nand U6498 (N_6498,N_5345,N_5898);
and U6499 (N_6499,N_5725,N_5989);
nor U6500 (N_6500,N_5282,N_5279);
or U6501 (N_6501,N_5970,N_5666);
and U6502 (N_6502,N_5486,N_5771);
and U6503 (N_6503,N_5285,N_5797);
nor U6504 (N_6504,N_5733,N_5632);
or U6505 (N_6505,N_5106,N_5811);
and U6506 (N_6506,N_5187,N_5338);
nor U6507 (N_6507,N_5973,N_5546);
or U6508 (N_6508,N_5399,N_5756);
nor U6509 (N_6509,N_5831,N_5825);
and U6510 (N_6510,N_5157,N_5518);
nor U6511 (N_6511,N_5525,N_5309);
nor U6512 (N_6512,N_5018,N_5903);
nand U6513 (N_6513,N_5072,N_5548);
nand U6514 (N_6514,N_5095,N_5178);
nor U6515 (N_6515,N_5679,N_5840);
nand U6516 (N_6516,N_5103,N_5415);
nor U6517 (N_6517,N_5536,N_5807);
nor U6518 (N_6518,N_5655,N_5536);
or U6519 (N_6519,N_5575,N_5156);
nand U6520 (N_6520,N_5430,N_5886);
and U6521 (N_6521,N_5531,N_5278);
and U6522 (N_6522,N_5327,N_5053);
or U6523 (N_6523,N_5096,N_5020);
or U6524 (N_6524,N_5224,N_5821);
nand U6525 (N_6525,N_5619,N_5494);
or U6526 (N_6526,N_5622,N_5054);
nor U6527 (N_6527,N_5965,N_5649);
and U6528 (N_6528,N_5728,N_5997);
nand U6529 (N_6529,N_5845,N_5194);
nand U6530 (N_6530,N_5726,N_5984);
and U6531 (N_6531,N_5311,N_5953);
and U6532 (N_6532,N_5997,N_5501);
nor U6533 (N_6533,N_5802,N_5433);
and U6534 (N_6534,N_5162,N_5942);
and U6535 (N_6535,N_5496,N_5596);
nor U6536 (N_6536,N_5661,N_5772);
and U6537 (N_6537,N_5408,N_5626);
and U6538 (N_6538,N_5701,N_5453);
nor U6539 (N_6539,N_5065,N_5003);
nor U6540 (N_6540,N_5768,N_5476);
or U6541 (N_6541,N_5120,N_5536);
nor U6542 (N_6542,N_5358,N_5175);
and U6543 (N_6543,N_5989,N_5938);
and U6544 (N_6544,N_5275,N_5300);
nand U6545 (N_6545,N_5457,N_5470);
nand U6546 (N_6546,N_5387,N_5116);
or U6547 (N_6547,N_5109,N_5503);
and U6548 (N_6548,N_5638,N_5602);
or U6549 (N_6549,N_5771,N_5311);
xor U6550 (N_6550,N_5497,N_5068);
nand U6551 (N_6551,N_5013,N_5474);
or U6552 (N_6552,N_5783,N_5285);
and U6553 (N_6553,N_5598,N_5257);
or U6554 (N_6554,N_5980,N_5472);
or U6555 (N_6555,N_5583,N_5985);
or U6556 (N_6556,N_5794,N_5914);
nand U6557 (N_6557,N_5383,N_5259);
nand U6558 (N_6558,N_5920,N_5097);
nand U6559 (N_6559,N_5308,N_5372);
or U6560 (N_6560,N_5093,N_5288);
nand U6561 (N_6561,N_5716,N_5190);
and U6562 (N_6562,N_5657,N_5207);
or U6563 (N_6563,N_5341,N_5983);
or U6564 (N_6564,N_5093,N_5461);
and U6565 (N_6565,N_5879,N_5362);
and U6566 (N_6566,N_5019,N_5500);
nor U6567 (N_6567,N_5526,N_5191);
and U6568 (N_6568,N_5238,N_5179);
or U6569 (N_6569,N_5412,N_5392);
and U6570 (N_6570,N_5105,N_5112);
nor U6571 (N_6571,N_5105,N_5081);
nand U6572 (N_6572,N_5573,N_5591);
and U6573 (N_6573,N_5597,N_5909);
nand U6574 (N_6574,N_5771,N_5656);
nand U6575 (N_6575,N_5607,N_5170);
nor U6576 (N_6576,N_5844,N_5757);
or U6577 (N_6577,N_5375,N_5501);
nor U6578 (N_6578,N_5740,N_5676);
xnor U6579 (N_6579,N_5632,N_5041);
nor U6580 (N_6580,N_5575,N_5998);
xnor U6581 (N_6581,N_5512,N_5895);
nor U6582 (N_6582,N_5479,N_5872);
nand U6583 (N_6583,N_5586,N_5942);
nand U6584 (N_6584,N_5556,N_5635);
nand U6585 (N_6585,N_5937,N_5733);
nand U6586 (N_6586,N_5505,N_5333);
xor U6587 (N_6587,N_5212,N_5069);
xor U6588 (N_6588,N_5797,N_5247);
and U6589 (N_6589,N_5363,N_5154);
and U6590 (N_6590,N_5275,N_5556);
and U6591 (N_6591,N_5108,N_5600);
nor U6592 (N_6592,N_5705,N_5643);
nand U6593 (N_6593,N_5159,N_5434);
and U6594 (N_6594,N_5931,N_5302);
xnor U6595 (N_6595,N_5932,N_5859);
nor U6596 (N_6596,N_5294,N_5126);
or U6597 (N_6597,N_5201,N_5964);
nand U6598 (N_6598,N_5797,N_5279);
nor U6599 (N_6599,N_5031,N_5772);
xor U6600 (N_6600,N_5820,N_5224);
and U6601 (N_6601,N_5139,N_5060);
nor U6602 (N_6602,N_5171,N_5807);
or U6603 (N_6603,N_5351,N_5696);
and U6604 (N_6604,N_5149,N_5660);
nand U6605 (N_6605,N_5921,N_5430);
or U6606 (N_6606,N_5840,N_5587);
nand U6607 (N_6607,N_5353,N_5787);
and U6608 (N_6608,N_5884,N_5249);
nor U6609 (N_6609,N_5178,N_5476);
or U6610 (N_6610,N_5704,N_5662);
nand U6611 (N_6611,N_5422,N_5896);
nor U6612 (N_6612,N_5704,N_5653);
nand U6613 (N_6613,N_5477,N_5307);
or U6614 (N_6614,N_5230,N_5519);
nand U6615 (N_6615,N_5042,N_5633);
xor U6616 (N_6616,N_5994,N_5679);
xor U6617 (N_6617,N_5469,N_5925);
or U6618 (N_6618,N_5423,N_5389);
or U6619 (N_6619,N_5721,N_5434);
or U6620 (N_6620,N_5289,N_5277);
or U6621 (N_6621,N_5030,N_5379);
nand U6622 (N_6622,N_5986,N_5379);
or U6623 (N_6623,N_5735,N_5066);
nand U6624 (N_6624,N_5044,N_5007);
nor U6625 (N_6625,N_5738,N_5795);
xor U6626 (N_6626,N_5691,N_5140);
or U6627 (N_6627,N_5563,N_5233);
nand U6628 (N_6628,N_5772,N_5787);
nand U6629 (N_6629,N_5013,N_5835);
xnor U6630 (N_6630,N_5155,N_5779);
and U6631 (N_6631,N_5414,N_5284);
or U6632 (N_6632,N_5422,N_5258);
nand U6633 (N_6633,N_5505,N_5495);
nand U6634 (N_6634,N_5533,N_5728);
nor U6635 (N_6635,N_5908,N_5749);
nor U6636 (N_6636,N_5842,N_5530);
nor U6637 (N_6637,N_5955,N_5134);
nand U6638 (N_6638,N_5391,N_5161);
nor U6639 (N_6639,N_5524,N_5555);
nor U6640 (N_6640,N_5117,N_5295);
nor U6641 (N_6641,N_5207,N_5410);
and U6642 (N_6642,N_5650,N_5686);
nor U6643 (N_6643,N_5565,N_5226);
xnor U6644 (N_6644,N_5141,N_5210);
or U6645 (N_6645,N_5019,N_5847);
and U6646 (N_6646,N_5727,N_5858);
nand U6647 (N_6647,N_5095,N_5662);
nand U6648 (N_6648,N_5829,N_5611);
nand U6649 (N_6649,N_5845,N_5370);
nor U6650 (N_6650,N_5529,N_5983);
or U6651 (N_6651,N_5877,N_5551);
nand U6652 (N_6652,N_5753,N_5132);
nor U6653 (N_6653,N_5901,N_5082);
and U6654 (N_6654,N_5261,N_5950);
nor U6655 (N_6655,N_5347,N_5816);
and U6656 (N_6656,N_5949,N_5700);
xnor U6657 (N_6657,N_5939,N_5194);
or U6658 (N_6658,N_5250,N_5111);
or U6659 (N_6659,N_5854,N_5227);
nand U6660 (N_6660,N_5197,N_5849);
and U6661 (N_6661,N_5500,N_5156);
or U6662 (N_6662,N_5684,N_5326);
or U6663 (N_6663,N_5081,N_5495);
and U6664 (N_6664,N_5510,N_5142);
and U6665 (N_6665,N_5256,N_5485);
and U6666 (N_6666,N_5465,N_5195);
xor U6667 (N_6667,N_5160,N_5974);
and U6668 (N_6668,N_5747,N_5314);
nor U6669 (N_6669,N_5277,N_5367);
nand U6670 (N_6670,N_5017,N_5193);
nand U6671 (N_6671,N_5857,N_5966);
and U6672 (N_6672,N_5753,N_5350);
or U6673 (N_6673,N_5991,N_5600);
nor U6674 (N_6674,N_5001,N_5653);
xnor U6675 (N_6675,N_5794,N_5813);
and U6676 (N_6676,N_5462,N_5191);
nand U6677 (N_6677,N_5906,N_5298);
and U6678 (N_6678,N_5686,N_5323);
and U6679 (N_6679,N_5763,N_5501);
and U6680 (N_6680,N_5385,N_5796);
nor U6681 (N_6681,N_5618,N_5912);
nand U6682 (N_6682,N_5173,N_5617);
nor U6683 (N_6683,N_5040,N_5366);
and U6684 (N_6684,N_5652,N_5360);
xnor U6685 (N_6685,N_5402,N_5201);
nand U6686 (N_6686,N_5103,N_5259);
or U6687 (N_6687,N_5446,N_5631);
and U6688 (N_6688,N_5855,N_5339);
nand U6689 (N_6689,N_5922,N_5793);
and U6690 (N_6690,N_5803,N_5578);
and U6691 (N_6691,N_5616,N_5787);
or U6692 (N_6692,N_5952,N_5654);
nor U6693 (N_6693,N_5467,N_5615);
xnor U6694 (N_6694,N_5173,N_5583);
and U6695 (N_6695,N_5520,N_5220);
nand U6696 (N_6696,N_5026,N_5426);
and U6697 (N_6697,N_5428,N_5932);
or U6698 (N_6698,N_5487,N_5778);
nor U6699 (N_6699,N_5371,N_5972);
and U6700 (N_6700,N_5041,N_5226);
nor U6701 (N_6701,N_5551,N_5715);
or U6702 (N_6702,N_5138,N_5860);
or U6703 (N_6703,N_5516,N_5586);
nand U6704 (N_6704,N_5939,N_5970);
nor U6705 (N_6705,N_5194,N_5547);
and U6706 (N_6706,N_5776,N_5560);
nor U6707 (N_6707,N_5708,N_5685);
nor U6708 (N_6708,N_5846,N_5883);
or U6709 (N_6709,N_5963,N_5459);
or U6710 (N_6710,N_5234,N_5442);
nor U6711 (N_6711,N_5204,N_5712);
nor U6712 (N_6712,N_5710,N_5816);
and U6713 (N_6713,N_5707,N_5506);
nand U6714 (N_6714,N_5225,N_5345);
nand U6715 (N_6715,N_5512,N_5806);
xor U6716 (N_6716,N_5534,N_5177);
and U6717 (N_6717,N_5583,N_5975);
or U6718 (N_6718,N_5883,N_5807);
nand U6719 (N_6719,N_5747,N_5281);
nor U6720 (N_6720,N_5008,N_5529);
nand U6721 (N_6721,N_5025,N_5440);
and U6722 (N_6722,N_5655,N_5495);
nor U6723 (N_6723,N_5108,N_5060);
nor U6724 (N_6724,N_5896,N_5219);
nor U6725 (N_6725,N_5765,N_5707);
and U6726 (N_6726,N_5407,N_5450);
and U6727 (N_6727,N_5500,N_5520);
nand U6728 (N_6728,N_5540,N_5352);
and U6729 (N_6729,N_5498,N_5958);
or U6730 (N_6730,N_5748,N_5453);
or U6731 (N_6731,N_5751,N_5862);
xor U6732 (N_6732,N_5627,N_5189);
nor U6733 (N_6733,N_5545,N_5166);
or U6734 (N_6734,N_5963,N_5268);
nand U6735 (N_6735,N_5992,N_5130);
and U6736 (N_6736,N_5272,N_5749);
nand U6737 (N_6737,N_5612,N_5924);
and U6738 (N_6738,N_5081,N_5068);
and U6739 (N_6739,N_5891,N_5613);
nor U6740 (N_6740,N_5757,N_5991);
and U6741 (N_6741,N_5922,N_5943);
nor U6742 (N_6742,N_5676,N_5813);
nand U6743 (N_6743,N_5593,N_5657);
nor U6744 (N_6744,N_5628,N_5475);
or U6745 (N_6745,N_5496,N_5400);
nand U6746 (N_6746,N_5780,N_5643);
and U6747 (N_6747,N_5091,N_5819);
and U6748 (N_6748,N_5966,N_5386);
nand U6749 (N_6749,N_5431,N_5366);
and U6750 (N_6750,N_5735,N_5364);
and U6751 (N_6751,N_5559,N_5306);
or U6752 (N_6752,N_5312,N_5535);
nor U6753 (N_6753,N_5966,N_5170);
or U6754 (N_6754,N_5823,N_5709);
and U6755 (N_6755,N_5103,N_5775);
and U6756 (N_6756,N_5742,N_5676);
or U6757 (N_6757,N_5955,N_5500);
or U6758 (N_6758,N_5532,N_5813);
or U6759 (N_6759,N_5839,N_5416);
nor U6760 (N_6760,N_5945,N_5021);
nand U6761 (N_6761,N_5668,N_5586);
nand U6762 (N_6762,N_5640,N_5673);
or U6763 (N_6763,N_5885,N_5950);
xnor U6764 (N_6764,N_5802,N_5724);
and U6765 (N_6765,N_5615,N_5375);
or U6766 (N_6766,N_5724,N_5500);
nor U6767 (N_6767,N_5679,N_5099);
and U6768 (N_6768,N_5665,N_5730);
or U6769 (N_6769,N_5521,N_5410);
nor U6770 (N_6770,N_5784,N_5320);
nor U6771 (N_6771,N_5754,N_5225);
nor U6772 (N_6772,N_5703,N_5157);
xor U6773 (N_6773,N_5180,N_5291);
xnor U6774 (N_6774,N_5181,N_5570);
nor U6775 (N_6775,N_5623,N_5956);
nand U6776 (N_6776,N_5099,N_5729);
nor U6777 (N_6777,N_5357,N_5520);
nand U6778 (N_6778,N_5786,N_5745);
nand U6779 (N_6779,N_5475,N_5292);
xor U6780 (N_6780,N_5538,N_5467);
nand U6781 (N_6781,N_5841,N_5049);
xor U6782 (N_6782,N_5161,N_5352);
xnor U6783 (N_6783,N_5163,N_5072);
or U6784 (N_6784,N_5046,N_5226);
or U6785 (N_6785,N_5305,N_5779);
nor U6786 (N_6786,N_5386,N_5284);
and U6787 (N_6787,N_5252,N_5704);
xor U6788 (N_6788,N_5098,N_5982);
nand U6789 (N_6789,N_5329,N_5560);
nor U6790 (N_6790,N_5168,N_5756);
nand U6791 (N_6791,N_5906,N_5507);
or U6792 (N_6792,N_5185,N_5742);
or U6793 (N_6793,N_5732,N_5696);
xor U6794 (N_6794,N_5503,N_5867);
or U6795 (N_6795,N_5604,N_5587);
xor U6796 (N_6796,N_5609,N_5521);
or U6797 (N_6797,N_5548,N_5095);
and U6798 (N_6798,N_5905,N_5260);
nor U6799 (N_6799,N_5142,N_5878);
nor U6800 (N_6800,N_5391,N_5346);
nor U6801 (N_6801,N_5788,N_5393);
and U6802 (N_6802,N_5304,N_5385);
nand U6803 (N_6803,N_5862,N_5994);
nor U6804 (N_6804,N_5384,N_5874);
or U6805 (N_6805,N_5689,N_5674);
nand U6806 (N_6806,N_5803,N_5892);
nand U6807 (N_6807,N_5990,N_5199);
nor U6808 (N_6808,N_5196,N_5700);
or U6809 (N_6809,N_5105,N_5418);
xor U6810 (N_6810,N_5501,N_5383);
or U6811 (N_6811,N_5013,N_5807);
or U6812 (N_6812,N_5959,N_5390);
xor U6813 (N_6813,N_5504,N_5178);
xnor U6814 (N_6814,N_5443,N_5648);
nand U6815 (N_6815,N_5466,N_5726);
or U6816 (N_6816,N_5591,N_5428);
nand U6817 (N_6817,N_5329,N_5262);
nor U6818 (N_6818,N_5997,N_5996);
and U6819 (N_6819,N_5270,N_5312);
and U6820 (N_6820,N_5105,N_5119);
and U6821 (N_6821,N_5164,N_5954);
and U6822 (N_6822,N_5042,N_5458);
nor U6823 (N_6823,N_5335,N_5527);
nor U6824 (N_6824,N_5938,N_5770);
nor U6825 (N_6825,N_5865,N_5709);
xor U6826 (N_6826,N_5350,N_5260);
nor U6827 (N_6827,N_5752,N_5925);
xnor U6828 (N_6828,N_5702,N_5333);
and U6829 (N_6829,N_5980,N_5883);
nand U6830 (N_6830,N_5455,N_5602);
or U6831 (N_6831,N_5051,N_5016);
nor U6832 (N_6832,N_5203,N_5425);
nor U6833 (N_6833,N_5131,N_5910);
nand U6834 (N_6834,N_5800,N_5153);
xor U6835 (N_6835,N_5586,N_5221);
or U6836 (N_6836,N_5424,N_5580);
and U6837 (N_6837,N_5978,N_5918);
xor U6838 (N_6838,N_5438,N_5789);
or U6839 (N_6839,N_5531,N_5049);
nand U6840 (N_6840,N_5684,N_5557);
and U6841 (N_6841,N_5661,N_5233);
or U6842 (N_6842,N_5156,N_5762);
or U6843 (N_6843,N_5704,N_5900);
nor U6844 (N_6844,N_5088,N_5034);
or U6845 (N_6845,N_5374,N_5682);
or U6846 (N_6846,N_5834,N_5630);
nor U6847 (N_6847,N_5257,N_5443);
nor U6848 (N_6848,N_5497,N_5353);
and U6849 (N_6849,N_5599,N_5185);
or U6850 (N_6850,N_5207,N_5399);
or U6851 (N_6851,N_5006,N_5516);
or U6852 (N_6852,N_5979,N_5125);
nand U6853 (N_6853,N_5126,N_5448);
xnor U6854 (N_6854,N_5947,N_5347);
or U6855 (N_6855,N_5984,N_5274);
and U6856 (N_6856,N_5112,N_5304);
and U6857 (N_6857,N_5304,N_5231);
and U6858 (N_6858,N_5033,N_5115);
or U6859 (N_6859,N_5831,N_5019);
nand U6860 (N_6860,N_5935,N_5503);
nand U6861 (N_6861,N_5446,N_5705);
nand U6862 (N_6862,N_5138,N_5113);
nand U6863 (N_6863,N_5837,N_5517);
nand U6864 (N_6864,N_5207,N_5361);
and U6865 (N_6865,N_5225,N_5523);
and U6866 (N_6866,N_5318,N_5352);
and U6867 (N_6867,N_5788,N_5928);
or U6868 (N_6868,N_5567,N_5159);
or U6869 (N_6869,N_5278,N_5026);
nor U6870 (N_6870,N_5894,N_5464);
nor U6871 (N_6871,N_5294,N_5107);
and U6872 (N_6872,N_5478,N_5581);
or U6873 (N_6873,N_5092,N_5667);
or U6874 (N_6874,N_5469,N_5485);
nor U6875 (N_6875,N_5200,N_5966);
and U6876 (N_6876,N_5113,N_5263);
nor U6877 (N_6877,N_5843,N_5317);
or U6878 (N_6878,N_5381,N_5683);
nand U6879 (N_6879,N_5478,N_5760);
nor U6880 (N_6880,N_5656,N_5956);
or U6881 (N_6881,N_5208,N_5710);
xor U6882 (N_6882,N_5052,N_5939);
nor U6883 (N_6883,N_5773,N_5212);
nand U6884 (N_6884,N_5868,N_5242);
or U6885 (N_6885,N_5274,N_5600);
xor U6886 (N_6886,N_5113,N_5086);
nand U6887 (N_6887,N_5477,N_5725);
nor U6888 (N_6888,N_5893,N_5184);
xnor U6889 (N_6889,N_5397,N_5897);
xor U6890 (N_6890,N_5831,N_5263);
and U6891 (N_6891,N_5033,N_5915);
or U6892 (N_6892,N_5727,N_5437);
nand U6893 (N_6893,N_5634,N_5690);
and U6894 (N_6894,N_5519,N_5644);
nor U6895 (N_6895,N_5671,N_5002);
nor U6896 (N_6896,N_5234,N_5383);
xor U6897 (N_6897,N_5516,N_5038);
nand U6898 (N_6898,N_5415,N_5041);
or U6899 (N_6899,N_5867,N_5692);
nand U6900 (N_6900,N_5048,N_5948);
and U6901 (N_6901,N_5936,N_5011);
and U6902 (N_6902,N_5568,N_5255);
and U6903 (N_6903,N_5887,N_5215);
nor U6904 (N_6904,N_5314,N_5344);
or U6905 (N_6905,N_5108,N_5502);
nand U6906 (N_6906,N_5706,N_5759);
nor U6907 (N_6907,N_5704,N_5199);
and U6908 (N_6908,N_5169,N_5222);
and U6909 (N_6909,N_5843,N_5809);
nand U6910 (N_6910,N_5899,N_5229);
and U6911 (N_6911,N_5549,N_5756);
nor U6912 (N_6912,N_5586,N_5096);
nor U6913 (N_6913,N_5153,N_5841);
nor U6914 (N_6914,N_5490,N_5556);
or U6915 (N_6915,N_5303,N_5584);
or U6916 (N_6916,N_5540,N_5740);
nand U6917 (N_6917,N_5473,N_5854);
xor U6918 (N_6918,N_5348,N_5261);
or U6919 (N_6919,N_5501,N_5164);
and U6920 (N_6920,N_5029,N_5373);
nand U6921 (N_6921,N_5389,N_5682);
or U6922 (N_6922,N_5475,N_5681);
nor U6923 (N_6923,N_5171,N_5665);
and U6924 (N_6924,N_5067,N_5398);
nand U6925 (N_6925,N_5053,N_5869);
or U6926 (N_6926,N_5502,N_5438);
nand U6927 (N_6927,N_5763,N_5347);
xor U6928 (N_6928,N_5427,N_5210);
and U6929 (N_6929,N_5803,N_5026);
or U6930 (N_6930,N_5332,N_5738);
nor U6931 (N_6931,N_5424,N_5487);
nor U6932 (N_6932,N_5151,N_5541);
nor U6933 (N_6933,N_5532,N_5215);
nor U6934 (N_6934,N_5598,N_5994);
nor U6935 (N_6935,N_5751,N_5281);
nor U6936 (N_6936,N_5583,N_5417);
or U6937 (N_6937,N_5267,N_5058);
and U6938 (N_6938,N_5535,N_5166);
nor U6939 (N_6939,N_5052,N_5205);
nand U6940 (N_6940,N_5529,N_5469);
xor U6941 (N_6941,N_5319,N_5182);
and U6942 (N_6942,N_5674,N_5362);
nor U6943 (N_6943,N_5695,N_5487);
and U6944 (N_6944,N_5294,N_5917);
nor U6945 (N_6945,N_5272,N_5155);
or U6946 (N_6946,N_5873,N_5123);
nor U6947 (N_6947,N_5094,N_5959);
nand U6948 (N_6948,N_5322,N_5756);
and U6949 (N_6949,N_5667,N_5104);
nor U6950 (N_6950,N_5341,N_5952);
or U6951 (N_6951,N_5291,N_5671);
or U6952 (N_6952,N_5931,N_5606);
nand U6953 (N_6953,N_5201,N_5308);
and U6954 (N_6954,N_5561,N_5312);
nand U6955 (N_6955,N_5212,N_5828);
nand U6956 (N_6956,N_5144,N_5262);
or U6957 (N_6957,N_5845,N_5703);
nand U6958 (N_6958,N_5838,N_5091);
or U6959 (N_6959,N_5367,N_5787);
or U6960 (N_6960,N_5594,N_5611);
and U6961 (N_6961,N_5639,N_5218);
and U6962 (N_6962,N_5886,N_5825);
or U6963 (N_6963,N_5418,N_5657);
nand U6964 (N_6964,N_5589,N_5561);
xor U6965 (N_6965,N_5565,N_5526);
nand U6966 (N_6966,N_5145,N_5786);
nand U6967 (N_6967,N_5366,N_5839);
and U6968 (N_6968,N_5350,N_5938);
and U6969 (N_6969,N_5622,N_5577);
nand U6970 (N_6970,N_5293,N_5700);
and U6971 (N_6971,N_5594,N_5342);
or U6972 (N_6972,N_5808,N_5176);
xor U6973 (N_6973,N_5796,N_5474);
and U6974 (N_6974,N_5170,N_5044);
xnor U6975 (N_6975,N_5541,N_5851);
xor U6976 (N_6976,N_5784,N_5743);
nor U6977 (N_6977,N_5205,N_5280);
nor U6978 (N_6978,N_5296,N_5638);
and U6979 (N_6979,N_5590,N_5811);
nand U6980 (N_6980,N_5254,N_5981);
nor U6981 (N_6981,N_5926,N_5399);
nand U6982 (N_6982,N_5146,N_5215);
or U6983 (N_6983,N_5172,N_5687);
nor U6984 (N_6984,N_5156,N_5810);
and U6985 (N_6985,N_5807,N_5293);
or U6986 (N_6986,N_5687,N_5521);
nand U6987 (N_6987,N_5050,N_5569);
nand U6988 (N_6988,N_5452,N_5889);
and U6989 (N_6989,N_5252,N_5622);
nor U6990 (N_6990,N_5332,N_5803);
nor U6991 (N_6991,N_5529,N_5425);
and U6992 (N_6992,N_5774,N_5966);
nor U6993 (N_6993,N_5553,N_5290);
nor U6994 (N_6994,N_5635,N_5350);
nand U6995 (N_6995,N_5973,N_5458);
xnor U6996 (N_6996,N_5858,N_5595);
and U6997 (N_6997,N_5844,N_5947);
nor U6998 (N_6998,N_5956,N_5405);
or U6999 (N_6999,N_5525,N_5555);
xor U7000 (N_7000,N_6443,N_6785);
nor U7001 (N_7001,N_6930,N_6351);
nor U7002 (N_7002,N_6190,N_6433);
nand U7003 (N_7003,N_6715,N_6383);
and U7004 (N_7004,N_6006,N_6671);
and U7005 (N_7005,N_6928,N_6487);
nor U7006 (N_7006,N_6011,N_6838);
or U7007 (N_7007,N_6848,N_6600);
or U7008 (N_7008,N_6696,N_6770);
xor U7009 (N_7009,N_6081,N_6924);
or U7010 (N_7010,N_6140,N_6989);
nor U7011 (N_7011,N_6742,N_6650);
and U7012 (N_7012,N_6904,N_6853);
and U7013 (N_7013,N_6029,N_6907);
xnor U7014 (N_7014,N_6633,N_6297);
nor U7015 (N_7015,N_6075,N_6423);
nand U7016 (N_7016,N_6911,N_6656);
nand U7017 (N_7017,N_6083,N_6273);
nor U7018 (N_7018,N_6200,N_6969);
or U7019 (N_7019,N_6408,N_6660);
and U7020 (N_7020,N_6221,N_6304);
nand U7021 (N_7021,N_6606,N_6258);
or U7022 (N_7022,N_6227,N_6166);
or U7023 (N_7023,N_6105,N_6553);
or U7024 (N_7024,N_6177,N_6555);
and U7025 (N_7025,N_6595,N_6894);
nand U7026 (N_7026,N_6941,N_6461);
and U7027 (N_7027,N_6816,N_6758);
nand U7028 (N_7028,N_6243,N_6126);
and U7029 (N_7029,N_6264,N_6797);
or U7030 (N_7030,N_6840,N_6254);
nand U7031 (N_7031,N_6976,N_6024);
nor U7032 (N_7032,N_6991,N_6884);
or U7033 (N_7033,N_6512,N_6145);
and U7034 (N_7034,N_6057,N_6452);
and U7035 (N_7035,N_6953,N_6438);
xor U7036 (N_7036,N_6677,N_6144);
nor U7037 (N_7037,N_6034,N_6617);
nor U7038 (N_7038,N_6730,N_6886);
or U7039 (N_7039,N_6966,N_6726);
nand U7040 (N_7040,N_6196,N_6870);
nand U7041 (N_7041,N_6073,N_6442);
nand U7042 (N_7042,N_6855,N_6475);
and U7043 (N_7043,N_6516,N_6471);
nand U7044 (N_7044,N_6546,N_6245);
and U7045 (N_7045,N_6421,N_6635);
nand U7046 (N_7046,N_6044,N_6535);
or U7047 (N_7047,N_6988,N_6026);
nand U7048 (N_7048,N_6468,N_6990);
nor U7049 (N_7049,N_6422,N_6756);
or U7050 (N_7050,N_6967,N_6532);
or U7051 (N_7051,N_6001,N_6672);
and U7052 (N_7052,N_6306,N_6776);
or U7053 (N_7053,N_6753,N_6813);
nand U7054 (N_7054,N_6128,N_6049);
or U7055 (N_7055,N_6932,N_6184);
nor U7056 (N_7056,N_6322,N_6665);
nand U7057 (N_7057,N_6880,N_6836);
and U7058 (N_7058,N_6141,N_6181);
or U7059 (N_7059,N_6565,N_6523);
nand U7060 (N_7060,N_6873,N_6241);
xor U7061 (N_7061,N_6805,N_6581);
nor U7062 (N_7062,N_6159,N_6385);
xor U7063 (N_7063,N_6288,N_6788);
and U7064 (N_7064,N_6927,N_6342);
or U7065 (N_7065,N_6175,N_6440);
or U7066 (N_7066,N_6333,N_6249);
or U7067 (N_7067,N_6768,N_6416);
xnor U7068 (N_7068,N_6667,N_6179);
and U7069 (N_7069,N_6301,N_6214);
and U7070 (N_7070,N_6389,N_6291);
nor U7071 (N_7071,N_6220,N_6998);
and U7072 (N_7072,N_6624,N_6290);
and U7073 (N_7073,N_6729,N_6920);
nor U7074 (N_7074,N_6231,N_6088);
or U7075 (N_7075,N_6474,N_6067);
xor U7076 (N_7076,N_6939,N_6430);
nor U7077 (N_7077,N_6154,N_6843);
and U7078 (N_7078,N_6626,N_6051);
or U7079 (N_7079,N_6335,N_6670);
nand U7080 (N_7080,N_6913,N_6480);
nor U7081 (N_7081,N_6597,N_6815);
nor U7082 (N_7082,N_6419,N_6089);
or U7083 (N_7083,N_6640,N_6217);
and U7084 (N_7084,N_6528,N_6109);
nand U7085 (N_7085,N_6136,N_6881);
or U7086 (N_7086,N_6348,N_6708);
xor U7087 (N_7087,N_6634,N_6686);
and U7088 (N_7088,N_6501,N_6395);
xor U7089 (N_7089,N_6142,N_6058);
xor U7090 (N_7090,N_6082,N_6275);
or U7091 (N_7091,N_6035,N_6949);
xor U7092 (N_7092,N_6513,N_6446);
nor U7093 (N_7093,N_6725,N_6601);
nor U7094 (N_7094,N_6917,N_6467);
nor U7095 (N_7095,N_6733,N_6820);
nand U7096 (N_7096,N_6460,N_6347);
or U7097 (N_7097,N_6219,N_6627);
or U7098 (N_7098,N_6394,N_6379);
or U7099 (N_7099,N_6208,N_6203);
and U7100 (N_7100,N_6874,N_6530);
nor U7101 (N_7101,N_6312,N_6673);
nand U7102 (N_7102,N_6132,N_6361);
nand U7103 (N_7103,N_6618,N_6269);
nor U7104 (N_7104,N_6596,N_6127);
nor U7105 (N_7105,N_6387,N_6902);
and U7106 (N_7106,N_6786,N_6824);
and U7107 (N_7107,N_6548,N_6028);
or U7108 (N_7108,N_6534,N_6977);
nand U7109 (N_7109,N_6915,N_6228);
or U7110 (N_7110,N_6226,N_6091);
or U7111 (N_7111,N_6518,N_6524);
or U7112 (N_7112,N_6586,N_6294);
and U7113 (N_7113,N_6162,N_6499);
or U7114 (N_7114,N_6683,N_6278);
or U7115 (N_7115,N_6102,N_6212);
nor U7116 (N_7116,N_6502,N_6354);
nand U7117 (N_7117,N_6774,N_6336);
and U7118 (N_7118,N_6974,N_6591);
or U7119 (N_7119,N_6092,N_6148);
nor U7120 (N_7120,N_6357,N_6772);
nor U7121 (N_7121,N_6572,N_6731);
nor U7122 (N_7122,N_6018,N_6038);
or U7123 (N_7123,N_6345,N_6852);
nor U7124 (N_7124,N_6434,N_6234);
nor U7125 (N_7125,N_6340,N_6527);
or U7126 (N_7126,N_6779,N_6752);
nor U7127 (N_7127,N_6699,N_6317);
or U7128 (N_7128,N_6666,N_6641);
nand U7129 (N_7129,N_6959,N_6537);
and U7130 (N_7130,N_6791,N_6380);
nor U7131 (N_7131,N_6116,N_6687);
nor U7132 (N_7132,N_6084,N_6149);
and U7133 (N_7133,N_6465,N_6946);
nand U7134 (N_7134,N_6093,N_6248);
nor U7135 (N_7135,N_6266,N_6777);
and U7136 (N_7136,N_6839,N_6255);
and U7137 (N_7137,N_6426,N_6503);
nor U7138 (N_7138,N_6287,N_6661);
and U7139 (N_7139,N_6644,N_6372);
or U7140 (N_7140,N_6935,N_6074);
nand U7141 (N_7141,N_6962,N_6384);
or U7142 (N_7142,N_6923,N_6152);
or U7143 (N_7143,N_6482,N_6504);
nand U7144 (N_7144,N_6114,N_6188);
or U7145 (N_7145,N_6303,N_6020);
and U7146 (N_7146,N_6302,N_6204);
or U7147 (N_7147,N_6519,N_6113);
or U7148 (N_7148,N_6763,N_6103);
or U7149 (N_7149,N_6106,N_6186);
nand U7150 (N_7150,N_6251,N_6605);
nand U7151 (N_7151,N_6849,N_6887);
nand U7152 (N_7152,N_6210,N_6013);
nand U7153 (N_7153,N_6701,N_6391);
nand U7154 (N_7154,N_6201,N_6439);
and U7155 (N_7155,N_6522,N_6858);
nor U7156 (N_7156,N_6578,N_6500);
or U7157 (N_7157,N_6560,N_6403);
and U7158 (N_7158,N_6846,N_6330);
and U7159 (N_7159,N_6065,N_6580);
nor U7160 (N_7160,N_6174,N_6331);
nand U7161 (N_7161,N_6736,N_6889);
and U7162 (N_7162,N_6579,N_6589);
and U7163 (N_7163,N_6005,N_6968);
nand U7164 (N_7164,N_6986,N_6137);
nand U7165 (N_7165,N_6897,N_6015);
and U7166 (N_7166,N_6134,N_6632);
nand U7167 (N_7167,N_6664,N_6495);
nor U7168 (N_7168,N_6329,N_6750);
nor U7169 (N_7169,N_6775,N_6246);
xor U7170 (N_7170,N_6676,N_6649);
and U7171 (N_7171,N_6030,N_6794);
nand U7172 (N_7172,N_6541,N_6451);
or U7173 (N_7173,N_6270,N_6021);
nor U7174 (N_7174,N_6994,N_6574);
nor U7175 (N_7175,N_6233,N_6163);
or U7176 (N_7176,N_6222,N_6636);
nor U7177 (N_7177,N_6765,N_6497);
and U7178 (N_7178,N_6762,N_6740);
nor U7179 (N_7179,N_6703,N_6926);
nor U7180 (N_7180,N_6436,N_6515);
and U7181 (N_7181,N_6053,N_6232);
nand U7182 (N_7182,N_6224,N_6898);
and U7183 (N_7183,N_6808,N_6691);
nor U7184 (N_7184,N_6412,N_6124);
nand U7185 (N_7185,N_6450,N_6801);
and U7186 (N_7186,N_6280,N_6704);
or U7187 (N_7187,N_6713,N_6047);
and U7188 (N_7188,N_6257,N_6033);
or U7189 (N_7189,N_6842,N_6919);
nand U7190 (N_7190,N_6993,N_6397);
nand U7191 (N_7191,N_6947,N_6984);
nor U7192 (N_7192,N_6400,N_6071);
xor U7193 (N_7193,N_6469,N_6638);
nor U7194 (N_7194,N_6300,N_6864);
or U7195 (N_7195,N_6476,N_6526);
and U7196 (N_7196,N_6909,N_6749);
nor U7197 (N_7197,N_6823,N_6645);
xnor U7198 (N_7198,N_6925,N_6378);
xor U7199 (N_7199,N_6646,N_6879);
or U7200 (N_7200,N_6707,N_6025);
nand U7201 (N_7201,N_6193,N_6027);
nand U7202 (N_7202,N_6343,N_6238);
or U7203 (N_7203,N_6334,N_6392);
nand U7204 (N_7204,N_6458,N_6800);
nand U7205 (N_7205,N_6374,N_6867);
xor U7206 (N_7206,N_6934,N_6971);
nor U7207 (N_7207,N_6680,N_6888);
and U7208 (N_7208,N_6050,N_6857);
nor U7209 (N_7209,N_6206,N_6851);
nor U7210 (N_7210,N_6484,N_6738);
nor U7211 (N_7211,N_6783,N_6751);
nand U7212 (N_7212,N_6960,N_6260);
nor U7213 (N_7213,N_6658,N_6054);
or U7214 (N_7214,N_6985,N_6337);
or U7215 (N_7215,N_6265,N_6895);
nand U7216 (N_7216,N_6160,N_6358);
and U7217 (N_7217,N_6097,N_6517);
xnor U7218 (N_7218,N_6830,N_6135);
nand U7219 (N_7219,N_6622,N_6556);
nand U7220 (N_7220,N_6016,N_6017);
and U7221 (N_7221,N_6723,N_6583);
nor U7222 (N_7222,N_6529,N_6414);
xor U7223 (N_7223,N_6316,N_6428);
or U7224 (N_7224,N_6720,N_6009);
nor U7225 (N_7225,N_6908,N_6724);
or U7226 (N_7226,N_6259,N_6183);
and U7227 (N_7227,N_6545,N_6138);
xnor U7228 (N_7228,N_6496,N_6975);
xnor U7229 (N_7229,N_6663,N_6295);
nor U7230 (N_7230,N_6153,N_6042);
or U7231 (N_7231,N_6236,N_6271);
or U7232 (N_7232,N_6916,N_6684);
and U7233 (N_7233,N_6115,N_6956);
nor U7234 (N_7234,N_6070,N_6420);
nand U7235 (N_7235,N_6061,N_6566);
nand U7236 (N_7236,N_6445,N_6767);
or U7237 (N_7237,N_6623,N_6628);
nor U7238 (N_7238,N_6931,N_6215);
nand U7239 (N_7239,N_6675,N_6229);
xnor U7240 (N_7240,N_6662,N_6702);
and U7241 (N_7241,N_6488,N_6004);
nor U7242 (N_7242,N_6818,N_6741);
nor U7243 (N_7243,N_6299,N_6182);
and U7244 (N_7244,N_6274,N_6388);
nor U7245 (N_7245,N_6178,N_6764);
nor U7246 (N_7246,N_6790,N_6856);
and U7247 (N_7247,N_6173,N_6120);
nor U7248 (N_7248,N_6697,N_6804);
or U7249 (N_7249,N_6877,N_6032);
and U7250 (N_7250,N_6454,N_6814);
or U7251 (N_7251,N_6958,N_6905);
and U7252 (N_7252,N_6463,N_6747);
or U7253 (N_7253,N_6401,N_6360);
nor U7254 (N_7254,N_6509,N_6709);
nand U7255 (N_7255,N_6043,N_6914);
nor U7256 (N_7256,N_6614,N_6890);
and U7257 (N_7257,N_6315,N_6950);
nor U7258 (N_7258,N_6377,N_6678);
or U7259 (N_7259,N_6368,N_6119);
and U7260 (N_7260,N_6798,N_6320);
and U7261 (N_7261,N_6826,N_6539);
or U7262 (N_7262,N_6418,N_6036);
nor U7263 (N_7263,N_6037,N_6230);
nor U7264 (N_7264,N_6883,N_6111);
nand U7265 (N_7265,N_6064,N_6668);
nor U7266 (N_7266,N_6938,N_6802);
nor U7267 (N_7267,N_6878,N_6531);
xnor U7268 (N_7268,N_6079,N_6659);
and U7269 (N_7269,N_6987,N_6817);
nor U7270 (N_7270,N_6373,N_6252);
nand U7271 (N_7271,N_6121,N_6171);
xor U7272 (N_7272,N_6462,N_6407);
or U7273 (N_7273,N_6072,N_6078);
nand U7274 (N_7274,N_6933,N_6326);
nand U7275 (N_7275,N_6746,N_6411);
nor U7276 (N_7276,N_6778,N_6899);
and U7277 (N_7277,N_6435,N_6940);
xor U7278 (N_7278,N_6429,N_6757);
xor U7279 (N_7279,N_6955,N_6608);
or U7280 (N_7280,N_6457,N_6540);
and U7281 (N_7281,N_6486,N_6716);
xor U7282 (N_7282,N_6982,N_6364);
and U7283 (N_7283,N_6854,N_6155);
nand U7284 (N_7284,N_6821,N_6191);
nor U7285 (N_7285,N_6570,N_6008);
or U7286 (N_7286,N_6584,N_6281);
nor U7287 (N_7287,N_6567,N_6900);
or U7288 (N_7288,N_6240,N_6737);
or U7289 (N_7289,N_6732,N_6727);
nand U7290 (N_7290,N_6076,N_6307);
or U7291 (N_7291,N_6789,N_6787);
or U7292 (N_7292,N_6748,N_6339);
nand U7293 (N_7293,N_6963,N_6399);
nor U7294 (N_7294,N_6272,N_6549);
or U7295 (N_7295,N_6314,N_6822);
and U7296 (N_7296,N_6937,N_6970);
nand U7297 (N_7297,N_6313,N_6328);
nand U7298 (N_7298,N_6755,N_6449);
or U7299 (N_7299,N_6261,N_6344);
and U7300 (N_7300,N_6353,N_6951);
and U7301 (N_7301,N_6189,N_6225);
or U7302 (N_7302,N_6912,N_6685);
or U7303 (N_7303,N_6045,N_6211);
or U7304 (N_7304,N_6041,N_6505);
nor U7305 (N_7305,N_6453,N_6616);
nor U7306 (N_7306,N_6356,N_6485);
and U7307 (N_7307,N_6594,N_6809);
or U7308 (N_7308,N_6615,N_6194);
nor U7309 (N_7309,N_6056,N_6533);
nand U7310 (N_7310,N_6376,N_6022);
xor U7311 (N_7311,N_6007,N_6803);
nand U7312 (N_7312,N_6352,N_6781);
or U7313 (N_7313,N_6557,N_6285);
and U7314 (N_7314,N_6305,N_6000);
and U7315 (N_7315,N_6810,N_6961);
xnor U7316 (N_7316,N_6620,N_6256);
or U7317 (N_7317,N_6850,N_6604);
nand U7318 (N_7318,N_6483,N_6263);
and U7319 (N_7319,N_6996,N_6719);
and U7320 (N_7320,N_6031,N_6997);
nand U7321 (N_7321,N_6631,N_6139);
or U7322 (N_7322,N_6172,N_6048);
or U7323 (N_7323,N_6865,N_6216);
nor U7324 (N_7324,N_6390,N_6866);
xnor U7325 (N_7325,N_6477,N_6157);
nand U7326 (N_7326,N_6739,N_6444);
xor U7327 (N_7327,N_6655,N_6169);
and U7328 (N_7328,N_6359,N_6478);
or U7329 (N_7329,N_6046,N_6369);
nand U7330 (N_7330,N_6382,N_6694);
or U7331 (N_7331,N_6718,N_6795);
nand U7332 (N_7332,N_6055,N_6643);
and U7333 (N_7333,N_6324,N_6187);
or U7334 (N_7334,N_6413,N_6362);
or U7335 (N_7335,N_6828,N_6619);
or U7336 (N_7336,N_6611,N_6068);
and U7337 (N_7337,N_6332,N_6875);
and U7338 (N_7338,N_6479,N_6829);
or U7339 (N_7339,N_6609,N_6693);
and U7340 (N_7340,N_6151,N_6207);
nor U7341 (N_7341,N_6455,N_6761);
and U7342 (N_7342,N_6965,N_6639);
and U7343 (N_7343,N_6393,N_6094);
and U7344 (N_7344,N_6972,N_6648);
nor U7345 (N_7345,N_6327,N_6575);
xnor U7346 (N_7346,N_6223,N_6101);
nor U7347 (N_7347,N_6587,N_6296);
or U7348 (N_7348,N_6003,N_6784);
nand U7349 (N_7349,N_6590,N_6863);
nor U7350 (N_7350,N_6247,N_6573);
xnor U7351 (N_7351,N_6613,N_6277);
or U7352 (N_7352,N_6876,N_6835);
or U7353 (N_7353,N_6095,N_6695);
nor U7354 (N_7354,N_6321,N_6610);
nor U7355 (N_7355,N_6323,N_6250);
nand U7356 (N_7356,N_6404,N_6447);
nand U7357 (N_7357,N_6869,N_6728);
or U7358 (N_7358,N_6481,N_6692);
and U7359 (N_7359,N_6346,N_6921);
nor U7360 (N_7360,N_6712,N_6367);
and U7361 (N_7361,N_6406,N_6122);
and U7362 (N_7362,N_6242,N_6576);
and U7363 (N_7363,N_6492,N_6398);
and U7364 (N_7364,N_6002,N_6493);
nor U7365 (N_7365,N_6559,N_6688);
xor U7366 (N_7366,N_6819,N_6896);
and U7367 (N_7367,N_6466,N_6366);
and U7368 (N_7368,N_6637,N_6903);
nand U7369 (N_7369,N_6812,N_6833);
nand U7370 (N_7370,N_6437,N_6213);
and U7371 (N_7371,N_6218,N_6780);
and U7372 (N_7372,N_6652,N_6268);
nor U7373 (N_7373,N_6284,N_6370);
nand U7374 (N_7374,N_6063,N_6341);
xor U7375 (N_7375,N_6396,N_6860);
nor U7376 (N_7376,N_6981,N_6629);
and U7377 (N_7377,N_6543,N_6156);
or U7378 (N_7378,N_6253,N_6536);
or U7379 (N_7379,N_6521,N_6470);
or U7380 (N_7380,N_6375,N_6918);
and U7381 (N_7381,N_6602,N_6040);
and U7382 (N_7382,N_6592,N_6562);
nor U7383 (N_7383,N_6150,N_6309);
nand U7384 (N_7384,N_6807,N_6992);
and U7385 (N_7385,N_6510,N_6973);
xnor U7386 (N_7386,N_6237,N_6131);
or U7387 (N_7387,N_6554,N_6847);
or U7388 (N_7388,N_6039,N_6859);
nand U7389 (N_7389,N_6901,N_6561);
nor U7390 (N_7390,N_6607,N_6612);
nor U7391 (N_7391,N_6205,N_6490);
or U7392 (N_7392,N_6796,N_6197);
nor U7393 (N_7393,N_6459,N_6711);
nor U7394 (N_7394,N_6117,N_6355);
nor U7395 (N_7395,N_6841,N_6773);
nor U7396 (N_7396,N_6811,N_6577);
nand U7397 (N_7397,N_6170,N_6472);
nand U7398 (N_7398,N_6892,N_6133);
nand U7399 (N_7399,N_6598,N_6432);
or U7400 (N_7400,N_6062,N_6948);
and U7401 (N_7401,N_6603,N_6180);
and U7402 (N_7402,N_6099,N_6569);
nor U7403 (N_7403,N_6410,N_6325);
nor U7404 (N_7404,N_6100,N_6571);
nand U7405 (N_7405,N_6464,N_6110);
and U7406 (N_7406,N_6882,N_6945);
nand U7407 (N_7407,N_6494,N_6276);
nand U7408 (N_7408,N_6108,N_6922);
and U7409 (N_7409,N_6125,N_6585);
nor U7410 (N_7410,N_6087,N_6161);
or U7411 (N_7411,N_6298,N_6832);
nand U7412 (N_7412,N_6621,N_6706);
nand U7413 (N_7413,N_6409,N_6402);
nand U7414 (N_7414,N_6754,N_6090);
nor U7415 (N_7415,N_6386,N_6743);
and U7416 (N_7416,N_6417,N_6999);
nand U7417 (N_7417,N_6674,N_6837);
nand U7418 (N_7418,N_6311,N_6593);
and U7419 (N_7419,N_6944,N_6568);
nor U7420 (N_7420,N_6292,N_6349);
nor U7421 (N_7421,N_6654,N_6086);
nand U7422 (N_7422,N_6168,N_6929);
xor U7423 (N_7423,N_6862,N_6441);
nand U7424 (N_7424,N_6793,N_6167);
nand U7425 (N_7425,N_6995,N_6514);
nor U7426 (N_7426,N_6363,N_6319);
and U7427 (N_7427,N_6957,N_6192);
or U7428 (N_7428,N_6371,N_6165);
nor U7429 (N_7429,N_6952,N_6844);
or U7430 (N_7430,N_6744,N_6698);
nor U7431 (N_7431,N_6456,N_6262);
nor U7432 (N_7432,N_6769,N_6282);
and U7433 (N_7433,N_6980,N_6415);
or U7434 (N_7434,N_6085,N_6158);
nor U7435 (N_7435,N_6508,N_6176);
or U7436 (N_7436,N_6146,N_6279);
nor U7437 (N_7437,N_6538,N_6520);
or U7438 (N_7438,N_6547,N_6112);
xor U7439 (N_7439,N_6118,N_6983);
nand U7440 (N_7440,N_6381,N_6489);
nand U7441 (N_7441,N_6782,N_6845);
xnor U7442 (N_7442,N_6338,N_6542);
nor U7443 (N_7443,N_6080,N_6283);
nor U7444 (N_7444,N_6143,N_6717);
and U7445 (N_7445,N_6424,N_6498);
or U7446 (N_7446,N_6310,N_6511);
and U7447 (N_7447,N_6129,N_6551);
xnor U7448 (N_7448,N_6653,N_6427);
nand U7449 (N_7449,N_6077,N_6104);
and U7450 (N_7450,N_6123,N_6365);
nor U7451 (N_7451,N_6198,N_6199);
xor U7452 (N_7452,N_6681,N_6964);
nand U7453 (N_7453,N_6491,N_6202);
nor U7454 (N_7454,N_6289,N_6164);
and U7455 (N_7455,N_6936,N_6023);
and U7456 (N_7456,N_6235,N_6760);
nor U7457 (N_7457,N_6893,N_6014);
nor U7458 (N_7458,N_6834,N_6979);
and U7459 (N_7459,N_6098,N_6588);
xnor U7460 (N_7460,N_6771,N_6318);
nand U7461 (N_7461,N_6147,N_6792);
nor U7462 (N_7462,N_6558,N_6431);
nand U7463 (N_7463,N_6052,N_6942);
nand U7464 (N_7464,N_6891,N_6550);
or U7465 (N_7465,N_6906,N_6642);
or U7466 (N_7466,N_6735,N_6871);
nand U7467 (N_7467,N_6599,N_6831);
nand U7468 (N_7468,N_6525,N_6868);
and U7469 (N_7469,N_6019,N_6107);
nand U7470 (N_7470,N_6059,N_6657);
xor U7471 (N_7471,N_6722,N_6244);
and U7472 (N_7472,N_6766,N_6564);
nor U7473 (N_7473,N_6425,N_6679);
nand U7474 (N_7474,N_6630,N_6647);
nand U7475 (N_7475,N_6745,N_6405);
nand U7476 (N_7476,N_6872,N_6714);
or U7477 (N_7477,N_6195,N_6705);
nand U7478 (N_7478,N_6069,N_6563);
nand U7479 (N_7479,N_6721,N_6978);
or U7480 (N_7480,N_6734,N_6827);
nor U7481 (N_7481,N_6625,N_6293);
and U7482 (N_7482,N_6286,N_6066);
nor U7483 (N_7483,N_6910,N_6759);
nor U7484 (N_7484,N_6012,N_6473);
or U7485 (N_7485,N_6885,N_6682);
nor U7486 (N_7486,N_6552,N_6689);
and U7487 (N_7487,N_6185,N_6651);
nand U7488 (N_7488,N_6861,N_6507);
nand U7489 (N_7489,N_6506,N_6806);
and U7490 (N_7490,N_6582,N_6308);
xnor U7491 (N_7491,N_6350,N_6130);
nor U7492 (N_7492,N_6096,N_6669);
nor U7493 (N_7493,N_6267,N_6448);
xnor U7494 (N_7494,N_6239,N_6209);
nor U7495 (N_7495,N_6825,N_6710);
nand U7496 (N_7496,N_6010,N_6954);
xor U7497 (N_7497,N_6943,N_6799);
nand U7498 (N_7498,N_6700,N_6060);
nor U7499 (N_7499,N_6690,N_6544);
nand U7500 (N_7500,N_6118,N_6021);
or U7501 (N_7501,N_6022,N_6222);
nor U7502 (N_7502,N_6346,N_6203);
nand U7503 (N_7503,N_6024,N_6736);
and U7504 (N_7504,N_6261,N_6768);
or U7505 (N_7505,N_6586,N_6295);
or U7506 (N_7506,N_6542,N_6816);
nor U7507 (N_7507,N_6317,N_6709);
or U7508 (N_7508,N_6171,N_6499);
and U7509 (N_7509,N_6532,N_6622);
nand U7510 (N_7510,N_6344,N_6214);
nor U7511 (N_7511,N_6926,N_6033);
xor U7512 (N_7512,N_6943,N_6500);
and U7513 (N_7513,N_6486,N_6274);
nor U7514 (N_7514,N_6254,N_6975);
xor U7515 (N_7515,N_6802,N_6555);
and U7516 (N_7516,N_6880,N_6841);
or U7517 (N_7517,N_6749,N_6666);
nor U7518 (N_7518,N_6079,N_6611);
nand U7519 (N_7519,N_6560,N_6524);
nand U7520 (N_7520,N_6820,N_6553);
nand U7521 (N_7521,N_6421,N_6863);
and U7522 (N_7522,N_6138,N_6911);
nand U7523 (N_7523,N_6762,N_6478);
nand U7524 (N_7524,N_6734,N_6442);
and U7525 (N_7525,N_6355,N_6366);
nand U7526 (N_7526,N_6645,N_6722);
nand U7527 (N_7527,N_6186,N_6756);
or U7528 (N_7528,N_6103,N_6359);
nor U7529 (N_7529,N_6091,N_6443);
nand U7530 (N_7530,N_6046,N_6408);
nor U7531 (N_7531,N_6367,N_6966);
nand U7532 (N_7532,N_6837,N_6976);
and U7533 (N_7533,N_6249,N_6913);
nor U7534 (N_7534,N_6549,N_6727);
or U7535 (N_7535,N_6046,N_6400);
or U7536 (N_7536,N_6024,N_6931);
or U7537 (N_7537,N_6217,N_6737);
nor U7538 (N_7538,N_6051,N_6635);
nor U7539 (N_7539,N_6933,N_6759);
or U7540 (N_7540,N_6460,N_6818);
and U7541 (N_7541,N_6334,N_6020);
nor U7542 (N_7542,N_6523,N_6765);
xor U7543 (N_7543,N_6448,N_6177);
nand U7544 (N_7544,N_6475,N_6927);
or U7545 (N_7545,N_6295,N_6135);
nor U7546 (N_7546,N_6615,N_6417);
xor U7547 (N_7547,N_6810,N_6147);
nor U7548 (N_7548,N_6246,N_6484);
and U7549 (N_7549,N_6148,N_6598);
or U7550 (N_7550,N_6556,N_6372);
xor U7551 (N_7551,N_6038,N_6816);
nor U7552 (N_7552,N_6031,N_6154);
nand U7553 (N_7553,N_6731,N_6904);
or U7554 (N_7554,N_6573,N_6925);
nand U7555 (N_7555,N_6321,N_6485);
or U7556 (N_7556,N_6874,N_6603);
and U7557 (N_7557,N_6903,N_6299);
and U7558 (N_7558,N_6951,N_6354);
nor U7559 (N_7559,N_6261,N_6686);
nand U7560 (N_7560,N_6116,N_6830);
nor U7561 (N_7561,N_6835,N_6445);
nand U7562 (N_7562,N_6300,N_6976);
nand U7563 (N_7563,N_6686,N_6045);
and U7564 (N_7564,N_6270,N_6259);
and U7565 (N_7565,N_6372,N_6636);
or U7566 (N_7566,N_6715,N_6623);
nor U7567 (N_7567,N_6265,N_6022);
nor U7568 (N_7568,N_6981,N_6536);
and U7569 (N_7569,N_6936,N_6219);
nor U7570 (N_7570,N_6645,N_6513);
nor U7571 (N_7571,N_6691,N_6759);
or U7572 (N_7572,N_6989,N_6337);
nor U7573 (N_7573,N_6896,N_6031);
nand U7574 (N_7574,N_6422,N_6384);
or U7575 (N_7575,N_6293,N_6918);
nor U7576 (N_7576,N_6661,N_6898);
or U7577 (N_7577,N_6005,N_6163);
nand U7578 (N_7578,N_6075,N_6144);
and U7579 (N_7579,N_6326,N_6834);
nor U7580 (N_7580,N_6616,N_6003);
nor U7581 (N_7581,N_6211,N_6629);
nand U7582 (N_7582,N_6659,N_6228);
or U7583 (N_7583,N_6872,N_6039);
nand U7584 (N_7584,N_6576,N_6655);
or U7585 (N_7585,N_6218,N_6407);
and U7586 (N_7586,N_6738,N_6259);
nor U7587 (N_7587,N_6052,N_6564);
nor U7588 (N_7588,N_6349,N_6342);
nand U7589 (N_7589,N_6446,N_6569);
and U7590 (N_7590,N_6432,N_6877);
nor U7591 (N_7591,N_6956,N_6727);
nor U7592 (N_7592,N_6810,N_6278);
nor U7593 (N_7593,N_6877,N_6027);
or U7594 (N_7594,N_6134,N_6753);
and U7595 (N_7595,N_6606,N_6711);
or U7596 (N_7596,N_6339,N_6196);
or U7597 (N_7597,N_6212,N_6959);
and U7598 (N_7598,N_6958,N_6401);
and U7599 (N_7599,N_6022,N_6937);
nand U7600 (N_7600,N_6305,N_6020);
and U7601 (N_7601,N_6675,N_6726);
nand U7602 (N_7602,N_6523,N_6853);
xor U7603 (N_7603,N_6633,N_6079);
nor U7604 (N_7604,N_6990,N_6827);
nor U7605 (N_7605,N_6342,N_6224);
xor U7606 (N_7606,N_6696,N_6354);
nand U7607 (N_7607,N_6452,N_6705);
nor U7608 (N_7608,N_6483,N_6848);
xnor U7609 (N_7609,N_6380,N_6397);
xnor U7610 (N_7610,N_6397,N_6894);
nand U7611 (N_7611,N_6829,N_6791);
nand U7612 (N_7612,N_6603,N_6643);
or U7613 (N_7613,N_6995,N_6435);
nand U7614 (N_7614,N_6037,N_6401);
and U7615 (N_7615,N_6898,N_6527);
xor U7616 (N_7616,N_6585,N_6877);
xnor U7617 (N_7617,N_6057,N_6558);
xor U7618 (N_7618,N_6090,N_6330);
or U7619 (N_7619,N_6492,N_6614);
xnor U7620 (N_7620,N_6420,N_6141);
nor U7621 (N_7621,N_6706,N_6858);
and U7622 (N_7622,N_6946,N_6728);
nor U7623 (N_7623,N_6047,N_6967);
nor U7624 (N_7624,N_6970,N_6631);
nand U7625 (N_7625,N_6485,N_6508);
xnor U7626 (N_7626,N_6738,N_6004);
nor U7627 (N_7627,N_6664,N_6089);
nor U7628 (N_7628,N_6397,N_6528);
or U7629 (N_7629,N_6911,N_6671);
or U7630 (N_7630,N_6883,N_6199);
or U7631 (N_7631,N_6840,N_6674);
nand U7632 (N_7632,N_6341,N_6596);
and U7633 (N_7633,N_6304,N_6482);
and U7634 (N_7634,N_6107,N_6573);
nor U7635 (N_7635,N_6905,N_6869);
xnor U7636 (N_7636,N_6227,N_6161);
and U7637 (N_7637,N_6617,N_6345);
nand U7638 (N_7638,N_6040,N_6973);
and U7639 (N_7639,N_6128,N_6072);
nand U7640 (N_7640,N_6146,N_6502);
or U7641 (N_7641,N_6459,N_6172);
nand U7642 (N_7642,N_6639,N_6816);
nand U7643 (N_7643,N_6625,N_6070);
xor U7644 (N_7644,N_6342,N_6521);
nand U7645 (N_7645,N_6689,N_6057);
and U7646 (N_7646,N_6042,N_6766);
and U7647 (N_7647,N_6569,N_6110);
nor U7648 (N_7648,N_6348,N_6563);
nand U7649 (N_7649,N_6295,N_6060);
nor U7650 (N_7650,N_6341,N_6517);
nor U7651 (N_7651,N_6253,N_6211);
nand U7652 (N_7652,N_6784,N_6508);
and U7653 (N_7653,N_6886,N_6326);
and U7654 (N_7654,N_6083,N_6121);
or U7655 (N_7655,N_6274,N_6330);
nor U7656 (N_7656,N_6266,N_6496);
nor U7657 (N_7657,N_6123,N_6764);
nor U7658 (N_7658,N_6242,N_6241);
nor U7659 (N_7659,N_6201,N_6749);
and U7660 (N_7660,N_6402,N_6972);
or U7661 (N_7661,N_6149,N_6197);
nor U7662 (N_7662,N_6020,N_6621);
nand U7663 (N_7663,N_6044,N_6528);
nor U7664 (N_7664,N_6402,N_6036);
or U7665 (N_7665,N_6348,N_6286);
xnor U7666 (N_7666,N_6049,N_6110);
nor U7667 (N_7667,N_6082,N_6152);
or U7668 (N_7668,N_6476,N_6252);
xnor U7669 (N_7669,N_6777,N_6730);
and U7670 (N_7670,N_6388,N_6893);
nor U7671 (N_7671,N_6403,N_6408);
nand U7672 (N_7672,N_6027,N_6874);
nand U7673 (N_7673,N_6509,N_6283);
and U7674 (N_7674,N_6479,N_6007);
nor U7675 (N_7675,N_6995,N_6035);
nor U7676 (N_7676,N_6246,N_6908);
nand U7677 (N_7677,N_6127,N_6267);
and U7678 (N_7678,N_6525,N_6860);
nand U7679 (N_7679,N_6324,N_6700);
and U7680 (N_7680,N_6408,N_6132);
or U7681 (N_7681,N_6565,N_6671);
and U7682 (N_7682,N_6147,N_6598);
and U7683 (N_7683,N_6179,N_6452);
and U7684 (N_7684,N_6481,N_6564);
or U7685 (N_7685,N_6833,N_6388);
nor U7686 (N_7686,N_6165,N_6020);
nor U7687 (N_7687,N_6574,N_6657);
and U7688 (N_7688,N_6978,N_6005);
or U7689 (N_7689,N_6335,N_6986);
nand U7690 (N_7690,N_6482,N_6253);
or U7691 (N_7691,N_6815,N_6865);
nor U7692 (N_7692,N_6233,N_6998);
and U7693 (N_7693,N_6813,N_6776);
nand U7694 (N_7694,N_6998,N_6884);
and U7695 (N_7695,N_6054,N_6793);
nor U7696 (N_7696,N_6429,N_6549);
xor U7697 (N_7697,N_6190,N_6720);
or U7698 (N_7698,N_6655,N_6280);
xnor U7699 (N_7699,N_6673,N_6548);
or U7700 (N_7700,N_6075,N_6430);
and U7701 (N_7701,N_6615,N_6682);
nor U7702 (N_7702,N_6643,N_6910);
xnor U7703 (N_7703,N_6425,N_6542);
xor U7704 (N_7704,N_6807,N_6630);
or U7705 (N_7705,N_6737,N_6980);
or U7706 (N_7706,N_6484,N_6261);
nand U7707 (N_7707,N_6149,N_6200);
and U7708 (N_7708,N_6591,N_6592);
nand U7709 (N_7709,N_6072,N_6448);
nor U7710 (N_7710,N_6477,N_6966);
nand U7711 (N_7711,N_6912,N_6041);
and U7712 (N_7712,N_6615,N_6909);
nand U7713 (N_7713,N_6199,N_6961);
or U7714 (N_7714,N_6086,N_6688);
or U7715 (N_7715,N_6533,N_6563);
and U7716 (N_7716,N_6503,N_6756);
nor U7717 (N_7717,N_6595,N_6749);
nor U7718 (N_7718,N_6687,N_6112);
and U7719 (N_7719,N_6249,N_6458);
nand U7720 (N_7720,N_6586,N_6361);
nor U7721 (N_7721,N_6829,N_6041);
nor U7722 (N_7722,N_6248,N_6166);
and U7723 (N_7723,N_6315,N_6575);
and U7724 (N_7724,N_6785,N_6505);
and U7725 (N_7725,N_6922,N_6498);
nand U7726 (N_7726,N_6783,N_6483);
nor U7727 (N_7727,N_6452,N_6100);
xnor U7728 (N_7728,N_6139,N_6883);
nor U7729 (N_7729,N_6072,N_6100);
and U7730 (N_7730,N_6356,N_6098);
nor U7731 (N_7731,N_6919,N_6890);
or U7732 (N_7732,N_6303,N_6893);
or U7733 (N_7733,N_6733,N_6512);
or U7734 (N_7734,N_6919,N_6714);
nor U7735 (N_7735,N_6150,N_6571);
and U7736 (N_7736,N_6047,N_6999);
or U7737 (N_7737,N_6410,N_6685);
or U7738 (N_7738,N_6654,N_6109);
and U7739 (N_7739,N_6568,N_6830);
nand U7740 (N_7740,N_6384,N_6086);
nor U7741 (N_7741,N_6083,N_6267);
or U7742 (N_7742,N_6645,N_6402);
or U7743 (N_7743,N_6881,N_6773);
or U7744 (N_7744,N_6743,N_6987);
nor U7745 (N_7745,N_6790,N_6723);
nor U7746 (N_7746,N_6962,N_6700);
nand U7747 (N_7747,N_6784,N_6464);
xor U7748 (N_7748,N_6352,N_6856);
nor U7749 (N_7749,N_6456,N_6323);
nand U7750 (N_7750,N_6866,N_6548);
and U7751 (N_7751,N_6722,N_6214);
xor U7752 (N_7752,N_6273,N_6222);
or U7753 (N_7753,N_6574,N_6178);
or U7754 (N_7754,N_6616,N_6421);
nor U7755 (N_7755,N_6804,N_6351);
nor U7756 (N_7756,N_6324,N_6373);
nand U7757 (N_7757,N_6449,N_6334);
and U7758 (N_7758,N_6483,N_6901);
nand U7759 (N_7759,N_6821,N_6533);
nor U7760 (N_7760,N_6975,N_6952);
xor U7761 (N_7761,N_6230,N_6488);
nor U7762 (N_7762,N_6715,N_6123);
or U7763 (N_7763,N_6087,N_6273);
nor U7764 (N_7764,N_6291,N_6996);
or U7765 (N_7765,N_6226,N_6198);
nand U7766 (N_7766,N_6969,N_6746);
xor U7767 (N_7767,N_6656,N_6279);
nor U7768 (N_7768,N_6798,N_6257);
and U7769 (N_7769,N_6204,N_6409);
or U7770 (N_7770,N_6839,N_6089);
xor U7771 (N_7771,N_6144,N_6389);
or U7772 (N_7772,N_6422,N_6895);
or U7773 (N_7773,N_6494,N_6497);
nand U7774 (N_7774,N_6972,N_6464);
xor U7775 (N_7775,N_6970,N_6839);
nor U7776 (N_7776,N_6369,N_6515);
nor U7777 (N_7777,N_6468,N_6170);
nand U7778 (N_7778,N_6352,N_6253);
nand U7779 (N_7779,N_6784,N_6466);
and U7780 (N_7780,N_6765,N_6037);
nor U7781 (N_7781,N_6682,N_6152);
or U7782 (N_7782,N_6812,N_6186);
nor U7783 (N_7783,N_6049,N_6133);
xnor U7784 (N_7784,N_6856,N_6653);
nor U7785 (N_7785,N_6149,N_6445);
and U7786 (N_7786,N_6420,N_6398);
nor U7787 (N_7787,N_6497,N_6445);
and U7788 (N_7788,N_6528,N_6486);
nand U7789 (N_7789,N_6481,N_6868);
and U7790 (N_7790,N_6303,N_6961);
nor U7791 (N_7791,N_6208,N_6631);
nor U7792 (N_7792,N_6739,N_6563);
or U7793 (N_7793,N_6345,N_6703);
and U7794 (N_7794,N_6913,N_6983);
xor U7795 (N_7795,N_6160,N_6165);
nand U7796 (N_7796,N_6581,N_6000);
nand U7797 (N_7797,N_6277,N_6734);
nor U7798 (N_7798,N_6234,N_6363);
and U7799 (N_7799,N_6090,N_6440);
and U7800 (N_7800,N_6978,N_6204);
nor U7801 (N_7801,N_6958,N_6061);
and U7802 (N_7802,N_6470,N_6535);
nand U7803 (N_7803,N_6845,N_6694);
xnor U7804 (N_7804,N_6413,N_6654);
and U7805 (N_7805,N_6933,N_6234);
or U7806 (N_7806,N_6194,N_6830);
and U7807 (N_7807,N_6971,N_6594);
or U7808 (N_7808,N_6462,N_6421);
or U7809 (N_7809,N_6271,N_6498);
or U7810 (N_7810,N_6561,N_6449);
nand U7811 (N_7811,N_6268,N_6962);
nand U7812 (N_7812,N_6061,N_6372);
or U7813 (N_7813,N_6013,N_6226);
nand U7814 (N_7814,N_6757,N_6319);
nor U7815 (N_7815,N_6932,N_6380);
or U7816 (N_7816,N_6580,N_6669);
nor U7817 (N_7817,N_6437,N_6641);
xor U7818 (N_7818,N_6300,N_6124);
nand U7819 (N_7819,N_6095,N_6355);
nand U7820 (N_7820,N_6887,N_6418);
and U7821 (N_7821,N_6704,N_6921);
and U7822 (N_7822,N_6087,N_6355);
or U7823 (N_7823,N_6277,N_6345);
xor U7824 (N_7824,N_6836,N_6650);
nor U7825 (N_7825,N_6670,N_6369);
nor U7826 (N_7826,N_6240,N_6923);
nor U7827 (N_7827,N_6304,N_6021);
nor U7828 (N_7828,N_6436,N_6569);
xnor U7829 (N_7829,N_6929,N_6369);
or U7830 (N_7830,N_6446,N_6614);
nor U7831 (N_7831,N_6970,N_6049);
nand U7832 (N_7832,N_6632,N_6494);
and U7833 (N_7833,N_6847,N_6659);
and U7834 (N_7834,N_6997,N_6532);
and U7835 (N_7835,N_6702,N_6931);
xor U7836 (N_7836,N_6253,N_6569);
and U7837 (N_7837,N_6521,N_6487);
nor U7838 (N_7838,N_6612,N_6876);
nand U7839 (N_7839,N_6517,N_6524);
nand U7840 (N_7840,N_6638,N_6264);
nand U7841 (N_7841,N_6976,N_6435);
or U7842 (N_7842,N_6147,N_6331);
or U7843 (N_7843,N_6439,N_6223);
nand U7844 (N_7844,N_6181,N_6923);
xnor U7845 (N_7845,N_6874,N_6648);
or U7846 (N_7846,N_6036,N_6027);
nand U7847 (N_7847,N_6986,N_6624);
nor U7848 (N_7848,N_6571,N_6016);
and U7849 (N_7849,N_6044,N_6718);
nand U7850 (N_7850,N_6771,N_6968);
nor U7851 (N_7851,N_6127,N_6914);
or U7852 (N_7852,N_6452,N_6037);
nand U7853 (N_7853,N_6895,N_6052);
xor U7854 (N_7854,N_6433,N_6536);
and U7855 (N_7855,N_6673,N_6421);
nor U7856 (N_7856,N_6207,N_6514);
and U7857 (N_7857,N_6499,N_6278);
nand U7858 (N_7858,N_6737,N_6313);
or U7859 (N_7859,N_6197,N_6915);
nand U7860 (N_7860,N_6660,N_6601);
nand U7861 (N_7861,N_6103,N_6170);
or U7862 (N_7862,N_6764,N_6271);
and U7863 (N_7863,N_6525,N_6296);
xnor U7864 (N_7864,N_6968,N_6850);
and U7865 (N_7865,N_6322,N_6990);
nor U7866 (N_7866,N_6553,N_6337);
or U7867 (N_7867,N_6159,N_6215);
nor U7868 (N_7868,N_6742,N_6714);
or U7869 (N_7869,N_6314,N_6833);
nand U7870 (N_7870,N_6920,N_6994);
or U7871 (N_7871,N_6517,N_6199);
nand U7872 (N_7872,N_6154,N_6943);
or U7873 (N_7873,N_6216,N_6197);
nor U7874 (N_7874,N_6694,N_6158);
nand U7875 (N_7875,N_6190,N_6278);
nand U7876 (N_7876,N_6753,N_6030);
nor U7877 (N_7877,N_6663,N_6040);
or U7878 (N_7878,N_6802,N_6644);
xor U7879 (N_7879,N_6646,N_6690);
or U7880 (N_7880,N_6805,N_6688);
and U7881 (N_7881,N_6333,N_6342);
or U7882 (N_7882,N_6489,N_6424);
or U7883 (N_7883,N_6906,N_6118);
nand U7884 (N_7884,N_6051,N_6015);
and U7885 (N_7885,N_6083,N_6647);
nor U7886 (N_7886,N_6546,N_6476);
and U7887 (N_7887,N_6727,N_6780);
nor U7888 (N_7888,N_6024,N_6016);
nor U7889 (N_7889,N_6790,N_6301);
or U7890 (N_7890,N_6747,N_6679);
nand U7891 (N_7891,N_6588,N_6671);
nor U7892 (N_7892,N_6754,N_6145);
nor U7893 (N_7893,N_6239,N_6993);
nand U7894 (N_7894,N_6164,N_6657);
and U7895 (N_7895,N_6957,N_6840);
and U7896 (N_7896,N_6980,N_6792);
nand U7897 (N_7897,N_6240,N_6134);
and U7898 (N_7898,N_6641,N_6111);
and U7899 (N_7899,N_6156,N_6007);
or U7900 (N_7900,N_6140,N_6459);
nand U7901 (N_7901,N_6637,N_6264);
nand U7902 (N_7902,N_6699,N_6033);
or U7903 (N_7903,N_6206,N_6359);
nand U7904 (N_7904,N_6692,N_6898);
nor U7905 (N_7905,N_6566,N_6164);
or U7906 (N_7906,N_6849,N_6463);
or U7907 (N_7907,N_6727,N_6347);
nand U7908 (N_7908,N_6826,N_6239);
nand U7909 (N_7909,N_6520,N_6915);
nand U7910 (N_7910,N_6501,N_6253);
or U7911 (N_7911,N_6405,N_6563);
nand U7912 (N_7912,N_6268,N_6688);
nand U7913 (N_7913,N_6770,N_6566);
nand U7914 (N_7914,N_6072,N_6034);
nor U7915 (N_7915,N_6669,N_6805);
nand U7916 (N_7916,N_6782,N_6006);
xnor U7917 (N_7917,N_6698,N_6803);
or U7918 (N_7918,N_6933,N_6309);
nor U7919 (N_7919,N_6540,N_6130);
nor U7920 (N_7920,N_6352,N_6726);
nor U7921 (N_7921,N_6639,N_6061);
or U7922 (N_7922,N_6293,N_6195);
nand U7923 (N_7923,N_6386,N_6649);
or U7924 (N_7924,N_6583,N_6750);
nand U7925 (N_7925,N_6554,N_6737);
nand U7926 (N_7926,N_6382,N_6145);
or U7927 (N_7927,N_6299,N_6426);
xor U7928 (N_7928,N_6872,N_6621);
nor U7929 (N_7929,N_6633,N_6743);
nand U7930 (N_7930,N_6770,N_6792);
xnor U7931 (N_7931,N_6555,N_6244);
nand U7932 (N_7932,N_6070,N_6165);
xnor U7933 (N_7933,N_6292,N_6112);
nor U7934 (N_7934,N_6187,N_6749);
nand U7935 (N_7935,N_6885,N_6144);
nor U7936 (N_7936,N_6963,N_6722);
and U7937 (N_7937,N_6247,N_6785);
xor U7938 (N_7938,N_6372,N_6898);
or U7939 (N_7939,N_6209,N_6900);
nand U7940 (N_7940,N_6825,N_6192);
nor U7941 (N_7941,N_6008,N_6200);
nor U7942 (N_7942,N_6881,N_6475);
or U7943 (N_7943,N_6053,N_6340);
nand U7944 (N_7944,N_6031,N_6123);
and U7945 (N_7945,N_6820,N_6176);
and U7946 (N_7946,N_6574,N_6613);
or U7947 (N_7947,N_6976,N_6801);
nor U7948 (N_7948,N_6567,N_6909);
xor U7949 (N_7949,N_6274,N_6658);
xnor U7950 (N_7950,N_6121,N_6840);
and U7951 (N_7951,N_6351,N_6535);
or U7952 (N_7952,N_6161,N_6965);
and U7953 (N_7953,N_6660,N_6716);
and U7954 (N_7954,N_6588,N_6566);
nand U7955 (N_7955,N_6399,N_6124);
nor U7956 (N_7956,N_6100,N_6255);
and U7957 (N_7957,N_6416,N_6833);
or U7958 (N_7958,N_6571,N_6466);
xor U7959 (N_7959,N_6702,N_6552);
nor U7960 (N_7960,N_6823,N_6784);
or U7961 (N_7961,N_6761,N_6960);
xnor U7962 (N_7962,N_6460,N_6123);
nor U7963 (N_7963,N_6493,N_6020);
and U7964 (N_7964,N_6328,N_6756);
and U7965 (N_7965,N_6768,N_6679);
and U7966 (N_7966,N_6623,N_6349);
xor U7967 (N_7967,N_6145,N_6066);
and U7968 (N_7968,N_6698,N_6998);
and U7969 (N_7969,N_6766,N_6225);
nor U7970 (N_7970,N_6238,N_6295);
nor U7971 (N_7971,N_6445,N_6137);
or U7972 (N_7972,N_6045,N_6842);
and U7973 (N_7973,N_6329,N_6028);
nor U7974 (N_7974,N_6853,N_6578);
nor U7975 (N_7975,N_6543,N_6066);
and U7976 (N_7976,N_6414,N_6577);
nand U7977 (N_7977,N_6854,N_6903);
nor U7978 (N_7978,N_6803,N_6016);
or U7979 (N_7979,N_6277,N_6438);
or U7980 (N_7980,N_6650,N_6806);
nand U7981 (N_7981,N_6479,N_6509);
and U7982 (N_7982,N_6441,N_6417);
nor U7983 (N_7983,N_6119,N_6882);
nand U7984 (N_7984,N_6834,N_6267);
nand U7985 (N_7985,N_6147,N_6282);
and U7986 (N_7986,N_6582,N_6862);
nor U7987 (N_7987,N_6656,N_6678);
nand U7988 (N_7988,N_6745,N_6750);
nand U7989 (N_7989,N_6703,N_6382);
nor U7990 (N_7990,N_6958,N_6596);
and U7991 (N_7991,N_6666,N_6473);
nor U7992 (N_7992,N_6191,N_6415);
nor U7993 (N_7993,N_6464,N_6064);
or U7994 (N_7994,N_6606,N_6075);
and U7995 (N_7995,N_6573,N_6448);
xnor U7996 (N_7996,N_6609,N_6820);
nand U7997 (N_7997,N_6806,N_6085);
or U7998 (N_7998,N_6447,N_6193);
and U7999 (N_7999,N_6614,N_6898);
nand U8000 (N_8000,N_7768,N_7147);
and U8001 (N_8001,N_7360,N_7200);
nand U8002 (N_8002,N_7625,N_7807);
nor U8003 (N_8003,N_7624,N_7653);
nand U8004 (N_8004,N_7158,N_7494);
and U8005 (N_8005,N_7443,N_7307);
nand U8006 (N_8006,N_7791,N_7611);
and U8007 (N_8007,N_7867,N_7887);
or U8008 (N_8008,N_7501,N_7640);
nor U8009 (N_8009,N_7765,N_7094);
nand U8010 (N_8010,N_7272,N_7236);
nand U8011 (N_8011,N_7415,N_7164);
nor U8012 (N_8012,N_7603,N_7239);
or U8013 (N_8013,N_7974,N_7652);
nor U8014 (N_8014,N_7851,N_7278);
or U8015 (N_8015,N_7519,N_7295);
nor U8016 (N_8016,N_7071,N_7479);
nor U8017 (N_8017,N_7952,N_7476);
nand U8018 (N_8018,N_7026,N_7133);
or U8019 (N_8019,N_7915,N_7602);
and U8020 (N_8020,N_7448,N_7840);
xnor U8021 (N_8021,N_7771,N_7464);
nor U8022 (N_8022,N_7811,N_7642);
and U8023 (N_8023,N_7114,N_7357);
nand U8024 (N_8024,N_7496,N_7341);
or U8025 (N_8025,N_7097,N_7676);
or U8026 (N_8026,N_7857,N_7264);
nor U8027 (N_8027,N_7474,N_7530);
nor U8028 (N_8028,N_7293,N_7763);
or U8029 (N_8029,N_7810,N_7886);
and U8030 (N_8030,N_7794,N_7711);
and U8031 (N_8031,N_7113,N_7121);
or U8032 (N_8032,N_7186,N_7358);
nand U8033 (N_8033,N_7673,N_7505);
nand U8034 (N_8034,N_7140,N_7083);
or U8035 (N_8035,N_7990,N_7368);
or U8036 (N_8036,N_7480,N_7724);
nand U8037 (N_8037,N_7224,N_7416);
or U8038 (N_8038,N_7498,N_7646);
xor U8039 (N_8039,N_7214,N_7924);
nand U8040 (N_8040,N_7234,N_7754);
or U8041 (N_8041,N_7271,N_7594);
nor U8042 (N_8042,N_7539,N_7165);
nand U8043 (N_8043,N_7403,N_7981);
nand U8044 (N_8044,N_7367,N_7363);
xnor U8045 (N_8045,N_7407,N_7418);
nand U8046 (N_8046,N_7824,N_7864);
nor U8047 (N_8047,N_7093,N_7662);
and U8048 (N_8048,N_7958,N_7375);
and U8049 (N_8049,N_7412,N_7347);
xor U8050 (N_8050,N_7232,N_7792);
or U8051 (N_8051,N_7637,N_7552);
nor U8052 (N_8052,N_7061,N_7429);
nor U8053 (N_8053,N_7090,N_7377);
and U8054 (N_8054,N_7329,N_7457);
or U8055 (N_8055,N_7134,N_7524);
nor U8056 (N_8056,N_7287,N_7683);
and U8057 (N_8057,N_7021,N_7720);
nor U8058 (N_8058,N_7593,N_7491);
nor U8059 (N_8059,N_7331,N_7571);
nand U8060 (N_8060,N_7332,N_7562);
nor U8061 (N_8061,N_7283,N_7649);
or U8062 (N_8062,N_7170,N_7199);
nand U8063 (N_8063,N_7806,N_7863);
or U8064 (N_8064,N_7832,N_7905);
xnor U8065 (N_8065,N_7439,N_7903);
xor U8066 (N_8066,N_7082,N_7871);
and U8067 (N_8067,N_7931,N_7175);
nand U8068 (N_8068,N_7639,N_7813);
nor U8069 (N_8069,N_7786,N_7553);
nor U8070 (N_8070,N_7010,N_7176);
and U8071 (N_8071,N_7185,N_7678);
nand U8072 (N_8072,N_7091,N_7188);
nand U8073 (N_8073,N_7411,N_7390);
nand U8074 (N_8074,N_7945,N_7233);
and U8075 (N_8075,N_7155,N_7019);
nor U8076 (N_8076,N_7627,N_7056);
nand U8077 (N_8077,N_7127,N_7294);
nand U8078 (N_8078,N_7353,N_7323);
xnor U8079 (N_8079,N_7219,N_7761);
and U8080 (N_8080,N_7537,N_7733);
nand U8081 (N_8081,N_7482,N_7364);
and U8082 (N_8082,N_7522,N_7405);
and U8083 (N_8083,N_7401,N_7752);
or U8084 (N_8084,N_7349,N_7820);
nor U8085 (N_8085,N_7535,N_7421);
xnor U8086 (N_8086,N_7260,N_7896);
and U8087 (N_8087,N_7115,N_7477);
or U8088 (N_8088,N_7462,N_7555);
or U8089 (N_8089,N_7445,N_7848);
or U8090 (N_8090,N_7668,N_7050);
nor U8091 (N_8091,N_7174,N_7317);
or U8092 (N_8092,N_7618,N_7104);
or U8093 (N_8093,N_7684,N_7354);
or U8094 (N_8094,N_7858,N_7167);
and U8095 (N_8095,N_7769,N_7612);
and U8096 (N_8096,N_7069,N_7959);
nor U8097 (N_8097,N_7849,N_7723);
or U8098 (N_8098,N_7687,N_7073);
and U8099 (N_8099,N_7484,N_7850);
xnor U8100 (N_8100,N_7085,N_7217);
nor U8101 (N_8101,N_7690,N_7833);
and U8102 (N_8102,N_7128,N_7731);
nand U8103 (N_8103,N_7345,N_7610);
nand U8104 (N_8104,N_7102,N_7322);
and U8105 (N_8105,N_7240,N_7879);
nor U8106 (N_8106,N_7275,N_7351);
or U8107 (N_8107,N_7413,N_7191);
and U8108 (N_8108,N_7468,N_7670);
and U8109 (N_8109,N_7576,N_7921);
nand U8110 (N_8110,N_7311,N_7695);
or U8111 (N_8111,N_7992,N_7908);
and U8112 (N_8112,N_7045,N_7805);
nand U8113 (N_8113,N_7098,N_7265);
and U8114 (N_8114,N_7744,N_7118);
and U8115 (N_8115,N_7528,N_7846);
and U8116 (N_8116,N_7961,N_7554);
nor U8117 (N_8117,N_7038,N_7187);
nor U8118 (N_8118,N_7635,N_7054);
nand U8119 (N_8119,N_7573,N_7391);
nor U8120 (N_8120,N_7614,N_7316);
xor U8121 (N_8121,N_7916,N_7772);
nor U8122 (N_8122,N_7526,N_7398);
and U8123 (N_8123,N_7551,N_7395);
or U8124 (N_8124,N_7031,N_7369);
or U8125 (N_8125,N_7606,N_7545);
or U8126 (N_8126,N_7297,N_7025);
and U8127 (N_8127,N_7760,N_7163);
nand U8128 (N_8128,N_7835,N_7587);
or U8129 (N_8129,N_7937,N_7304);
nand U8130 (N_8130,N_7953,N_7388);
nand U8131 (N_8131,N_7111,N_7737);
nand U8132 (N_8132,N_7490,N_7561);
or U8133 (N_8133,N_7386,N_7719);
nor U8134 (N_8134,N_7276,N_7067);
and U8135 (N_8135,N_7302,N_7968);
nand U8136 (N_8136,N_7036,N_7117);
or U8137 (N_8137,N_7116,N_7076);
or U8138 (N_8138,N_7325,N_7352);
nor U8139 (N_8139,N_7320,N_7617);
nor U8140 (N_8140,N_7201,N_7366);
xnor U8141 (N_8141,N_7442,N_7248);
nor U8142 (N_8142,N_7667,N_7856);
nand U8143 (N_8143,N_7099,N_7972);
nor U8144 (N_8144,N_7438,N_7842);
and U8145 (N_8145,N_7534,N_7204);
and U8146 (N_8146,N_7142,N_7310);
nand U8147 (N_8147,N_7862,N_7874);
nor U8148 (N_8148,N_7447,N_7762);
or U8149 (N_8149,N_7712,N_7507);
xnor U8150 (N_8150,N_7651,N_7566);
and U8151 (N_8151,N_7253,N_7256);
and U8152 (N_8152,N_7558,N_7735);
nand U8153 (N_8153,N_7657,N_7816);
nor U8154 (N_8154,N_7106,N_7120);
and U8155 (N_8155,N_7827,N_7515);
or U8156 (N_8156,N_7124,N_7060);
nand U8157 (N_8157,N_7909,N_7800);
or U8158 (N_8158,N_7773,N_7514);
and U8159 (N_8159,N_7984,N_7556);
and U8160 (N_8160,N_7081,N_7198);
and U8161 (N_8161,N_7801,N_7729);
or U8162 (N_8162,N_7630,N_7699);
nand U8163 (N_8163,N_7608,N_7343);
or U8164 (N_8164,N_7425,N_7444);
and U8165 (N_8165,N_7680,N_7394);
xnor U8166 (N_8166,N_7847,N_7006);
nand U8167 (N_8167,N_7892,N_7714);
nor U8168 (N_8168,N_7169,N_7095);
nand U8169 (N_8169,N_7437,N_7280);
nor U8170 (N_8170,N_7237,N_7975);
nor U8171 (N_8171,N_7956,N_7138);
nand U8172 (N_8172,N_7454,N_7957);
xor U8173 (N_8173,N_7231,N_7826);
nand U8174 (N_8174,N_7273,N_7802);
nor U8175 (N_8175,N_7725,N_7179);
nor U8176 (N_8176,N_7011,N_7033);
or U8177 (N_8177,N_7641,N_7891);
nand U8178 (N_8178,N_7020,N_7075);
xnor U8179 (N_8179,N_7289,N_7463);
nand U8180 (N_8180,N_7225,N_7334);
and U8181 (N_8181,N_7902,N_7694);
xnor U8182 (N_8182,N_7563,N_7404);
or U8183 (N_8183,N_7532,N_7852);
nor U8184 (N_8184,N_7796,N_7266);
nand U8185 (N_8185,N_7035,N_7718);
nand U8186 (N_8186,N_7930,N_7540);
nor U8187 (N_8187,N_7279,N_7172);
or U8188 (N_8188,N_7628,N_7255);
or U8189 (N_8189,N_7359,N_7277);
nor U8190 (N_8190,N_7578,N_7742);
xor U8191 (N_8191,N_7313,N_7478);
nand U8192 (N_8192,N_7135,N_7793);
or U8193 (N_8193,N_7977,N_7192);
nand U8194 (N_8194,N_7638,N_7440);
or U8195 (N_8195,N_7570,N_7782);
or U8196 (N_8196,N_7997,N_7597);
nor U8197 (N_8197,N_7985,N_7195);
nand U8198 (N_8198,N_7516,N_7986);
nand U8199 (N_8199,N_7103,N_7979);
nand U8200 (N_8200,N_7854,N_7643);
nand U8201 (N_8201,N_7636,N_7453);
nand U8202 (N_8202,N_7235,N_7065);
nand U8203 (N_8203,N_7929,N_7942);
nor U8204 (N_8204,N_7938,N_7845);
nand U8205 (N_8205,N_7586,N_7679);
or U8206 (N_8206,N_7365,N_7427);
nor U8207 (N_8207,N_7621,N_7456);
or U8208 (N_8208,N_7868,N_7092);
nand U8209 (N_8209,N_7243,N_7108);
or U8210 (N_8210,N_7549,N_7839);
nand U8211 (N_8211,N_7865,N_7876);
nand U8212 (N_8212,N_7631,N_7348);
and U8213 (N_8213,N_7296,N_7205);
nor U8214 (N_8214,N_7434,N_7996);
nand U8215 (N_8215,N_7966,N_7654);
xnor U8216 (N_8216,N_7809,N_7321);
and U8217 (N_8217,N_7947,N_7776);
xor U8218 (N_8218,N_7568,N_7126);
or U8219 (N_8219,N_7105,N_7130);
nand U8220 (N_8220,N_7898,N_7890);
or U8221 (N_8221,N_7202,N_7346);
and U8222 (N_8222,N_7184,N_7301);
nor U8223 (N_8223,N_7873,N_7764);
and U8224 (N_8224,N_7557,N_7546);
nor U8225 (N_8225,N_7923,N_7156);
and U8226 (N_8226,N_7223,N_7692);
and U8227 (N_8227,N_7181,N_7143);
nand U8228 (N_8228,N_7250,N_7601);
nand U8229 (N_8229,N_7843,N_7564);
nand U8230 (N_8230,N_7604,N_7221);
or U8231 (N_8231,N_7356,N_7086);
nor U8232 (N_8232,N_7433,N_7918);
nand U8233 (N_8233,N_7954,N_7647);
or U8234 (N_8234,N_7877,N_7748);
and U8235 (N_8235,N_7982,N_7666);
nand U8236 (N_8236,N_7312,N_7702);
and U8237 (N_8237,N_7072,N_7978);
or U8238 (N_8238,N_7932,N_7605);
or U8239 (N_8239,N_7686,N_7517);
nand U8240 (N_8240,N_7860,N_7663);
or U8241 (N_8241,N_7671,N_7971);
xor U8242 (N_8242,N_7770,N_7007);
and U8243 (N_8243,N_7987,N_7378);
nand U8244 (N_8244,N_7339,N_7465);
nor U8245 (N_8245,N_7585,N_7577);
nand U8246 (N_8246,N_7788,N_7338);
and U8247 (N_8247,N_7907,N_7922);
nand U8248 (N_8248,N_7241,N_7913);
and U8249 (N_8249,N_7706,N_7327);
nor U8250 (N_8250,N_7672,N_7344);
or U8251 (N_8251,N_7989,N_7910);
nor U8252 (N_8252,N_7335,N_7151);
nand U8253 (N_8253,N_7376,N_7789);
nor U8254 (N_8254,N_7410,N_7125);
nand U8255 (N_8255,N_7177,N_7728);
or U8256 (N_8256,N_7459,N_7944);
nor U8257 (N_8257,N_7661,N_7542);
nand U8258 (N_8258,N_7137,N_7658);
or U8259 (N_8259,N_7077,N_7100);
nor U8260 (N_8260,N_7374,N_7489);
nand U8261 (N_8261,N_7935,N_7159);
nor U8262 (N_8262,N_7052,N_7426);
and U8263 (N_8263,N_7051,N_7467);
nand U8264 (N_8264,N_7853,N_7973);
or U8265 (N_8265,N_7251,N_7591);
or U8266 (N_8266,N_7436,N_7029);
nor U8267 (N_8267,N_7626,N_7965);
nor U8268 (N_8268,N_7392,N_7709);
nand U8269 (N_8269,N_7040,N_7506);
or U8270 (N_8270,N_7584,N_7780);
and U8271 (N_8271,N_7660,N_7139);
nand U8272 (N_8272,N_7084,N_7999);
or U8273 (N_8273,N_7252,N_7834);
and U8274 (N_8274,N_7629,N_7057);
nor U8275 (N_8275,N_7161,N_7715);
or U8276 (N_8276,N_7209,N_7967);
nand U8277 (N_8277,N_7032,N_7449);
nor U8278 (N_8278,N_7948,N_7087);
or U8279 (N_8279,N_7904,N_7939);
and U8280 (N_8280,N_7567,N_7513);
or U8281 (N_8281,N_7227,N_7001);
nand U8282 (N_8282,N_7767,N_7207);
or U8283 (N_8283,N_7408,N_7337);
and U8284 (N_8284,N_7704,N_7218);
nand U8285 (N_8285,N_7895,N_7582);
and U8286 (N_8286,N_7633,N_7815);
nand U8287 (N_8287,N_7122,N_7983);
and U8288 (N_8288,N_7171,N_7998);
nand U8289 (N_8289,N_7046,N_7609);
nand U8290 (N_8290,N_7423,N_7180);
nand U8291 (N_8291,N_7194,N_7037);
and U8292 (N_8292,N_7373,N_7245);
nand U8293 (N_8293,N_7544,N_7785);
nor U8294 (N_8294,N_7149,N_7732);
nor U8295 (N_8295,N_7028,N_7677);
nor U8296 (N_8296,N_7370,N_7005);
nand U8297 (N_8297,N_7875,N_7096);
or U8298 (N_8298,N_7914,N_7736);
nand U8299 (N_8299,N_7166,N_7306);
xor U8300 (N_8300,N_7016,N_7615);
or U8301 (N_8301,N_7299,N_7964);
and U8302 (N_8302,N_7379,N_7705);
or U8303 (N_8303,N_7043,N_7648);
xor U8304 (N_8304,N_7784,N_7995);
nand U8305 (N_8305,N_7825,N_7689);
and U8306 (N_8306,N_7291,N_7009);
or U8307 (N_8307,N_7520,N_7015);
nor U8308 (N_8308,N_7855,N_7074);
nor U8309 (N_8309,N_7281,N_7308);
or U8310 (N_8310,N_7211,N_7483);
nand U8311 (N_8311,N_7027,N_7745);
nor U8312 (N_8312,N_7698,N_7812);
or U8313 (N_8313,N_7883,N_7970);
nor U8314 (N_8314,N_7685,N_7583);
and U8315 (N_8315,N_7927,N_7716);
nand U8316 (N_8316,N_7216,N_7326);
or U8317 (N_8317,N_7389,N_7330);
and U8318 (N_8318,N_7962,N_7538);
xnor U8319 (N_8319,N_7512,N_7779);
nor U8320 (N_8320,N_7747,N_7417);
or U8321 (N_8321,N_7881,N_7814);
or U8322 (N_8322,N_7665,N_7949);
nor U8323 (N_8323,N_7422,N_7249);
nor U8324 (N_8324,N_7047,N_7596);
nand U8325 (N_8325,N_7795,N_7936);
nor U8326 (N_8326,N_7196,N_7844);
nor U8327 (N_8327,N_7409,N_7878);
and U8328 (N_8328,N_7469,N_7925);
or U8329 (N_8329,N_7829,N_7472);
and U8330 (N_8330,N_7220,N_7148);
and U8331 (N_8331,N_7708,N_7645);
and U8332 (N_8332,N_7002,N_7523);
and U8333 (N_8333,N_7870,N_7920);
and U8334 (N_8334,N_7955,N_7059);
nor U8335 (N_8335,N_7739,N_7473);
or U8336 (N_8336,N_7861,N_7541);
nand U8337 (N_8337,N_7088,N_7940);
and U8338 (N_8338,N_7525,N_7527);
xor U8339 (N_8339,N_7384,N_7397);
nor U8340 (N_8340,N_7682,N_7675);
and U8341 (N_8341,N_7778,N_7178);
xor U8342 (N_8342,N_7136,N_7753);
xor U8343 (N_8343,N_7650,N_7058);
or U8344 (N_8344,N_7655,N_7109);
nand U8345 (N_8345,N_7536,N_7432);
xor U8346 (N_8346,N_7722,N_7361);
and U8347 (N_8347,N_7153,N_7182);
xor U8348 (N_8348,N_7493,N_7701);
or U8349 (N_8349,N_7048,N_7589);
and U8350 (N_8350,N_7696,N_7034);
nor U8351 (N_8351,N_7740,N_7828);
and U8352 (N_8352,N_7548,N_7560);
and U8353 (N_8353,N_7014,N_7497);
nor U8354 (N_8354,N_7466,N_7831);
and U8355 (N_8355,N_7242,N_7288);
nand U8356 (N_8356,N_7492,N_7681);
and U8357 (N_8357,N_7580,N_7836);
nor U8358 (N_8358,N_7822,N_7818);
nand U8359 (N_8359,N_7424,N_7726);
nand U8360 (N_8360,N_7414,N_7934);
and U8361 (N_8361,N_7619,N_7509);
nand U8362 (N_8362,N_7495,N_7960);
and U8363 (N_8363,N_7912,N_7309);
nor U8364 (N_8364,N_7215,N_7688);
nor U8365 (N_8365,N_7141,N_7656);
xor U8366 (N_8366,N_7707,N_7980);
nand U8367 (N_8367,N_7906,N_7888);
xnor U8368 (N_8368,N_7503,N_7229);
nand U8369 (N_8369,N_7254,N_7994);
or U8370 (N_8370,N_7743,N_7068);
or U8371 (N_8371,N_7766,N_7441);
nor U8372 (N_8372,N_7008,N_7481);
nand U8373 (N_8373,N_7697,N_7933);
nor U8374 (N_8374,N_7044,N_7168);
nor U8375 (N_8375,N_7446,N_7777);
nand U8376 (N_8376,N_7659,N_7119);
and U8377 (N_8377,N_7838,N_7790);
or U8378 (N_8378,N_7713,N_7882);
nor U8379 (N_8379,N_7669,N_7969);
xnor U8380 (N_8380,N_7259,N_7372);
xnor U8381 (N_8381,N_7926,N_7529);
nand U8382 (N_8382,N_7599,N_7285);
and U8383 (N_8383,N_7144,N_7460);
nor U8384 (N_8384,N_7268,N_7470);
and U8385 (N_8385,N_7774,N_7559);
and U8386 (N_8386,N_7362,N_7450);
and U8387 (N_8387,N_7055,N_7226);
or U8388 (N_8388,N_7230,N_7703);
nand U8389 (N_8389,N_7623,N_7350);
or U8390 (N_8390,N_7502,N_7521);
and U8391 (N_8391,N_7292,N_7080);
nor U8392 (N_8392,N_7004,N_7160);
and U8393 (N_8393,N_7132,N_7943);
nor U8394 (N_8394,N_7588,N_7799);
and U8395 (N_8395,N_7393,N_7693);
nor U8396 (N_8396,N_7569,N_7872);
nand U8397 (N_8397,N_7262,N_7064);
nor U8398 (N_8398,N_7017,N_7721);
and U8399 (N_8399,N_7193,N_7951);
nand U8400 (N_8400,N_7428,N_7157);
or U8401 (N_8401,N_7565,N_7808);
nand U8402 (N_8402,N_7941,N_7257);
nor U8403 (N_8403,N_7821,N_7324);
and U8404 (N_8404,N_7859,N_7823);
and U8405 (N_8405,N_7162,N_7781);
and U8406 (N_8406,N_7717,N_7632);
nand U8407 (N_8407,N_7189,N_7804);
nand U8408 (N_8408,N_7018,N_7210);
or U8409 (N_8409,N_7146,N_7664);
nand U8410 (N_8410,N_7042,N_7003);
nand U8411 (N_8411,N_7066,N_7475);
xnor U8412 (N_8412,N_7183,N_7575);
nand U8413 (N_8413,N_7798,N_7458);
nand U8414 (N_8414,N_7900,N_7487);
xnor U8415 (N_8415,N_7885,N_7893);
and U8416 (N_8416,N_7261,N_7590);
or U8417 (N_8417,N_7270,N_7727);
or U8418 (N_8418,N_7620,N_7817);
and U8419 (N_8419,N_7290,N_7471);
xnor U8420 (N_8420,N_7328,N_7284);
and U8421 (N_8421,N_7298,N_7543);
xnor U8422 (N_8422,N_7598,N_7381);
nor U8423 (N_8423,N_7592,N_7547);
and U8424 (N_8424,N_7371,N_7510);
xor U8425 (N_8425,N_7741,N_7282);
nor U8426 (N_8426,N_7616,N_7129);
nand U8427 (N_8427,N_7755,N_7738);
and U8428 (N_8428,N_7382,N_7451);
nor U8429 (N_8429,N_7746,N_7511);
nor U8430 (N_8430,N_7333,N_7000);
and U8431 (N_8431,N_7600,N_7644);
nor U8432 (N_8432,N_7899,N_7244);
or U8433 (N_8433,N_7756,N_7634);
nor U8434 (N_8434,N_7247,N_7110);
nor U8435 (N_8435,N_7894,N_7819);
and U8436 (N_8436,N_7579,N_7355);
nor U8437 (N_8437,N_7988,N_7691);
and U8438 (N_8438,N_7206,N_7734);
or U8439 (N_8439,N_7783,N_7504);
and U8440 (N_8440,N_7246,N_7315);
xor U8441 (N_8441,N_7123,N_7749);
and U8442 (N_8442,N_7710,N_7500);
xor U8443 (N_8443,N_7595,N_7751);
and U8444 (N_8444,N_7213,N_7112);
nor U8445 (N_8445,N_7869,N_7336);
and U8446 (N_8446,N_7550,N_7730);
nand U8447 (N_8447,N_7101,N_7622);
or U8448 (N_8448,N_7486,N_7488);
nor U8449 (N_8449,N_7078,N_7203);
or U8450 (N_8450,N_7228,N_7340);
nand U8451 (N_8451,N_7039,N_7318);
nand U8452 (N_8452,N_7430,N_7107);
nor U8453 (N_8453,N_7797,N_7062);
nor U8454 (N_8454,N_7190,N_7841);
xnor U8455 (N_8455,N_7917,N_7607);
or U8456 (N_8456,N_7574,N_7837);
nor U8457 (N_8457,N_7173,N_7884);
nor U8458 (N_8458,N_7435,N_7267);
xor U8459 (N_8459,N_7012,N_7387);
nand U8460 (N_8460,N_7775,N_7303);
nor U8461 (N_8461,N_7385,N_7803);
nor U8462 (N_8462,N_7830,N_7946);
nor U8463 (N_8463,N_7499,N_7757);
nand U8464 (N_8464,N_7399,N_7222);
or U8465 (N_8465,N_7053,N_7485);
nor U8466 (N_8466,N_7396,N_7238);
and U8467 (N_8467,N_7269,N_7022);
nor U8468 (N_8468,N_7208,N_7518);
xnor U8469 (N_8469,N_7919,N_7452);
nor U8470 (N_8470,N_7897,N_7150);
and U8471 (N_8471,N_7041,N_7089);
or U8472 (N_8472,N_7420,N_7911);
nor U8473 (N_8473,N_7419,N_7063);
or U8474 (N_8474,N_7880,N_7145);
nor U8475 (N_8475,N_7197,N_7131);
nand U8476 (N_8476,N_7286,N_7400);
or U8477 (N_8477,N_7079,N_7152);
xor U8478 (N_8478,N_7963,N_7976);
nand U8479 (N_8479,N_7508,N_7674);
or U8480 (N_8480,N_7928,N_7750);
nand U8481 (N_8481,N_7314,N_7431);
or U8482 (N_8482,N_7319,N_7049);
nand U8483 (N_8483,N_7342,N_7154);
or U8484 (N_8484,N_7406,N_7300);
nor U8485 (N_8485,N_7866,N_7402);
and U8486 (N_8486,N_7991,N_7993);
or U8487 (N_8487,N_7070,N_7758);
or U8488 (N_8488,N_7700,N_7889);
nand U8489 (N_8489,N_7024,N_7787);
or U8490 (N_8490,N_7461,N_7258);
nor U8491 (N_8491,N_7023,N_7212);
nand U8492 (N_8492,N_7305,N_7901);
or U8493 (N_8493,N_7263,N_7533);
or U8494 (N_8494,N_7030,N_7274);
xor U8495 (N_8495,N_7531,N_7013);
nand U8496 (N_8496,N_7380,N_7759);
and U8497 (N_8497,N_7572,N_7613);
nand U8498 (N_8498,N_7383,N_7581);
and U8499 (N_8499,N_7455,N_7950);
nor U8500 (N_8500,N_7327,N_7045);
nand U8501 (N_8501,N_7559,N_7832);
or U8502 (N_8502,N_7607,N_7145);
and U8503 (N_8503,N_7609,N_7116);
and U8504 (N_8504,N_7421,N_7792);
or U8505 (N_8505,N_7870,N_7104);
or U8506 (N_8506,N_7914,N_7754);
nand U8507 (N_8507,N_7596,N_7626);
nor U8508 (N_8508,N_7919,N_7950);
nor U8509 (N_8509,N_7069,N_7965);
nand U8510 (N_8510,N_7076,N_7313);
nand U8511 (N_8511,N_7352,N_7964);
nor U8512 (N_8512,N_7852,N_7226);
xor U8513 (N_8513,N_7957,N_7894);
nor U8514 (N_8514,N_7406,N_7542);
nor U8515 (N_8515,N_7696,N_7689);
nand U8516 (N_8516,N_7595,N_7172);
and U8517 (N_8517,N_7351,N_7377);
nor U8518 (N_8518,N_7053,N_7473);
xnor U8519 (N_8519,N_7499,N_7273);
and U8520 (N_8520,N_7272,N_7113);
and U8521 (N_8521,N_7207,N_7611);
nor U8522 (N_8522,N_7143,N_7170);
or U8523 (N_8523,N_7953,N_7632);
and U8524 (N_8524,N_7194,N_7869);
nand U8525 (N_8525,N_7329,N_7037);
nor U8526 (N_8526,N_7751,N_7291);
xor U8527 (N_8527,N_7568,N_7525);
or U8528 (N_8528,N_7167,N_7828);
or U8529 (N_8529,N_7622,N_7700);
nor U8530 (N_8530,N_7675,N_7140);
nand U8531 (N_8531,N_7224,N_7062);
nor U8532 (N_8532,N_7295,N_7800);
nand U8533 (N_8533,N_7717,N_7807);
nor U8534 (N_8534,N_7998,N_7155);
or U8535 (N_8535,N_7427,N_7824);
and U8536 (N_8536,N_7581,N_7010);
xor U8537 (N_8537,N_7102,N_7273);
or U8538 (N_8538,N_7404,N_7361);
nand U8539 (N_8539,N_7700,N_7469);
and U8540 (N_8540,N_7982,N_7447);
nand U8541 (N_8541,N_7557,N_7010);
and U8542 (N_8542,N_7402,N_7547);
or U8543 (N_8543,N_7978,N_7525);
xor U8544 (N_8544,N_7856,N_7255);
or U8545 (N_8545,N_7681,N_7487);
or U8546 (N_8546,N_7899,N_7239);
xor U8547 (N_8547,N_7986,N_7726);
and U8548 (N_8548,N_7465,N_7414);
nor U8549 (N_8549,N_7821,N_7398);
or U8550 (N_8550,N_7982,N_7043);
or U8551 (N_8551,N_7668,N_7838);
nor U8552 (N_8552,N_7580,N_7485);
nor U8553 (N_8553,N_7652,N_7044);
nand U8554 (N_8554,N_7762,N_7501);
or U8555 (N_8555,N_7901,N_7838);
or U8556 (N_8556,N_7695,N_7670);
xnor U8557 (N_8557,N_7601,N_7935);
nor U8558 (N_8558,N_7754,N_7477);
nand U8559 (N_8559,N_7720,N_7267);
and U8560 (N_8560,N_7500,N_7610);
nand U8561 (N_8561,N_7393,N_7997);
nand U8562 (N_8562,N_7166,N_7745);
nand U8563 (N_8563,N_7436,N_7051);
and U8564 (N_8564,N_7207,N_7133);
or U8565 (N_8565,N_7453,N_7830);
nor U8566 (N_8566,N_7237,N_7841);
nand U8567 (N_8567,N_7778,N_7712);
nor U8568 (N_8568,N_7666,N_7519);
and U8569 (N_8569,N_7777,N_7752);
nand U8570 (N_8570,N_7721,N_7951);
nand U8571 (N_8571,N_7295,N_7185);
or U8572 (N_8572,N_7977,N_7041);
or U8573 (N_8573,N_7833,N_7769);
nor U8574 (N_8574,N_7295,N_7056);
nand U8575 (N_8575,N_7800,N_7339);
xor U8576 (N_8576,N_7877,N_7984);
nand U8577 (N_8577,N_7667,N_7085);
nor U8578 (N_8578,N_7435,N_7017);
or U8579 (N_8579,N_7215,N_7903);
or U8580 (N_8580,N_7590,N_7522);
xor U8581 (N_8581,N_7071,N_7990);
nor U8582 (N_8582,N_7978,N_7628);
and U8583 (N_8583,N_7773,N_7140);
and U8584 (N_8584,N_7100,N_7333);
xor U8585 (N_8585,N_7975,N_7722);
nor U8586 (N_8586,N_7736,N_7154);
and U8587 (N_8587,N_7168,N_7317);
and U8588 (N_8588,N_7863,N_7837);
or U8589 (N_8589,N_7661,N_7933);
nand U8590 (N_8590,N_7686,N_7398);
or U8591 (N_8591,N_7956,N_7674);
nor U8592 (N_8592,N_7158,N_7809);
and U8593 (N_8593,N_7503,N_7677);
nand U8594 (N_8594,N_7049,N_7083);
or U8595 (N_8595,N_7096,N_7012);
or U8596 (N_8596,N_7459,N_7429);
and U8597 (N_8597,N_7712,N_7609);
and U8598 (N_8598,N_7140,N_7620);
nor U8599 (N_8599,N_7690,N_7363);
or U8600 (N_8600,N_7604,N_7741);
nor U8601 (N_8601,N_7483,N_7013);
xor U8602 (N_8602,N_7856,N_7914);
and U8603 (N_8603,N_7610,N_7703);
and U8604 (N_8604,N_7753,N_7015);
nand U8605 (N_8605,N_7223,N_7932);
nor U8606 (N_8606,N_7077,N_7613);
xnor U8607 (N_8607,N_7267,N_7555);
nor U8608 (N_8608,N_7455,N_7879);
or U8609 (N_8609,N_7738,N_7014);
nor U8610 (N_8610,N_7926,N_7658);
and U8611 (N_8611,N_7667,N_7624);
or U8612 (N_8612,N_7631,N_7514);
nor U8613 (N_8613,N_7124,N_7265);
or U8614 (N_8614,N_7324,N_7577);
and U8615 (N_8615,N_7367,N_7076);
nand U8616 (N_8616,N_7162,N_7310);
nand U8617 (N_8617,N_7343,N_7250);
nor U8618 (N_8618,N_7943,N_7771);
nand U8619 (N_8619,N_7745,N_7065);
and U8620 (N_8620,N_7248,N_7409);
and U8621 (N_8621,N_7124,N_7236);
nand U8622 (N_8622,N_7320,N_7853);
nand U8623 (N_8623,N_7504,N_7419);
xor U8624 (N_8624,N_7397,N_7091);
nor U8625 (N_8625,N_7613,N_7419);
nand U8626 (N_8626,N_7302,N_7369);
nand U8627 (N_8627,N_7904,N_7468);
and U8628 (N_8628,N_7814,N_7607);
nand U8629 (N_8629,N_7336,N_7648);
and U8630 (N_8630,N_7514,N_7264);
or U8631 (N_8631,N_7301,N_7250);
xnor U8632 (N_8632,N_7795,N_7154);
and U8633 (N_8633,N_7258,N_7595);
nand U8634 (N_8634,N_7634,N_7919);
nand U8635 (N_8635,N_7751,N_7603);
or U8636 (N_8636,N_7937,N_7195);
xnor U8637 (N_8637,N_7307,N_7519);
nand U8638 (N_8638,N_7918,N_7543);
nand U8639 (N_8639,N_7887,N_7348);
nor U8640 (N_8640,N_7234,N_7459);
and U8641 (N_8641,N_7548,N_7316);
xnor U8642 (N_8642,N_7866,N_7936);
nor U8643 (N_8643,N_7769,N_7670);
or U8644 (N_8644,N_7119,N_7981);
or U8645 (N_8645,N_7043,N_7544);
nand U8646 (N_8646,N_7353,N_7245);
xor U8647 (N_8647,N_7004,N_7797);
nor U8648 (N_8648,N_7183,N_7082);
xnor U8649 (N_8649,N_7308,N_7616);
nor U8650 (N_8650,N_7264,N_7068);
nand U8651 (N_8651,N_7926,N_7498);
xor U8652 (N_8652,N_7769,N_7108);
nor U8653 (N_8653,N_7886,N_7762);
xnor U8654 (N_8654,N_7328,N_7535);
and U8655 (N_8655,N_7573,N_7832);
nand U8656 (N_8656,N_7356,N_7798);
and U8657 (N_8657,N_7301,N_7524);
and U8658 (N_8658,N_7721,N_7466);
nor U8659 (N_8659,N_7058,N_7192);
or U8660 (N_8660,N_7736,N_7316);
nor U8661 (N_8661,N_7228,N_7323);
nor U8662 (N_8662,N_7219,N_7757);
nor U8663 (N_8663,N_7802,N_7419);
and U8664 (N_8664,N_7450,N_7337);
nand U8665 (N_8665,N_7157,N_7704);
or U8666 (N_8666,N_7703,N_7783);
and U8667 (N_8667,N_7842,N_7090);
or U8668 (N_8668,N_7779,N_7780);
nor U8669 (N_8669,N_7335,N_7797);
or U8670 (N_8670,N_7363,N_7496);
nor U8671 (N_8671,N_7028,N_7916);
or U8672 (N_8672,N_7366,N_7607);
nor U8673 (N_8673,N_7977,N_7221);
nand U8674 (N_8674,N_7220,N_7155);
nand U8675 (N_8675,N_7139,N_7439);
nor U8676 (N_8676,N_7915,N_7289);
nor U8677 (N_8677,N_7512,N_7876);
or U8678 (N_8678,N_7437,N_7426);
or U8679 (N_8679,N_7037,N_7727);
nor U8680 (N_8680,N_7321,N_7379);
or U8681 (N_8681,N_7637,N_7287);
and U8682 (N_8682,N_7465,N_7806);
or U8683 (N_8683,N_7084,N_7647);
nand U8684 (N_8684,N_7987,N_7520);
and U8685 (N_8685,N_7011,N_7150);
nor U8686 (N_8686,N_7547,N_7336);
nor U8687 (N_8687,N_7432,N_7214);
or U8688 (N_8688,N_7269,N_7538);
or U8689 (N_8689,N_7242,N_7038);
xnor U8690 (N_8690,N_7013,N_7923);
and U8691 (N_8691,N_7579,N_7029);
and U8692 (N_8692,N_7922,N_7350);
or U8693 (N_8693,N_7170,N_7107);
xnor U8694 (N_8694,N_7928,N_7964);
nand U8695 (N_8695,N_7822,N_7689);
nor U8696 (N_8696,N_7307,N_7327);
or U8697 (N_8697,N_7465,N_7216);
and U8698 (N_8698,N_7686,N_7801);
nand U8699 (N_8699,N_7519,N_7589);
or U8700 (N_8700,N_7289,N_7686);
and U8701 (N_8701,N_7462,N_7962);
nor U8702 (N_8702,N_7184,N_7198);
nor U8703 (N_8703,N_7400,N_7262);
nand U8704 (N_8704,N_7148,N_7907);
nor U8705 (N_8705,N_7422,N_7543);
and U8706 (N_8706,N_7836,N_7377);
nor U8707 (N_8707,N_7191,N_7627);
xnor U8708 (N_8708,N_7525,N_7660);
nor U8709 (N_8709,N_7987,N_7786);
and U8710 (N_8710,N_7412,N_7776);
or U8711 (N_8711,N_7363,N_7428);
and U8712 (N_8712,N_7575,N_7639);
nor U8713 (N_8713,N_7469,N_7199);
and U8714 (N_8714,N_7336,N_7343);
or U8715 (N_8715,N_7503,N_7728);
nand U8716 (N_8716,N_7057,N_7645);
nand U8717 (N_8717,N_7912,N_7828);
nor U8718 (N_8718,N_7321,N_7640);
nand U8719 (N_8719,N_7045,N_7649);
nand U8720 (N_8720,N_7215,N_7604);
and U8721 (N_8721,N_7414,N_7117);
nor U8722 (N_8722,N_7565,N_7006);
and U8723 (N_8723,N_7491,N_7589);
or U8724 (N_8724,N_7033,N_7042);
nor U8725 (N_8725,N_7735,N_7967);
nand U8726 (N_8726,N_7305,N_7805);
nor U8727 (N_8727,N_7248,N_7679);
nor U8728 (N_8728,N_7044,N_7445);
xnor U8729 (N_8729,N_7295,N_7518);
nand U8730 (N_8730,N_7154,N_7700);
nor U8731 (N_8731,N_7491,N_7288);
and U8732 (N_8732,N_7318,N_7245);
and U8733 (N_8733,N_7368,N_7636);
and U8734 (N_8734,N_7307,N_7898);
or U8735 (N_8735,N_7360,N_7247);
and U8736 (N_8736,N_7107,N_7491);
nor U8737 (N_8737,N_7511,N_7470);
nor U8738 (N_8738,N_7963,N_7396);
nand U8739 (N_8739,N_7931,N_7646);
nand U8740 (N_8740,N_7147,N_7365);
and U8741 (N_8741,N_7652,N_7770);
or U8742 (N_8742,N_7486,N_7048);
nor U8743 (N_8743,N_7943,N_7925);
xnor U8744 (N_8744,N_7024,N_7621);
nand U8745 (N_8745,N_7610,N_7861);
and U8746 (N_8746,N_7458,N_7914);
nand U8747 (N_8747,N_7907,N_7468);
nand U8748 (N_8748,N_7813,N_7573);
nand U8749 (N_8749,N_7764,N_7003);
and U8750 (N_8750,N_7079,N_7998);
or U8751 (N_8751,N_7826,N_7901);
or U8752 (N_8752,N_7212,N_7029);
nor U8753 (N_8753,N_7196,N_7430);
and U8754 (N_8754,N_7605,N_7136);
nand U8755 (N_8755,N_7624,N_7134);
nor U8756 (N_8756,N_7987,N_7035);
nand U8757 (N_8757,N_7051,N_7344);
nor U8758 (N_8758,N_7806,N_7324);
nand U8759 (N_8759,N_7900,N_7620);
nor U8760 (N_8760,N_7324,N_7366);
nor U8761 (N_8761,N_7255,N_7539);
and U8762 (N_8762,N_7894,N_7498);
or U8763 (N_8763,N_7769,N_7478);
and U8764 (N_8764,N_7855,N_7176);
xnor U8765 (N_8765,N_7585,N_7628);
nor U8766 (N_8766,N_7224,N_7370);
and U8767 (N_8767,N_7949,N_7151);
or U8768 (N_8768,N_7184,N_7837);
or U8769 (N_8769,N_7296,N_7872);
and U8770 (N_8770,N_7456,N_7514);
and U8771 (N_8771,N_7937,N_7814);
or U8772 (N_8772,N_7044,N_7385);
nor U8773 (N_8773,N_7552,N_7019);
and U8774 (N_8774,N_7649,N_7398);
and U8775 (N_8775,N_7080,N_7082);
or U8776 (N_8776,N_7434,N_7395);
or U8777 (N_8777,N_7003,N_7851);
nor U8778 (N_8778,N_7096,N_7050);
and U8779 (N_8779,N_7318,N_7563);
nor U8780 (N_8780,N_7307,N_7181);
nand U8781 (N_8781,N_7373,N_7202);
nor U8782 (N_8782,N_7956,N_7383);
and U8783 (N_8783,N_7439,N_7257);
nor U8784 (N_8784,N_7150,N_7513);
or U8785 (N_8785,N_7466,N_7468);
nand U8786 (N_8786,N_7213,N_7659);
and U8787 (N_8787,N_7649,N_7305);
and U8788 (N_8788,N_7604,N_7538);
or U8789 (N_8789,N_7169,N_7671);
xor U8790 (N_8790,N_7859,N_7748);
and U8791 (N_8791,N_7214,N_7028);
nor U8792 (N_8792,N_7223,N_7260);
xnor U8793 (N_8793,N_7723,N_7175);
nand U8794 (N_8794,N_7210,N_7722);
or U8795 (N_8795,N_7221,N_7863);
nand U8796 (N_8796,N_7257,N_7790);
nand U8797 (N_8797,N_7614,N_7689);
nand U8798 (N_8798,N_7554,N_7452);
and U8799 (N_8799,N_7228,N_7689);
or U8800 (N_8800,N_7910,N_7784);
and U8801 (N_8801,N_7215,N_7812);
nor U8802 (N_8802,N_7949,N_7595);
xnor U8803 (N_8803,N_7848,N_7181);
or U8804 (N_8804,N_7821,N_7269);
nand U8805 (N_8805,N_7473,N_7643);
xor U8806 (N_8806,N_7677,N_7785);
nor U8807 (N_8807,N_7654,N_7171);
nor U8808 (N_8808,N_7781,N_7799);
or U8809 (N_8809,N_7556,N_7242);
nand U8810 (N_8810,N_7153,N_7902);
xor U8811 (N_8811,N_7808,N_7241);
nand U8812 (N_8812,N_7325,N_7438);
and U8813 (N_8813,N_7787,N_7121);
nand U8814 (N_8814,N_7740,N_7933);
nand U8815 (N_8815,N_7623,N_7735);
nor U8816 (N_8816,N_7814,N_7317);
nor U8817 (N_8817,N_7126,N_7816);
nand U8818 (N_8818,N_7915,N_7797);
nand U8819 (N_8819,N_7809,N_7619);
nand U8820 (N_8820,N_7303,N_7307);
nor U8821 (N_8821,N_7725,N_7751);
or U8822 (N_8822,N_7775,N_7652);
nor U8823 (N_8823,N_7843,N_7061);
and U8824 (N_8824,N_7957,N_7139);
or U8825 (N_8825,N_7049,N_7266);
and U8826 (N_8826,N_7059,N_7158);
and U8827 (N_8827,N_7943,N_7118);
nor U8828 (N_8828,N_7035,N_7515);
nor U8829 (N_8829,N_7467,N_7548);
or U8830 (N_8830,N_7626,N_7819);
or U8831 (N_8831,N_7406,N_7331);
nand U8832 (N_8832,N_7266,N_7488);
and U8833 (N_8833,N_7000,N_7652);
or U8834 (N_8834,N_7886,N_7637);
nand U8835 (N_8835,N_7359,N_7532);
or U8836 (N_8836,N_7885,N_7541);
and U8837 (N_8837,N_7034,N_7202);
and U8838 (N_8838,N_7081,N_7060);
nor U8839 (N_8839,N_7396,N_7303);
and U8840 (N_8840,N_7348,N_7269);
and U8841 (N_8841,N_7136,N_7573);
nand U8842 (N_8842,N_7144,N_7439);
or U8843 (N_8843,N_7388,N_7806);
nand U8844 (N_8844,N_7437,N_7940);
nor U8845 (N_8845,N_7990,N_7678);
and U8846 (N_8846,N_7990,N_7091);
and U8847 (N_8847,N_7224,N_7105);
nand U8848 (N_8848,N_7713,N_7022);
and U8849 (N_8849,N_7363,N_7165);
nand U8850 (N_8850,N_7445,N_7868);
nand U8851 (N_8851,N_7612,N_7136);
nand U8852 (N_8852,N_7267,N_7689);
and U8853 (N_8853,N_7401,N_7359);
or U8854 (N_8854,N_7444,N_7236);
or U8855 (N_8855,N_7314,N_7241);
nand U8856 (N_8856,N_7075,N_7025);
and U8857 (N_8857,N_7036,N_7596);
and U8858 (N_8858,N_7801,N_7243);
nand U8859 (N_8859,N_7792,N_7484);
nor U8860 (N_8860,N_7552,N_7435);
nand U8861 (N_8861,N_7202,N_7093);
or U8862 (N_8862,N_7879,N_7428);
nand U8863 (N_8863,N_7064,N_7315);
or U8864 (N_8864,N_7404,N_7120);
nand U8865 (N_8865,N_7629,N_7645);
xor U8866 (N_8866,N_7023,N_7573);
nand U8867 (N_8867,N_7052,N_7569);
nand U8868 (N_8868,N_7756,N_7575);
nor U8869 (N_8869,N_7526,N_7978);
xor U8870 (N_8870,N_7892,N_7131);
xnor U8871 (N_8871,N_7161,N_7616);
nand U8872 (N_8872,N_7606,N_7256);
nor U8873 (N_8873,N_7346,N_7698);
nor U8874 (N_8874,N_7168,N_7127);
xor U8875 (N_8875,N_7352,N_7601);
nor U8876 (N_8876,N_7438,N_7632);
nand U8877 (N_8877,N_7575,N_7969);
nor U8878 (N_8878,N_7298,N_7280);
nand U8879 (N_8879,N_7336,N_7970);
and U8880 (N_8880,N_7349,N_7346);
nand U8881 (N_8881,N_7908,N_7320);
nand U8882 (N_8882,N_7290,N_7214);
and U8883 (N_8883,N_7561,N_7536);
nand U8884 (N_8884,N_7994,N_7573);
xnor U8885 (N_8885,N_7749,N_7608);
nand U8886 (N_8886,N_7315,N_7800);
and U8887 (N_8887,N_7976,N_7458);
nand U8888 (N_8888,N_7498,N_7002);
nand U8889 (N_8889,N_7820,N_7738);
nor U8890 (N_8890,N_7692,N_7724);
nor U8891 (N_8891,N_7275,N_7785);
xnor U8892 (N_8892,N_7996,N_7484);
or U8893 (N_8893,N_7573,N_7869);
and U8894 (N_8894,N_7620,N_7353);
nor U8895 (N_8895,N_7528,N_7667);
nand U8896 (N_8896,N_7461,N_7219);
and U8897 (N_8897,N_7067,N_7525);
xnor U8898 (N_8898,N_7319,N_7538);
nor U8899 (N_8899,N_7867,N_7916);
or U8900 (N_8900,N_7415,N_7623);
nor U8901 (N_8901,N_7680,N_7726);
nor U8902 (N_8902,N_7602,N_7301);
nand U8903 (N_8903,N_7667,N_7665);
nand U8904 (N_8904,N_7356,N_7973);
nand U8905 (N_8905,N_7392,N_7456);
nor U8906 (N_8906,N_7868,N_7651);
or U8907 (N_8907,N_7408,N_7859);
or U8908 (N_8908,N_7644,N_7173);
and U8909 (N_8909,N_7510,N_7126);
and U8910 (N_8910,N_7303,N_7820);
nor U8911 (N_8911,N_7655,N_7210);
and U8912 (N_8912,N_7159,N_7470);
nor U8913 (N_8913,N_7504,N_7949);
nand U8914 (N_8914,N_7197,N_7150);
and U8915 (N_8915,N_7700,N_7567);
xor U8916 (N_8916,N_7142,N_7834);
nand U8917 (N_8917,N_7792,N_7294);
xor U8918 (N_8918,N_7662,N_7975);
nand U8919 (N_8919,N_7339,N_7499);
and U8920 (N_8920,N_7462,N_7086);
nor U8921 (N_8921,N_7083,N_7558);
or U8922 (N_8922,N_7981,N_7379);
xor U8923 (N_8923,N_7167,N_7861);
xor U8924 (N_8924,N_7889,N_7683);
nor U8925 (N_8925,N_7469,N_7176);
or U8926 (N_8926,N_7803,N_7167);
and U8927 (N_8927,N_7716,N_7617);
or U8928 (N_8928,N_7142,N_7012);
nor U8929 (N_8929,N_7973,N_7256);
and U8930 (N_8930,N_7281,N_7605);
nand U8931 (N_8931,N_7721,N_7014);
and U8932 (N_8932,N_7262,N_7093);
nand U8933 (N_8933,N_7927,N_7761);
nand U8934 (N_8934,N_7605,N_7263);
and U8935 (N_8935,N_7851,N_7991);
xor U8936 (N_8936,N_7595,N_7531);
or U8937 (N_8937,N_7117,N_7736);
nand U8938 (N_8938,N_7979,N_7108);
nand U8939 (N_8939,N_7089,N_7129);
and U8940 (N_8940,N_7101,N_7751);
or U8941 (N_8941,N_7822,N_7231);
nand U8942 (N_8942,N_7167,N_7450);
and U8943 (N_8943,N_7054,N_7537);
and U8944 (N_8944,N_7249,N_7111);
and U8945 (N_8945,N_7262,N_7580);
or U8946 (N_8946,N_7169,N_7557);
and U8947 (N_8947,N_7446,N_7473);
xor U8948 (N_8948,N_7163,N_7338);
nor U8949 (N_8949,N_7852,N_7580);
xor U8950 (N_8950,N_7430,N_7598);
nand U8951 (N_8951,N_7906,N_7689);
nor U8952 (N_8952,N_7152,N_7963);
nand U8953 (N_8953,N_7414,N_7658);
nand U8954 (N_8954,N_7208,N_7060);
nand U8955 (N_8955,N_7048,N_7322);
or U8956 (N_8956,N_7612,N_7662);
nand U8957 (N_8957,N_7226,N_7000);
xnor U8958 (N_8958,N_7003,N_7201);
nand U8959 (N_8959,N_7818,N_7412);
and U8960 (N_8960,N_7514,N_7007);
xor U8961 (N_8961,N_7311,N_7788);
nor U8962 (N_8962,N_7221,N_7388);
nand U8963 (N_8963,N_7877,N_7764);
or U8964 (N_8964,N_7787,N_7014);
nor U8965 (N_8965,N_7927,N_7709);
nor U8966 (N_8966,N_7531,N_7025);
and U8967 (N_8967,N_7437,N_7331);
nor U8968 (N_8968,N_7077,N_7285);
nand U8969 (N_8969,N_7265,N_7350);
nand U8970 (N_8970,N_7270,N_7623);
nor U8971 (N_8971,N_7794,N_7481);
and U8972 (N_8972,N_7183,N_7564);
nor U8973 (N_8973,N_7073,N_7430);
and U8974 (N_8974,N_7912,N_7845);
or U8975 (N_8975,N_7639,N_7475);
or U8976 (N_8976,N_7520,N_7413);
or U8977 (N_8977,N_7918,N_7012);
nor U8978 (N_8978,N_7791,N_7607);
nor U8979 (N_8979,N_7262,N_7430);
nand U8980 (N_8980,N_7495,N_7955);
nor U8981 (N_8981,N_7706,N_7153);
or U8982 (N_8982,N_7474,N_7454);
and U8983 (N_8983,N_7867,N_7236);
xnor U8984 (N_8984,N_7658,N_7472);
and U8985 (N_8985,N_7976,N_7460);
nand U8986 (N_8986,N_7748,N_7784);
nor U8987 (N_8987,N_7652,N_7344);
and U8988 (N_8988,N_7469,N_7763);
nor U8989 (N_8989,N_7410,N_7170);
nor U8990 (N_8990,N_7189,N_7965);
and U8991 (N_8991,N_7549,N_7512);
or U8992 (N_8992,N_7472,N_7674);
nand U8993 (N_8993,N_7913,N_7357);
or U8994 (N_8994,N_7796,N_7578);
nand U8995 (N_8995,N_7888,N_7518);
and U8996 (N_8996,N_7728,N_7386);
nor U8997 (N_8997,N_7315,N_7465);
nand U8998 (N_8998,N_7845,N_7859);
nand U8999 (N_8999,N_7985,N_7227);
or U9000 (N_9000,N_8915,N_8218);
nand U9001 (N_9001,N_8246,N_8573);
or U9002 (N_9002,N_8873,N_8383);
xnor U9003 (N_9003,N_8385,N_8020);
xnor U9004 (N_9004,N_8286,N_8179);
xnor U9005 (N_9005,N_8474,N_8240);
nor U9006 (N_9006,N_8697,N_8559);
nand U9007 (N_9007,N_8431,N_8751);
xor U9008 (N_9008,N_8794,N_8323);
or U9009 (N_9009,N_8106,N_8967);
nand U9010 (N_9010,N_8144,N_8761);
or U9011 (N_9011,N_8226,N_8622);
and U9012 (N_9012,N_8931,N_8128);
nand U9013 (N_9013,N_8613,N_8419);
and U9014 (N_9014,N_8355,N_8594);
nand U9015 (N_9015,N_8919,N_8845);
nand U9016 (N_9016,N_8554,N_8148);
or U9017 (N_9017,N_8305,N_8508);
and U9018 (N_9018,N_8036,N_8909);
or U9019 (N_9019,N_8839,N_8781);
or U9020 (N_9020,N_8718,N_8347);
or U9021 (N_9021,N_8985,N_8177);
nor U9022 (N_9022,N_8009,N_8297);
nor U9023 (N_9023,N_8166,N_8171);
or U9024 (N_9024,N_8170,N_8512);
nor U9025 (N_9025,N_8889,N_8662);
xor U9026 (N_9026,N_8247,N_8844);
or U9027 (N_9027,N_8363,N_8068);
nor U9028 (N_9028,N_8417,N_8534);
nor U9029 (N_9029,N_8397,N_8441);
nand U9030 (N_9030,N_8436,N_8969);
nand U9031 (N_9031,N_8760,N_8610);
nor U9032 (N_9032,N_8167,N_8414);
nor U9033 (N_9033,N_8310,N_8567);
nand U9034 (N_9034,N_8540,N_8536);
or U9035 (N_9035,N_8766,N_8852);
or U9036 (N_9036,N_8913,N_8388);
nand U9037 (N_9037,N_8618,N_8731);
and U9038 (N_9038,N_8014,N_8461);
xor U9039 (N_9039,N_8937,N_8335);
or U9040 (N_9040,N_8425,N_8269);
nand U9041 (N_9041,N_8409,N_8819);
nor U9042 (N_9042,N_8306,N_8619);
nor U9043 (N_9043,N_8550,N_8309);
nor U9044 (N_9044,N_8719,N_8152);
or U9045 (N_9045,N_8423,N_8894);
or U9046 (N_9046,N_8392,N_8198);
and U9047 (N_9047,N_8353,N_8445);
nand U9048 (N_9048,N_8139,N_8565);
nand U9049 (N_9049,N_8292,N_8365);
and U9050 (N_9050,N_8447,N_8214);
nand U9051 (N_9051,N_8614,N_8775);
or U9052 (N_9052,N_8968,N_8261);
nand U9053 (N_9053,N_8245,N_8348);
or U9054 (N_9054,N_8216,N_8377);
nor U9055 (N_9055,N_8782,N_8429);
and U9056 (N_9056,N_8859,N_8635);
nor U9057 (N_9057,N_8394,N_8548);
nand U9058 (N_9058,N_8869,N_8552);
nor U9059 (N_9059,N_8453,N_8225);
xnor U9060 (N_9060,N_8814,N_8189);
or U9061 (N_9061,N_8283,N_8603);
nor U9062 (N_9062,N_8346,N_8136);
nand U9063 (N_9063,N_8007,N_8910);
nor U9064 (N_9064,N_8497,N_8091);
or U9065 (N_9065,N_8290,N_8041);
or U9066 (N_9066,N_8588,N_8275);
nor U9067 (N_9067,N_8026,N_8024);
or U9068 (N_9068,N_8812,N_8750);
nor U9069 (N_9069,N_8285,N_8800);
or U9070 (N_9070,N_8126,N_8174);
and U9071 (N_9071,N_8176,N_8475);
nor U9072 (N_9072,N_8288,N_8786);
and U9073 (N_9073,N_8119,N_8015);
and U9074 (N_9074,N_8195,N_8252);
or U9075 (N_9075,N_8090,N_8244);
or U9076 (N_9076,N_8890,N_8639);
and U9077 (N_9077,N_8974,N_8096);
or U9078 (N_9078,N_8021,N_8955);
and U9079 (N_9079,N_8029,N_8851);
nand U9080 (N_9080,N_8455,N_8138);
or U9081 (N_9081,N_8607,N_8510);
and U9082 (N_9082,N_8746,N_8878);
or U9083 (N_9083,N_8975,N_8145);
nand U9084 (N_9084,N_8696,N_8713);
or U9085 (N_9085,N_8884,N_8666);
nand U9086 (N_9086,N_8287,N_8577);
nand U9087 (N_9087,N_8542,N_8608);
nand U9088 (N_9088,N_8316,N_8075);
xor U9089 (N_9089,N_8291,N_8893);
nor U9090 (N_9090,N_8952,N_8998);
or U9091 (N_9091,N_8242,N_8105);
and U9092 (N_9092,N_8059,N_8277);
nor U9093 (N_9093,N_8575,N_8169);
nor U9094 (N_9094,N_8768,N_8787);
nand U9095 (N_9095,N_8232,N_8949);
or U9096 (N_9096,N_8100,N_8725);
nor U9097 (N_9097,N_8935,N_8204);
nor U9098 (N_9098,N_8518,N_8591);
nor U9099 (N_9099,N_8837,N_8531);
nand U9100 (N_9100,N_8324,N_8446);
nor U9101 (N_9101,N_8081,N_8156);
or U9102 (N_9102,N_8328,N_8048);
or U9103 (N_9103,N_8765,N_8127);
and U9104 (N_9104,N_8574,N_8272);
or U9105 (N_9105,N_8063,N_8143);
nand U9106 (N_9106,N_8582,N_8856);
nand U9107 (N_9107,N_8891,N_8898);
nand U9108 (N_9108,N_8535,N_8354);
and U9109 (N_9109,N_8117,N_8399);
nand U9110 (N_9110,N_8281,N_8071);
nor U9111 (N_9111,N_8403,N_8107);
nor U9112 (N_9112,N_8312,N_8074);
nand U9113 (N_9113,N_8759,N_8338);
or U9114 (N_9114,N_8407,N_8861);
xnor U9115 (N_9115,N_8589,N_8359);
nor U9116 (N_9116,N_8192,N_8317);
nand U9117 (N_9117,N_8378,N_8122);
nor U9118 (N_9118,N_8572,N_8904);
and U9119 (N_9119,N_8430,N_8806);
and U9120 (N_9120,N_8838,N_8989);
nor U9121 (N_9121,N_8815,N_8372);
xnor U9122 (N_9122,N_8146,N_8903);
and U9123 (N_9123,N_8331,N_8154);
and U9124 (N_9124,N_8595,N_8767);
nand U9125 (N_9125,N_8628,N_8830);
and U9126 (N_9126,N_8108,N_8736);
nand U9127 (N_9127,N_8279,N_8080);
and U9128 (N_9128,N_8289,N_8871);
and U9129 (N_9129,N_8978,N_8769);
nand U9130 (N_9130,N_8630,N_8433);
xnor U9131 (N_9131,N_8957,N_8992);
or U9132 (N_9132,N_8771,N_8562);
nor U9133 (N_9133,N_8185,N_8911);
nor U9134 (N_9134,N_8853,N_8868);
xnor U9135 (N_9135,N_8817,N_8360);
xor U9136 (N_9136,N_8202,N_8364);
or U9137 (N_9137,N_8712,N_8113);
and U9138 (N_9138,N_8458,N_8660);
xor U9139 (N_9139,N_8069,N_8468);
and U9140 (N_9140,N_8165,N_8327);
nand U9141 (N_9141,N_8141,N_8592);
nor U9142 (N_9142,N_8566,N_8135);
and U9143 (N_9143,N_8930,N_8568);
xor U9144 (N_9144,N_8263,N_8197);
nand U9145 (N_9145,N_8717,N_8473);
or U9146 (N_9146,N_8857,N_8877);
nor U9147 (N_9147,N_8023,N_8914);
and U9148 (N_9148,N_8503,N_8631);
and U9149 (N_9149,N_8270,N_8236);
or U9150 (N_9150,N_8826,N_8017);
nor U9151 (N_9151,N_8991,N_8368);
and U9152 (N_9152,N_8576,N_8428);
and U9153 (N_9153,N_8326,N_8657);
nand U9154 (N_9154,N_8448,N_8744);
xnor U9155 (N_9155,N_8304,N_8078);
and U9156 (N_9156,N_8370,N_8563);
nand U9157 (N_9157,N_8895,N_8386);
and U9158 (N_9158,N_8033,N_8502);
or U9159 (N_9159,N_8945,N_8778);
or U9160 (N_9160,N_8284,N_8703);
nand U9161 (N_9161,N_8587,N_8757);
xor U9162 (N_9162,N_8454,N_8175);
or U9163 (N_9163,N_8130,N_8381);
xnor U9164 (N_9164,N_8770,N_8557);
and U9165 (N_9165,N_8537,N_8382);
xor U9166 (N_9166,N_8708,N_8229);
or U9167 (N_9167,N_8209,N_8104);
nor U9168 (N_9168,N_8186,N_8808);
xnor U9169 (N_9169,N_8132,N_8711);
or U9170 (N_9170,N_8199,N_8350);
nand U9171 (N_9171,N_8450,N_8402);
nand U9172 (N_9172,N_8439,N_8529);
or U9173 (N_9173,N_8584,N_8371);
xor U9174 (N_9174,N_8656,N_8042);
xnor U9175 (N_9175,N_8694,N_8401);
xnor U9176 (N_9176,N_8494,N_8564);
nand U9177 (N_9177,N_8161,N_8016);
nand U9178 (N_9178,N_8823,N_8274);
and U9179 (N_9179,N_8267,N_8066);
nand U9180 (N_9180,N_8001,N_8626);
or U9181 (N_9181,N_8493,N_8031);
nand U9182 (N_9182,N_8466,N_8905);
or U9183 (N_9183,N_8341,N_8940);
or U9184 (N_9184,N_8013,N_8996);
nand U9185 (N_9185,N_8956,N_8487);
xor U9186 (N_9186,N_8089,N_8469);
nor U9187 (N_9187,N_8203,N_8602);
and U9188 (N_9188,N_8298,N_8410);
nand U9189 (N_9189,N_8411,N_8999);
xnor U9190 (N_9190,N_8748,N_8065);
nand U9191 (N_9191,N_8791,N_8926);
and U9192 (N_9192,N_8490,N_8387);
nor U9193 (N_9193,N_8389,N_8253);
and U9194 (N_9194,N_8881,N_8665);
nor U9195 (N_9195,N_8349,N_8037);
nand U9196 (N_9196,N_8351,N_8231);
and U9197 (N_9197,N_8040,N_8221);
nand U9198 (N_9198,N_8783,N_8743);
and U9199 (N_9199,N_8390,N_8586);
or U9200 (N_9200,N_8982,N_8738);
nor U9201 (N_9201,N_8633,N_8432);
and U9202 (N_9202,N_8732,N_8959);
or U9203 (N_9203,N_8848,N_8046);
nor U9204 (N_9204,N_8964,N_8963);
nor U9205 (N_9205,N_8380,N_8239);
nand U9206 (N_9206,N_8051,N_8832);
nand U9207 (N_9207,N_8028,N_8282);
and U9208 (N_9208,N_8444,N_8803);
nor U9209 (N_9209,N_8879,N_8793);
nand U9210 (N_9210,N_8836,N_8649);
nand U9211 (N_9211,N_8524,N_8627);
nand U9212 (N_9212,N_8934,N_8249);
and U9213 (N_9213,N_8276,N_8661);
or U9214 (N_9214,N_8673,N_8506);
and U9215 (N_9215,N_8375,N_8958);
nand U9216 (N_9216,N_8257,N_8337);
or U9217 (N_9217,N_8867,N_8753);
or U9218 (N_9218,N_8084,N_8965);
nor U9219 (N_9219,N_8435,N_8217);
or U9220 (N_9220,N_8303,N_8483);
and U9221 (N_9221,N_8509,N_8313);
and U9222 (N_9222,N_8621,N_8311);
xnor U9223 (N_9223,N_8343,N_8356);
nand U9224 (N_9224,N_8440,N_8646);
and U9225 (N_9225,N_8593,N_8082);
nor U9226 (N_9226,N_8211,N_8296);
or U9227 (N_9227,N_8067,N_8034);
nand U9228 (N_9228,N_8155,N_8465);
nand U9229 (N_9229,N_8482,N_8943);
nand U9230 (N_9230,N_8669,N_8115);
xor U9231 (N_9231,N_8319,N_8230);
nand U9232 (N_9232,N_8342,N_8019);
nand U9233 (N_9233,N_8684,N_8809);
or U9234 (N_9234,N_8530,N_8336);
nand U9235 (N_9235,N_8682,N_8097);
and U9236 (N_9236,N_8302,N_8625);
nor U9237 (N_9237,N_8828,N_8056);
and U9238 (N_9238,N_8295,N_8561);
nand U9239 (N_9239,N_8609,N_8874);
and U9240 (N_9240,N_8526,N_8443);
and U9241 (N_9241,N_8058,N_8521);
nor U9242 (N_9242,N_8818,N_8032);
xor U9243 (N_9243,N_8792,N_8971);
and U9244 (N_9244,N_8514,N_8882);
or U9245 (N_9245,N_8413,N_8095);
nor U9246 (N_9246,N_8495,N_8332);
nand U9247 (N_9247,N_8896,N_8396);
or U9248 (N_9248,N_8087,N_8352);
and U9249 (N_9249,N_8228,N_8426);
nand U9250 (N_9250,N_8980,N_8578);
nor U9251 (N_9251,N_8273,N_8266);
or U9252 (N_9252,N_8504,N_8271);
or U9253 (N_9253,N_8695,N_8099);
nand U9254 (N_9254,N_8908,N_8715);
nand U9255 (N_9255,N_8570,N_8671);
nand U9256 (N_9256,N_8194,N_8841);
and U9257 (N_9257,N_8864,N_8123);
and U9258 (N_9258,N_8357,N_8412);
or U9259 (N_9259,N_8667,N_8278);
xor U9260 (N_9260,N_8484,N_8004);
nand U9261 (N_9261,N_8842,N_8102);
xor U9262 (N_9262,N_8654,N_8709);
nand U9263 (N_9263,N_8103,N_8796);
or U9264 (N_9264,N_8234,N_8057);
nand U9265 (N_9265,N_8072,N_8973);
xnor U9266 (N_9266,N_8422,N_8318);
nand U9267 (N_9267,N_8116,N_8520);
nor U9268 (N_9268,N_8917,N_8688);
or U9269 (N_9269,N_8345,N_8358);
or U9270 (N_9270,N_8062,N_8233);
and U9271 (N_9271,N_8047,N_8724);
or U9272 (N_9272,N_8749,N_8339);
nand U9273 (N_9273,N_8551,N_8824);
nand U9274 (N_9274,N_8600,N_8259);
nand U9275 (N_9275,N_8611,N_8693);
or U9276 (N_9276,N_8515,N_8039);
or U9277 (N_9277,N_8979,N_8936);
nand U9278 (N_9278,N_8164,N_8044);
nand U9279 (N_9279,N_8083,N_8449);
or U9280 (N_9280,N_8994,N_8404);
nor U9281 (N_9281,N_8705,N_8799);
nand U9282 (N_9282,N_8367,N_8110);
or U9283 (N_9283,N_8710,N_8801);
nor U9284 (N_9284,N_8962,N_8321);
nor U9285 (N_9285,N_8804,N_8953);
nand U9286 (N_9286,N_8686,N_8846);
and U9287 (N_9287,N_8320,N_8716);
nor U9288 (N_9288,N_8816,N_8672);
nand U9289 (N_9289,N_8183,N_8650);
and U9290 (N_9290,N_8597,N_8870);
nand U9291 (N_9291,N_8157,N_8325);
nor U9292 (N_9292,N_8920,N_8137);
nor U9293 (N_9293,N_8172,N_8981);
nand U9294 (N_9294,N_8901,N_8772);
xor U9295 (N_9295,N_8735,N_8706);
and U9296 (N_9296,N_8250,N_8191);
and U9297 (N_9297,N_8220,N_8254);
nand U9298 (N_9298,N_8022,N_8617);
or U9299 (N_9299,N_8109,N_8741);
and U9300 (N_9300,N_8664,N_8427);
and U9301 (N_9301,N_8789,N_8605);
nand U9302 (N_9302,N_8076,N_8843);
xor U9303 (N_9303,N_8027,N_8210);
nand U9304 (N_9304,N_8012,N_8553);
nand U9305 (N_9305,N_8235,N_8742);
xor U9306 (N_9306,N_8866,N_8714);
and U9307 (N_9307,N_8590,N_8580);
nor U9308 (N_9308,N_8018,N_8632);
and U9309 (N_9309,N_8322,N_8173);
xnor U9310 (N_9310,N_8835,N_8984);
or U9311 (N_9311,N_8681,N_8215);
and U9312 (N_9312,N_8050,N_8685);
or U9313 (N_9313,N_8928,N_8299);
nand U9314 (N_9314,N_8112,N_8213);
and U9315 (N_9315,N_8834,N_8142);
xnor U9316 (N_9316,N_8807,N_8798);
or U9317 (N_9317,N_8262,N_8492);
and U9318 (N_9318,N_8049,N_8053);
or U9319 (N_9319,N_8615,N_8970);
nand U9320 (N_9320,N_8636,N_8993);
nand U9321 (N_9321,N_8523,N_8147);
and U9322 (N_9322,N_8481,N_8912);
nor U9323 (N_9323,N_8498,N_8424);
or U9324 (N_9324,N_8923,N_8902);
and U9325 (N_9325,N_8038,N_8129);
xor U9326 (N_9326,N_8476,N_8865);
or U9327 (N_9327,N_8227,N_8527);
and U9328 (N_9328,N_8692,N_8315);
xnor U9329 (N_9329,N_8641,N_8002);
nor U9330 (N_9330,N_8925,N_8733);
nand U9331 (N_9331,N_8361,N_8241);
and U9332 (N_9332,N_8188,N_8690);
and U9333 (N_9333,N_8932,N_8942);
or U9334 (N_9334,N_8256,N_8088);
or U9335 (N_9335,N_8212,N_8206);
and U9336 (N_9336,N_8634,N_8379);
nor U9337 (N_9337,N_8488,N_8612);
or U9338 (N_9338,N_8479,N_8764);
nor U9339 (N_9339,N_8196,N_8223);
nand U9340 (N_9340,N_8820,N_8885);
and U9341 (N_9341,N_8120,N_8092);
or U9342 (N_9342,N_8011,N_8831);
or U9343 (N_9343,N_8960,N_8421);
nand U9344 (N_9344,N_8929,N_8079);
nor U9345 (N_9345,N_8140,N_8875);
nand U9346 (N_9346,N_8391,N_8663);
nand U9347 (N_9347,N_8511,N_8077);
nand U9348 (N_9348,N_8900,N_8976);
nand U9349 (N_9349,N_8307,N_8500);
or U9350 (N_9350,N_8585,N_8677);
and U9351 (N_9351,N_8645,N_8810);
or U9352 (N_9352,N_8747,N_8707);
nand U9353 (N_9353,N_8121,N_8651);
xnor U9354 (N_9354,N_8599,N_8420);
or U9355 (N_9355,N_8933,N_8921);
xnor U9356 (N_9356,N_8948,N_8545);
nand U9357 (N_9357,N_8480,N_8774);
nand U9358 (N_9358,N_8085,N_8549);
nor U9359 (N_9359,N_8457,N_8679);
nand U9360 (N_9360,N_8726,N_8111);
and U9361 (N_9361,N_8187,N_8918);
nor U9362 (N_9362,N_8642,N_8797);
or U9363 (N_9363,N_8862,N_8528);
and U9364 (N_9364,N_8168,N_8437);
or U9365 (N_9365,N_8193,N_8517);
and U9366 (N_9366,N_8485,N_8604);
nor U9367 (N_9367,N_8855,N_8163);
nand U9368 (N_9368,N_8003,N_8652);
and U9369 (N_9369,N_8616,N_8777);
nand U9370 (N_9370,N_8434,N_8539);
or U9371 (N_9371,N_8060,N_8972);
nor U9372 (N_9372,N_8525,N_8655);
or U9373 (N_9373,N_8308,N_8045);
nand U9374 (N_9374,N_8237,N_8405);
or U9375 (N_9375,N_8334,N_8883);
or U9376 (N_9376,N_8456,N_8471);
nand U9377 (N_9377,N_8486,N_8704);
or U9378 (N_9378,N_8093,N_8010);
nand U9379 (N_9379,N_8734,N_8073);
xnor U9380 (N_9380,N_8990,N_8569);
or U9381 (N_9381,N_8008,N_8653);
nor U9382 (N_9382,N_8125,N_8762);
or U9383 (N_9383,N_8000,N_8055);
and U9384 (N_9384,N_8406,N_8064);
nand U9385 (N_9385,N_8727,N_8648);
nand U9386 (N_9386,N_8344,N_8670);
nand U9387 (N_9387,N_8238,N_8675);
nor U9388 (N_9388,N_8847,N_8647);
or U9389 (N_9389,N_8314,N_8880);
or U9390 (N_9390,N_8416,N_8756);
nand U9391 (N_9391,N_8678,N_8938);
nor U9392 (N_9392,N_8395,N_8698);
nor U9393 (N_9393,N_8776,N_8556);
nor U9394 (N_9394,N_8030,N_8532);
nand U9395 (N_9395,N_8153,N_8598);
or U9396 (N_9396,N_8854,N_8086);
xnor U9397 (N_9397,N_8637,N_8489);
nor U9398 (N_9398,N_8888,N_8330);
nor U9399 (N_9399,N_8795,N_8384);
or U9400 (N_9400,N_8268,N_8101);
and U9401 (N_9401,N_8644,N_8983);
nand U9402 (N_9402,N_8802,N_8219);
nand U9403 (N_9403,N_8373,N_8683);
and U9404 (N_9404,N_8638,N_8477);
nand U9405 (N_9405,N_8374,N_8516);
nand U9406 (N_9406,N_8547,N_8462);
xor U9407 (N_9407,N_8442,N_8555);
xor U9408 (N_9408,N_8987,N_8522);
xnor U9409 (N_9409,N_8150,N_8151);
nand U9410 (N_9410,N_8745,N_8916);
nor U9411 (N_9411,N_8546,N_8755);
and U9412 (N_9412,N_8790,N_8581);
and U9413 (N_9413,N_8950,N_8620);
nor U9414 (N_9414,N_8505,N_8947);
or U9415 (N_9415,N_8721,N_8850);
or U9416 (N_9416,N_8927,N_8451);
and U9417 (N_9417,N_8222,N_8114);
nor U9418 (N_9418,N_8583,N_8366);
nor U9419 (N_9419,N_8779,N_8758);
xor U9420 (N_9420,N_8723,N_8460);
or U9421 (N_9421,N_8533,N_8643);
nand U9422 (N_9422,N_8813,N_8702);
or U9423 (N_9423,N_8944,N_8181);
nand U9424 (N_9424,N_8729,N_8408);
nor U9425 (N_9425,N_8501,N_8728);
or U9426 (N_9426,N_8763,N_8624);
and U9427 (N_9427,N_8264,N_8251);
xor U9428 (N_9428,N_8393,N_8398);
nand U9429 (N_9429,N_8376,N_8201);
and U9430 (N_9430,N_8571,N_8739);
and U9431 (N_9431,N_8329,N_8159);
and U9432 (N_9432,N_8301,N_8025);
nand U9433 (N_9433,N_8182,N_8070);
nor U9434 (N_9434,N_8260,N_8676);
or U9435 (N_9435,N_8689,N_8785);
nor U9436 (N_9436,N_8265,N_8208);
and U9437 (N_9437,N_8300,N_8467);
nor U9438 (N_9438,N_8596,N_8640);
or U9439 (N_9439,N_8369,N_8255);
or U9440 (N_9440,N_8700,N_8054);
or U9441 (N_9441,N_8752,N_8773);
nor U9442 (N_9442,N_8519,N_8496);
and U9443 (N_9443,N_8863,N_8939);
nor U9444 (N_9444,N_8098,N_8941);
xor U9445 (N_9445,N_8513,N_8200);
nand U9446 (N_9446,N_8452,N_8623);
xnor U9447 (N_9447,N_8558,N_8924);
or U9448 (N_9448,N_8205,N_8543);
nand U9449 (N_9449,N_8829,N_8780);
xnor U9450 (N_9450,N_8180,N_8951);
and U9451 (N_9451,N_8858,N_8658);
or U9452 (N_9452,N_8158,N_8438);
nor U9453 (N_9453,N_8400,N_8997);
and U9454 (N_9454,N_8966,N_8131);
nand U9455 (N_9455,N_8872,N_8899);
or U9456 (N_9456,N_8886,N_8833);
xor U9457 (N_9457,N_8118,N_8740);
nand U9458 (N_9458,N_8876,N_8207);
xor U9459 (N_9459,N_8340,N_8629);
xnor U9460 (N_9460,N_8472,N_8892);
nand U9461 (N_9461,N_8124,N_8579);
and U9462 (N_9462,N_8184,N_8293);
or U9463 (N_9463,N_8988,N_8907);
and U9464 (N_9464,N_8668,N_8720);
or U9465 (N_9465,N_8840,N_8094);
xor U9466 (N_9466,N_8160,N_8248);
nand U9467 (N_9467,N_8463,N_8995);
and U9468 (N_9468,N_8687,N_8897);
or U9469 (N_9469,N_8961,N_8258);
and U9470 (N_9470,N_8821,N_8470);
nor U9471 (N_9471,N_8294,N_8977);
or U9472 (N_9472,N_8860,N_8224);
nand U9473 (N_9473,N_8052,N_8680);
and U9474 (N_9474,N_8499,N_8280);
or U9475 (N_9475,N_8507,N_8005);
nand U9476 (N_9476,N_8825,N_8544);
nor U9477 (N_9477,N_8178,N_8415);
and U9478 (N_9478,N_8459,N_8788);
nor U9479 (N_9479,N_8333,N_8133);
and U9480 (N_9480,N_8784,N_8827);
or U9481 (N_9481,N_8006,N_8464);
or U9482 (N_9482,N_8906,N_8190);
and U9483 (N_9483,N_8043,N_8922);
and U9484 (N_9484,N_8986,N_8418);
nand U9485 (N_9485,N_8035,N_8730);
and U9486 (N_9486,N_8601,N_8805);
and U9487 (N_9487,N_8541,N_8560);
nand U9488 (N_9488,N_8061,N_8362);
nor U9489 (N_9489,N_8811,N_8887);
or U9490 (N_9490,N_8701,N_8822);
nand U9491 (N_9491,N_8954,N_8691);
or U9492 (N_9492,N_8699,N_8946);
nor U9493 (N_9493,N_8659,N_8674);
nor U9494 (N_9494,N_8722,N_8162);
nand U9495 (N_9495,N_8478,N_8606);
and U9496 (N_9496,N_8134,N_8243);
nand U9497 (N_9497,N_8491,N_8538);
nor U9498 (N_9498,N_8737,N_8754);
or U9499 (N_9499,N_8149,N_8849);
nand U9500 (N_9500,N_8039,N_8139);
or U9501 (N_9501,N_8294,N_8031);
and U9502 (N_9502,N_8752,N_8282);
or U9503 (N_9503,N_8754,N_8834);
or U9504 (N_9504,N_8716,N_8270);
or U9505 (N_9505,N_8151,N_8621);
nand U9506 (N_9506,N_8466,N_8793);
and U9507 (N_9507,N_8908,N_8574);
or U9508 (N_9508,N_8858,N_8319);
and U9509 (N_9509,N_8164,N_8788);
or U9510 (N_9510,N_8060,N_8057);
and U9511 (N_9511,N_8015,N_8488);
nand U9512 (N_9512,N_8385,N_8560);
nand U9513 (N_9513,N_8653,N_8181);
nand U9514 (N_9514,N_8058,N_8216);
nand U9515 (N_9515,N_8902,N_8551);
or U9516 (N_9516,N_8275,N_8118);
nor U9517 (N_9517,N_8229,N_8768);
and U9518 (N_9518,N_8887,N_8544);
nor U9519 (N_9519,N_8674,N_8150);
nor U9520 (N_9520,N_8584,N_8315);
nor U9521 (N_9521,N_8628,N_8529);
or U9522 (N_9522,N_8680,N_8879);
nor U9523 (N_9523,N_8336,N_8579);
and U9524 (N_9524,N_8755,N_8117);
nand U9525 (N_9525,N_8519,N_8969);
nor U9526 (N_9526,N_8119,N_8132);
nand U9527 (N_9527,N_8150,N_8018);
xnor U9528 (N_9528,N_8779,N_8783);
nand U9529 (N_9529,N_8138,N_8074);
and U9530 (N_9530,N_8755,N_8041);
or U9531 (N_9531,N_8578,N_8842);
nor U9532 (N_9532,N_8592,N_8319);
nor U9533 (N_9533,N_8994,N_8442);
nor U9534 (N_9534,N_8395,N_8617);
nor U9535 (N_9535,N_8651,N_8566);
or U9536 (N_9536,N_8934,N_8501);
nor U9537 (N_9537,N_8142,N_8992);
xnor U9538 (N_9538,N_8095,N_8058);
or U9539 (N_9539,N_8632,N_8388);
and U9540 (N_9540,N_8960,N_8149);
xnor U9541 (N_9541,N_8524,N_8924);
nand U9542 (N_9542,N_8111,N_8064);
nand U9543 (N_9543,N_8562,N_8095);
nand U9544 (N_9544,N_8837,N_8788);
or U9545 (N_9545,N_8886,N_8982);
nor U9546 (N_9546,N_8496,N_8841);
or U9547 (N_9547,N_8038,N_8903);
nor U9548 (N_9548,N_8983,N_8728);
nor U9549 (N_9549,N_8975,N_8075);
and U9550 (N_9550,N_8310,N_8407);
nor U9551 (N_9551,N_8362,N_8021);
or U9552 (N_9552,N_8180,N_8279);
nand U9553 (N_9553,N_8527,N_8305);
nor U9554 (N_9554,N_8527,N_8454);
xor U9555 (N_9555,N_8393,N_8739);
or U9556 (N_9556,N_8318,N_8293);
or U9557 (N_9557,N_8300,N_8357);
nor U9558 (N_9558,N_8518,N_8207);
and U9559 (N_9559,N_8784,N_8500);
and U9560 (N_9560,N_8994,N_8121);
nor U9561 (N_9561,N_8424,N_8815);
nor U9562 (N_9562,N_8444,N_8017);
nand U9563 (N_9563,N_8227,N_8429);
and U9564 (N_9564,N_8745,N_8153);
or U9565 (N_9565,N_8983,N_8592);
nor U9566 (N_9566,N_8710,N_8422);
and U9567 (N_9567,N_8875,N_8306);
or U9568 (N_9568,N_8608,N_8538);
nand U9569 (N_9569,N_8093,N_8855);
or U9570 (N_9570,N_8946,N_8940);
nand U9571 (N_9571,N_8045,N_8271);
xor U9572 (N_9572,N_8805,N_8533);
nand U9573 (N_9573,N_8565,N_8206);
and U9574 (N_9574,N_8481,N_8882);
and U9575 (N_9575,N_8414,N_8939);
nand U9576 (N_9576,N_8548,N_8397);
or U9577 (N_9577,N_8106,N_8718);
or U9578 (N_9578,N_8595,N_8377);
xnor U9579 (N_9579,N_8610,N_8495);
and U9580 (N_9580,N_8498,N_8822);
nand U9581 (N_9581,N_8852,N_8097);
nand U9582 (N_9582,N_8803,N_8928);
or U9583 (N_9583,N_8310,N_8719);
nor U9584 (N_9584,N_8064,N_8169);
nor U9585 (N_9585,N_8837,N_8126);
or U9586 (N_9586,N_8230,N_8488);
and U9587 (N_9587,N_8315,N_8296);
or U9588 (N_9588,N_8949,N_8446);
nand U9589 (N_9589,N_8241,N_8808);
or U9590 (N_9590,N_8967,N_8773);
nand U9591 (N_9591,N_8612,N_8373);
nand U9592 (N_9592,N_8037,N_8733);
nor U9593 (N_9593,N_8377,N_8641);
and U9594 (N_9594,N_8680,N_8413);
and U9595 (N_9595,N_8657,N_8960);
nor U9596 (N_9596,N_8075,N_8344);
nor U9597 (N_9597,N_8240,N_8271);
or U9598 (N_9598,N_8869,N_8788);
and U9599 (N_9599,N_8373,N_8904);
or U9600 (N_9600,N_8458,N_8181);
nor U9601 (N_9601,N_8781,N_8008);
or U9602 (N_9602,N_8481,N_8511);
and U9603 (N_9603,N_8769,N_8308);
nand U9604 (N_9604,N_8074,N_8516);
or U9605 (N_9605,N_8601,N_8357);
nor U9606 (N_9606,N_8708,N_8920);
and U9607 (N_9607,N_8603,N_8327);
nor U9608 (N_9608,N_8075,N_8262);
nor U9609 (N_9609,N_8031,N_8638);
nor U9610 (N_9610,N_8500,N_8866);
xnor U9611 (N_9611,N_8416,N_8776);
xnor U9612 (N_9612,N_8116,N_8238);
nor U9613 (N_9613,N_8704,N_8246);
and U9614 (N_9614,N_8919,N_8638);
and U9615 (N_9615,N_8066,N_8331);
nor U9616 (N_9616,N_8292,N_8174);
nor U9617 (N_9617,N_8701,N_8973);
or U9618 (N_9618,N_8909,N_8868);
or U9619 (N_9619,N_8278,N_8296);
or U9620 (N_9620,N_8363,N_8177);
or U9621 (N_9621,N_8359,N_8057);
and U9622 (N_9622,N_8762,N_8794);
or U9623 (N_9623,N_8214,N_8301);
and U9624 (N_9624,N_8185,N_8245);
nand U9625 (N_9625,N_8095,N_8681);
nand U9626 (N_9626,N_8805,N_8864);
xnor U9627 (N_9627,N_8199,N_8567);
nor U9628 (N_9628,N_8308,N_8780);
and U9629 (N_9629,N_8675,N_8817);
nand U9630 (N_9630,N_8663,N_8182);
and U9631 (N_9631,N_8371,N_8804);
or U9632 (N_9632,N_8567,N_8661);
and U9633 (N_9633,N_8220,N_8457);
xnor U9634 (N_9634,N_8320,N_8785);
nor U9635 (N_9635,N_8501,N_8157);
nor U9636 (N_9636,N_8619,N_8204);
and U9637 (N_9637,N_8349,N_8792);
xor U9638 (N_9638,N_8111,N_8086);
xor U9639 (N_9639,N_8493,N_8465);
nor U9640 (N_9640,N_8778,N_8248);
nand U9641 (N_9641,N_8248,N_8984);
and U9642 (N_9642,N_8289,N_8658);
nor U9643 (N_9643,N_8887,N_8321);
and U9644 (N_9644,N_8575,N_8027);
and U9645 (N_9645,N_8487,N_8446);
nand U9646 (N_9646,N_8779,N_8688);
nor U9647 (N_9647,N_8909,N_8125);
or U9648 (N_9648,N_8751,N_8029);
nand U9649 (N_9649,N_8118,N_8474);
nor U9650 (N_9650,N_8119,N_8665);
nand U9651 (N_9651,N_8176,N_8613);
or U9652 (N_9652,N_8803,N_8866);
or U9653 (N_9653,N_8854,N_8719);
xnor U9654 (N_9654,N_8762,N_8246);
nor U9655 (N_9655,N_8675,N_8072);
or U9656 (N_9656,N_8296,N_8270);
and U9657 (N_9657,N_8861,N_8205);
nor U9658 (N_9658,N_8869,N_8366);
xnor U9659 (N_9659,N_8375,N_8298);
or U9660 (N_9660,N_8377,N_8033);
nand U9661 (N_9661,N_8320,N_8729);
nand U9662 (N_9662,N_8084,N_8973);
nand U9663 (N_9663,N_8358,N_8156);
nor U9664 (N_9664,N_8468,N_8203);
nand U9665 (N_9665,N_8171,N_8915);
nor U9666 (N_9666,N_8919,N_8591);
xnor U9667 (N_9667,N_8237,N_8567);
or U9668 (N_9668,N_8281,N_8628);
nand U9669 (N_9669,N_8295,N_8674);
nand U9670 (N_9670,N_8461,N_8040);
nand U9671 (N_9671,N_8271,N_8842);
nand U9672 (N_9672,N_8382,N_8723);
nand U9673 (N_9673,N_8211,N_8401);
and U9674 (N_9674,N_8032,N_8705);
and U9675 (N_9675,N_8042,N_8980);
and U9676 (N_9676,N_8082,N_8257);
or U9677 (N_9677,N_8959,N_8399);
and U9678 (N_9678,N_8941,N_8727);
or U9679 (N_9679,N_8058,N_8817);
nor U9680 (N_9680,N_8367,N_8150);
or U9681 (N_9681,N_8280,N_8552);
or U9682 (N_9682,N_8545,N_8483);
or U9683 (N_9683,N_8258,N_8584);
nand U9684 (N_9684,N_8610,N_8386);
and U9685 (N_9685,N_8930,N_8070);
or U9686 (N_9686,N_8867,N_8131);
nor U9687 (N_9687,N_8393,N_8654);
nand U9688 (N_9688,N_8132,N_8163);
nand U9689 (N_9689,N_8522,N_8400);
nor U9690 (N_9690,N_8535,N_8012);
and U9691 (N_9691,N_8272,N_8887);
nor U9692 (N_9692,N_8939,N_8513);
and U9693 (N_9693,N_8962,N_8474);
nor U9694 (N_9694,N_8773,N_8762);
or U9695 (N_9695,N_8603,N_8782);
xor U9696 (N_9696,N_8226,N_8155);
nand U9697 (N_9697,N_8361,N_8900);
nand U9698 (N_9698,N_8821,N_8639);
nor U9699 (N_9699,N_8378,N_8924);
nor U9700 (N_9700,N_8693,N_8265);
or U9701 (N_9701,N_8699,N_8992);
xor U9702 (N_9702,N_8771,N_8919);
xor U9703 (N_9703,N_8129,N_8384);
xnor U9704 (N_9704,N_8020,N_8440);
nand U9705 (N_9705,N_8584,N_8455);
or U9706 (N_9706,N_8833,N_8512);
nor U9707 (N_9707,N_8147,N_8859);
and U9708 (N_9708,N_8617,N_8934);
nor U9709 (N_9709,N_8834,N_8020);
nor U9710 (N_9710,N_8887,N_8530);
or U9711 (N_9711,N_8705,N_8685);
and U9712 (N_9712,N_8994,N_8247);
nand U9713 (N_9713,N_8487,N_8100);
nor U9714 (N_9714,N_8651,N_8188);
nor U9715 (N_9715,N_8503,N_8064);
and U9716 (N_9716,N_8791,N_8534);
nor U9717 (N_9717,N_8334,N_8335);
and U9718 (N_9718,N_8887,N_8624);
nand U9719 (N_9719,N_8564,N_8733);
or U9720 (N_9720,N_8531,N_8384);
nor U9721 (N_9721,N_8713,N_8187);
or U9722 (N_9722,N_8327,N_8881);
nand U9723 (N_9723,N_8702,N_8666);
and U9724 (N_9724,N_8836,N_8129);
nor U9725 (N_9725,N_8932,N_8375);
nor U9726 (N_9726,N_8585,N_8054);
nor U9727 (N_9727,N_8799,N_8566);
and U9728 (N_9728,N_8682,N_8041);
nand U9729 (N_9729,N_8055,N_8150);
nor U9730 (N_9730,N_8696,N_8003);
and U9731 (N_9731,N_8807,N_8182);
or U9732 (N_9732,N_8130,N_8682);
or U9733 (N_9733,N_8842,N_8749);
or U9734 (N_9734,N_8310,N_8969);
nor U9735 (N_9735,N_8200,N_8694);
or U9736 (N_9736,N_8396,N_8407);
nand U9737 (N_9737,N_8433,N_8157);
xor U9738 (N_9738,N_8464,N_8927);
nor U9739 (N_9739,N_8106,N_8981);
nand U9740 (N_9740,N_8044,N_8196);
and U9741 (N_9741,N_8624,N_8325);
nor U9742 (N_9742,N_8891,N_8762);
nor U9743 (N_9743,N_8761,N_8550);
nand U9744 (N_9744,N_8815,N_8285);
or U9745 (N_9745,N_8370,N_8467);
nand U9746 (N_9746,N_8598,N_8489);
or U9747 (N_9747,N_8285,N_8219);
xnor U9748 (N_9748,N_8786,N_8724);
and U9749 (N_9749,N_8815,N_8366);
nand U9750 (N_9750,N_8301,N_8578);
or U9751 (N_9751,N_8060,N_8205);
or U9752 (N_9752,N_8932,N_8002);
nand U9753 (N_9753,N_8290,N_8657);
and U9754 (N_9754,N_8254,N_8845);
nor U9755 (N_9755,N_8547,N_8929);
and U9756 (N_9756,N_8415,N_8452);
nand U9757 (N_9757,N_8356,N_8628);
nand U9758 (N_9758,N_8626,N_8069);
or U9759 (N_9759,N_8811,N_8357);
nand U9760 (N_9760,N_8748,N_8004);
nand U9761 (N_9761,N_8172,N_8610);
nor U9762 (N_9762,N_8147,N_8371);
nand U9763 (N_9763,N_8160,N_8988);
nor U9764 (N_9764,N_8205,N_8445);
nand U9765 (N_9765,N_8314,N_8771);
and U9766 (N_9766,N_8815,N_8848);
xnor U9767 (N_9767,N_8322,N_8467);
nor U9768 (N_9768,N_8053,N_8057);
or U9769 (N_9769,N_8931,N_8107);
nor U9770 (N_9770,N_8511,N_8360);
nor U9771 (N_9771,N_8567,N_8952);
xnor U9772 (N_9772,N_8975,N_8247);
nand U9773 (N_9773,N_8039,N_8523);
and U9774 (N_9774,N_8009,N_8726);
and U9775 (N_9775,N_8472,N_8376);
nor U9776 (N_9776,N_8334,N_8425);
or U9777 (N_9777,N_8120,N_8634);
and U9778 (N_9778,N_8386,N_8899);
and U9779 (N_9779,N_8505,N_8444);
or U9780 (N_9780,N_8776,N_8117);
nand U9781 (N_9781,N_8340,N_8634);
nor U9782 (N_9782,N_8139,N_8121);
or U9783 (N_9783,N_8449,N_8154);
and U9784 (N_9784,N_8082,N_8752);
xnor U9785 (N_9785,N_8955,N_8074);
nand U9786 (N_9786,N_8175,N_8381);
and U9787 (N_9787,N_8630,N_8424);
and U9788 (N_9788,N_8009,N_8910);
nor U9789 (N_9789,N_8144,N_8681);
and U9790 (N_9790,N_8757,N_8737);
nor U9791 (N_9791,N_8652,N_8899);
and U9792 (N_9792,N_8503,N_8914);
or U9793 (N_9793,N_8948,N_8705);
nor U9794 (N_9794,N_8774,N_8609);
nand U9795 (N_9795,N_8271,N_8412);
or U9796 (N_9796,N_8971,N_8715);
nand U9797 (N_9797,N_8004,N_8405);
nor U9798 (N_9798,N_8647,N_8452);
nor U9799 (N_9799,N_8827,N_8141);
or U9800 (N_9800,N_8415,N_8244);
nor U9801 (N_9801,N_8819,N_8402);
xnor U9802 (N_9802,N_8022,N_8573);
and U9803 (N_9803,N_8489,N_8103);
xnor U9804 (N_9804,N_8228,N_8160);
nor U9805 (N_9805,N_8853,N_8527);
nand U9806 (N_9806,N_8353,N_8863);
nand U9807 (N_9807,N_8248,N_8166);
nand U9808 (N_9808,N_8048,N_8463);
nand U9809 (N_9809,N_8424,N_8473);
nand U9810 (N_9810,N_8137,N_8755);
and U9811 (N_9811,N_8929,N_8912);
nand U9812 (N_9812,N_8704,N_8019);
nand U9813 (N_9813,N_8761,N_8907);
nand U9814 (N_9814,N_8500,N_8176);
and U9815 (N_9815,N_8901,N_8553);
nand U9816 (N_9816,N_8495,N_8970);
xnor U9817 (N_9817,N_8235,N_8816);
or U9818 (N_9818,N_8152,N_8073);
and U9819 (N_9819,N_8928,N_8100);
xnor U9820 (N_9820,N_8959,N_8729);
nand U9821 (N_9821,N_8724,N_8169);
or U9822 (N_9822,N_8806,N_8091);
or U9823 (N_9823,N_8671,N_8459);
nor U9824 (N_9824,N_8054,N_8574);
nor U9825 (N_9825,N_8688,N_8031);
or U9826 (N_9826,N_8063,N_8002);
nand U9827 (N_9827,N_8554,N_8634);
nor U9828 (N_9828,N_8977,N_8071);
nand U9829 (N_9829,N_8680,N_8402);
or U9830 (N_9830,N_8048,N_8618);
nand U9831 (N_9831,N_8002,N_8087);
nor U9832 (N_9832,N_8581,N_8707);
and U9833 (N_9833,N_8669,N_8780);
or U9834 (N_9834,N_8267,N_8042);
nor U9835 (N_9835,N_8264,N_8988);
nor U9836 (N_9836,N_8592,N_8725);
xor U9837 (N_9837,N_8899,N_8779);
nand U9838 (N_9838,N_8748,N_8577);
nand U9839 (N_9839,N_8875,N_8087);
nor U9840 (N_9840,N_8730,N_8026);
and U9841 (N_9841,N_8990,N_8958);
or U9842 (N_9842,N_8601,N_8184);
nand U9843 (N_9843,N_8621,N_8167);
nand U9844 (N_9844,N_8049,N_8054);
nor U9845 (N_9845,N_8517,N_8383);
or U9846 (N_9846,N_8407,N_8604);
nand U9847 (N_9847,N_8304,N_8122);
nand U9848 (N_9848,N_8399,N_8823);
nand U9849 (N_9849,N_8818,N_8704);
nor U9850 (N_9850,N_8832,N_8569);
and U9851 (N_9851,N_8150,N_8352);
nand U9852 (N_9852,N_8774,N_8519);
nor U9853 (N_9853,N_8633,N_8453);
nor U9854 (N_9854,N_8593,N_8185);
and U9855 (N_9855,N_8777,N_8746);
nand U9856 (N_9856,N_8639,N_8565);
nand U9857 (N_9857,N_8162,N_8053);
nand U9858 (N_9858,N_8541,N_8831);
or U9859 (N_9859,N_8467,N_8079);
or U9860 (N_9860,N_8781,N_8754);
nor U9861 (N_9861,N_8117,N_8386);
or U9862 (N_9862,N_8403,N_8301);
and U9863 (N_9863,N_8994,N_8262);
and U9864 (N_9864,N_8709,N_8048);
or U9865 (N_9865,N_8518,N_8640);
nand U9866 (N_9866,N_8452,N_8468);
nor U9867 (N_9867,N_8270,N_8290);
nand U9868 (N_9868,N_8976,N_8129);
and U9869 (N_9869,N_8807,N_8256);
nor U9870 (N_9870,N_8845,N_8335);
or U9871 (N_9871,N_8025,N_8927);
nor U9872 (N_9872,N_8346,N_8876);
nand U9873 (N_9873,N_8661,N_8100);
nand U9874 (N_9874,N_8025,N_8259);
nor U9875 (N_9875,N_8319,N_8837);
or U9876 (N_9876,N_8582,N_8085);
nand U9877 (N_9877,N_8326,N_8265);
and U9878 (N_9878,N_8751,N_8150);
nor U9879 (N_9879,N_8561,N_8838);
xor U9880 (N_9880,N_8271,N_8332);
and U9881 (N_9881,N_8504,N_8498);
or U9882 (N_9882,N_8024,N_8583);
and U9883 (N_9883,N_8341,N_8863);
nor U9884 (N_9884,N_8862,N_8406);
nor U9885 (N_9885,N_8382,N_8657);
xnor U9886 (N_9886,N_8165,N_8675);
nand U9887 (N_9887,N_8839,N_8905);
or U9888 (N_9888,N_8817,N_8144);
nor U9889 (N_9889,N_8378,N_8678);
or U9890 (N_9890,N_8856,N_8620);
and U9891 (N_9891,N_8112,N_8542);
and U9892 (N_9892,N_8813,N_8912);
nand U9893 (N_9893,N_8395,N_8625);
and U9894 (N_9894,N_8781,N_8984);
or U9895 (N_9895,N_8413,N_8555);
nand U9896 (N_9896,N_8979,N_8001);
and U9897 (N_9897,N_8665,N_8323);
nor U9898 (N_9898,N_8000,N_8328);
nor U9899 (N_9899,N_8649,N_8301);
or U9900 (N_9900,N_8691,N_8993);
nand U9901 (N_9901,N_8474,N_8808);
xor U9902 (N_9902,N_8166,N_8479);
or U9903 (N_9903,N_8840,N_8179);
nor U9904 (N_9904,N_8928,N_8043);
or U9905 (N_9905,N_8520,N_8257);
and U9906 (N_9906,N_8430,N_8226);
and U9907 (N_9907,N_8073,N_8450);
nor U9908 (N_9908,N_8630,N_8184);
and U9909 (N_9909,N_8956,N_8831);
nand U9910 (N_9910,N_8062,N_8770);
or U9911 (N_9911,N_8837,N_8950);
nand U9912 (N_9912,N_8199,N_8776);
xor U9913 (N_9913,N_8536,N_8912);
nor U9914 (N_9914,N_8946,N_8824);
or U9915 (N_9915,N_8247,N_8001);
or U9916 (N_9916,N_8047,N_8629);
and U9917 (N_9917,N_8122,N_8147);
nor U9918 (N_9918,N_8319,N_8308);
and U9919 (N_9919,N_8894,N_8715);
nand U9920 (N_9920,N_8024,N_8950);
or U9921 (N_9921,N_8621,N_8158);
nand U9922 (N_9922,N_8020,N_8755);
or U9923 (N_9923,N_8263,N_8107);
and U9924 (N_9924,N_8231,N_8034);
and U9925 (N_9925,N_8976,N_8181);
nor U9926 (N_9926,N_8670,N_8694);
xnor U9927 (N_9927,N_8249,N_8710);
nor U9928 (N_9928,N_8377,N_8730);
or U9929 (N_9929,N_8770,N_8410);
nor U9930 (N_9930,N_8944,N_8799);
or U9931 (N_9931,N_8043,N_8074);
or U9932 (N_9932,N_8244,N_8332);
nand U9933 (N_9933,N_8487,N_8879);
nor U9934 (N_9934,N_8372,N_8299);
or U9935 (N_9935,N_8560,N_8532);
or U9936 (N_9936,N_8629,N_8559);
nand U9937 (N_9937,N_8358,N_8216);
and U9938 (N_9938,N_8158,N_8518);
and U9939 (N_9939,N_8263,N_8560);
and U9940 (N_9940,N_8777,N_8779);
or U9941 (N_9941,N_8722,N_8091);
or U9942 (N_9942,N_8524,N_8688);
and U9943 (N_9943,N_8853,N_8641);
or U9944 (N_9944,N_8410,N_8523);
xnor U9945 (N_9945,N_8028,N_8011);
nor U9946 (N_9946,N_8160,N_8252);
nor U9947 (N_9947,N_8633,N_8945);
xnor U9948 (N_9948,N_8801,N_8707);
nor U9949 (N_9949,N_8947,N_8456);
or U9950 (N_9950,N_8875,N_8912);
or U9951 (N_9951,N_8527,N_8955);
and U9952 (N_9952,N_8301,N_8874);
nand U9953 (N_9953,N_8961,N_8473);
xor U9954 (N_9954,N_8672,N_8620);
nor U9955 (N_9955,N_8953,N_8609);
nor U9956 (N_9956,N_8454,N_8229);
or U9957 (N_9957,N_8997,N_8869);
xnor U9958 (N_9958,N_8772,N_8186);
and U9959 (N_9959,N_8782,N_8131);
nor U9960 (N_9960,N_8912,N_8320);
and U9961 (N_9961,N_8491,N_8855);
or U9962 (N_9962,N_8912,N_8666);
nor U9963 (N_9963,N_8219,N_8016);
and U9964 (N_9964,N_8427,N_8630);
nor U9965 (N_9965,N_8325,N_8283);
nand U9966 (N_9966,N_8499,N_8713);
nor U9967 (N_9967,N_8731,N_8683);
or U9968 (N_9968,N_8179,N_8077);
or U9969 (N_9969,N_8089,N_8027);
nor U9970 (N_9970,N_8601,N_8686);
nor U9971 (N_9971,N_8696,N_8578);
or U9972 (N_9972,N_8780,N_8859);
and U9973 (N_9973,N_8062,N_8535);
xor U9974 (N_9974,N_8054,N_8386);
xnor U9975 (N_9975,N_8588,N_8249);
and U9976 (N_9976,N_8327,N_8308);
nor U9977 (N_9977,N_8338,N_8147);
xor U9978 (N_9978,N_8168,N_8505);
nand U9979 (N_9979,N_8236,N_8596);
and U9980 (N_9980,N_8085,N_8555);
and U9981 (N_9981,N_8073,N_8576);
nor U9982 (N_9982,N_8907,N_8488);
xor U9983 (N_9983,N_8344,N_8058);
or U9984 (N_9984,N_8677,N_8178);
xnor U9985 (N_9985,N_8171,N_8465);
and U9986 (N_9986,N_8102,N_8529);
and U9987 (N_9987,N_8734,N_8950);
nand U9988 (N_9988,N_8169,N_8545);
nand U9989 (N_9989,N_8898,N_8018);
nor U9990 (N_9990,N_8053,N_8195);
and U9991 (N_9991,N_8235,N_8132);
and U9992 (N_9992,N_8094,N_8006);
nor U9993 (N_9993,N_8299,N_8814);
and U9994 (N_9994,N_8311,N_8161);
nand U9995 (N_9995,N_8387,N_8304);
nand U9996 (N_9996,N_8924,N_8730);
xor U9997 (N_9997,N_8509,N_8506);
and U9998 (N_9998,N_8578,N_8542);
nand U9999 (N_9999,N_8190,N_8581);
nand U10000 (N_10000,N_9186,N_9393);
or U10001 (N_10001,N_9665,N_9468);
and U10002 (N_10002,N_9419,N_9832);
or U10003 (N_10003,N_9926,N_9081);
xor U10004 (N_10004,N_9127,N_9739);
xor U10005 (N_10005,N_9734,N_9959);
or U10006 (N_10006,N_9196,N_9449);
xor U10007 (N_10007,N_9376,N_9292);
nand U10008 (N_10008,N_9314,N_9110);
and U10009 (N_10009,N_9350,N_9705);
and U10010 (N_10010,N_9256,N_9299);
and U10011 (N_10011,N_9581,N_9029);
nor U10012 (N_10012,N_9202,N_9509);
and U10013 (N_10013,N_9593,N_9652);
and U10014 (N_10014,N_9451,N_9444);
or U10015 (N_10015,N_9436,N_9975);
or U10016 (N_10016,N_9093,N_9637);
nand U10017 (N_10017,N_9058,N_9427);
or U10018 (N_10018,N_9609,N_9426);
or U10019 (N_10019,N_9464,N_9620);
nand U10020 (N_10020,N_9332,N_9895);
or U10021 (N_10021,N_9813,N_9987);
nand U10022 (N_10022,N_9657,N_9692);
nor U10023 (N_10023,N_9401,N_9709);
or U10024 (N_10024,N_9381,N_9302);
nand U10025 (N_10025,N_9452,N_9828);
xnor U10026 (N_10026,N_9375,N_9741);
or U10027 (N_10027,N_9659,N_9224);
nand U10028 (N_10028,N_9954,N_9598);
and U10029 (N_10029,N_9803,N_9364);
nand U10030 (N_10030,N_9486,N_9011);
and U10031 (N_10031,N_9320,N_9726);
nand U10032 (N_10032,N_9586,N_9841);
or U10033 (N_10033,N_9238,N_9974);
nand U10034 (N_10034,N_9520,N_9372);
nand U10035 (N_10035,N_9856,N_9365);
nand U10036 (N_10036,N_9465,N_9596);
nor U10037 (N_10037,N_9570,N_9024);
or U10038 (N_10038,N_9924,N_9909);
or U10039 (N_10039,N_9453,N_9119);
nand U10040 (N_10040,N_9074,N_9807);
and U10041 (N_10041,N_9958,N_9099);
nand U10042 (N_10042,N_9893,N_9335);
or U10043 (N_10043,N_9086,N_9795);
xnor U10044 (N_10044,N_9358,N_9274);
xor U10045 (N_10045,N_9404,N_9773);
and U10046 (N_10046,N_9138,N_9215);
or U10047 (N_10047,N_9928,N_9675);
nor U10048 (N_10048,N_9471,N_9680);
nor U10049 (N_10049,N_9346,N_9548);
nor U10050 (N_10050,N_9148,N_9681);
nand U10051 (N_10051,N_9085,N_9027);
nor U10052 (N_10052,N_9658,N_9176);
nor U10053 (N_10053,N_9245,N_9382);
and U10054 (N_10054,N_9206,N_9319);
and U10055 (N_10055,N_9949,N_9757);
or U10056 (N_10056,N_9446,N_9062);
nand U10057 (N_10057,N_9740,N_9566);
or U10058 (N_10058,N_9904,N_9748);
or U10059 (N_10059,N_9247,N_9802);
or U10060 (N_10060,N_9158,N_9778);
nor U10061 (N_10061,N_9535,N_9950);
or U10062 (N_10062,N_9666,N_9122);
nand U10063 (N_10063,N_9023,N_9971);
xor U10064 (N_10064,N_9736,N_9996);
and U10065 (N_10065,N_9738,N_9756);
nor U10066 (N_10066,N_9050,N_9435);
nor U10067 (N_10067,N_9445,N_9525);
and U10068 (N_10068,N_9687,N_9617);
nor U10069 (N_10069,N_9012,N_9569);
and U10070 (N_10070,N_9685,N_9183);
xnor U10071 (N_10071,N_9283,N_9897);
nor U10072 (N_10072,N_9155,N_9106);
nand U10073 (N_10073,N_9036,N_9549);
and U10074 (N_10074,N_9615,N_9216);
and U10075 (N_10075,N_9330,N_9338);
and U10076 (N_10076,N_9053,N_9785);
or U10077 (N_10077,N_9955,N_9174);
nand U10078 (N_10078,N_9817,N_9339);
nor U10079 (N_10079,N_9069,N_9266);
and U10080 (N_10080,N_9990,N_9994);
nor U10081 (N_10081,N_9398,N_9510);
and U10082 (N_10082,N_9920,N_9530);
or U10083 (N_10083,N_9575,N_9234);
nand U10084 (N_10084,N_9661,N_9422);
nand U10085 (N_10085,N_9275,N_9821);
xor U10086 (N_10086,N_9706,N_9745);
and U10087 (N_10087,N_9839,N_9639);
nand U10088 (N_10088,N_9041,N_9852);
nand U10089 (N_10089,N_9628,N_9386);
nor U10090 (N_10090,N_9348,N_9116);
nor U10091 (N_10091,N_9491,N_9260);
and U10092 (N_10092,N_9564,N_9582);
nor U10093 (N_10093,N_9316,N_9084);
nor U10094 (N_10094,N_9013,N_9560);
nand U10095 (N_10095,N_9290,N_9295);
and U10096 (N_10096,N_9945,N_9503);
or U10097 (N_10097,N_9363,N_9134);
xnor U10098 (N_10098,N_9887,N_9908);
and U10099 (N_10099,N_9577,N_9166);
and U10100 (N_10100,N_9618,N_9989);
nor U10101 (N_10101,N_9480,N_9825);
and U10102 (N_10102,N_9496,N_9699);
or U10103 (N_10103,N_9656,N_9132);
nand U10104 (N_10104,N_9875,N_9285);
nor U10105 (N_10105,N_9834,N_9860);
nand U10106 (N_10106,N_9703,N_9727);
or U10107 (N_10107,N_9653,N_9001);
or U10108 (N_10108,N_9812,N_9595);
nand U10109 (N_10109,N_9667,N_9884);
nor U10110 (N_10110,N_9109,N_9991);
nor U10111 (N_10111,N_9101,N_9447);
nor U10112 (N_10112,N_9967,N_9353);
nand U10113 (N_10113,N_9291,N_9562);
nand U10114 (N_10114,N_9787,N_9563);
or U10115 (N_10115,N_9087,N_9208);
xnor U10116 (N_10116,N_9755,N_9482);
nor U10117 (N_10117,N_9218,N_9052);
or U10118 (N_10118,N_9108,N_9157);
nor U10119 (N_10119,N_9823,N_9307);
nand U10120 (N_10120,N_9673,N_9677);
nor U10121 (N_10121,N_9272,N_9630);
nor U10122 (N_10122,N_9671,N_9540);
and U10123 (N_10123,N_9645,N_9125);
and U10124 (N_10124,N_9054,N_9523);
nand U10125 (N_10125,N_9670,N_9051);
xor U10126 (N_10126,N_9801,N_9017);
and U10127 (N_10127,N_9182,N_9409);
nor U10128 (N_10128,N_9941,N_9288);
nand U10129 (N_10129,N_9889,N_9842);
xnor U10130 (N_10130,N_9693,N_9818);
and U10131 (N_10131,N_9221,N_9475);
nor U10132 (N_10132,N_9059,N_9168);
or U10133 (N_10133,N_9229,N_9819);
and U10134 (N_10134,N_9254,N_9883);
or U10135 (N_10135,N_9980,N_9160);
or U10136 (N_10136,N_9995,N_9690);
and U10137 (N_10137,N_9175,N_9321);
xor U10138 (N_10138,N_9370,N_9402);
and U10139 (N_10139,N_9988,N_9809);
or U10140 (N_10140,N_9406,N_9642);
nor U10141 (N_10141,N_9118,N_9930);
or U10142 (N_10142,N_9746,N_9697);
nor U10143 (N_10143,N_9120,N_9131);
nand U10144 (N_10144,N_9629,N_9483);
xor U10145 (N_10145,N_9002,N_9973);
nor U10146 (N_10146,N_9499,N_9905);
nand U10147 (N_10147,N_9105,N_9205);
or U10148 (N_10148,N_9682,N_9911);
or U10149 (N_10149,N_9416,N_9289);
or U10150 (N_10150,N_9711,N_9635);
nand U10151 (N_10151,N_9064,N_9870);
nor U10152 (N_10152,N_9646,N_9421);
nand U10153 (N_10153,N_9760,N_9729);
nand U10154 (N_10154,N_9579,N_9783);
nand U10155 (N_10155,N_9651,N_9144);
or U10156 (N_10156,N_9458,N_9481);
nand U10157 (N_10157,N_9648,N_9150);
or U10158 (N_10158,N_9223,N_9898);
or U10159 (N_10159,N_9572,N_9679);
nand U10160 (N_10160,N_9797,N_9297);
and U10161 (N_10161,N_9810,N_9534);
nor U10162 (N_10162,N_9932,N_9301);
nand U10163 (N_10163,N_9322,N_9312);
or U10164 (N_10164,N_9325,N_9360);
nand U10165 (N_10165,N_9261,N_9149);
nor U10166 (N_10166,N_9268,N_9391);
and U10167 (N_10167,N_9390,N_9284);
or U10168 (N_10168,N_9318,N_9805);
and U10169 (N_10169,N_9907,N_9777);
xor U10170 (N_10170,N_9235,N_9696);
nor U10171 (N_10171,N_9559,N_9032);
nor U10172 (N_10172,N_9811,N_9347);
nand U10173 (N_10173,N_9923,N_9672);
or U10174 (N_10174,N_9603,N_9177);
or U10175 (N_10175,N_9478,N_9669);
or U10176 (N_10176,N_9878,N_9015);
nor U10177 (N_10177,N_9356,N_9063);
nand U10178 (N_10178,N_9145,N_9749);
nand U10179 (N_10179,N_9425,N_9497);
nand U10180 (N_10180,N_9820,N_9104);
nor U10181 (N_10181,N_9660,N_9913);
nand U10182 (N_10182,N_9487,N_9914);
nand U10183 (N_10183,N_9018,N_9713);
and U10184 (N_10184,N_9663,N_9143);
nor U10185 (N_10185,N_9972,N_9009);
nand U10186 (N_10186,N_9886,N_9798);
or U10187 (N_10187,N_9257,N_9744);
and U10188 (N_10188,N_9373,N_9583);
or U10189 (N_10189,N_9964,N_9770);
nor U10190 (N_10190,N_9936,N_9126);
or U10191 (N_10191,N_9624,N_9599);
nand U10192 (N_10192,N_9121,N_9374);
nand U10193 (N_10193,N_9858,N_9430);
nand U10194 (N_10194,N_9243,N_9394);
or U10195 (N_10195,N_9529,N_9007);
nor U10196 (N_10196,N_9742,N_9644);
or U10197 (N_10197,N_9846,N_9781);
xor U10198 (N_10198,N_9873,N_9837);
and U10199 (N_10199,N_9429,N_9668);
xnor U10200 (N_10200,N_9537,N_9517);
or U10201 (N_10201,N_9743,N_9005);
or U10202 (N_10202,N_9655,N_9249);
nor U10203 (N_10203,N_9606,N_9782);
and U10204 (N_10204,N_9197,N_9279);
nor U10205 (N_10205,N_9733,N_9953);
and U10206 (N_10206,N_9031,N_9040);
nand U10207 (N_10207,N_9198,N_9396);
and U10208 (N_10208,N_9894,N_9488);
nor U10209 (N_10209,N_9721,N_9367);
nand U10210 (N_10210,N_9042,N_9688);
and U10211 (N_10211,N_9490,N_9986);
xor U10212 (N_10212,N_9650,N_9047);
or U10213 (N_10213,N_9546,N_9210);
nor U10214 (N_10214,N_9890,N_9413);
nor U10215 (N_10215,N_9576,N_9207);
nand U10216 (N_10216,N_9255,N_9233);
and U10217 (N_10217,N_9754,N_9985);
and U10218 (N_10218,N_9361,N_9385);
or U10219 (N_10219,N_9849,N_9872);
and U10220 (N_10220,N_9112,N_9766);
nor U10221 (N_10221,N_9474,N_9647);
and U10222 (N_10222,N_9512,N_9800);
xor U10223 (N_10223,N_9379,N_9891);
nand U10224 (N_10224,N_9146,N_9351);
nand U10225 (N_10225,N_9035,N_9469);
nand U10226 (N_10226,N_9824,N_9225);
nand U10227 (N_10227,N_9558,N_9702);
and U10228 (N_10228,N_9951,N_9184);
xor U10229 (N_10229,N_9280,N_9431);
nor U10230 (N_10230,N_9850,N_9181);
or U10231 (N_10231,N_9264,N_9683);
or U10232 (N_10232,N_9078,N_9336);
nand U10233 (N_10233,N_9056,N_9942);
xor U10234 (N_10234,N_9979,N_9762);
or U10235 (N_10235,N_9489,N_9355);
nand U10236 (N_10236,N_9626,N_9792);
or U10237 (N_10237,N_9129,N_9484);
or U10238 (N_10238,N_9424,N_9287);
nor U10239 (N_10239,N_9567,N_9293);
nand U10240 (N_10240,N_9442,N_9730);
nor U10241 (N_10241,N_9270,N_9060);
and U10242 (N_10242,N_9165,N_9956);
or U10243 (N_10243,N_9432,N_9326);
nor U10244 (N_10244,N_9940,N_9133);
nand U10245 (N_10245,N_9113,N_9075);
or U10246 (N_10246,N_9173,N_9296);
or U10247 (N_10247,N_9830,N_9412);
and U10248 (N_10248,N_9585,N_9384);
nand U10249 (N_10249,N_9498,N_9328);
or U10250 (N_10250,N_9764,N_9269);
and U10251 (N_10251,N_9095,N_9551);
nor U10252 (N_10252,N_9259,N_9354);
nor U10253 (N_10253,N_9357,N_9854);
nand U10254 (N_10254,N_9128,N_9248);
and U10255 (N_10255,N_9506,N_9039);
nand U10256 (N_10256,N_9840,N_9044);
nand U10257 (N_10257,N_9935,N_9731);
or U10258 (N_10258,N_9403,N_9934);
xor U10259 (N_10259,N_9966,N_9494);
nand U10260 (N_10260,N_9055,N_9674);
and U10261 (N_10261,N_9737,N_9070);
and U10262 (N_10262,N_9508,N_9473);
nor U10263 (N_10263,N_9010,N_9578);
nand U10264 (N_10264,N_9392,N_9377);
or U10265 (N_10265,N_9789,N_9467);
or U10266 (N_10266,N_9072,N_9507);
nor U10267 (N_10267,N_9045,N_9371);
or U10268 (N_10268,N_9545,N_9278);
or U10269 (N_10269,N_9418,N_9957);
nand U10270 (N_10270,N_9978,N_9536);
or U10271 (N_10271,N_9169,N_9750);
or U10272 (N_10272,N_9796,N_9759);
nand U10273 (N_10273,N_9747,N_9306);
nor U10274 (N_10274,N_9107,N_9619);
nand U10275 (N_10275,N_9008,N_9389);
nor U10276 (N_10276,N_9794,N_9833);
nand U10277 (N_10277,N_9231,N_9485);
or U10278 (N_10278,N_9822,N_9241);
nand U10279 (N_10279,N_9201,N_9772);
and U10280 (N_10280,N_9541,N_9139);
and U10281 (N_10281,N_9879,N_9092);
or U10282 (N_10282,N_9410,N_9862);
or U10283 (N_10283,N_9542,N_9098);
nor U10284 (N_10284,N_9843,N_9701);
nand U10285 (N_10285,N_9788,N_9547);
nand U10286 (N_10286,N_9686,N_9882);
or U10287 (N_10287,N_9917,N_9610);
nor U10288 (N_10288,N_9969,N_9874);
and U10289 (N_10289,N_9641,N_9901);
and U10290 (N_10290,N_9511,N_9030);
or U10291 (N_10291,N_9947,N_9455);
and U10292 (N_10292,N_9405,N_9970);
nand U10293 (N_10293,N_9147,N_9019);
or U10294 (N_10294,N_9597,N_9526);
nand U10295 (N_10295,N_9689,N_9034);
nor U10296 (N_10296,N_9992,N_9694);
nand U10297 (N_10297,N_9171,N_9433);
or U10298 (N_10298,N_9865,N_9876);
and U10299 (N_10299,N_9561,N_9152);
nor U10300 (N_10300,N_9538,N_9938);
nand U10301 (N_10301,N_9505,N_9999);
nor U10302 (N_10302,N_9790,N_9303);
or U10303 (N_10303,N_9340,N_9472);
and U10304 (N_10304,N_9162,N_9925);
and U10305 (N_10305,N_9501,N_9252);
nor U10306 (N_10306,N_9869,N_9910);
nor U10307 (N_10307,N_9179,N_9466);
nand U10308 (N_10308,N_9998,N_9775);
nor U10309 (N_10309,N_9151,N_9903);
or U10310 (N_10310,N_9720,N_9804);
or U10311 (N_10311,N_9604,N_9723);
and U10312 (N_10312,N_9057,N_9004);
and U10313 (N_10313,N_9698,N_9808);
nor U10314 (N_10314,N_9033,N_9944);
nor U10315 (N_10315,N_9153,N_9344);
or U10316 (N_10316,N_9187,N_9571);
nor U10317 (N_10317,N_9912,N_9902);
and U10318 (N_10318,N_9929,N_9415);
and U10319 (N_10319,N_9997,N_9049);
or U10320 (N_10320,N_9724,N_9477);
nand U10321 (N_10321,N_9317,N_9163);
or U10322 (N_10322,N_9456,N_9533);
nand U10323 (N_10323,N_9281,N_9515);
and U10324 (N_10324,N_9199,N_9067);
nor U10325 (N_10325,N_9844,N_9799);
nor U10326 (N_10326,N_9352,N_9459);
nand U10327 (N_10327,N_9282,N_9123);
nand U10328 (N_10328,N_9826,N_9142);
nand U10329 (N_10329,N_9211,N_9388);
and U10330 (N_10330,N_9786,N_9554);
or U10331 (N_10331,N_9963,N_9079);
or U10332 (N_10332,N_9073,N_9791);
nor U10333 (N_10333,N_9141,N_9753);
nor U10334 (N_10334,N_9094,N_9000);
or U10335 (N_10335,N_9359,N_9632);
nor U10336 (N_10336,N_9984,N_9190);
nor U10337 (N_10337,N_9440,N_9065);
nor U10338 (N_10338,N_9622,N_9922);
xnor U10339 (N_10339,N_9025,N_9500);
nor U10340 (N_10340,N_9020,N_9276);
and U10341 (N_10341,N_9779,N_9423);
and U10342 (N_10342,N_9140,N_9568);
xnor U10343 (N_10343,N_9717,N_9514);
nand U10344 (N_10344,N_9977,N_9961);
nor U10345 (N_10345,N_9111,N_9634);
or U10346 (N_10346,N_9752,N_9532);
and U10347 (N_10347,N_9845,N_9960);
nor U10348 (N_10348,N_9704,N_9308);
nand U10349 (N_10349,N_9919,N_9868);
xor U10350 (N_10350,N_9605,N_9495);
nor U10351 (N_10351,N_9838,N_9294);
nand U10352 (N_10352,N_9556,N_9851);
or U10353 (N_10353,N_9937,N_9470);
nor U10354 (N_10354,N_9083,N_9776);
and U10355 (N_10355,N_9993,N_9881);
and U10356 (N_10356,N_9918,N_9200);
xor U10357 (N_10357,N_9968,N_9209);
or U10358 (N_10358,N_9513,N_9071);
nor U10359 (N_10359,N_9885,N_9311);
and U10360 (N_10360,N_9366,N_9780);
and U10361 (N_10361,N_9521,N_9691);
nand U10362 (N_10362,N_9708,N_9414);
nor U10363 (N_10363,N_9531,N_9304);
and U10364 (N_10364,N_9028,N_9082);
or U10365 (N_10365,N_9476,N_9089);
or U10366 (N_10366,N_9298,N_9965);
or U10367 (N_10367,N_9806,N_9100);
xor U10368 (N_10368,N_9277,N_9172);
and U10369 (N_10369,N_9715,N_9387);
nand U10370 (N_10370,N_9649,N_9204);
or U10371 (N_10371,N_9203,N_9719);
or U10372 (N_10372,N_9115,N_9921);
or U10373 (N_10373,N_9528,N_9156);
or U10374 (N_10374,N_9076,N_9349);
nor U10375 (N_10375,N_9616,N_9716);
or U10376 (N_10376,N_9263,N_9627);
or U10377 (N_10377,N_9608,N_9237);
xnor U10378 (N_10378,N_9952,N_9006);
nor U10379 (N_10379,N_9369,N_9022);
nor U10380 (N_10380,N_9601,N_9591);
nand U10381 (N_10381,N_9976,N_9417);
and U10382 (N_10382,N_9315,N_9625);
or U10383 (N_10383,N_9867,N_9983);
or U10384 (N_10384,N_9038,N_9220);
nand U10385 (N_10385,N_9592,N_9342);
nand U10386 (N_10386,N_9130,N_9195);
nand U10387 (N_10387,N_9946,N_9899);
and U10388 (N_10388,N_9916,N_9258);
nor U10389 (N_10389,N_9552,N_9262);
nor U10390 (N_10390,N_9021,N_9539);
or U10391 (N_10391,N_9827,N_9219);
nand U10392 (N_10392,N_9573,N_9265);
nand U10393 (N_10393,N_9518,N_9253);
nand U10394 (N_10394,N_9271,N_9584);
xnor U10395 (N_10395,N_9273,N_9300);
xnor U10396 (N_10396,N_9829,N_9454);
nand U10397 (N_10397,N_9324,N_9343);
nor U10398 (N_10398,N_9714,N_9154);
or U10399 (N_10399,N_9565,N_9927);
nand U10400 (N_10400,N_9502,N_9161);
or U10401 (N_10401,N_9103,N_9493);
xnor U10402 (N_10402,N_9728,N_9438);
and U10403 (N_10403,N_9814,N_9333);
and U10404 (N_10404,N_9088,N_9981);
nand U10405 (N_10405,N_9185,N_9188);
nor U10406 (N_10406,N_9222,N_9461);
and U10407 (N_10407,N_9240,N_9864);
nor U10408 (N_10408,N_9191,N_9479);
and U10409 (N_10409,N_9189,N_9068);
nor U10410 (N_10410,N_9544,N_9411);
xor U10411 (N_10411,N_9136,N_9815);
and U10412 (N_10412,N_9962,N_9077);
nand U10413 (N_10413,N_9710,N_9250);
nand U10414 (N_10414,N_9114,N_9439);
nor U10415 (N_10415,N_9091,N_9492);
and U10416 (N_10416,N_9448,N_9016);
or U10417 (N_10417,N_9117,N_9242);
xnor U10418 (N_10418,N_9246,N_9137);
or U10419 (N_10419,N_9066,N_9732);
nand U10420 (N_10420,N_9310,N_9574);
or U10421 (N_10421,N_9758,N_9135);
nand U10422 (N_10422,N_9640,N_9607);
nand U10423 (N_10423,N_9323,N_9654);
or U10424 (N_10424,N_9003,N_9880);
and U10425 (N_10425,N_9124,N_9861);
nor U10426 (N_10426,N_9167,N_9866);
or U10427 (N_10427,N_9313,N_9621);
and U10428 (N_10428,N_9192,N_9228);
nand U10429 (N_10429,N_9847,N_9048);
nor U10430 (N_10430,N_9345,N_9676);
nor U10431 (N_10431,N_9631,N_9037);
nor U10432 (N_10432,N_9588,N_9768);
nand U10433 (N_10433,N_9587,N_9580);
and U10434 (N_10434,N_9329,N_9848);
or U10435 (N_10435,N_9636,N_9457);
nand U10436 (N_10436,N_9305,N_9722);
nand U10437 (N_10437,N_9589,N_9437);
nor U10438 (N_10438,N_9543,N_9217);
nand U10439 (N_10439,N_9982,N_9769);
xnor U10440 (N_10440,N_9831,N_9193);
nand U10441 (N_10441,N_9550,N_9892);
nor U10442 (N_10442,N_9853,N_9286);
nor U10443 (N_10443,N_9395,N_9164);
or U10444 (N_10444,N_9232,N_9463);
or U10445 (N_10445,N_9227,N_9614);
and U10446 (N_10446,N_9043,N_9662);
nor U10447 (N_10447,N_9516,N_9718);
and U10448 (N_10448,N_9519,N_9871);
or U10449 (N_10449,N_9612,N_9767);
and U10450 (N_10450,N_9180,N_9524);
nor U10451 (N_10451,N_9080,N_9341);
or U10452 (N_10452,N_9751,N_9600);
and U10453 (N_10453,N_9836,N_9400);
nor U10454 (N_10454,N_9443,N_9420);
nor U10455 (N_10455,N_9707,N_9097);
or U10456 (N_10456,N_9362,N_9900);
nand U10457 (N_10457,N_9327,N_9337);
nor U10458 (N_10458,N_9915,N_9061);
and U10459 (N_10459,N_9236,N_9765);
or U10460 (N_10460,N_9026,N_9784);
nand U10461 (N_10461,N_9735,N_9933);
xor U10462 (N_10462,N_9613,N_9712);
or U10463 (N_10463,N_9793,N_9906);
or U10464 (N_10464,N_9943,N_9212);
nand U10465 (N_10465,N_9504,N_9014);
xnor U10466 (N_10466,N_9331,N_9590);
and U10467 (N_10467,N_9368,N_9434);
and U10468 (N_10468,N_9888,N_9214);
nor U10469 (N_10469,N_9527,N_9159);
xor U10470 (N_10470,N_9602,N_9380);
nand U10471 (N_10471,N_9623,N_9460);
nor U10472 (N_10472,N_9877,N_9557);
and U10473 (N_10473,N_9383,N_9643);
nand U10474 (N_10474,N_9678,N_9664);
or U10475 (N_10475,N_9230,N_9896);
and U10476 (N_10476,N_9102,N_9553);
and U10477 (N_10477,N_9857,N_9695);
nor U10478 (N_10478,N_9684,N_9939);
and U10479 (N_10479,N_9725,N_9816);
nand U10480 (N_10480,N_9441,N_9863);
and U10481 (N_10481,N_9178,N_9397);
nor U10482 (N_10482,N_9244,N_9251);
nand U10483 (N_10483,N_9334,N_9633);
or U10484 (N_10484,N_9450,N_9428);
and U10485 (N_10485,N_9763,N_9859);
nor U10486 (N_10486,N_9771,N_9555);
or U10487 (N_10487,N_9267,N_9408);
or U10488 (N_10488,N_9213,N_9700);
or U10489 (N_10489,N_9611,N_9638);
nor U10490 (N_10490,N_9835,N_9239);
xor U10491 (N_10491,N_9378,N_9948);
or U10492 (N_10492,N_9046,N_9761);
nor U10493 (N_10493,N_9309,N_9399);
or U10494 (N_10494,N_9522,N_9407);
nor U10495 (N_10495,N_9855,N_9194);
and U10496 (N_10496,N_9594,N_9170);
nand U10497 (N_10497,N_9096,N_9931);
xor U10498 (N_10498,N_9226,N_9090);
xnor U10499 (N_10499,N_9462,N_9774);
or U10500 (N_10500,N_9337,N_9338);
and U10501 (N_10501,N_9917,N_9095);
or U10502 (N_10502,N_9416,N_9777);
and U10503 (N_10503,N_9115,N_9983);
or U10504 (N_10504,N_9747,N_9812);
or U10505 (N_10505,N_9120,N_9213);
or U10506 (N_10506,N_9894,N_9800);
or U10507 (N_10507,N_9549,N_9291);
nand U10508 (N_10508,N_9745,N_9273);
nand U10509 (N_10509,N_9453,N_9089);
nor U10510 (N_10510,N_9158,N_9427);
xnor U10511 (N_10511,N_9450,N_9210);
and U10512 (N_10512,N_9040,N_9774);
or U10513 (N_10513,N_9332,N_9419);
nand U10514 (N_10514,N_9421,N_9319);
xor U10515 (N_10515,N_9454,N_9879);
and U10516 (N_10516,N_9916,N_9613);
or U10517 (N_10517,N_9326,N_9307);
and U10518 (N_10518,N_9467,N_9169);
nor U10519 (N_10519,N_9335,N_9003);
or U10520 (N_10520,N_9689,N_9952);
xnor U10521 (N_10521,N_9768,N_9665);
and U10522 (N_10522,N_9497,N_9736);
nor U10523 (N_10523,N_9596,N_9436);
nand U10524 (N_10524,N_9834,N_9240);
nor U10525 (N_10525,N_9335,N_9282);
or U10526 (N_10526,N_9794,N_9554);
nand U10527 (N_10527,N_9346,N_9551);
nand U10528 (N_10528,N_9644,N_9367);
and U10529 (N_10529,N_9850,N_9955);
or U10530 (N_10530,N_9330,N_9161);
or U10531 (N_10531,N_9585,N_9575);
nand U10532 (N_10532,N_9854,N_9921);
and U10533 (N_10533,N_9460,N_9749);
nand U10534 (N_10534,N_9198,N_9230);
and U10535 (N_10535,N_9912,N_9736);
or U10536 (N_10536,N_9990,N_9828);
nand U10537 (N_10537,N_9584,N_9576);
xor U10538 (N_10538,N_9432,N_9069);
or U10539 (N_10539,N_9490,N_9530);
nand U10540 (N_10540,N_9131,N_9716);
nand U10541 (N_10541,N_9638,N_9069);
and U10542 (N_10542,N_9319,N_9825);
nand U10543 (N_10543,N_9675,N_9373);
or U10544 (N_10544,N_9478,N_9747);
or U10545 (N_10545,N_9573,N_9223);
nand U10546 (N_10546,N_9999,N_9078);
or U10547 (N_10547,N_9169,N_9571);
nor U10548 (N_10548,N_9275,N_9103);
or U10549 (N_10549,N_9528,N_9728);
nand U10550 (N_10550,N_9576,N_9909);
and U10551 (N_10551,N_9234,N_9723);
nand U10552 (N_10552,N_9777,N_9929);
nor U10553 (N_10553,N_9827,N_9872);
nand U10554 (N_10554,N_9458,N_9631);
and U10555 (N_10555,N_9714,N_9806);
and U10556 (N_10556,N_9126,N_9633);
nand U10557 (N_10557,N_9025,N_9986);
nand U10558 (N_10558,N_9307,N_9111);
or U10559 (N_10559,N_9956,N_9402);
or U10560 (N_10560,N_9224,N_9909);
xor U10561 (N_10561,N_9059,N_9343);
nor U10562 (N_10562,N_9878,N_9040);
and U10563 (N_10563,N_9813,N_9023);
nor U10564 (N_10564,N_9624,N_9950);
or U10565 (N_10565,N_9255,N_9569);
nor U10566 (N_10566,N_9150,N_9975);
nand U10567 (N_10567,N_9353,N_9876);
nand U10568 (N_10568,N_9877,N_9242);
and U10569 (N_10569,N_9727,N_9534);
or U10570 (N_10570,N_9692,N_9367);
nand U10571 (N_10571,N_9829,N_9430);
xor U10572 (N_10572,N_9357,N_9117);
nor U10573 (N_10573,N_9004,N_9928);
nor U10574 (N_10574,N_9164,N_9463);
nand U10575 (N_10575,N_9801,N_9591);
nand U10576 (N_10576,N_9594,N_9390);
nor U10577 (N_10577,N_9773,N_9473);
nor U10578 (N_10578,N_9502,N_9348);
xor U10579 (N_10579,N_9995,N_9018);
and U10580 (N_10580,N_9448,N_9864);
or U10581 (N_10581,N_9710,N_9459);
or U10582 (N_10582,N_9207,N_9536);
xor U10583 (N_10583,N_9047,N_9752);
nand U10584 (N_10584,N_9861,N_9975);
and U10585 (N_10585,N_9168,N_9740);
nand U10586 (N_10586,N_9572,N_9849);
nor U10587 (N_10587,N_9983,N_9970);
xnor U10588 (N_10588,N_9418,N_9598);
and U10589 (N_10589,N_9409,N_9194);
and U10590 (N_10590,N_9572,N_9635);
or U10591 (N_10591,N_9400,N_9611);
nor U10592 (N_10592,N_9732,N_9069);
or U10593 (N_10593,N_9366,N_9319);
or U10594 (N_10594,N_9004,N_9044);
nor U10595 (N_10595,N_9372,N_9561);
nand U10596 (N_10596,N_9483,N_9568);
and U10597 (N_10597,N_9575,N_9009);
nand U10598 (N_10598,N_9854,N_9110);
nor U10599 (N_10599,N_9782,N_9753);
or U10600 (N_10600,N_9154,N_9614);
and U10601 (N_10601,N_9525,N_9701);
or U10602 (N_10602,N_9175,N_9826);
nor U10603 (N_10603,N_9675,N_9414);
or U10604 (N_10604,N_9570,N_9955);
nand U10605 (N_10605,N_9930,N_9964);
xor U10606 (N_10606,N_9805,N_9609);
and U10607 (N_10607,N_9284,N_9425);
xor U10608 (N_10608,N_9346,N_9104);
and U10609 (N_10609,N_9482,N_9169);
nor U10610 (N_10610,N_9810,N_9877);
xor U10611 (N_10611,N_9973,N_9841);
or U10612 (N_10612,N_9759,N_9411);
nand U10613 (N_10613,N_9836,N_9558);
nand U10614 (N_10614,N_9771,N_9072);
nor U10615 (N_10615,N_9585,N_9854);
nand U10616 (N_10616,N_9631,N_9088);
nand U10617 (N_10617,N_9102,N_9851);
nand U10618 (N_10618,N_9755,N_9804);
or U10619 (N_10619,N_9741,N_9895);
nand U10620 (N_10620,N_9414,N_9324);
nand U10621 (N_10621,N_9280,N_9053);
or U10622 (N_10622,N_9087,N_9038);
or U10623 (N_10623,N_9900,N_9718);
or U10624 (N_10624,N_9478,N_9659);
nand U10625 (N_10625,N_9543,N_9233);
xor U10626 (N_10626,N_9201,N_9712);
xor U10627 (N_10627,N_9454,N_9095);
nand U10628 (N_10628,N_9292,N_9896);
and U10629 (N_10629,N_9480,N_9842);
nand U10630 (N_10630,N_9608,N_9099);
nand U10631 (N_10631,N_9059,N_9044);
and U10632 (N_10632,N_9319,N_9434);
xnor U10633 (N_10633,N_9315,N_9529);
or U10634 (N_10634,N_9059,N_9345);
xnor U10635 (N_10635,N_9167,N_9761);
and U10636 (N_10636,N_9845,N_9541);
nand U10637 (N_10637,N_9491,N_9193);
or U10638 (N_10638,N_9928,N_9213);
nand U10639 (N_10639,N_9164,N_9413);
nor U10640 (N_10640,N_9158,N_9580);
nor U10641 (N_10641,N_9137,N_9092);
or U10642 (N_10642,N_9047,N_9448);
and U10643 (N_10643,N_9583,N_9357);
or U10644 (N_10644,N_9856,N_9047);
or U10645 (N_10645,N_9773,N_9163);
nor U10646 (N_10646,N_9003,N_9971);
nor U10647 (N_10647,N_9479,N_9847);
and U10648 (N_10648,N_9142,N_9324);
xor U10649 (N_10649,N_9653,N_9783);
nand U10650 (N_10650,N_9530,N_9713);
and U10651 (N_10651,N_9370,N_9638);
and U10652 (N_10652,N_9000,N_9020);
nand U10653 (N_10653,N_9438,N_9259);
nand U10654 (N_10654,N_9886,N_9551);
nor U10655 (N_10655,N_9930,N_9622);
nand U10656 (N_10656,N_9128,N_9841);
nor U10657 (N_10657,N_9948,N_9786);
xnor U10658 (N_10658,N_9436,N_9081);
nor U10659 (N_10659,N_9104,N_9239);
or U10660 (N_10660,N_9919,N_9160);
nor U10661 (N_10661,N_9611,N_9493);
nand U10662 (N_10662,N_9672,N_9586);
nor U10663 (N_10663,N_9106,N_9712);
xnor U10664 (N_10664,N_9863,N_9903);
or U10665 (N_10665,N_9736,N_9001);
and U10666 (N_10666,N_9884,N_9186);
and U10667 (N_10667,N_9585,N_9303);
nand U10668 (N_10668,N_9929,N_9967);
xnor U10669 (N_10669,N_9588,N_9677);
and U10670 (N_10670,N_9025,N_9085);
or U10671 (N_10671,N_9281,N_9065);
and U10672 (N_10672,N_9633,N_9921);
or U10673 (N_10673,N_9690,N_9640);
nor U10674 (N_10674,N_9170,N_9267);
xnor U10675 (N_10675,N_9407,N_9787);
and U10676 (N_10676,N_9587,N_9537);
nor U10677 (N_10677,N_9062,N_9824);
nor U10678 (N_10678,N_9404,N_9871);
nand U10679 (N_10679,N_9935,N_9365);
nand U10680 (N_10680,N_9294,N_9226);
nand U10681 (N_10681,N_9857,N_9448);
or U10682 (N_10682,N_9195,N_9750);
xor U10683 (N_10683,N_9940,N_9346);
nand U10684 (N_10684,N_9034,N_9171);
nor U10685 (N_10685,N_9710,N_9900);
nand U10686 (N_10686,N_9287,N_9109);
nor U10687 (N_10687,N_9674,N_9631);
or U10688 (N_10688,N_9551,N_9072);
nand U10689 (N_10689,N_9199,N_9170);
nor U10690 (N_10690,N_9488,N_9387);
xnor U10691 (N_10691,N_9302,N_9798);
nand U10692 (N_10692,N_9059,N_9692);
and U10693 (N_10693,N_9398,N_9946);
xor U10694 (N_10694,N_9588,N_9761);
nand U10695 (N_10695,N_9416,N_9908);
or U10696 (N_10696,N_9902,N_9195);
nor U10697 (N_10697,N_9129,N_9953);
or U10698 (N_10698,N_9406,N_9635);
nand U10699 (N_10699,N_9617,N_9864);
or U10700 (N_10700,N_9262,N_9159);
nor U10701 (N_10701,N_9976,N_9972);
or U10702 (N_10702,N_9065,N_9081);
xnor U10703 (N_10703,N_9453,N_9557);
xnor U10704 (N_10704,N_9313,N_9452);
nor U10705 (N_10705,N_9662,N_9289);
xor U10706 (N_10706,N_9246,N_9807);
and U10707 (N_10707,N_9328,N_9351);
nand U10708 (N_10708,N_9546,N_9306);
nand U10709 (N_10709,N_9085,N_9697);
nor U10710 (N_10710,N_9229,N_9172);
nor U10711 (N_10711,N_9444,N_9973);
xor U10712 (N_10712,N_9780,N_9461);
and U10713 (N_10713,N_9416,N_9015);
or U10714 (N_10714,N_9602,N_9240);
xor U10715 (N_10715,N_9715,N_9329);
nor U10716 (N_10716,N_9362,N_9347);
or U10717 (N_10717,N_9822,N_9315);
and U10718 (N_10718,N_9939,N_9409);
nand U10719 (N_10719,N_9693,N_9252);
or U10720 (N_10720,N_9674,N_9062);
or U10721 (N_10721,N_9283,N_9990);
xnor U10722 (N_10722,N_9956,N_9679);
and U10723 (N_10723,N_9026,N_9718);
and U10724 (N_10724,N_9435,N_9915);
or U10725 (N_10725,N_9242,N_9815);
or U10726 (N_10726,N_9687,N_9973);
nor U10727 (N_10727,N_9423,N_9023);
nor U10728 (N_10728,N_9598,N_9157);
xnor U10729 (N_10729,N_9903,N_9673);
xor U10730 (N_10730,N_9396,N_9158);
or U10731 (N_10731,N_9333,N_9063);
and U10732 (N_10732,N_9813,N_9384);
or U10733 (N_10733,N_9911,N_9890);
and U10734 (N_10734,N_9579,N_9033);
nor U10735 (N_10735,N_9469,N_9316);
nand U10736 (N_10736,N_9576,N_9647);
or U10737 (N_10737,N_9064,N_9511);
or U10738 (N_10738,N_9240,N_9700);
nand U10739 (N_10739,N_9057,N_9372);
or U10740 (N_10740,N_9454,N_9223);
nor U10741 (N_10741,N_9302,N_9309);
and U10742 (N_10742,N_9436,N_9940);
and U10743 (N_10743,N_9588,N_9068);
xor U10744 (N_10744,N_9259,N_9323);
nor U10745 (N_10745,N_9953,N_9646);
and U10746 (N_10746,N_9363,N_9894);
or U10747 (N_10747,N_9710,N_9375);
or U10748 (N_10748,N_9727,N_9519);
nand U10749 (N_10749,N_9835,N_9806);
xor U10750 (N_10750,N_9231,N_9063);
or U10751 (N_10751,N_9960,N_9260);
and U10752 (N_10752,N_9843,N_9160);
nor U10753 (N_10753,N_9817,N_9893);
nor U10754 (N_10754,N_9825,N_9698);
nand U10755 (N_10755,N_9414,N_9809);
and U10756 (N_10756,N_9078,N_9459);
nor U10757 (N_10757,N_9614,N_9312);
or U10758 (N_10758,N_9508,N_9877);
and U10759 (N_10759,N_9725,N_9706);
nand U10760 (N_10760,N_9919,N_9479);
and U10761 (N_10761,N_9366,N_9291);
or U10762 (N_10762,N_9773,N_9442);
nor U10763 (N_10763,N_9194,N_9349);
or U10764 (N_10764,N_9217,N_9101);
and U10765 (N_10765,N_9700,N_9451);
and U10766 (N_10766,N_9756,N_9308);
and U10767 (N_10767,N_9124,N_9654);
and U10768 (N_10768,N_9309,N_9961);
nand U10769 (N_10769,N_9873,N_9633);
or U10770 (N_10770,N_9484,N_9272);
nand U10771 (N_10771,N_9550,N_9437);
nand U10772 (N_10772,N_9963,N_9264);
nor U10773 (N_10773,N_9482,N_9663);
or U10774 (N_10774,N_9538,N_9964);
or U10775 (N_10775,N_9695,N_9743);
xnor U10776 (N_10776,N_9332,N_9658);
xor U10777 (N_10777,N_9588,N_9908);
or U10778 (N_10778,N_9270,N_9184);
or U10779 (N_10779,N_9574,N_9022);
nand U10780 (N_10780,N_9717,N_9954);
and U10781 (N_10781,N_9290,N_9104);
nand U10782 (N_10782,N_9478,N_9431);
nor U10783 (N_10783,N_9264,N_9953);
nand U10784 (N_10784,N_9082,N_9757);
nand U10785 (N_10785,N_9579,N_9163);
and U10786 (N_10786,N_9153,N_9880);
and U10787 (N_10787,N_9804,N_9190);
xnor U10788 (N_10788,N_9846,N_9955);
nand U10789 (N_10789,N_9362,N_9554);
and U10790 (N_10790,N_9994,N_9751);
nand U10791 (N_10791,N_9308,N_9171);
and U10792 (N_10792,N_9537,N_9442);
and U10793 (N_10793,N_9347,N_9380);
or U10794 (N_10794,N_9937,N_9085);
nand U10795 (N_10795,N_9889,N_9628);
nor U10796 (N_10796,N_9547,N_9880);
nand U10797 (N_10797,N_9161,N_9100);
and U10798 (N_10798,N_9922,N_9405);
and U10799 (N_10799,N_9123,N_9419);
nor U10800 (N_10800,N_9623,N_9796);
or U10801 (N_10801,N_9900,N_9242);
nand U10802 (N_10802,N_9794,N_9281);
or U10803 (N_10803,N_9839,N_9277);
or U10804 (N_10804,N_9358,N_9351);
or U10805 (N_10805,N_9013,N_9812);
or U10806 (N_10806,N_9202,N_9112);
xor U10807 (N_10807,N_9545,N_9328);
or U10808 (N_10808,N_9387,N_9864);
or U10809 (N_10809,N_9682,N_9948);
nor U10810 (N_10810,N_9601,N_9496);
nor U10811 (N_10811,N_9308,N_9520);
or U10812 (N_10812,N_9042,N_9088);
nand U10813 (N_10813,N_9626,N_9574);
and U10814 (N_10814,N_9788,N_9346);
or U10815 (N_10815,N_9245,N_9749);
or U10816 (N_10816,N_9600,N_9906);
and U10817 (N_10817,N_9798,N_9646);
nor U10818 (N_10818,N_9036,N_9847);
and U10819 (N_10819,N_9324,N_9073);
or U10820 (N_10820,N_9218,N_9981);
nor U10821 (N_10821,N_9896,N_9510);
or U10822 (N_10822,N_9842,N_9832);
and U10823 (N_10823,N_9810,N_9454);
xor U10824 (N_10824,N_9707,N_9408);
or U10825 (N_10825,N_9135,N_9010);
and U10826 (N_10826,N_9360,N_9141);
nand U10827 (N_10827,N_9391,N_9051);
nor U10828 (N_10828,N_9995,N_9861);
nor U10829 (N_10829,N_9706,N_9473);
nand U10830 (N_10830,N_9421,N_9759);
and U10831 (N_10831,N_9303,N_9439);
nand U10832 (N_10832,N_9602,N_9587);
xor U10833 (N_10833,N_9275,N_9254);
and U10834 (N_10834,N_9662,N_9178);
or U10835 (N_10835,N_9876,N_9846);
or U10836 (N_10836,N_9131,N_9286);
or U10837 (N_10837,N_9236,N_9368);
or U10838 (N_10838,N_9188,N_9502);
nor U10839 (N_10839,N_9984,N_9484);
nor U10840 (N_10840,N_9137,N_9607);
nand U10841 (N_10841,N_9818,N_9045);
nor U10842 (N_10842,N_9573,N_9087);
nor U10843 (N_10843,N_9581,N_9147);
nand U10844 (N_10844,N_9482,N_9876);
nand U10845 (N_10845,N_9736,N_9519);
or U10846 (N_10846,N_9758,N_9561);
nand U10847 (N_10847,N_9873,N_9534);
and U10848 (N_10848,N_9059,N_9071);
and U10849 (N_10849,N_9794,N_9999);
and U10850 (N_10850,N_9401,N_9297);
nand U10851 (N_10851,N_9855,N_9955);
or U10852 (N_10852,N_9613,N_9179);
or U10853 (N_10853,N_9491,N_9068);
and U10854 (N_10854,N_9147,N_9817);
or U10855 (N_10855,N_9215,N_9548);
nand U10856 (N_10856,N_9556,N_9445);
or U10857 (N_10857,N_9770,N_9012);
and U10858 (N_10858,N_9249,N_9625);
or U10859 (N_10859,N_9520,N_9234);
nor U10860 (N_10860,N_9298,N_9271);
and U10861 (N_10861,N_9829,N_9979);
and U10862 (N_10862,N_9077,N_9220);
and U10863 (N_10863,N_9331,N_9485);
and U10864 (N_10864,N_9800,N_9604);
and U10865 (N_10865,N_9468,N_9844);
nand U10866 (N_10866,N_9487,N_9962);
or U10867 (N_10867,N_9284,N_9179);
xor U10868 (N_10868,N_9624,N_9014);
nand U10869 (N_10869,N_9335,N_9810);
nand U10870 (N_10870,N_9654,N_9332);
and U10871 (N_10871,N_9409,N_9899);
and U10872 (N_10872,N_9436,N_9591);
and U10873 (N_10873,N_9478,N_9721);
and U10874 (N_10874,N_9341,N_9664);
or U10875 (N_10875,N_9117,N_9302);
and U10876 (N_10876,N_9981,N_9222);
nand U10877 (N_10877,N_9528,N_9890);
or U10878 (N_10878,N_9660,N_9741);
nand U10879 (N_10879,N_9739,N_9446);
xnor U10880 (N_10880,N_9929,N_9403);
and U10881 (N_10881,N_9493,N_9988);
or U10882 (N_10882,N_9310,N_9904);
and U10883 (N_10883,N_9679,N_9427);
or U10884 (N_10884,N_9728,N_9576);
nor U10885 (N_10885,N_9786,N_9117);
or U10886 (N_10886,N_9973,N_9834);
and U10887 (N_10887,N_9427,N_9257);
xnor U10888 (N_10888,N_9110,N_9420);
nor U10889 (N_10889,N_9340,N_9805);
nor U10890 (N_10890,N_9445,N_9165);
nand U10891 (N_10891,N_9700,N_9612);
nand U10892 (N_10892,N_9221,N_9645);
xnor U10893 (N_10893,N_9245,N_9176);
xnor U10894 (N_10894,N_9666,N_9445);
and U10895 (N_10895,N_9369,N_9141);
and U10896 (N_10896,N_9383,N_9706);
and U10897 (N_10897,N_9160,N_9027);
nand U10898 (N_10898,N_9363,N_9223);
nor U10899 (N_10899,N_9017,N_9949);
nand U10900 (N_10900,N_9992,N_9119);
or U10901 (N_10901,N_9459,N_9660);
nor U10902 (N_10902,N_9087,N_9258);
or U10903 (N_10903,N_9574,N_9970);
nor U10904 (N_10904,N_9748,N_9176);
nor U10905 (N_10905,N_9343,N_9090);
nor U10906 (N_10906,N_9326,N_9706);
and U10907 (N_10907,N_9401,N_9951);
or U10908 (N_10908,N_9603,N_9837);
or U10909 (N_10909,N_9053,N_9317);
nand U10910 (N_10910,N_9522,N_9784);
and U10911 (N_10911,N_9042,N_9254);
or U10912 (N_10912,N_9498,N_9013);
nor U10913 (N_10913,N_9852,N_9542);
or U10914 (N_10914,N_9920,N_9371);
or U10915 (N_10915,N_9897,N_9483);
and U10916 (N_10916,N_9389,N_9138);
xor U10917 (N_10917,N_9113,N_9151);
or U10918 (N_10918,N_9904,N_9155);
nand U10919 (N_10919,N_9130,N_9626);
nand U10920 (N_10920,N_9239,N_9375);
or U10921 (N_10921,N_9578,N_9337);
nor U10922 (N_10922,N_9260,N_9891);
and U10923 (N_10923,N_9066,N_9929);
or U10924 (N_10924,N_9176,N_9968);
and U10925 (N_10925,N_9651,N_9293);
and U10926 (N_10926,N_9771,N_9338);
and U10927 (N_10927,N_9614,N_9836);
xnor U10928 (N_10928,N_9609,N_9033);
and U10929 (N_10929,N_9756,N_9753);
nand U10930 (N_10930,N_9423,N_9367);
and U10931 (N_10931,N_9435,N_9561);
nand U10932 (N_10932,N_9478,N_9170);
and U10933 (N_10933,N_9263,N_9196);
or U10934 (N_10934,N_9501,N_9601);
nand U10935 (N_10935,N_9924,N_9105);
and U10936 (N_10936,N_9034,N_9005);
nor U10937 (N_10937,N_9991,N_9687);
nand U10938 (N_10938,N_9712,N_9887);
or U10939 (N_10939,N_9225,N_9797);
and U10940 (N_10940,N_9043,N_9577);
or U10941 (N_10941,N_9760,N_9171);
xnor U10942 (N_10942,N_9581,N_9621);
nand U10943 (N_10943,N_9360,N_9842);
and U10944 (N_10944,N_9214,N_9364);
nor U10945 (N_10945,N_9808,N_9323);
nand U10946 (N_10946,N_9817,N_9804);
nand U10947 (N_10947,N_9262,N_9912);
nor U10948 (N_10948,N_9262,N_9453);
and U10949 (N_10949,N_9053,N_9494);
nor U10950 (N_10950,N_9615,N_9561);
or U10951 (N_10951,N_9424,N_9989);
or U10952 (N_10952,N_9477,N_9190);
nor U10953 (N_10953,N_9064,N_9470);
or U10954 (N_10954,N_9828,N_9594);
and U10955 (N_10955,N_9708,N_9261);
nor U10956 (N_10956,N_9769,N_9322);
nand U10957 (N_10957,N_9184,N_9638);
or U10958 (N_10958,N_9584,N_9846);
nor U10959 (N_10959,N_9328,N_9458);
or U10960 (N_10960,N_9618,N_9411);
nand U10961 (N_10961,N_9576,N_9531);
nand U10962 (N_10962,N_9493,N_9529);
and U10963 (N_10963,N_9182,N_9156);
or U10964 (N_10964,N_9275,N_9391);
or U10965 (N_10965,N_9137,N_9542);
nor U10966 (N_10966,N_9715,N_9714);
xor U10967 (N_10967,N_9903,N_9505);
xor U10968 (N_10968,N_9521,N_9466);
nor U10969 (N_10969,N_9065,N_9135);
nor U10970 (N_10970,N_9822,N_9398);
or U10971 (N_10971,N_9252,N_9995);
or U10972 (N_10972,N_9603,N_9962);
and U10973 (N_10973,N_9675,N_9861);
and U10974 (N_10974,N_9193,N_9771);
or U10975 (N_10975,N_9742,N_9286);
or U10976 (N_10976,N_9141,N_9819);
and U10977 (N_10977,N_9304,N_9196);
nor U10978 (N_10978,N_9542,N_9600);
and U10979 (N_10979,N_9834,N_9463);
xnor U10980 (N_10980,N_9914,N_9860);
and U10981 (N_10981,N_9094,N_9347);
or U10982 (N_10982,N_9060,N_9944);
nor U10983 (N_10983,N_9131,N_9478);
nor U10984 (N_10984,N_9305,N_9118);
and U10985 (N_10985,N_9940,N_9403);
nand U10986 (N_10986,N_9115,N_9534);
nor U10987 (N_10987,N_9382,N_9260);
or U10988 (N_10988,N_9184,N_9995);
nand U10989 (N_10989,N_9331,N_9255);
and U10990 (N_10990,N_9545,N_9601);
or U10991 (N_10991,N_9897,N_9358);
nor U10992 (N_10992,N_9808,N_9951);
or U10993 (N_10993,N_9565,N_9131);
xnor U10994 (N_10994,N_9473,N_9292);
nand U10995 (N_10995,N_9058,N_9856);
nand U10996 (N_10996,N_9197,N_9624);
nor U10997 (N_10997,N_9219,N_9740);
nor U10998 (N_10998,N_9375,N_9469);
nor U10999 (N_10999,N_9417,N_9020);
or U11000 (N_11000,N_10066,N_10765);
and U11001 (N_11001,N_10146,N_10950);
nor U11002 (N_11002,N_10505,N_10311);
nor U11003 (N_11003,N_10323,N_10745);
or U11004 (N_11004,N_10751,N_10973);
nor U11005 (N_11005,N_10432,N_10251);
nor U11006 (N_11006,N_10707,N_10279);
or U11007 (N_11007,N_10641,N_10747);
or U11008 (N_11008,N_10955,N_10150);
nand U11009 (N_11009,N_10832,N_10770);
nor U11010 (N_11010,N_10133,N_10103);
and U11011 (N_11011,N_10424,N_10224);
nand U11012 (N_11012,N_10781,N_10607);
nor U11013 (N_11013,N_10276,N_10377);
nand U11014 (N_11014,N_10847,N_10665);
nor U11015 (N_11015,N_10797,N_10867);
nor U11016 (N_11016,N_10392,N_10697);
or U11017 (N_11017,N_10637,N_10417);
or U11018 (N_11018,N_10004,N_10910);
nand U11019 (N_11019,N_10318,N_10236);
and U11020 (N_11020,N_10099,N_10698);
nor U11021 (N_11021,N_10828,N_10678);
xor U11022 (N_11022,N_10442,N_10443);
nand U11023 (N_11023,N_10151,N_10932);
or U11024 (N_11024,N_10605,N_10299);
and U11025 (N_11025,N_10568,N_10750);
or U11026 (N_11026,N_10541,N_10295);
or U11027 (N_11027,N_10499,N_10886);
nor U11028 (N_11028,N_10724,N_10209);
and U11029 (N_11029,N_10170,N_10595);
or U11030 (N_11030,N_10701,N_10575);
or U11031 (N_11031,N_10100,N_10971);
nor U11032 (N_11032,N_10135,N_10264);
nand U11033 (N_11033,N_10018,N_10769);
nor U11034 (N_11034,N_10438,N_10455);
xnor U11035 (N_11035,N_10997,N_10090);
or U11036 (N_11036,N_10598,N_10578);
or U11037 (N_11037,N_10487,N_10016);
and U11038 (N_11038,N_10091,N_10996);
or U11039 (N_11039,N_10001,N_10901);
nand U11040 (N_11040,N_10591,N_10364);
and U11041 (N_11041,N_10760,N_10310);
nand U11042 (N_11042,N_10109,N_10457);
xor U11043 (N_11043,N_10241,N_10243);
nand U11044 (N_11044,N_10611,N_10190);
nor U11045 (N_11045,N_10385,N_10929);
nand U11046 (N_11046,N_10835,N_10511);
nor U11047 (N_11047,N_10970,N_10218);
nor U11048 (N_11048,N_10551,N_10705);
nor U11049 (N_11049,N_10221,N_10708);
or U11050 (N_11050,N_10720,N_10566);
or U11051 (N_11051,N_10275,N_10362);
nor U11052 (N_11052,N_10830,N_10391);
xnor U11053 (N_11053,N_10069,N_10040);
or U11054 (N_11054,N_10853,N_10126);
and U11055 (N_11055,N_10723,N_10137);
and U11056 (N_11056,N_10005,N_10922);
nor U11057 (N_11057,N_10683,N_10301);
nor U11058 (N_11058,N_10784,N_10262);
or U11059 (N_11059,N_10968,N_10848);
nor U11060 (N_11060,N_10608,N_10493);
nand U11061 (N_11061,N_10398,N_10967);
xor U11062 (N_11062,N_10987,N_10246);
or U11063 (N_11063,N_10829,N_10325);
nor U11064 (N_11064,N_10521,N_10002);
nand U11065 (N_11065,N_10051,N_10673);
and U11066 (N_11066,N_10397,N_10703);
or U11067 (N_11067,N_10143,N_10702);
nand U11068 (N_11068,N_10721,N_10649);
and U11069 (N_11069,N_10658,N_10532);
nand U11070 (N_11070,N_10490,N_10237);
nor U11071 (N_11071,N_10643,N_10184);
nor U11072 (N_11072,N_10677,N_10865);
and U11073 (N_11073,N_10125,N_10336);
nand U11074 (N_11074,N_10523,N_10934);
or U11075 (N_11075,N_10817,N_10918);
or U11076 (N_11076,N_10020,N_10925);
and U11077 (N_11077,N_10909,N_10947);
or U11078 (N_11078,N_10902,N_10851);
and U11079 (N_11079,N_10270,N_10895);
nor U11080 (N_11080,N_10429,N_10335);
or U11081 (N_11081,N_10104,N_10719);
nand U11082 (N_11082,N_10669,N_10965);
nor U11083 (N_11083,N_10743,N_10861);
nand U11084 (N_11084,N_10193,N_10489);
or U11085 (N_11085,N_10891,N_10175);
nand U11086 (N_11086,N_10360,N_10113);
or U11087 (N_11087,N_10194,N_10067);
or U11088 (N_11088,N_10794,N_10282);
nor U11089 (N_11089,N_10339,N_10988);
and U11090 (N_11090,N_10024,N_10261);
nand U11091 (N_11091,N_10186,N_10075);
nand U11092 (N_11092,N_10453,N_10802);
and U11093 (N_11093,N_10022,N_10727);
and U11094 (N_11094,N_10268,N_10889);
xnor U11095 (N_11095,N_10957,N_10783);
nor U11096 (N_11096,N_10000,N_10614);
xnor U11097 (N_11097,N_10728,N_10142);
nor U11098 (N_11098,N_10631,N_10687);
and U11099 (N_11099,N_10786,N_10920);
or U11100 (N_11100,N_10796,N_10624);
or U11101 (N_11101,N_10199,N_10804);
nand U11102 (N_11102,N_10448,N_10176);
nor U11103 (N_11103,N_10841,N_10880);
nor U11104 (N_11104,N_10191,N_10156);
and U11105 (N_11105,N_10418,N_10354);
nand U11106 (N_11106,N_10811,N_10500);
and U11107 (N_11107,N_10842,N_10297);
and U11108 (N_11108,N_10390,N_10820);
nor U11109 (N_11109,N_10250,N_10296);
nor U11110 (N_11110,N_10917,N_10451);
or U11111 (N_11111,N_10373,N_10612);
or U11112 (N_11112,N_10414,N_10138);
or U11113 (N_11113,N_10187,N_10228);
or U11114 (N_11114,N_10936,N_10182);
or U11115 (N_11115,N_10063,N_10473);
nor U11116 (N_11116,N_10277,N_10471);
nand U11117 (N_11117,N_10388,N_10862);
or U11118 (N_11118,N_10434,N_10904);
xor U11119 (N_11119,N_10494,N_10872);
or U11120 (N_11120,N_10452,N_10078);
or U11121 (N_11121,N_10634,N_10793);
nand U11122 (N_11122,N_10680,N_10736);
and U11123 (N_11123,N_10742,N_10030);
or U11124 (N_11124,N_10106,N_10128);
or U11125 (N_11125,N_10481,N_10361);
or U11126 (N_11126,N_10419,N_10546);
and U11127 (N_11127,N_10337,N_10771);
nor U11128 (N_11128,N_10038,N_10426);
and U11129 (N_11129,N_10626,N_10039);
or U11130 (N_11130,N_10327,N_10960);
or U11131 (N_11131,N_10839,N_10466);
nor U11132 (N_11132,N_10463,N_10510);
and U11133 (N_11133,N_10587,N_10502);
and U11134 (N_11134,N_10685,N_10795);
and U11135 (N_11135,N_10244,N_10780);
or U11136 (N_11136,N_10699,N_10376);
and U11137 (N_11137,N_10083,N_10164);
nand U11138 (N_11138,N_10633,N_10172);
or U11139 (N_11139,N_10691,N_10982);
and U11140 (N_11140,N_10632,N_10107);
and U11141 (N_11141,N_10343,N_10613);
xnor U11142 (N_11142,N_10435,N_10718);
xor U11143 (N_11143,N_10212,N_10342);
and U11144 (N_11144,N_10507,N_10827);
or U11145 (N_11145,N_10514,N_10476);
xor U11146 (N_11146,N_10704,N_10756);
xor U11147 (N_11147,N_10367,N_10401);
nand U11148 (N_11148,N_10378,N_10974);
and U11149 (N_11149,N_10402,N_10892);
nand U11150 (N_11150,N_10064,N_10203);
or U11151 (N_11151,N_10431,N_10215);
or U11152 (N_11152,N_10406,N_10287);
or U11153 (N_11153,N_10334,N_10615);
xnor U11154 (N_11154,N_10921,N_10580);
nand U11155 (N_11155,N_10084,N_10216);
nor U11156 (N_11156,N_10217,N_10055);
nand U11157 (N_11157,N_10710,N_10522);
nor U11158 (N_11158,N_10893,N_10530);
or U11159 (N_11159,N_10089,N_10010);
or U11160 (N_11160,N_10951,N_10630);
or U11161 (N_11161,N_10449,N_10877);
nor U11162 (N_11162,N_10171,N_10681);
and U11163 (N_11163,N_10948,N_10748);
or U11164 (N_11164,N_10396,N_10349);
nor U11165 (N_11165,N_10025,N_10700);
and U11166 (N_11166,N_10809,N_10110);
nor U11167 (N_11167,N_10445,N_10653);
nand U11168 (N_11168,N_10386,N_10374);
or U11169 (N_11169,N_10547,N_10539);
or U11170 (N_11170,N_10328,N_10846);
nor U11171 (N_11171,N_10450,N_10118);
or U11172 (N_11172,N_10468,N_10239);
nor U11173 (N_11173,N_10864,N_10593);
nor U11174 (N_11174,N_10283,N_10144);
and U11175 (N_11175,N_10651,N_10717);
nor U11176 (N_11176,N_10352,N_10280);
or U11177 (N_11177,N_10584,N_10253);
or U11178 (N_11178,N_10357,N_10200);
nand U11179 (N_11179,N_10588,N_10753);
xnor U11180 (N_11180,N_10806,N_10271);
nor U11181 (N_11181,N_10696,N_10715);
nor U11182 (N_11182,N_10488,N_10528);
nand U11183 (N_11183,N_10496,N_10117);
and U11184 (N_11184,N_10625,N_10792);
or U11185 (N_11185,N_10101,N_10709);
and U11186 (N_11186,N_10870,N_10542);
and U11187 (N_11187,N_10787,N_10577);
or U11188 (N_11188,N_10824,N_10088);
or U11189 (N_11189,N_10459,N_10814);
and U11190 (N_11190,N_10223,N_10197);
or U11191 (N_11191,N_10914,N_10790);
or U11192 (N_11192,N_10731,N_10854);
nand U11193 (N_11193,N_10169,N_10694);
nor U11194 (N_11194,N_10706,N_10121);
nand U11195 (N_11195,N_10482,N_10884);
nor U11196 (N_11196,N_10778,N_10400);
or U11197 (N_11197,N_10458,N_10945);
or U11198 (N_11198,N_10013,N_10245);
nand U11199 (N_11199,N_10729,N_10267);
and U11200 (N_11200,N_10603,N_10671);
and U11201 (N_11201,N_10874,N_10585);
or U11202 (N_11202,N_10887,N_10382);
nand U11203 (N_11203,N_10056,N_10622);
or U11204 (N_11204,N_10561,N_10883);
nand U11205 (N_11205,N_10928,N_10387);
and U11206 (N_11206,N_10211,N_10368);
and U11207 (N_11207,N_10439,N_10008);
nor U11208 (N_11208,N_10474,N_10646);
xor U11209 (N_11209,N_10062,N_10610);
or U11210 (N_11210,N_10773,N_10559);
xnor U11211 (N_11211,N_10776,N_10141);
nor U11212 (N_11212,N_10119,N_10554);
nor U11213 (N_11213,N_10185,N_10423);
nor U11214 (N_11214,N_10105,N_10043);
nor U11215 (N_11215,N_10042,N_10356);
xnor U11216 (N_11216,N_10157,N_10695);
nand U11217 (N_11217,N_10550,N_10739);
xnor U11218 (N_11218,N_10120,N_10938);
or U11219 (N_11219,N_10816,N_10518);
and U11220 (N_11220,N_10755,N_10956);
and U11221 (N_11221,N_10491,N_10220);
and U11222 (N_11222,N_10659,N_10949);
nand U11223 (N_11223,N_10322,N_10531);
or U11224 (N_11224,N_10340,N_10111);
and U11225 (N_11225,N_10412,N_10962);
and U11226 (N_11226,N_10462,N_10574);
nand U11227 (N_11227,N_10077,N_10799);
and U11228 (N_11228,N_10616,N_10980);
nor U11229 (N_11229,N_10810,N_10095);
nand U11230 (N_11230,N_10140,N_10549);
nor U11231 (N_11231,N_10319,N_10272);
or U11232 (N_11232,N_10619,N_10158);
nor U11233 (N_11233,N_10281,N_10353);
nand U11234 (N_11234,N_10876,N_10300);
nand U11235 (N_11235,N_10399,N_10623);
nor U11236 (N_11236,N_10991,N_10512);
or U11237 (N_11237,N_10347,N_10366);
and U11238 (N_11238,N_10079,N_10684);
or U11239 (N_11239,N_10746,N_10636);
nor U11240 (N_11240,N_10969,N_10341);
nor U11241 (N_11241,N_10871,N_10249);
xor U11242 (N_11242,N_10690,N_10782);
and U11243 (N_11243,N_10907,N_10779);
nor U11244 (N_11244,N_10394,N_10456);
nand U11245 (N_11245,N_10682,N_10534);
xor U11246 (N_11246,N_10210,N_10898);
nor U11247 (N_11247,N_10330,N_10447);
or U11248 (N_11248,N_10427,N_10978);
and U11249 (N_11249,N_10933,N_10831);
and U11250 (N_11250,N_10308,N_10213);
xor U11251 (N_11251,N_10201,N_10940);
and U11252 (N_11252,N_10660,N_10007);
nor U11253 (N_11253,N_10127,N_10420);
nand U11254 (N_11254,N_10048,N_10766);
nand U11255 (N_11255,N_10284,N_10053);
or U11256 (N_11256,N_10037,N_10915);
or U11257 (N_11257,N_10526,N_10102);
and U11258 (N_11258,N_10302,N_10744);
or U11259 (N_11259,N_10233,N_10881);
nand U11260 (N_11260,N_10291,N_10761);
and U11261 (N_11261,N_10012,N_10358);
and U11262 (N_11262,N_10321,N_10017);
or U11263 (N_11263,N_10097,N_10207);
or U11264 (N_11264,N_10560,N_10122);
nand U11265 (N_11265,N_10548,N_10467);
or U11266 (N_11266,N_10805,N_10732);
nor U11267 (N_11267,N_10942,N_10441);
or U11268 (N_11268,N_10312,N_10028);
and U11269 (N_11269,N_10994,N_10617);
and U11270 (N_11270,N_10734,N_10259);
nand U11271 (N_11271,N_10768,N_10344);
and U11272 (N_11272,N_10826,N_10843);
nand U11273 (N_11273,N_10219,N_10019);
or U11274 (N_11274,N_10324,N_10285);
nand U11275 (N_11275,N_10908,N_10757);
and U11276 (N_11276,N_10981,N_10911);
or U11277 (N_11277,N_10508,N_10214);
nor U11278 (N_11278,N_10989,N_10676);
and U11279 (N_11279,N_10403,N_10014);
or U11280 (N_11280,N_10808,N_10258);
nand U11281 (N_11281,N_10189,N_10672);
xor U11282 (N_11282,N_10475,N_10029);
or U11283 (N_11283,N_10803,N_10894);
and U11284 (N_11284,N_10556,N_10430);
nand U11285 (N_11285,N_10993,N_10903);
or U11286 (N_11286,N_10562,N_10509);
or U11287 (N_11287,N_10538,N_10527);
nor U11288 (N_11288,N_10195,N_10576);
or U11289 (N_11289,N_10639,N_10317);
or U11290 (N_11290,N_10305,N_10517);
nor U11291 (N_11291,N_10320,N_10477);
and U11292 (N_11292,N_10492,N_10134);
and U11293 (N_11293,N_10080,N_10912);
nor U11294 (N_11294,N_10979,N_10712);
nor U11295 (N_11295,N_10073,N_10713);
nor U11296 (N_11296,N_10057,N_10404);
and U11297 (N_11297,N_10147,N_10260);
nand U11298 (N_11298,N_10196,N_10306);
and U11299 (N_11299,N_10229,N_10293);
nand U11300 (N_11300,N_10966,N_10597);
or U11301 (N_11301,N_10177,N_10206);
nand U11302 (N_11302,N_10174,N_10995);
nand U11303 (N_11303,N_10085,N_10759);
or U11304 (N_11304,N_10944,N_10621);
and U11305 (N_11305,N_10304,N_10529);
nor U11306 (N_11306,N_10648,N_10166);
or U11307 (N_11307,N_10180,N_10976);
nand U11308 (N_11308,N_10906,N_10274);
and U11309 (N_11309,N_10823,N_10885);
nor U11310 (N_11310,N_10844,N_10946);
or U11311 (N_11311,N_10015,N_10555);
or U11312 (N_11312,N_10592,N_10045);
nor U11313 (N_11313,N_10655,N_10036);
or U11314 (N_11314,N_10266,N_10112);
nor U11315 (N_11315,N_10952,N_10983);
or U11316 (N_11316,N_10941,N_10294);
nor U11317 (N_11317,N_10202,N_10192);
nand U11318 (N_11318,N_10225,N_10931);
nand U11319 (N_11319,N_10689,N_10963);
or U11320 (N_11320,N_10762,N_10572);
nor U11321 (N_11321,N_10054,N_10645);
or U11322 (N_11322,N_10178,N_10834);
nor U11323 (N_11323,N_10638,N_10332);
nand U11324 (N_11324,N_10035,N_10092);
and U11325 (N_11325,N_10818,N_10383);
nand U11326 (N_11326,N_10813,N_10837);
or U11327 (N_11327,N_10647,N_10533);
nand U11328 (N_11328,N_10389,N_10984);
and U11329 (N_11329,N_10800,N_10860);
xnor U11330 (N_11330,N_10596,N_10132);
and U11331 (N_11331,N_10875,N_10372);
nand U11332 (N_11332,N_10565,N_10772);
nor U11333 (N_11333,N_10888,N_10384);
xnor U11334 (N_11334,N_10571,N_10044);
or U11335 (N_11335,N_10858,N_10628);
nand U11336 (N_11336,N_10975,N_10663);
nor U11337 (N_11337,N_10298,N_10838);
nor U11338 (N_11338,N_10433,N_10031);
xor U11339 (N_11339,N_10081,N_10850);
nor U11340 (N_11340,N_10849,N_10254);
nor U11341 (N_11341,N_10620,N_10937);
nand U11342 (N_11342,N_10670,N_10930);
xor U11343 (N_11343,N_10856,N_10599);
nor U11344 (N_11344,N_10136,N_10600);
or U11345 (N_11345,N_10812,N_10232);
nor U11346 (N_11346,N_10845,N_10520);
nor U11347 (N_11347,N_10640,N_10365);
nand U11348 (N_11348,N_10752,N_10954);
and U11349 (N_11349,N_10540,N_10722);
and U11350 (N_11350,N_10819,N_10086);
xor U11351 (N_11351,N_10869,N_10393);
nor U11352 (N_11352,N_10290,N_10205);
nand U11353 (N_11353,N_10131,N_10924);
and U11354 (N_11354,N_10737,N_10011);
nand U11355 (N_11355,N_10506,N_10058);
or U11356 (N_11356,N_10240,N_10798);
nand U11357 (N_11357,N_10428,N_10286);
or U11358 (N_11358,N_10758,N_10208);
xor U11359 (N_11359,N_10879,N_10654);
or U11360 (N_11360,N_10569,N_10198);
and U11361 (N_11361,N_10992,N_10686);
xnor U11362 (N_11362,N_10338,N_10943);
and U11363 (N_11363,N_10155,N_10405);
nor U11364 (N_11364,N_10033,N_10740);
and U11365 (N_11365,N_10461,N_10986);
or U11366 (N_11366,N_10688,N_10935);
or U11367 (N_11367,N_10789,N_10047);
nor U11368 (N_11368,N_10315,N_10469);
nor U11369 (N_11369,N_10153,N_10098);
nor U11370 (N_11370,N_10149,N_10375);
nand U11371 (N_11371,N_10307,N_10152);
and U11372 (N_11372,N_10160,N_10552);
nand U11373 (N_11373,N_10730,N_10242);
and U11374 (N_11374,N_10775,N_10168);
or U11375 (N_11375,N_10878,N_10049);
nand U11376 (N_11376,N_10582,N_10525);
and U11377 (N_11377,N_10788,N_10657);
or U11378 (N_11378,N_10093,N_10733);
nor U11379 (N_11379,N_10503,N_10407);
nand U11380 (N_11380,N_10679,N_10557);
or U11381 (N_11381,N_10256,N_10873);
nand U11382 (N_11382,N_10618,N_10183);
nor U11383 (N_11383,N_10961,N_10741);
nand U11384 (N_11384,N_10919,N_10825);
and U11385 (N_11385,N_10668,N_10333);
nand U11386 (N_11386,N_10923,N_10667);
nor U11387 (N_11387,N_10501,N_10009);
nor U11388 (N_11388,N_10791,N_10822);
nand U11389 (N_11389,N_10905,N_10515);
nor U11390 (N_11390,N_10583,N_10479);
nand U11391 (N_11391,N_10999,N_10716);
or U11392 (N_11392,N_10913,N_10454);
and U11393 (N_11393,N_10032,N_10263);
and U11394 (N_11394,N_10484,N_10958);
nand U11395 (N_11395,N_10927,N_10711);
nor U11396 (N_11396,N_10238,N_10543);
or U11397 (N_11397,N_10519,N_10807);
or U11398 (N_11398,N_10188,N_10114);
xor U11399 (N_11399,N_10470,N_10411);
or U11400 (N_11400,N_10558,N_10278);
and U11401 (N_11401,N_10478,N_10693);
or U11402 (N_11402,N_10725,N_10345);
nor U11403 (N_11403,N_10348,N_10662);
nand U11404 (N_11404,N_10094,N_10351);
or U11405 (N_11405,N_10159,N_10675);
and U11406 (N_11406,N_10774,N_10859);
or U11407 (N_11407,N_10785,N_10777);
or U11408 (N_11408,N_10897,N_10460);
nor U11409 (N_11409,N_10065,N_10006);
nor U11410 (N_11410,N_10735,N_10269);
xnor U11411 (N_11411,N_10313,N_10714);
or U11412 (N_11412,N_10052,N_10537);
or U11413 (N_11413,N_10738,N_10674);
or U11414 (N_11414,N_10154,N_10754);
nand U11415 (N_11415,N_10590,N_10900);
xnor U11416 (N_11416,N_10444,N_10369);
or U11417 (N_11417,N_10939,N_10464);
nand U11418 (N_11418,N_10570,N_10265);
or U11419 (N_11419,N_10314,N_10288);
or U11420 (N_11420,N_10370,N_10034);
and U11421 (N_11421,N_10497,N_10553);
and U11422 (N_11422,N_10896,N_10495);
nand U11423 (N_11423,N_10204,N_10763);
or U11424 (N_11424,N_10027,N_10567);
or U11425 (N_11425,N_10326,N_10642);
nand U11426 (N_11426,N_10959,N_10129);
nand U11427 (N_11427,N_10363,N_10222);
or U11428 (N_11428,N_10379,N_10627);
nor U11429 (N_11429,N_10235,N_10465);
or U11430 (N_11430,N_10666,N_10486);
nor U11431 (N_11431,N_10070,N_10380);
nand U11432 (N_11432,N_10564,N_10899);
nand U11433 (N_11433,N_10726,N_10664);
xor U11434 (N_11434,N_10485,N_10162);
nor U11435 (N_11435,N_10041,N_10139);
nand U11436 (N_11436,N_10059,N_10609);
nor U11437 (N_11437,N_10573,N_10329);
nor U11438 (N_11438,N_10161,N_10226);
xnor U11439 (N_11439,N_10586,N_10292);
or U11440 (N_11440,N_10446,N_10108);
and U11441 (N_11441,N_10026,N_10413);
xor U11442 (N_11442,N_10355,N_10504);
or U11443 (N_11443,N_10123,N_10046);
nor U11444 (N_11444,N_10359,N_10227);
and U11445 (N_11445,N_10309,N_10255);
nand U11446 (N_11446,N_10833,N_10516);
or U11447 (N_11447,N_10248,N_10953);
or U11448 (N_11448,N_10408,N_10247);
or U11449 (N_11449,N_10273,N_10395);
nand U11450 (N_11450,N_10998,N_10231);
nor U11451 (N_11451,N_10440,N_10563);
or U11452 (N_11452,N_10425,N_10331);
or U11453 (N_11453,N_10868,N_10076);
or U11454 (N_11454,N_10289,N_10116);
or U11455 (N_11455,N_10436,N_10252);
or U11456 (N_11456,N_10589,N_10074);
or U11457 (N_11457,N_10115,N_10230);
nand U11458 (N_11458,N_10749,N_10257);
nand U11459 (N_11459,N_10821,N_10023);
and U11460 (N_11460,N_10416,N_10179);
nand U11461 (N_11461,N_10985,N_10072);
or U11462 (N_11462,N_10480,N_10087);
or U11463 (N_11463,N_10371,N_10606);
nor U11464 (N_11464,N_10173,N_10060);
nor U11465 (N_11465,N_10003,N_10472);
nand U11466 (N_11466,N_10890,N_10852);
or U11467 (N_11467,N_10635,N_10524);
and U11468 (N_11468,N_10855,N_10483);
nor U11469 (N_11469,N_10165,N_10840);
or U11470 (N_11470,N_10167,N_10124);
nand U11471 (N_11471,N_10346,N_10421);
nor U11472 (N_11472,N_10650,N_10234);
nor U11473 (N_11473,N_10303,N_10661);
nor U11474 (N_11474,N_10579,N_10581);
xnor U11475 (N_11475,N_10021,N_10437);
and U11476 (N_11476,N_10130,N_10145);
nor U11477 (N_11477,N_10409,N_10602);
or U11478 (N_11478,N_10536,N_10882);
nor U11479 (N_11479,N_10801,N_10863);
xnor U11480 (N_11480,N_10972,N_10163);
nor U11481 (N_11481,N_10350,N_10857);
and U11482 (N_11482,N_10866,N_10422);
or U11483 (N_11483,N_10977,N_10656);
nand U11484 (N_11484,N_10692,N_10545);
nor U11485 (N_11485,N_10415,N_10316);
and U11486 (N_11486,N_10071,N_10652);
nand U11487 (N_11487,N_10990,N_10644);
nor U11488 (N_11488,N_10410,N_10604);
and U11489 (N_11489,N_10148,N_10535);
and U11490 (N_11490,N_10629,N_10964);
or U11491 (N_11491,N_10544,N_10815);
or U11492 (N_11492,N_10601,N_10050);
or U11493 (N_11493,N_10836,N_10513);
and U11494 (N_11494,N_10096,N_10068);
and U11495 (N_11495,N_10082,N_10498);
xnor U11496 (N_11496,N_10764,N_10767);
nor U11497 (N_11497,N_10061,N_10381);
nand U11498 (N_11498,N_10916,N_10926);
nand U11499 (N_11499,N_10594,N_10181);
and U11500 (N_11500,N_10905,N_10875);
or U11501 (N_11501,N_10925,N_10451);
or U11502 (N_11502,N_10774,N_10256);
and U11503 (N_11503,N_10326,N_10293);
nand U11504 (N_11504,N_10492,N_10031);
nand U11505 (N_11505,N_10406,N_10002);
xor U11506 (N_11506,N_10499,N_10077);
xnor U11507 (N_11507,N_10778,N_10263);
xnor U11508 (N_11508,N_10334,N_10648);
nor U11509 (N_11509,N_10333,N_10304);
or U11510 (N_11510,N_10456,N_10879);
or U11511 (N_11511,N_10637,N_10831);
or U11512 (N_11512,N_10887,N_10089);
and U11513 (N_11513,N_10686,N_10291);
nor U11514 (N_11514,N_10284,N_10945);
nor U11515 (N_11515,N_10912,N_10976);
and U11516 (N_11516,N_10324,N_10230);
or U11517 (N_11517,N_10444,N_10052);
nand U11518 (N_11518,N_10223,N_10244);
xnor U11519 (N_11519,N_10468,N_10071);
xnor U11520 (N_11520,N_10567,N_10868);
nor U11521 (N_11521,N_10973,N_10949);
nor U11522 (N_11522,N_10409,N_10057);
and U11523 (N_11523,N_10654,N_10471);
or U11524 (N_11524,N_10436,N_10685);
nand U11525 (N_11525,N_10912,N_10847);
or U11526 (N_11526,N_10335,N_10522);
xor U11527 (N_11527,N_10892,N_10383);
and U11528 (N_11528,N_10200,N_10270);
nor U11529 (N_11529,N_10608,N_10807);
or U11530 (N_11530,N_10571,N_10457);
or U11531 (N_11531,N_10138,N_10918);
nor U11532 (N_11532,N_10061,N_10441);
and U11533 (N_11533,N_10067,N_10851);
or U11534 (N_11534,N_10026,N_10009);
xor U11535 (N_11535,N_10368,N_10463);
nor U11536 (N_11536,N_10264,N_10973);
nor U11537 (N_11537,N_10255,N_10936);
and U11538 (N_11538,N_10515,N_10326);
and U11539 (N_11539,N_10930,N_10803);
or U11540 (N_11540,N_10873,N_10056);
and U11541 (N_11541,N_10640,N_10309);
and U11542 (N_11542,N_10448,N_10898);
nand U11543 (N_11543,N_10191,N_10687);
and U11544 (N_11544,N_10568,N_10369);
nand U11545 (N_11545,N_10983,N_10851);
or U11546 (N_11546,N_10567,N_10571);
nand U11547 (N_11547,N_10725,N_10258);
or U11548 (N_11548,N_10563,N_10027);
nor U11549 (N_11549,N_10532,N_10602);
xor U11550 (N_11550,N_10182,N_10575);
and U11551 (N_11551,N_10306,N_10867);
xnor U11552 (N_11552,N_10260,N_10484);
nand U11553 (N_11553,N_10654,N_10283);
and U11554 (N_11554,N_10439,N_10481);
xnor U11555 (N_11555,N_10144,N_10987);
or U11556 (N_11556,N_10501,N_10785);
or U11557 (N_11557,N_10138,N_10833);
or U11558 (N_11558,N_10830,N_10811);
and U11559 (N_11559,N_10521,N_10630);
and U11560 (N_11560,N_10056,N_10738);
nor U11561 (N_11561,N_10410,N_10577);
nand U11562 (N_11562,N_10875,N_10651);
nor U11563 (N_11563,N_10756,N_10775);
or U11564 (N_11564,N_10979,N_10024);
or U11565 (N_11565,N_10137,N_10894);
or U11566 (N_11566,N_10748,N_10356);
nand U11567 (N_11567,N_10863,N_10091);
and U11568 (N_11568,N_10864,N_10476);
nand U11569 (N_11569,N_10615,N_10343);
or U11570 (N_11570,N_10336,N_10988);
or U11571 (N_11571,N_10116,N_10628);
and U11572 (N_11572,N_10023,N_10615);
or U11573 (N_11573,N_10128,N_10728);
nor U11574 (N_11574,N_10941,N_10495);
or U11575 (N_11575,N_10756,N_10721);
or U11576 (N_11576,N_10152,N_10681);
or U11577 (N_11577,N_10794,N_10869);
or U11578 (N_11578,N_10780,N_10656);
nor U11579 (N_11579,N_10730,N_10792);
nand U11580 (N_11580,N_10875,N_10954);
and U11581 (N_11581,N_10526,N_10456);
or U11582 (N_11582,N_10028,N_10482);
or U11583 (N_11583,N_10402,N_10266);
and U11584 (N_11584,N_10082,N_10292);
nor U11585 (N_11585,N_10396,N_10696);
nand U11586 (N_11586,N_10809,N_10575);
and U11587 (N_11587,N_10240,N_10402);
and U11588 (N_11588,N_10878,N_10524);
and U11589 (N_11589,N_10633,N_10354);
and U11590 (N_11590,N_10191,N_10142);
nand U11591 (N_11591,N_10559,N_10719);
nand U11592 (N_11592,N_10835,N_10959);
nor U11593 (N_11593,N_10277,N_10814);
and U11594 (N_11594,N_10841,N_10770);
nor U11595 (N_11595,N_10269,N_10792);
nor U11596 (N_11596,N_10339,N_10860);
or U11597 (N_11597,N_10768,N_10703);
and U11598 (N_11598,N_10042,N_10616);
and U11599 (N_11599,N_10216,N_10245);
nor U11600 (N_11600,N_10284,N_10585);
or U11601 (N_11601,N_10606,N_10746);
nand U11602 (N_11602,N_10446,N_10393);
and U11603 (N_11603,N_10169,N_10568);
and U11604 (N_11604,N_10375,N_10796);
and U11605 (N_11605,N_10149,N_10813);
nor U11606 (N_11606,N_10709,N_10840);
and U11607 (N_11607,N_10493,N_10829);
and U11608 (N_11608,N_10694,N_10346);
xor U11609 (N_11609,N_10641,N_10366);
or U11610 (N_11610,N_10481,N_10511);
and U11611 (N_11611,N_10460,N_10515);
xnor U11612 (N_11612,N_10797,N_10047);
and U11613 (N_11613,N_10941,N_10704);
and U11614 (N_11614,N_10691,N_10554);
nand U11615 (N_11615,N_10786,N_10257);
xnor U11616 (N_11616,N_10790,N_10870);
nor U11617 (N_11617,N_10313,N_10088);
or U11618 (N_11618,N_10722,N_10780);
nor U11619 (N_11619,N_10852,N_10554);
or U11620 (N_11620,N_10035,N_10615);
nor U11621 (N_11621,N_10232,N_10312);
nor U11622 (N_11622,N_10777,N_10539);
xor U11623 (N_11623,N_10708,N_10458);
nand U11624 (N_11624,N_10266,N_10967);
and U11625 (N_11625,N_10666,N_10191);
xnor U11626 (N_11626,N_10444,N_10021);
or U11627 (N_11627,N_10424,N_10233);
nor U11628 (N_11628,N_10099,N_10213);
nor U11629 (N_11629,N_10728,N_10203);
nor U11630 (N_11630,N_10714,N_10829);
nor U11631 (N_11631,N_10969,N_10918);
or U11632 (N_11632,N_10551,N_10619);
and U11633 (N_11633,N_10706,N_10852);
or U11634 (N_11634,N_10004,N_10289);
nand U11635 (N_11635,N_10949,N_10554);
nor U11636 (N_11636,N_10242,N_10024);
nor U11637 (N_11637,N_10064,N_10687);
and U11638 (N_11638,N_10183,N_10307);
nand U11639 (N_11639,N_10305,N_10337);
and U11640 (N_11640,N_10961,N_10958);
and U11641 (N_11641,N_10068,N_10964);
or U11642 (N_11642,N_10105,N_10080);
nand U11643 (N_11643,N_10336,N_10006);
nand U11644 (N_11644,N_10982,N_10195);
and U11645 (N_11645,N_10018,N_10464);
nand U11646 (N_11646,N_10721,N_10659);
and U11647 (N_11647,N_10269,N_10971);
nand U11648 (N_11648,N_10073,N_10765);
nor U11649 (N_11649,N_10889,N_10370);
nand U11650 (N_11650,N_10853,N_10069);
nand U11651 (N_11651,N_10746,N_10408);
and U11652 (N_11652,N_10353,N_10708);
or U11653 (N_11653,N_10756,N_10724);
and U11654 (N_11654,N_10678,N_10280);
xnor U11655 (N_11655,N_10146,N_10489);
or U11656 (N_11656,N_10576,N_10233);
and U11657 (N_11657,N_10123,N_10775);
or U11658 (N_11658,N_10081,N_10119);
nand U11659 (N_11659,N_10460,N_10534);
xnor U11660 (N_11660,N_10979,N_10392);
and U11661 (N_11661,N_10562,N_10768);
or U11662 (N_11662,N_10350,N_10744);
or U11663 (N_11663,N_10422,N_10473);
nand U11664 (N_11664,N_10402,N_10437);
and U11665 (N_11665,N_10113,N_10034);
and U11666 (N_11666,N_10527,N_10053);
and U11667 (N_11667,N_10460,N_10071);
nor U11668 (N_11668,N_10755,N_10186);
or U11669 (N_11669,N_10426,N_10721);
nand U11670 (N_11670,N_10916,N_10186);
nor U11671 (N_11671,N_10154,N_10906);
nor U11672 (N_11672,N_10222,N_10353);
nor U11673 (N_11673,N_10302,N_10004);
nor U11674 (N_11674,N_10598,N_10252);
or U11675 (N_11675,N_10830,N_10271);
nand U11676 (N_11676,N_10835,N_10132);
and U11677 (N_11677,N_10667,N_10408);
or U11678 (N_11678,N_10701,N_10385);
or U11679 (N_11679,N_10913,N_10941);
nand U11680 (N_11680,N_10450,N_10985);
xor U11681 (N_11681,N_10316,N_10468);
or U11682 (N_11682,N_10645,N_10832);
xnor U11683 (N_11683,N_10937,N_10379);
nor U11684 (N_11684,N_10167,N_10874);
nor U11685 (N_11685,N_10840,N_10762);
nand U11686 (N_11686,N_10202,N_10263);
and U11687 (N_11687,N_10503,N_10130);
nor U11688 (N_11688,N_10851,N_10199);
and U11689 (N_11689,N_10816,N_10807);
and U11690 (N_11690,N_10612,N_10356);
nor U11691 (N_11691,N_10084,N_10935);
and U11692 (N_11692,N_10928,N_10555);
nor U11693 (N_11693,N_10826,N_10334);
and U11694 (N_11694,N_10831,N_10276);
and U11695 (N_11695,N_10211,N_10953);
xor U11696 (N_11696,N_10266,N_10028);
nand U11697 (N_11697,N_10432,N_10794);
nand U11698 (N_11698,N_10264,N_10246);
nor U11699 (N_11699,N_10701,N_10845);
or U11700 (N_11700,N_10730,N_10608);
and U11701 (N_11701,N_10827,N_10147);
nor U11702 (N_11702,N_10011,N_10865);
xor U11703 (N_11703,N_10264,N_10752);
or U11704 (N_11704,N_10149,N_10640);
nor U11705 (N_11705,N_10078,N_10397);
nor U11706 (N_11706,N_10918,N_10409);
and U11707 (N_11707,N_10849,N_10479);
nand U11708 (N_11708,N_10835,N_10204);
or U11709 (N_11709,N_10115,N_10409);
nor U11710 (N_11710,N_10839,N_10174);
or U11711 (N_11711,N_10103,N_10504);
nand U11712 (N_11712,N_10475,N_10088);
or U11713 (N_11713,N_10312,N_10176);
or U11714 (N_11714,N_10600,N_10919);
and U11715 (N_11715,N_10249,N_10831);
nand U11716 (N_11716,N_10257,N_10706);
or U11717 (N_11717,N_10228,N_10392);
nor U11718 (N_11718,N_10200,N_10943);
nand U11719 (N_11719,N_10298,N_10867);
or U11720 (N_11720,N_10317,N_10440);
and U11721 (N_11721,N_10331,N_10337);
nor U11722 (N_11722,N_10716,N_10052);
and U11723 (N_11723,N_10567,N_10484);
nor U11724 (N_11724,N_10311,N_10887);
or U11725 (N_11725,N_10912,N_10716);
and U11726 (N_11726,N_10532,N_10150);
nand U11727 (N_11727,N_10620,N_10278);
or U11728 (N_11728,N_10375,N_10668);
or U11729 (N_11729,N_10115,N_10860);
or U11730 (N_11730,N_10181,N_10643);
and U11731 (N_11731,N_10423,N_10078);
nand U11732 (N_11732,N_10241,N_10672);
xor U11733 (N_11733,N_10552,N_10790);
nor U11734 (N_11734,N_10997,N_10563);
and U11735 (N_11735,N_10569,N_10455);
nor U11736 (N_11736,N_10041,N_10040);
xnor U11737 (N_11737,N_10156,N_10577);
nor U11738 (N_11738,N_10561,N_10949);
nor U11739 (N_11739,N_10761,N_10630);
or U11740 (N_11740,N_10165,N_10953);
xnor U11741 (N_11741,N_10944,N_10075);
and U11742 (N_11742,N_10179,N_10866);
and U11743 (N_11743,N_10251,N_10825);
nand U11744 (N_11744,N_10510,N_10424);
and U11745 (N_11745,N_10831,N_10550);
or U11746 (N_11746,N_10863,N_10439);
nor U11747 (N_11747,N_10623,N_10279);
xnor U11748 (N_11748,N_10836,N_10082);
nor U11749 (N_11749,N_10459,N_10238);
and U11750 (N_11750,N_10637,N_10155);
nor U11751 (N_11751,N_10034,N_10654);
nor U11752 (N_11752,N_10035,N_10626);
or U11753 (N_11753,N_10224,N_10320);
nand U11754 (N_11754,N_10183,N_10462);
nor U11755 (N_11755,N_10971,N_10120);
nand U11756 (N_11756,N_10445,N_10652);
or U11757 (N_11757,N_10204,N_10081);
or U11758 (N_11758,N_10016,N_10287);
and U11759 (N_11759,N_10971,N_10355);
nand U11760 (N_11760,N_10529,N_10653);
nor U11761 (N_11761,N_10591,N_10924);
nand U11762 (N_11762,N_10592,N_10698);
nand U11763 (N_11763,N_10364,N_10281);
nand U11764 (N_11764,N_10933,N_10949);
nor U11765 (N_11765,N_10847,N_10075);
xor U11766 (N_11766,N_10999,N_10255);
or U11767 (N_11767,N_10579,N_10422);
xnor U11768 (N_11768,N_10951,N_10152);
nand U11769 (N_11769,N_10035,N_10883);
nor U11770 (N_11770,N_10109,N_10892);
or U11771 (N_11771,N_10744,N_10793);
or U11772 (N_11772,N_10734,N_10814);
nand U11773 (N_11773,N_10499,N_10789);
and U11774 (N_11774,N_10725,N_10276);
nand U11775 (N_11775,N_10317,N_10396);
nor U11776 (N_11776,N_10565,N_10985);
nor U11777 (N_11777,N_10628,N_10390);
nor U11778 (N_11778,N_10610,N_10499);
or U11779 (N_11779,N_10203,N_10304);
and U11780 (N_11780,N_10155,N_10353);
nor U11781 (N_11781,N_10296,N_10824);
and U11782 (N_11782,N_10168,N_10462);
nand U11783 (N_11783,N_10033,N_10450);
xor U11784 (N_11784,N_10663,N_10351);
nor U11785 (N_11785,N_10064,N_10810);
nand U11786 (N_11786,N_10682,N_10662);
nand U11787 (N_11787,N_10326,N_10224);
xnor U11788 (N_11788,N_10268,N_10401);
and U11789 (N_11789,N_10154,N_10846);
and U11790 (N_11790,N_10708,N_10947);
nand U11791 (N_11791,N_10310,N_10629);
or U11792 (N_11792,N_10679,N_10230);
nand U11793 (N_11793,N_10629,N_10920);
nand U11794 (N_11794,N_10782,N_10812);
and U11795 (N_11795,N_10196,N_10605);
or U11796 (N_11796,N_10423,N_10262);
nor U11797 (N_11797,N_10593,N_10325);
and U11798 (N_11798,N_10825,N_10449);
and U11799 (N_11799,N_10607,N_10537);
nor U11800 (N_11800,N_10213,N_10049);
xor U11801 (N_11801,N_10533,N_10020);
or U11802 (N_11802,N_10263,N_10049);
nand U11803 (N_11803,N_10790,N_10937);
nor U11804 (N_11804,N_10255,N_10953);
nor U11805 (N_11805,N_10145,N_10529);
nand U11806 (N_11806,N_10658,N_10586);
or U11807 (N_11807,N_10626,N_10511);
nand U11808 (N_11808,N_10038,N_10765);
nand U11809 (N_11809,N_10666,N_10665);
and U11810 (N_11810,N_10712,N_10144);
and U11811 (N_11811,N_10653,N_10919);
nand U11812 (N_11812,N_10470,N_10763);
or U11813 (N_11813,N_10737,N_10745);
nand U11814 (N_11814,N_10935,N_10094);
or U11815 (N_11815,N_10541,N_10003);
xnor U11816 (N_11816,N_10696,N_10581);
nor U11817 (N_11817,N_10328,N_10023);
or U11818 (N_11818,N_10505,N_10357);
xor U11819 (N_11819,N_10297,N_10750);
nand U11820 (N_11820,N_10273,N_10471);
and U11821 (N_11821,N_10171,N_10353);
and U11822 (N_11822,N_10822,N_10736);
and U11823 (N_11823,N_10377,N_10754);
and U11824 (N_11824,N_10478,N_10118);
xnor U11825 (N_11825,N_10627,N_10131);
nand U11826 (N_11826,N_10290,N_10027);
nor U11827 (N_11827,N_10067,N_10622);
nor U11828 (N_11828,N_10004,N_10720);
nand U11829 (N_11829,N_10553,N_10656);
and U11830 (N_11830,N_10593,N_10505);
nor U11831 (N_11831,N_10162,N_10589);
nand U11832 (N_11832,N_10924,N_10498);
nor U11833 (N_11833,N_10550,N_10685);
nand U11834 (N_11834,N_10848,N_10086);
nor U11835 (N_11835,N_10521,N_10764);
nor U11836 (N_11836,N_10471,N_10368);
or U11837 (N_11837,N_10089,N_10631);
xnor U11838 (N_11838,N_10943,N_10055);
xor U11839 (N_11839,N_10659,N_10190);
nor U11840 (N_11840,N_10217,N_10499);
and U11841 (N_11841,N_10896,N_10035);
or U11842 (N_11842,N_10184,N_10936);
nor U11843 (N_11843,N_10383,N_10097);
and U11844 (N_11844,N_10097,N_10378);
and U11845 (N_11845,N_10266,N_10311);
xnor U11846 (N_11846,N_10909,N_10327);
nand U11847 (N_11847,N_10744,N_10984);
nand U11848 (N_11848,N_10700,N_10046);
or U11849 (N_11849,N_10303,N_10616);
and U11850 (N_11850,N_10912,N_10631);
or U11851 (N_11851,N_10947,N_10524);
nand U11852 (N_11852,N_10940,N_10964);
nor U11853 (N_11853,N_10760,N_10316);
nand U11854 (N_11854,N_10596,N_10294);
xor U11855 (N_11855,N_10964,N_10122);
nand U11856 (N_11856,N_10754,N_10694);
and U11857 (N_11857,N_10716,N_10531);
and U11858 (N_11858,N_10091,N_10335);
xor U11859 (N_11859,N_10660,N_10364);
nor U11860 (N_11860,N_10918,N_10434);
or U11861 (N_11861,N_10107,N_10539);
nand U11862 (N_11862,N_10766,N_10008);
nand U11863 (N_11863,N_10505,N_10240);
or U11864 (N_11864,N_10039,N_10100);
nand U11865 (N_11865,N_10576,N_10501);
nor U11866 (N_11866,N_10183,N_10426);
or U11867 (N_11867,N_10641,N_10566);
and U11868 (N_11868,N_10761,N_10414);
nor U11869 (N_11869,N_10996,N_10528);
nand U11870 (N_11870,N_10450,N_10089);
and U11871 (N_11871,N_10172,N_10205);
nor U11872 (N_11872,N_10081,N_10573);
or U11873 (N_11873,N_10589,N_10878);
or U11874 (N_11874,N_10142,N_10112);
or U11875 (N_11875,N_10425,N_10666);
and U11876 (N_11876,N_10972,N_10564);
nor U11877 (N_11877,N_10501,N_10166);
nor U11878 (N_11878,N_10040,N_10816);
and U11879 (N_11879,N_10512,N_10358);
nand U11880 (N_11880,N_10067,N_10198);
or U11881 (N_11881,N_10976,N_10809);
nor U11882 (N_11882,N_10516,N_10265);
or U11883 (N_11883,N_10305,N_10780);
or U11884 (N_11884,N_10772,N_10736);
nor U11885 (N_11885,N_10294,N_10318);
xor U11886 (N_11886,N_10247,N_10800);
and U11887 (N_11887,N_10925,N_10423);
or U11888 (N_11888,N_10598,N_10878);
nor U11889 (N_11889,N_10148,N_10829);
or U11890 (N_11890,N_10848,N_10919);
nand U11891 (N_11891,N_10923,N_10571);
xnor U11892 (N_11892,N_10170,N_10202);
nand U11893 (N_11893,N_10938,N_10351);
or U11894 (N_11894,N_10651,N_10691);
and U11895 (N_11895,N_10091,N_10127);
or U11896 (N_11896,N_10513,N_10820);
nand U11897 (N_11897,N_10548,N_10970);
and U11898 (N_11898,N_10653,N_10569);
or U11899 (N_11899,N_10093,N_10736);
nand U11900 (N_11900,N_10438,N_10561);
and U11901 (N_11901,N_10912,N_10942);
or U11902 (N_11902,N_10118,N_10125);
nor U11903 (N_11903,N_10375,N_10762);
nand U11904 (N_11904,N_10256,N_10268);
or U11905 (N_11905,N_10658,N_10505);
nand U11906 (N_11906,N_10301,N_10119);
and U11907 (N_11907,N_10488,N_10742);
nand U11908 (N_11908,N_10393,N_10814);
nand U11909 (N_11909,N_10210,N_10111);
nor U11910 (N_11910,N_10623,N_10162);
or U11911 (N_11911,N_10866,N_10521);
nand U11912 (N_11912,N_10114,N_10277);
nand U11913 (N_11913,N_10147,N_10521);
and U11914 (N_11914,N_10329,N_10609);
or U11915 (N_11915,N_10227,N_10040);
nand U11916 (N_11916,N_10497,N_10405);
and U11917 (N_11917,N_10471,N_10628);
nor U11918 (N_11918,N_10319,N_10696);
nand U11919 (N_11919,N_10610,N_10244);
nand U11920 (N_11920,N_10386,N_10411);
xnor U11921 (N_11921,N_10055,N_10985);
or U11922 (N_11922,N_10941,N_10185);
nor U11923 (N_11923,N_10736,N_10874);
xor U11924 (N_11924,N_10393,N_10741);
nor U11925 (N_11925,N_10639,N_10694);
xnor U11926 (N_11926,N_10558,N_10140);
nand U11927 (N_11927,N_10729,N_10427);
nor U11928 (N_11928,N_10197,N_10099);
nand U11929 (N_11929,N_10648,N_10366);
xor U11930 (N_11930,N_10491,N_10379);
or U11931 (N_11931,N_10733,N_10383);
nor U11932 (N_11932,N_10604,N_10596);
or U11933 (N_11933,N_10790,N_10581);
nor U11934 (N_11934,N_10678,N_10805);
or U11935 (N_11935,N_10731,N_10889);
and U11936 (N_11936,N_10828,N_10090);
nand U11937 (N_11937,N_10851,N_10049);
nor U11938 (N_11938,N_10848,N_10037);
nor U11939 (N_11939,N_10721,N_10879);
nor U11940 (N_11940,N_10720,N_10192);
and U11941 (N_11941,N_10583,N_10929);
xor U11942 (N_11942,N_10656,N_10226);
and U11943 (N_11943,N_10598,N_10911);
xnor U11944 (N_11944,N_10724,N_10387);
and U11945 (N_11945,N_10006,N_10158);
nand U11946 (N_11946,N_10317,N_10291);
and U11947 (N_11947,N_10161,N_10048);
and U11948 (N_11948,N_10286,N_10081);
or U11949 (N_11949,N_10114,N_10916);
nor U11950 (N_11950,N_10102,N_10796);
nand U11951 (N_11951,N_10889,N_10497);
nand U11952 (N_11952,N_10221,N_10164);
nor U11953 (N_11953,N_10341,N_10935);
or U11954 (N_11954,N_10313,N_10234);
and U11955 (N_11955,N_10935,N_10337);
or U11956 (N_11956,N_10157,N_10413);
nand U11957 (N_11957,N_10335,N_10694);
and U11958 (N_11958,N_10893,N_10946);
and U11959 (N_11959,N_10282,N_10369);
and U11960 (N_11960,N_10096,N_10033);
or U11961 (N_11961,N_10760,N_10649);
xor U11962 (N_11962,N_10755,N_10531);
and U11963 (N_11963,N_10741,N_10011);
nand U11964 (N_11964,N_10575,N_10187);
and U11965 (N_11965,N_10309,N_10558);
nor U11966 (N_11966,N_10434,N_10092);
and U11967 (N_11967,N_10775,N_10722);
or U11968 (N_11968,N_10122,N_10146);
or U11969 (N_11969,N_10883,N_10616);
xnor U11970 (N_11970,N_10504,N_10011);
or U11971 (N_11971,N_10398,N_10562);
nand U11972 (N_11972,N_10944,N_10905);
nor U11973 (N_11973,N_10418,N_10040);
or U11974 (N_11974,N_10801,N_10453);
nor U11975 (N_11975,N_10818,N_10871);
nor U11976 (N_11976,N_10281,N_10011);
or U11977 (N_11977,N_10441,N_10787);
and U11978 (N_11978,N_10633,N_10560);
or U11979 (N_11979,N_10473,N_10428);
and U11980 (N_11980,N_10875,N_10708);
nor U11981 (N_11981,N_10391,N_10032);
or U11982 (N_11982,N_10746,N_10385);
nand U11983 (N_11983,N_10827,N_10090);
or U11984 (N_11984,N_10166,N_10778);
xor U11985 (N_11985,N_10735,N_10703);
and U11986 (N_11986,N_10850,N_10241);
nor U11987 (N_11987,N_10846,N_10497);
nand U11988 (N_11988,N_10571,N_10495);
nand U11989 (N_11989,N_10313,N_10243);
or U11990 (N_11990,N_10431,N_10399);
and U11991 (N_11991,N_10129,N_10092);
or U11992 (N_11992,N_10087,N_10809);
xnor U11993 (N_11993,N_10313,N_10349);
or U11994 (N_11994,N_10159,N_10225);
and U11995 (N_11995,N_10580,N_10526);
or U11996 (N_11996,N_10519,N_10620);
nand U11997 (N_11997,N_10135,N_10708);
or U11998 (N_11998,N_10613,N_10640);
nand U11999 (N_11999,N_10939,N_10055);
or U12000 (N_12000,N_11721,N_11885);
nor U12001 (N_12001,N_11872,N_11334);
nor U12002 (N_12002,N_11296,N_11078);
nand U12003 (N_12003,N_11640,N_11681);
or U12004 (N_12004,N_11265,N_11268);
and U12005 (N_12005,N_11969,N_11896);
nand U12006 (N_12006,N_11856,N_11750);
nor U12007 (N_12007,N_11371,N_11395);
and U12008 (N_12008,N_11327,N_11238);
nand U12009 (N_12009,N_11911,N_11262);
nand U12010 (N_12010,N_11567,N_11445);
or U12011 (N_12011,N_11740,N_11847);
or U12012 (N_12012,N_11363,N_11093);
or U12013 (N_12013,N_11016,N_11424);
nor U12014 (N_12014,N_11696,N_11916);
or U12015 (N_12015,N_11904,N_11032);
nor U12016 (N_12016,N_11846,N_11170);
nor U12017 (N_12017,N_11633,N_11315);
or U12018 (N_12018,N_11050,N_11511);
and U12019 (N_12019,N_11760,N_11858);
and U12020 (N_12020,N_11456,N_11983);
and U12021 (N_12021,N_11678,N_11278);
nand U12022 (N_12022,N_11764,N_11831);
or U12023 (N_12023,N_11336,N_11018);
and U12024 (N_12024,N_11804,N_11042);
nand U12025 (N_12025,N_11167,N_11069);
nand U12026 (N_12026,N_11449,N_11840);
and U12027 (N_12027,N_11410,N_11746);
and U12028 (N_12028,N_11785,N_11477);
or U12029 (N_12029,N_11792,N_11534);
nor U12030 (N_12030,N_11544,N_11163);
or U12031 (N_12031,N_11903,N_11246);
nand U12032 (N_12032,N_11217,N_11564);
or U12033 (N_12033,N_11396,N_11450);
nor U12034 (N_12034,N_11063,N_11193);
xor U12035 (N_12035,N_11893,N_11062);
nand U12036 (N_12036,N_11214,N_11059);
nor U12037 (N_12037,N_11386,N_11144);
nor U12038 (N_12038,N_11512,N_11157);
nand U12039 (N_12039,N_11286,N_11457);
and U12040 (N_12040,N_11701,N_11699);
nand U12041 (N_12041,N_11291,N_11734);
nor U12042 (N_12042,N_11491,N_11022);
and U12043 (N_12043,N_11021,N_11901);
nor U12044 (N_12044,N_11087,N_11923);
nor U12045 (N_12045,N_11912,N_11761);
or U12046 (N_12046,N_11684,N_11254);
nand U12047 (N_12047,N_11680,N_11828);
nand U12048 (N_12048,N_11728,N_11049);
nor U12049 (N_12049,N_11682,N_11944);
nor U12050 (N_12050,N_11630,N_11955);
or U12051 (N_12051,N_11139,N_11810);
nor U12052 (N_12052,N_11205,N_11455);
or U12053 (N_12053,N_11460,N_11184);
nor U12054 (N_12054,N_11124,N_11624);
and U12055 (N_12055,N_11494,N_11741);
and U12056 (N_12056,N_11290,N_11434);
and U12057 (N_12057,N_11351,N_11462);
nor U12058 (N_12058,N_11580,N_11419);
nand U12059 (N_12059,N_11492,N_11578);
nand U12060 (N_12060,N_11694,N_11917);
nor U12061 (N_12061,N_11751,N_11364);
nand U12062 (N_12062,N_11322,N_11031);
xnor U12063 (N_12063,N_11418,N_11066);
nand U12064 (N_12064,N_11826,N_11835);
or U12065 (N_12065,N_11978,N_11388);
and U12066 (N_12066,N_11550,N_11498);
and U12067 (N_12067,N_11379,N_11330);
or U12068 (N_12068,N_11248,N_11256);
or U12069 (N_12069,N_11281,N_11987);
nand U12070 (N_12070,N_11754,N_11180);
or U12071 (N_12071,N_11933,N_11676);
nand U12072 (N_12072,N_11178,N_11739);
or U12073 (N_12073,N_11479,N_11894);
nor U12074 (N_12074,N_11713,N_11196);
nand U12075 (N_12075,N_11834,N_11801);
xor U12076 (N_12076,N_11710,N_11960);
or U12077 (N_12077,N_11165,N_11092);
xor U12078 (N_12078,N_11272,N_11690);
and U12079 (N_12079,N_11429,N_11487);
nand U12080 (N_12080,N_11519,N_11448);
or U12081 (N_12081,N_11639,N_11210);
nor U12082 (N_12082,N_11103,N_11697);
and U12083 (N_12083,N_11168,N_11907);
nor U12084 (N_12084,N_11202,N_11380);
xor U12085 (N_12085,N_11867,N_11602);
or U12086 (N_12086,N_11098,N_11158);
and U12087 (N_12087,N_11375,N_11558);
nand U12088 (N_12088,N_11687,N_11280);
and U12089 (N_12089,N_11535,N_11310);
or U12090 (N_12090,N_11902,N_11224);
or U12091 (N_12091,N_11360,N_11914);
nor U12092 (N_12092,N_11913,N_11725);
and U12093 (N_12093,N_11720,N_11161);
nand U12094 (N_12094,N_11313,N_11986);
xor U12095 (N_12095,N_11146,N_11890);
and U12096 (N_12096,N_11809,N_11897);
nor U12097 (N_12097,N_11669,N_11505);
and U12098 (N_12098,N_11420,N_11219);
or U12099 (N_12099,N_11179,N_11052);
and U12100 (N_12100,N_11467,N_11057);
nand U12101 (N_12101,N_11962,N_11811);
xor U12102 (N_12102,N_11077,N_11323);
nand U12103 (N_12103,N_11570,N_11166);
or U12104 (N_12104,N_11129,N_11878);
or U12105 (N_12105,N_11671,N_11007);
xnor U12106 (N_12106,N_11886,N_11372);
and U12107 (N_12107,N_11476,N_11316);
nor U12108 (N_12108,N_11159,N_11616);
or U12109 (N_12109,N_11083,N_11325);
xnor U12110 (N_12110,N_11125,N_11993);
xnor U12111 (N_12111,N_11777,N_11963);
and U12112 (N_12112,N_11403,N_11520);
xor U12113 (N_12113,N_11005,N_11150);
nand U12114 (N_12114,N_11939,N_11484);
and U12115 (N_12115,N_11392,N_11107);
xnor U12116 (N_12116,N_11892,N_11436);
and U12117 (N_12117,N_11156,N_11068);
nor U12118 (N_12118,N_11575,N_11645);
nand U12119 (N_12119,N_11688,N_11407);
nor U12120 (N_12120,N_11672,N_11938);
and U12121 (N_12121,N_11613,N_11474);
nor U12122 (N_12122,N_11752,N_11979);
nand U12123 (N_12123,N_11788,N_11258);
xor U12124 (N_12124,N_11096,N_11206);
and U12125 (N_12125,N_11628,N_11667);
nor U12126 (N_12126,N_11171,N_11590);
nor U12127 (N_12127,N_11047,N_11025);
and U12128 (N_12128,N_11433,N_11763);
xor U12129 (N_12129,N_11416,N_11112);
nand U12130 (N_12130,N_11757,N_11298);
nor U12131 (N_12131,N_11715,N_11515);
or U12132 (N_12132,N_11431,N_11230);
nor U12133 (N_12133,N_11413,N_11592);
nand U12134 (N_12134,N_11131,N_11088);
xor U12135 (N_12135,N_11686,N_11081);
nand U12136 (N_12136,N_11597,N_11382);
nand U12137 (N_12137,N_11441,N_11054);
and U12138 (N_12138,N_11399,N_11438);
and U12139 (N_12139,N_11880,N_11634);
xnor U12140 (N_12140,N_11173,N_11247);
nor U12141 (N_12141,N_11989,N_11461);
or U12142 (N_12142,N_11242,N_11709);
nand U12143 (N_12143,N_11612,N_11953);
and U12144 (N_12144,N_11321,N_11756);
nand U12145 (N_12145,N_11397,N_11342);
or U12146 (N_12146,N_11936,N_11727);
and U12147 (N_12147,N_11311,N_11530);
and U12148 (N_12148,N_11582,N_11120);
nand U12149 (N_12149,N_11865,N_11154);
and U12150 (N_12150,N_11666,N_11773);
nor U12151 (N_12151,N_11623,N_11164);
and U12152 (N_12152,N_11943,N_11776);
nand U12153 (N_12153,N_11390,N_11784);
and U12154 (N_12154,N_11506,N_11422);
nor U12155 (N_12155,N_11521,N_11350);
nand U12156 (N_12156,N_11931,N_11743);
xor U12157 (N_12157,N_11621,N_11266);
xnor U12158 (N_12158,N_11853,N_11679);
and U12159 (N_12159,N_11443,N_11584);
or U12160 (N_12160,N_11384,N_11961);
nand U12161 (N_12161,N_11394,N_11192);
or U12162 (N_12162,N_11502,N_11780);
nor U12163 (N_12163,N_11288,N_11444);
nand U12164 (N_12164,N_11646,N_11275);
nand U12165 (N_12165,N_11277,N_11860);
nand U12166 (N_12166,N_11004,N_11412);
and U12167 (N_12167,N_11080,N_11181);
nor U12168 (N_12168,N_11304,N_11928);
or U12169 (N_12169,N_11089,N_11562);
and U12170 (N_12170,N_11056,N_11114);
nand U12171 (N_12171,N_11825,N_11516);
nor U12172 (N_12172,N_11225,N_11653);
and U12173 (N_12173,N_11040,N_11620);
or U12174 (N_12174,N_11389,N_11329);
xnor U12175 (N_12175,N_11029,N_11373);
or U12176 (N_12176,N_11712,N_11815);
and U12177 (N_12177,N_11563,N_11947);
nor U12178 (N_12178,N_11117,N_11177);
nand U12179 (N_12179,N_11787,N_11798);
nor U12180 (N_12180,N_11014,N_11038);
and U12181 (N_12181,N_11489,N_11099);
nor U12182 (N_12182,N_11642,N_11768);
and U12183 (N_12183,N_11133,N_11400);
nor U12184 (N_12184,N_11997,N_11661);
or U12185 (N_12185,N_11340,N_11656);
or U12186 (N_12186,N_11585,N_11257);
nand U12187 (N_12187,N_11552,N_11453);
nor U12188 (N_12188,N_11898,N_11510);
xnor U12189 (N_12189,N_11331,N_11415);
nor U12190 (N_12190,N_11794,N_11465);
nand U12191 (N_12191,N_11932,N_11383);
and U12192 (N_12192,N_11952,N_11485);
and U12193 (N_12193,N_11941,N_11309);
and U12194 (N_12194,N_11097,N_11607);
or U12195 (N_12195,N_11283,N_11716);
nor U12196 (N_12196,N_11548,N_11358);
or U12197 (N_12197,N_11744,N_11660);
xor U12198 (N_12198,N_11188,N_11136);
and U12199 (N_12199,N_11946,N_11971);
or U12200 (N_12200,N_11199,N_11668);
nand U12201 (N_12201,N_11020,N_11104);
and U12202 (N_12202,N_11244,N_11176);
or U12203 (N_12203,N_11977,N_11499);
nand U12204 (N_12204,N_11920,N_11006);
nand U12205 (N_12205,N_11127,N_11724);
or U12206 (N_12206,N_11800,N_11102);
or U12207 (N_12207,N_11036,N_11027);
or U12208 (N_12208,N_11532,N_11749);
nand U12209 (N_12209,N_11837,N_11189);
nor U12210 (N_12210,N_11705,N_11355);
nand U12211 (N_12211,N_11733,N_11895);
or U12212 (N_12212,N_11204,N_11545);
nor U12213 (N_12213,N_11058,N_11200);
and U12214 (N_12214,N_11803,N_11755);
or U12215 (N_12215,N_11293,N_11393);
or U12216 (N_12216,N_11574,N_11560);
and U12217 (N_12217,N_11683,N_11781);
or U12218 (N_12218,N_11100,N_11387);
nor U12219 (N_12219,N_11033,N_11561);
nand U12220 (N_12220,N_11879,N_11013);
xnor U12221 (N_12221,N_11579,N_11041);
nor U12222 (N_12222,N_11536,N_11985);
nand U12223 (N_12223,N_11957,N_11859);
or U12224 (N_12224,N_11595,N_11748);
xor U12225 (N_12225,N_11354,N_11259);
nand U12226 (N_12226,N_11368,N_11113);
or U12227 (N_12227,N_11486,N_11269);
or U12228 (N_12228,N_11338,N_11875);
nand U12229 (N_12229,N_11593,N_11026);
nand U12230 (N_12230,N_11190,N_11786);
nor U12231 (N_12231,N_11588,N_11719);
nand U12232 (N_12232,N_11654,N_11411);
and U12233 (N_12233,N_11982,N_11201);
xor U12234 (N_12234,N_11421,N_11468);
and U12235 (N_12235,N_11542,N_11148);
or U12236 (N_12236,N_11480,N_11673);
or U12237 (N_12237,N_11111,N_11643);
or U12238 (N_12238,N_11974,N_11820);
xnor U12239 (N_12239,N_11182,N_11635);
or U12240 (N_12240,N_11430,N_11723);
or U12241 (N_12241,N_11629,N_11888);
nand U12242 (N_12242,N_11609,N_11874);
xnor U12243 (N_12243,N_11615,N_11263);
or U12244 (N_12244,N_11503,N_11600);
nand U12245 (N_12245,N_11228,N_11346);
nand U12246 (N_12246,N_11704,N_11866);
or U12247 (N_12247,N_11324,N_11990);
nand U12248 (N_12248,N_11626,N_11827);
nand U12249 (N_12249,N_11481,N_11958);
nor U12250 (N_12250,N_11848,N_11314);
nand U12251 (N_12251,N_11197,N_11814);
and U12252 (N_12252,N_11950,N_11547);
and U12253 (N_12253,N_11126,N_11900);
and U12254 (N_12254,N_11657,N_11121);
nor U12255 (N_12255,N_11599,N_11488);
xor U12256 (N_12256,N_11299,N_11402);
or U12257 (N_12257,N_11968,N_11589);
and U12258 (N_12258,N_11249,N_11398);
nor U12259 (N_12259,N_11935,N_11862);
and U12260 (N_12260,N_11861,N_11426);
nor U12261 (N_12261,N_11906,N_11769);
or U12262 (N_12262,N_11253,N_11638);
xor U12263 (N_12263,N_11789,N_11405);
or U12264 (N_12264,N_11128,N_11307);
or U12265 (N_12265,N_11352,N_11483);
and U12266 (N_12266,N_11348,N_11587);
or U12267 (N_12267,N_11135,N_11852);
and U12268 (N_12268,N_11401,N_11586);
nand U12269 (N_12269,N_11541,N_11658);
or U12270 (N_12270,N_11086,N_11425);
nand U12271 (N_12271,N_11142,N_11458);
and U12272 (N_12272,N_11915,N_11264);
or U12273 (N_12273,N_11849,N_11076);
or U12274 (N_12274,N_11300,N_11821);
xor U12275 (N_12275,N_11094,N_11791);
or U12276 (N_12276,N_11292,N_11767);
and U12277 (N_12277,N_11836,N_11353);
or U12278 (N_12278,N_11959,N_11965);
or U12279 (N_12279,N_11319,N_11707);
or U12280 (N_12280,N_11223,N_11326);
xor U12281 (N_12281,N_11910,N_11736);
or U12282 (N_12282,N_11137,N_11540);
or U12283 (N_12283,N_11366,N_11664);
or U12284 (N_12284,N_11212,N_11509);
nor U12285 (N_12285,N_11118,N_11030);
or U12286 (N_12286,N_11070,N_11140);
or U12287 (N_12287,N_11169,N_11617);
nand U12288 (N_12288,N_11537,N_11677);
or U12289 (N_12289,N_11122,N_11610);
and U12290 (N_12290,N_11863,N_11194);
and U12291 (N_12291,N_11447,N_11216);
nor U12292 (N_12292,N_11605,N_11162);
nand U12293 (N_12293,N_11970,N_11949);
and U12294 (N_12294,N_11344,N_11466);
or U12295 (N_12295,N_11706,N_11622);
and U12296 (N_12296,N_11691,N_11463);
and U12297 (N_12297,N_11877,N_11883);
nand U12298 (N_12298,N_11869,N_11546);
nor U12299 (N_12299,N_11708,N_11003);
and U12300 (N_12300,N_11925,N_11737);
and U12301 (N_12301,N_11497,N_11881);
or U12302 (N_12302,N_11591,N_11454);
nand U12303 (N_12303,N_11349,N_11374);
and U12304 (N_12304,N_11976,N_11339);
and U12305 (N_12305,N_11967,N_11566);
nand U12306 (N_12306,N_11842,N_11889);
and U12307 (N_12307,N_11034,N_11758);
xor U12308 (N_12308,N_11432,N_11260);
nand U12309 (N_12309,N_11115,N_11730);
nand U12310 (N_12310,N_11899,N_11064);
nor U12311 (N_12311,N_11328,N_11303);
nor U12312 (N_12312,N_11975,N_11844);
or U12313 (N_12313,N_11337,N_11215);
nand U12314 (N_12314,N_11237,N_11551);
xor U12315 (N_12315,N_11252,N_11318);
or U12316 (N_12316,N_11472,N_11294);
nand U12317 (N_12317,N_11700,N_11729);
or U12318 (N_12318,N_11555,N_11071);
nor U12319 (N_12319,N_11649,N_11608);
or U12320 (N_12320,N_11232,N_11009);
xnor U12321 (N_12321,N_11830,N_11945);
and U12322 (N_12322,N_11245,N_11981);
nor U12323 (N_12323,N_11475,N_11940);
xnor U12324 (N_12324,N_11221,N_11067);
nand U12325 (N_12325,N_11175,N_11464);
nand U12326 (N_12326,N_11060,N_11378);
xor U12327 (N_12327,N_11999,N_11045);
nand U12328 (N_12328,N_11583,N_11692);
nand U12329 (N_12329,N_11942,N_11377);
xor U12330 (N_12330,N_11948,N_11934);
nor U12331 (N_12331,N_11345,N_11408);
and U12332 (N_12332,N_11841,N_11854);
or U12333 (N_12333,N_11048,N_11569);
nor U12334 (N_12334,N_11251,N_11614);
and U12335 (N_12335,N_11183,N_11864);
and U12336 (N_12336,N_11085,N_11271);
and U12337 (N_12337,N_11601,N_11356);
nand U12338 (N_12338,N_11305,N_11195);
nand U12339 (N_12339,N_11731,N_11808);
nor U12340 (N_12340,N_11812,N_11236);
nand U12341 (N_12341,N_11153,N_11442);
and U12342 (N_12342,N_11665,N_11308);
nor U12343 (N_12343,N_11742,N_11797);
nor U12344 (N_12344,N_11851,N_11522);
or U12345 (N_12345,N_11250,N_11317);
or U12346 (N_12346,N_11529,N_11446);
and U12347 (N_12347,N_11526,N_11823);
or U12348 (N_12348,N_11527,N_11119);
and U12349 (N_12349,N_11650,N_11276);
nand U12350 (N_12350,N_11759,N_11839);
nand U12351 (N_12351,N_11270,N_11576);
xor U12352 (N_12352,N_11469,N_11651);
and U12353 (N_12353,N_11289,N_11500);
and U12354 (N_12354,N_11306,N_11010);
or U12355 (N_12355,N_11185,N_11929);
nor U12356 (N_12356,N_11722,N_11966);
or U12357 (N_12357,N_11627,N_11647);
or U12358 (N_12358,N_11972,N_11241);
nor U12359 (N_12359,N_11332,N_11106);
nor U12360 (N_12360,N_11095,N_11044);
xor U12361 (N_12361,N_11019,N_11980);
and U12362 (N_12362,N_11084,N_11648);
nor U12363 (N_12363,N_11641,N_11451);
and U12364 (N_12364,N_11817,N_11495);
or U12365 (N_12365,N_11905,N_11596);
xnor U12366 (N_12366,N_11011,N_11427);
or U12367 (N_12367,N_11130,N_11765);
xnor U12368 (N_12368,N_11922,N_11343);
nor U12369 (N_12369,N_11285,N_11652);
nor U12370 (N_12370,N_11984,N_11138);
and U12371 (N_12371,N_11783,N_11220);
or U12372 (N_12372,N_11818,N_11046);
and U12373 (N_12373,N_11132,N_11796);
nand U12374 (N_12374,N_11414,N_11015);
nor U12375 (N_12375,N_11134,N_11514);
nand U12376 (N_12376,N_11152,N_11341);
xnor U12377 (N_12377,N_11101,N_11274);
and U12378 (N_12378,N_11239,N_11908);
xor U12379 (N_12379,N_11793,N_11735);
nand U12380 (N_12380,N_11282,N_11284);
and U12381 (N_12381,N_11012,N_11771);
nand U12382 (N_12382,N_11822,N_11790);
and U12383 (N_12383,N_11229,N_11075);
nor U12384 (N_12384,N_11528,N_11919);
xnor U12385 (N_12385,N_11116,N_11659);
or U12386 (N_12386,N_11518,N_11838);
nor U12387 (N_12387,N_11008,N_11218);
nor U12388 (N_12388,N_11186,N_11747);
and U12389 (N_12389,N_11795,N_11061);
and U12390 (N_12390,N_11829,N_11110);
or U12391 (N_12391,N_11753,N_11235);
or U12392 (N_12392,N_11409,N_11553);
nand U12393 (N_12393,N_11816,N_11714);
nor U12394 (N_12394,N_11273,N_11297);
nor U12395 (N_12395,N_11850,N_11996);
or U12396 (N_12396,N_11000,N_11082);
nand U12397 (N_12397,N_11473,N_11452);
or U12398 (N_12398,N_11423,N_11577);
and U12399 (N_12399,N_11891,N_11039);
and U12400 (N_12400,N_11365,N_11573);
nor U12401 (N_12401,N_11857,N_11279);
nor U12402 (N_12402,N_11927,N_11774);
and U12403 (N_12403,N_11543,N_11361);
and U12404 (N_12404,N_11951,N_11833);
xor U12405 (N_12405,N_11956,N_11357);
nor U12406 (N_12406,N_11369,N_11718);
nand U12407 (N_12407,N_11782,N_11909);
nor U12408 (N_12408,N_11470,N_11240);
nand U12409 (N_12409,N_11698,N_11043);
and U12410 (N_12410,N_11203,N_11554);
nand U12411 (N_12411,N_11689,N_11227);
or U12412 (N_12412,N_11994,N_11772);
nor U12413 (N_12413,N_11998,N_11208);
and U12414 (N_12414,N_11151,N_11002);
and U12415 (N_12415,N_11604,N_11632);
or U12416 (N_12416,N_11995,N_11404);
nor U12417 (N_12417,N_11581,N_11770);
nand U12418 (N_12418,N_11711,N_11766);
nand U12419 (N_12419,N_11504,N_11918);
nand U12420 (N_12420,N_11367,N_11799);
or U12421 (N_12421,N_11559,N_11695);
or U12422 (N_12422,N_11988,N_11406);
or U12423 (N_12423,N_11090,N_11625);
nand U12424 (N_12424,N_11843,N_11105);
nor U12425 (N_12425,N_11073,N_11362);
nor U12426 (N_12426,N_11805,N_11637);
xor U12427 (N_12427,N_11233,N_11525);
nand U12428 (N_12428,N_11887,N_11209);
xor U12429 (N_12429,N_11053,N_11598);
and U12430 (N_12430,N_11147,N_11824);
nand U12431 (N_12431,N_11871,N_11556);
nand U12432 (N_12432,N_11644,N_11065);
nor U12433 (N_12433,N_11868,N_11035);
and U12434 (N_12434,N_11557,N_11762);
and U12435 (N_12435,N_11072,N_11370);
or U12436 (N_12436,N_11482,N_11172);
nor U12437 (N_12437,N_11802,N_11141);
or U12438 (N_12438,N_11191,N_11261);
and U12439 (N_12439,N_11693,N_11287);
nor U12440 (N_12440,N_11674,N_11611);
nor U12441 (N_12441,N_11149,N_11391);
nor U12442 (N_12442,N_11312,N_11517);
nor U12443 (N_12443,N_11631,N_11302);
xor U12444 (N_12444,N_11347,N_11539);
xor U12445 (N_12445,N_11655,N_11490);
or U12446 (N_12446,N_11493,N_11876);
nand U12447 (N_12447,N_11675,N_11670);
and U12448 (N_12448,N_11778,N_11496);
xor U12449 (N_12449,N_11603,N_11832);
nor U12450 (N_12450,N_11924,N_11779);
or U12451 (N_12451,N_11954,N_11813);
and U12452 (N_12452,N_11531,N_11381);
xor U12453 (N_12453,N_11618,N_11109);
and U12454 (N_12454,N_11301,N_11501);
nor U12455 (N_12455,N_11145,N_11471);
and U12456 (N_12456,N_11508,N_11775);
and U12457 (N_12457,N_11732,N_11538);
or U12458 (N_12458,N_11417,N_11459);
and U12459 (N_12459,N_11991,N_11187);
xnor U12460 (N_12460,N_11855,N_11222);
nand U12461 (N_12461,N_11143,N_11160);
and U12462 (N_12462,N_11845,N_11964);
nand U12463 (N_12463,N_11882,N_11079);
nand U12464 (N_12464,N_11685,N_11507);
and U12465 (N_12465,N_11523,N_11017);
xor U12466 (N_12466,N_11234,N_11662);
and U12467 (N_12467,N_11437,N_11295);
nor U12468 (N_12468,N_11930,N_11001);
xnor U12469 (N_12469,N_11513,N_11091);
nand U12470 (N_12470,N_11619,N_11385);
or U12471 (N_12471,N_11051,N_11594);
and U12472 (N_12472,N_11606,N_11376);
or U12473 (N_12473,N_11198,N_11726);
nand U12474 (N_12474,N_11870,N_11267);
or U12475 (N_12475,N_11335,N_11243);
nand U12476 (N_12476,N_11439,N_11211);
or U12477 (N_12477,N_11703,N_11359);
nand U12478 (N_12478,N_11565,N_11037);
nor U12479 (N_12479,N_11819,N_11636);
xor U12480 (N_12480,N_11926,N_11568);
nor U12481 (N_12481,N_11702,N_11174);
or U12482 (N_12482,N_11873,N_11921);
or U12483 (N_12483,N_11226,N_11108);
nor U12484 (N_12484,N_11806,N_11028);
or U12485 (N_12485,N_11738,N_11533);
and U12486 (N_12486,N_11992,N_11213);
xor U12487 (N_12487,N_11255,N_11973);
nand U12488 (N_12488,N_11435,N_11745);
and U12489 (N_12489,N_11155,N_11123);
nand U12490 (N_12490,N_11231,N_11549);
or U12491 (N_12491,N_11428,N_11524);
nor U12492 (N_12492,N_11440,N_11572);
or U12493 (N_12493,N_11717,N_11571);
or U12494 (N_12494,N_11663,N_11478);
and U12495 (N_12495,N_11074,N_11320);
xnor U12496 (N_12496,N_11884,N_11333);
and U12497 (N_12497,N_11937,N_11055);
nor U12498 (N_12498,N_11024,N_11023);
nand U12499 (N_12499,N_11207,N_11807);
or U12500 (N_12500,N_11693,N_11905);
or U12501 (N_12501,N_11056,N_11142);
and U12502 (N_12502,N_11950,N_11640);
and U12503 (N_12503,N_11383,N_11446);
nand U12504 (N_12504,N_11927,N_11670);
nand U12505 (N_12505,N_11308,N_11237);
and U12506 (N_12506,N_11904,N_11864);
nand U12507 (N_12507,N_11730,N_11299);
nor U12508 (N_12508,N_11171,N_11247);
nor U12509 (N_12509,N_11601,N_11547);
nand U12510 (N_12510,N_11857,N_11496);
nor U12511 (N_12511,N_11918,N_11842);
and U12512 (N_12512,N_11155,N_11160);
xor U12513 (N_12513,N_11955,N_11556);
xnor U12514 (N_12514,N_11467,N_11764);
nor U12515 (N_12515,N_11443,N_11342);
nand U12516 (N_12516,N_11538,N_11845);
nor U12517 (N_12517,N_11118,N_11161);
or U12518 (N_12518,N_11257,N_11692);
and U12519 (N_12519,N_11755,N_11499);
or U12520 (N_12520,N_11068,N_11427);
and U12521 (N_12521,N_11323,N_11454);
nor U12522 (N_12522,N_11544,N_11607);
nand U12523 (N_12523,N_11512,N_11650);
xor U12524 (N_12524,N_11705,N_11147);
xor U12525 (N_12525,N_11498,N_11834);
nor U12526 (N_12526,N_11840,N_11677);
nor U12527 (N_12527,N_11958,N_11251);
or U12528 (N_12528,N_11936,N_11442);
nor U12529 (N_12529,N_11066,N_11001);
nor U12530 (N_12530,N_11600,N_11134);
or U12531 (N_12531,N_11272,N_11418);
nor U12532 (N_12532,N_11556,N_11376);
or U12533 (N_12533,N_11098,N_11995);
nand U12534 (N_12534,N_11604,N_11379);
nand U12535 (N_12535,N_11350,N_11599);
or U12536 (N_12536,N_11935,N_11406);
and U12537 (N_12537,N_11592,N_11548);
and U12538 (N_12538,N_11782,N_11435);
and U12539 (N_12539,N_11187,N_11122);
nand U12540 (N_12540,N_11620,N_11352);
or U12541 (N_12541,N_11811,N_11877);
and U12542 (N_12542,N_11130,N_11850);
or U12543 (N_12543,N_11924,N_11339);
or U12544 (N_12544,N_11554,N_11865);
xnor U12545 (N_12545,N_11426,N_11729);
nor U12546 (N_12546,N_11609,N_11742);
nand U12547 (N_12547,N_11840,N_11855);
nand U12548 (N_12548,N_11340,N_11406);
nor U12549 (N_12549,N_11839,N_11391);
nand U12550 (N_12550,N_11084,N_11398);
nor U12551 (N_12551,N_11073,N_11327);
nand U12552 (N_12552,N_11074,N_11391);
xnor U12553 (N_12553,N_11967,N_11312);
xnor U12554 (N_12554,N_11143,N_11387);
nor U12555 (N_12555,N_11387,N_11734);
nor U12556 (N_12556,N_11105,N_11890);
nor U12557 (N_12557,N_11639,N_11648);
nand U12558 (N_12558,N_11331,N_11030);
nor U12559 (N_12559,N_11521,N_11378);
or U12560 (N_12560,N_11638,N_11839);
nand U12561 (N_12561,N_11324,N_11083);
nand U12562 (N_12562,N_11392,N_11277);
nand U12563 (N_12563,N_11776,N_11528);
nor U12564 (N_12564,N_11598,N_11871);
and U12565 (N_12565,N_11982,N_11425);
nor U12566 (N_12566,N_11395,N_11586);
and U12567 (N_12567,N_11654,N_11518);
and U12568 (N_12568,N_11463,N_11692);
nand U12569 (N_12569,N_11066,N_11493);
or U12570 (N_12570,N_11753,N_11936);
and U12571 (N_12571,N_11448,N_11682);
nand U12572 (N_12572,N_11117,N_11281);
and U12573 (N_12573,N_11189,N_11165);
and U12574 (N_12574,N_11713,N_11678);
and U12575 (N_12575,N_11917,N_11793);
nand U12576 (N_12576,N_11981,N_11634);
or U12577 (N_12577,N_11579,N_11778);
nor U12578 (N_12578,N_11619,N_11883);
and U12579 (N_12579,N_11214,N_11490);
or U12580 (N_12580,N_11050,N_11720);
xor U12581 (N_12581,N_11967,N_11727);
nor U12582 (N_12582,N_11617,N_11548);
and U12583 (N_12583,N_11780,N_11602);
and U12584 (N_12584,N_11512,N_11530);
and U12585 (N_12585,N_11379,N_11278);
nand U12586 (N_12586,N_11058,N_11762);
and U12587 (N_12587,N_11366,N_11225);
nor U12588 (N_12588,N_11521,N_11526);
and U12589 (N_12589,N_11738,N_11791);
nand U12590 (N_12590,N_11653,N_11423);
and U12591 (N_12591,N_11571,N_11995);
or U12592 (N_12592,N_11828,N_11056);
and U12593 (N_12593,N_11814,N_11191);
nand U12594 (N_12594,N_11850,N_11893);
nand U12595 (N_12595,N_11108,N_11737);
or U12596 (N_12596,N_11728,N_11201);
and U12597 (N_12597,N_11804,N_11375);
nor U12598 (N_12598,N_11472,N_11522);
and U12599 (N_12599,N_11762,N_11302);
xnor U12600 (N_12600,N_11742,N_11015);
nor U12601 (N_12601,N_11583,N_11010);
xnor U12602 (N_12602,N_11446,N_11501);
and U12603 (N_12603,N_11792,N_11162);
and U12604 (N_12604,N_11815,N_11694);
and U12605 (N_12605,N_11360,N_11080);
nor U12606 (N_12606,N_11110,N_11649);
nor U12607 (N_12607,N_11244,N_11017);
nand U12608 (N_12608,N_11516,N_11848);
and U12609 (N_12609,N_11822,N_11540);
or U12610 (N_12610,N_11437,N_11157);
nand U12611 (N_12611,N_11987,N_11980);
and U12612 (N_12612,N_11365,N_11510);
xor U12613 (N_12613,N_11788,N_11070);
nor U12614 (N_12614,N_11976,N_11437);
nor U12615 (N_12615,N_11883,N_11204);
nand U12616 (N_12616,N_11295,N_11770);
and U12617 (N_12617,N_11468,N_11008);
xnor U12618 (N_12618,N_11341,N_11211);
and U12619 (N_12619,N_11229,N_11162);
nand U12620 (N_12620,N_11132,N_11475);
nand U12621 (N_12621,N_11068,N_11738);
and U12622 (N_12622,N_11469,N_11633);
or U12623 (N_12623,N_11672,N_11009);
and U12624 (N_12624,N_11012,N_11296);
and U12625 (N_12625,N_11229,N_11855);
nand U12626 (N_12626,N_11792,N_11856);
and U12627 (N_12627,N_11690,N_11442);
or U12628 (N_12628,N_11253,N_11922);
or U12629 (N_12629,N_11608,N_11596);
nor U12630 (N_12630,N_11027,N_11809);
nor U12631 (N_12631,N_11271,N_11658);
xnor U12632 (N_12632,N_11813,N_11659);
and U12633 (N_12633,N_11932,N_11543);
or U12634 (N_12634,N_11194,N_11818);
nor U12635 (N_12635,N_11975,N_11286);
nor U12636 (N_12636,N_11043,N_11300);
and U12637 (N_12637,N_11555,N_11918);
nand U12638 (N_12638,N_11168,N_11071);
and U12639 (N_12639,N_11289,N_11364);
nand U12640 (N_12640,N_11372,N_11505);
xor U12641 (N_12641,N_11648,N_11517);
nor U12642 (N_12642,N_11702,N_11917);
and U12643 (N_12643,N_11400,N_11655);
and U12644 (N_12644,N_11185,N_11234);
and U12645 (N_12645,N_11892,N_11619);
and U12646 (N_12646,N_11604,N_11343);
nor U12647 (N_12647,N_11370,N_11253);
nand U12648 (N_12648,N_11735,N_11398);
and U12649 (N_12649,N_11149,N_11540);
nor U12650 (N_12650,N_11278,N_11812);
and U12651 (N_12651,N_11400,N_11085);
or U12652 (N_12652,N_11138,N_11019);
nor U12653 (N_12653,N_11573,N_11801);
nor U12654 (N_12654,N_11759,N_11965);
nor U12655 (N_12655,N_11683,N_11911);
xnor U12656 (N_12656,N_11986,N_11831);
or U12657 (N_12657,N_11026,N_11387);
or U12658 (N_12658,N_11337,N_11535);
and U12659 (N_12659,N_11616,N_11213);
and U12660 (N_12660,N_11360,N_11131);
xnor U12661 (N_12661,N_11596,N_11355);
or U12662 (N_12662,N_11018,N_11146);
or U12663 (N_12663,N_11735,N_11755);
or U12664 (N_12664,N_11151,N_11157);
and U12665 (N_12665,N_11006,N_11088);
nor U12666 (N_12666,N_11333,N_11578);
and U12667 (N_12667,N_11011,N_11865);
xor U12668 (N_12668,N_11685,N_11340);
or U12669 (N_12669,N_11341,N_11113);
nand U12670 (N_12670,N_11641,N_11397);
nor U12671 (N_12671,N_11829,N_11808);
and U12672 (N_12672,N_11454,N_11107);
nand U12673 (N_12673,N_11133,N_11943);
or U12674 (N_12674,N_11741,N_11598);
and U12675 (N_12675,N_11864,N_11002);
nand U12676 (N_12676,N_11127,N_11337);
nand U12677 (N_12677,N_11570,N_11307);
or U12678 (N_12678,N_11592,N_11468);
and U12679 (N_12679,N_11508,N_11350);
and U12680 (N_12680,N_11576,N_11874);
nor U12681 (N_12681,N_11150,N_11789);
nor U12682 (N_12682,N_11052,N_11397);
and U12683 (N_12683,N_11330,N_11503);
xor U12684 (N_12684,N_11708,N_11955);
or U12685 (N_12685,N_11643,N_11182);
or U12686 (N_12686,N_11092,N_11435);
nor U12687 (N_12687,N_11003,N_11046);
nor U12688 (N_12688,N_11781,N_11542);
or U12689 (N_12689,N_11992,N_11436);
nand U12690 (N_12690,N_11957,N_11096);
and U12691 (N_12691,N_11983,N_11803);
nor U12692 (N_12692,N_11605,N_11656);
or U12693 (N_12693,N_11942,N_11624);
and U12694 (N_12694,N_11051,N_11655);
and U12695 (N_12695,N_11314,N_11918);
and U12696 (N_12696,N_11056,N_11351);
xor U12697 (N_12697,N_11913,N_11797);
xor U12698 (N_12698,N_11364,N_11757);
or U12699 (N_12699,N_11426,N_11476);
nand U12700 (N_12700,N_11338,N_11050);
xor U12701 (N_12701,N_11572,N_11725);
nand U12702 (N_12702,N_11194,N_11877);
nand U12703 (N_12703,N_11690,N_11609);
xor U12704 (N_12704,N_11822,N_11171);
and U12705 (N_12705,N_11177,N_11902);
nand U12706 (N_12706,N_11148,N_11791);
xnor U12707 (N_12707,N_11589,N_11021);
and U12708 (N_12708,N_11774,N_11237);
nand U12709 (N_12709,N_11873,N_11832);
nor U12710 (N_12710,N_11837,N_11431);
xnor U12711 (N_12711,N_11180,N_11225);
nand U12712 (N_12712,N_11383,N_11933);
nor U12713 (N_12713,N_11199,N_11804);
nor U12714 (N_12714,N_11554,N_11984);
nand U12715 (N_12715,N_11258,N_11083);
nand U12716 (N_12716,N_11797,N_11945);
or U12717 (N_12717,N_11207,N_11330);
or U12718 (N_12718,N_11503,N_11022);
and U12719 (N_12719,N_11906,N_11136);
nand U12720 (N_12720,N_11141,N_11872);
nor U12721 (N_12721,N_11750,N_11025);
and U12722 (N_12722,N_11524,N_11376);
nand U12723 (N_12723,N_11672,N_11799);
or U12724 (N_12724,N_11566,N_11095);
nand U12725 (N_12725,N_11355,N_11288);
or U12726 (N_12726,N_11922,N_11994);
nor U12727 (N_12727,N_11723,N_11880);
or U12728 (N_12728,N_11988,N_11601);
nor U12729 (N_12729,N_11742,N_11645);
and U12730 (N_12730,N_11952,N_11279);
nand U12731 (N_12731,N_11792,N_11564);
or U12732 (N_12732,N_11908,N_11464);
nor U12733 (N_12733,N_11440,N_11002);
xor U12734 (N_12734,N_11706,N_11104);
nor U12735 (N_12735,N_11404,N_11151);
nand U12736 (N_12736,N_11232,N_11151);
or U12737 (N_12737,N_11931,N_11235);
or U12738 (N_12738,N_11208,N_11715);
and U12739 (N_12739,N_11923,N_11328);
and U12740 (N_12740,N_11575,N_11241);
and U12741 (N_12741,N_11158,N_11124);
and U12742 (N_12742,N_11943,N_11649);
xnor U12743 (N_12743,N_11147,N_11917);
and U12744 (N_12744,N_11431,N_11085);
nand U12745 (N_12745,N_11605,N_11007);
and U12746 (N_12746,N_11634,N_11553);
and U12747 (N_12747,N_11387,N_11382);
nor U12748 (N_12748,N_11738,N_11313);
or U12749 (N_12749,N_11753,N_11699);
nand U12750 (N_12750,N_11928,N_11964);
xor U12751 (N_12751,N_11593,N_11653);
and U12752 (N_12752,N_11890,N_11704);
or U12753 (N_12753,N_11031,N_11634);
or U12754 (N_12754,N_11960,N_11540);
or U12755 (N_12755,N_11616,N_11433);
nor U12756 (N_12756,N_11616,N_11400);
nand U12757 (N_12757,N_11397,N_11007);
nand U12758 (N_12758,N_11386,N_11567);
xnor U12759 (N_12759,N_11565,N_11345);
nor U12760 (N_12760,N_11931,N_11677);
and U12761 (N_12761,N_11993,N_11553);
nor U12762 (N_12762,N_11248,N_11540);
or U12763 (N_12763,N_11834,N_11049);
or U12764 (N_12764,N_11255,N_11367);
and U12765 (N_12765,N_11043,N_11847);
nor U12766 (N_12766,N_11502,N_11188);
or U12767 (N_12767,N_11438,N_11733);
nor U12768 (N_12768,N_11603,N_11403);
and U12769 (N_12769,N_11181,N_11991);
and U12770 (N_12770,N_11700,N_11703);
and U12771 (N_12771,N_11350,N_11471);
nand U12772 (N_12772,N_11268,N_11537);
xor U12773 (N_12773,N_11373,N_11370);
and U12774 (N_12774,N_11681,N_11368);
nor U12775 (N_12775,N_11698,N_11152);
and U12776 (N_12776,N_11250,N_11304);
and U12777 (N_12777,N_11177,N_11951);
or U12778 (N_12778,N_11760,N_11626);
xnor U12779 (N_12779,N_11127,N_11880);
and U12780 (N_12780,N_11248,N_11024);
and U12781 (N_12781,N_11918,N_11259);
or U12782 (N_12782,N_11587,N_11648);
nor U12783 (N_12783,N_11471,N_11814);
nor U12784 (N_12784,N_11942,N_11881);
nor U12785 (N_12785,N_11125,N_11688);
or U12786 (N_12786,N_11325,N_11512);
or U12787 (N_12787,N_11508,N_11910);
nor U12788 (N_12788,N_11772,N_11517);
nor U12789 (N_12789,N_11597,N_11621);
nor U12790 (N_12790,N_11709,N_11112);
nand U12791 (N_12791,N_11963,N_11786);
nand U12792 (N_12792,N_11436,N_11061);
nand U12793 (N_12793,N_11648,N_11130);
and U12794 (N_12794,N_11353,N_11010);
or U12795 (N_12795,N_11048,N_11410);
nand U12796 (N_12796,N_11816,N_11121);
or U12797 (N_12797,N_11070,N_11646);
and U12798 (N_12798,N_11502,N_11141);
xor U12799 (N_12799,N_11925,N_11871);
nor U12800 (N_12800,N_11541,N_11424);
nor U12801 (N_12801,N_11123,N_11269);
nor U12802 (N_12802,N_11134,N_11666);
or U12803 (N_12803,N_11088,N_11939);
nor U12804 (N_12804,N_11380,N_11658);
nand U12805 (N_12805,N_11197,N_11199);
or U12806 (N_12806,N_11591,N_11540);
and U12807 (N_12807,N_11898,N_11187);
nor U12808 (N_12808,N_11972,N_11585);
nand U12809 (N_12809,N_11474,N_11253);
nand U12810 (N_12810,N_11093,N_11372);
nand U12811 (N_12811,N_11063,N_11766);
nand U12812 (N_12812,N_11872,N_11042);
nor U12813 (N_12813,N_11162,N_11819);
nand U12814 (N_12814,N_11985,N_11499);
or U12815 (N_12815,N_11219,N_11651);
and U12816 (N_12816,N_11239,N_11326);
nand U12817 (N_12817,N_11964,N_11654);
nor U12818 (N_12818,N_11279,N_11699);
and U12819 (N_12819,N_11064,N_11443);
and U12820 (N_12820,N_11975,N_11572);
nor U12821 (N_12821,N_11313,N_11156);
nor U12822 (N_12822,N_11786,N_11675);
nor U12823 (N_12823,N_11559,N_11086);
or U12824 (N_12824,N_11402,N_11789);
nor U12825 (N_12825,N_11264,N_11551);
or U12826 (N_12826,N_11387,N_11140);
and U12827 (N_12827,N_11320,N_11468);
and U12828 (N_12828,N_11747,N_11229);
and U12829 (N_12829,N_11042,N_11114);
or U12830 (N_12830,N_11806,N_11920);
nand U12831 (N_12831,N_11369,N_11734);
and U12832 (N_12832,N_11591,N_11324);
or U12833 (N_12833,N_11281,N_11820);
and U12834 (N_12834,N_11927,N_11370);
nand U12835 (N_12835,N_11098,N_11629);
and U12836 (N_12836,N_11314,N_11602);
nand U12837 (N_12837,N_11543,N_11822);
nand U12838 (N_12838,N_11132,N_11713);
and U12839 (N_12839,N_11909,N_11225);
nand U12840 (N_12840,N_11241,N_11155);
nor U12841 (N_12841,N_11631,N_11119);
or U12842 (N_12842,N_11508,N_11271);
or U12843 (N_12843,N_11798,N_11628);
or U12844 (N_12844,N_11093,N_11825);
nor U12845 (N_12845,N_11411,N_11170);
xnor U12846 (N_12846,N_11263,N_11208);
nor U12847 (N_12847,N_11042,N_11600);
nor U12848 (N_12848,N_11363,N_11542);
or U12849 (N_12849,N_11780,N_11352);
or U12850 (N_12850,N_11962,N_11841);
and U12851 (N_12851,N_11062,N_11208);
nand U12852 (N_12852,N_11521,N_11208);
or U12853 (N_12853,N_11965,N_11423);
and U12854 (N_12854,N_11567,N_11857);
xor U12855 (N_12855,N_11369,N_11110);
nor U12856 (N_12856,N_11082,N_11133);
and U12857 (N_12857,N_11073,N_11274);
nand U12858 (N_12858,N_11152,N_11435);
or U12859 (N_12859,N_11641,N_11027);
or U12860 (N_12860,N_11780,N_11099);
nand U12861 (N_12861,N_11005,N_11855);
nor U12862 (N_12862,N_11187,N_11315);
nor U12863 (N_12863,N_11562,N_11334);
and U12864 (N_12864,N_11657,N_11525);
xnor U12865 (N_12865,N_11379,N_11386);
nand U12866 (N_12866,N_11755,N_11078);
and U12867 (N_12867,N_11358,N_11946);
or U12868 (N_12868,N_11638,N_11097);
nand U12869 (N_12869,N_11931,N_11357);
nand U12870 (N_12870,N_11183,N_11741);
or U12871 (N_12871,N_11632,N_11935);
nand U12872 (N_12872,N_11763,N_11130);
or U12873 (N_12873,N_11197,N_11843);
and U12874 (N_12874,N_11951,N_11334);
or U12875 (N_12875,N_11564,N_11981);
nor U12876 (N_12876,N_11078,N_11179);
nor U12877 (N_12877,N_11052,N_11040);
nor U12878 (N_12878,N_11532,N_11160);
and U12879 (N_12879,N_11409,N_11453);
nand U12880 (N_12880,N_11757,N_11634);
and U12881 (N_12881,N_11001,N_11087);
xnor U12882 (N_12882,N_11933,N_11800);
nor U12883 (N_12883,N_11219,N_11088);
and U12884 (N_12884,N_11620,N_11174);
nor U12885 (N_12885,N_11548,N_11195);
nand U12886 (N_12886,N_11888,N_11203);
or U12887 (N_12887,N_11364,N_11575);
or U12888 (N_12888,N_11655,N_11478);
or U12889 (N_12889,N_11707,N_11493);
nor U12890 (N_12890,N_11044,N_11567);
nor U12891 (N_12891,N_11925,N_11348);
and U12892 (N_12892,N_11184,N_11746);
nand U12893 (N_12893,N_11433,N_11404);
nand U12894 (N_12894,N_11191,N_11914);
nor U12895 (N_12895,N_11604,N_11964);
xor U12896 (N_12896,N_11455,N_11909);
nor U12897 (N_12897,N_11813,N_11838);
or U12898 (N_12898,N_11049,N_11982);
and U12899 (N_12899,N_11013,N_11415);
nand U12900 (N_12900,N_11836,N_11570);
or U12901 (N_12901,N_11561,N_11696);
and U12902 (N_12902,N_11208,N_11829);
nor U12903 (N_12903,N_11989,N_11183);
or U12904 (N_12904,N_11579,N_11809);
or U12905 (N_12905,N_11744,N_11332);
and U12906 (N_12906,N_11665,N_11792);
and U12907 (N_12907,N_11404,N_11999);
nor U12908 (N_12908,N_11967,N_11594);
nand U12909 (N_12909,N_11401,N_11358);
and U12910 (N_12910,N_11831,N_11653);
and U12911 (N_12911,N_11686,N_11806);
or U12912 (N_12912,N_11376,N_11073);
nor U12913 (N_12913,N_11468,N_11309);
nand U12914 (N_12914,N_11415,N_11829);
xor U12915 (N_12915,N_11291,N_11458);
nand U12916 (N_12916,N_11676,N_11375);
or U12917 (N_12917,N_11702,N_11175);
nor U12918 (N_12918,N_11907,N_11825);
xor U12919 (N_12919,N_11901,N_11572);
nor U12920 (N_12920,N_11893,N_11515);
and U12921 (N_12921,N_11099,N_11899);
and U12922 (N_12922,N_11246,N_11101);
or U12923 (N_12923,N_11970,N_11576);
xnor U12924 (N_12924,N_11415,N_11058);
nand U12925 (N_12925,N_11327,N_11297);
nand U12926 (N_12926,N_11375,N_11946);
nor U12927 (N_12927,N_11266,N_11834);
and U12928 (N_12928,N_11766,N_11911);
nand U12929 (N_12929,N_11203,N_11279);
xor U12930 (N_12930,N_11511,N_11487);
nor U12931 (N_12931,N_11088,N_11119);
xor U12932 (N_12932,N_11517,N_11940);
nand U12933 (N_12933,N_11842,N_11802);
xor U12934 (N_12934,N_11891,N_11562);
nand U12935 (N_12935,N_11125,N_11600);
and U12936 (N_12936,N_11800,N_11217);
xnor U12937 (N_12937,N_11142,N_11568);
nor U12938 (N_12938,N_11959,N_11384);
nor U12939 (N_12939,N_11079,N_11155);
xor U12940 (N_12940,N_11128,N_11767);
and U12941 (N_12941,N_11235,N_11124);
nor U12942 (N_12942,N_11069,N_11006);
nand U12943 (N_12943,N_11271,N_11679);
nor U12944 (N_12944,N_11818,N_11768);
or U12945 (N_12945,N_11172,N_11168);
and U12946 (N_12946,N_11392,N_11266);
and U12947 (N_12947,N_11888,N_11991);
nand U12948 (N_12948,N_11328,N_11850);
nor U12949 (N_12949,N_11025,N_11318);
nand U12950 (N_12950,N_11043,N_11271);
nor U12951 (N_12951,N_11681,N_11523);
nor U12952 (N_12952,N_11942,N_11665);
nand U12953 (N_12953,N_11957,N_11423);
nand U12954 (N_12954,N_11532,N_11839);
or U12955 (N_12955,N_11610,N_11464);
nand U12956 (N_12956,N_11678,N_11985);
and U12957 (N_12957,N_11293,N_11243);
and U12958 (N_12958,N_11540,N_11967);
or U12959 (N_12959,N_11616,N_11898);
nand U12960 (N_12960,N_11786,N_11898);
xor U12961 (N_12961,N_11249,N_11644);
and U12962 (N_12962,N_11961,N_11001);
nor U12963 (N_12963,N_11614,N_11731);
nand U12964 (N_12964,N_11893,N_11391);
or U12965 (N_12965,N_11680,N_11356);
nor U12966 (N_12966,N_11488,N_11167);
or U12967 (N_12967,N_11202,N_11767);
or U12968 (N_12968,N_11628,N_11142);
nand U12969 (N_12969,N_11775,N_11774);
nor U12970 (N_12970,N_11820,N_11105);
or U12971 (N_12971,N_11761,N_11049);
and U12972 (N_12972,N_11216,N_11599);
xnor U12973 (N_12973,N_11077,N_11982);
or U12974 (N_12974,N_11294,N_11420);
nand U12975 (N_12975,N_11497,N_11416);
nand U12976 (N_12976,N_11784,N_11442);
and U12977 (N_12977,N_11474,N_11667);
nor U12978 (N_12978,N_11675,N_11688);
and U12979 (N_12979,N_11877,N_11775);
xor U12980 (N_12980,N_11680,N_11531);
nor U12981 (N_12981,N_11267,N_11669);
nand U12982 (N_12982,N_11803,N_11788);
or U12983 (N_12983,N_11768,N_11986);
nor U12984 (N_12984,N_11753,N_11966);
and U12985 (N_12985,N_11229,N_11619);
nand U12986 (N_12986,N_11264,N_11624);
or U12987 (N_12987,N_11199,N_11932);
or U12988 (N_12988,N_11985,N_11986);
or U12989 (N_12989,N_11054,N_11216);
nor U12990 (N_12990,N_11706,N_11147);
nand U12991 (N_12991,N_11710,N_11640);
and U12992 (N_12992,N_11658,N_11871);
and U12993 (N_12993,N_11359,N_11184);
and U12994 (N_12994,N_11020,N_11688);
nand U12995 (N_12995,N_11824,N_11244);
nor U12996 (N_12996,N_11057,N_11926);
nor U12997 (N_12997,N_11028,N_11411);
xor U12998 (N_12998,N_11753,N_11346);
xor U12999 (N_12999,N_11072,N_11060);
nor U13000 (N_13000,N_12212,N_12464);
or U13001 (N_13001,N_12003,N_12164);
and U13002 (N_13002,N_12847,N_12161);
nand U13003 (N_13003,N_12248,N_12416);
or U13004 (N_13004,N_12724,N_12288);
xnor U13005 (N_13005,N_12691,N_12150);
nand U13006 (N_13006,N_12127,N_12110);
xnor U13007 (N_13007,N_12276,N_12129);
or U13008 (N_13008,N_12382,N_12094);
nand U13009 (N_13009,N_12014,N_12917);
and U13010 (N_13010,N_12759,N_12629);
or U13011 (N_13011,N_12045,N_12189);
nand U13012 (N_13012,N_12099,N_12031);
xnor U13013 (N_13013,N_12865,N_12067);
nand U13014 (N_13014,N_12651,N_12595);
nand U13015 (N_13015,N_12566,N_12412);
and U13016 (N_13016,N_12694,N_12295);
nand U13017 (N_13017,N_12763,N_12206);
or U13018 (N_13018,N_12444,N_12082);
or U13019 (N_13019,N_12916,N_12034);
and U13020 (N_13020,N_12618,N_12955);
nand U13021 (N_13021,N_12885,N_12365);
xnor U13022 (N_13022,N_12591,N_12088);
nand U13023 (N_13023,N_12216,N_12572);
nand U13024 (N_13024,N_12434,N_12509);
nand U13025 (N_13025,N_12390,N_12748);
nor U13026 (N_13026,N_12892,N_12035);
or U13027 (N_13027,N_12816,N_12745);
and U13028 (N_13028,N_12617,N_12689);
and U13029 (N_13029,N_12881,N_12484);
xor U13030 (N_13030,N_12645,N_12784);
and U13031 (N_13031,N_12404,N_12648);
or U13032 (N_13032,N_12729,N_12485);
or U13033 (N_13033,N_12450,N_12820);
and U13034 (N_13034,N_12793,N_12176);
xor U13035 (N_13035,N_12265,N_12534);
xor U13036 (N_13036,N_12733,N_12605);
nand U13037 (N_13037,N_12103,N_12918);
nand U13038 (N_13038,N_12050,N_12627);
nor U13039 (N_13039,N_12397,N_12941);
and U13040 (N_13040,N_12153,N_12079);
nand U13041 (N_13041,N_12077,N_12215);
and U13042 (N_13042,N_12321,N_12654);
or U13043 (N_13043,N_12155,N_12965);
or U13044 (N_13044,N_12315,N_12228);
nand U13045 (N_13045,N_12306,N_12561);
nor U13046 (N_13046,N_12564,N_12010);
nand U13047 (N_13047,N_12719,N_12197);
nor U13048 (N_13048,N_12953,N_12507);
nor U13049 (N_13049,N_12323,N_12089);
or U13050 (N_13050,N_12353,N_12779);
and U13051 (N_13051,N_12049,N_12500);
or U13052 (N_13052,N_12951,N_12557);
nor U13053 (N_13053,N_12300,N_12301);
and U13054 (N_13054,N_12979,N_12396);
nor U13055 (N_13055,N_12247,N_12123);
and U13056 (N_13056,N_12244,N_12961);
and U13057 (N_13057,N_12897,N_12125);
and U13058 (N_13058,N_12086,N_12144);
nor U13059 (N_13059,N_12170,N_12836);
nand U13060 (N_13060,N_12932,N_12738);
or U13061 (N_13061,N_12819,N_12436);
or U13062 (N_13062,N_12923,N_12322);
nor U13063 (N_13063,N_12347,N_12196);
nand U13064 (N_13064,N_12266,N_12976);
and U13065 (N_13065,N_12269,N_12672);
or U13066 (N_13066,N_12807,N_12024);
xnor U13067 (N_13067,N_12439,N_12281);
and U13068 (N_13068,N_12044,N_12324);
and U13069 (N_13069,N_12767,N_12180);
nand U13070 (N_13070,N_12379,N_12147);
nand U13071 (N_13071,N_12364,N_12590);
xor U13072 (N_13072,N_12194,N_12367);
or U13073 (N_13073,N_12752,N_12320);
and U13074 (N_13074,N_12853,N_12051);
nor U13075 (N_13075,N_12751,N_12895);
nor U13076 (N_13076,N_12805,N_12638);
nor U13077 (N_13077,N_12652,N_12234);
nand U13078 (N_13078,N_12934,N_12744);
and U13079 (N_13079,N_12523,N_12945);
and U13080 (N_13080,N_12204,N_12665);
and U13081 (N_13081,N_12866,N_12357);
xor U13082 (N_13082,N_12452,N_12690);
nor U13083 (N_13083,N_12877,N_12825);
xnor U13084 (N_13084,N_12880,N_12311);
or U13085 (N_13085,N_12407,N_12226);
and U13086 (N_13086,N_12019,N_12747);
or U13087 (N_13087,N_12810,N_12774);
nor U13088 (N_13088,N_12175,N_12644);
nor U13089 (N_13089,N_12373,N_12122);
and U13090 (N_13090,N_12526,N_12162);
and U13091 (N_13091,N_12947,N_12430);
nand U13092 (N_13092,N_12016,N_12984);
and U13093 (N_13093,N_12702,N_12706);
nor U13094 (N_13094,N_12701,N_12737);
or U13095 (N_13095,N_12531,N_12418);
nand U13096 (N_13096,N_12705,N_12355);
or U13097 (N_13097,N_12275,N_12427);
or U13098 (N_13098,N_12026,N_12878);
nor U13099 (N_13099,N_12402,N_12603);
nor U13100 (N_13100,N_12578,N_12312);
nand U13101 (N_13101,N_12548,N_12620);
and U13102 (N_13102,N_12375,N_12842);
nor U13103 (N_13103,N_12156,N_12078);
nand U13104 (N_13104,N_12195,N_12870);
or U13105 (N_13105,N_12616,N_12358);
nor U13106 (N_13106,N_12183,N_12341);
or U13107 (N_13107,N_12399,N_12208);
and U13108 (N_13108,N_12114,N_12891);
and U13109 (N_13109,N_12679,N_12827);
nor U13110 (N_13110,N_12915,N_12458);
xnor U13111 (N_13111,N_12210,N_12850);
or U13112 (N_13112,N_12108,N_12568);
nor U13113 (N_13113,N_12995,N_12801);
or U13114 (N_13114,N_12036,N_12506);
nor U13115 (N_13115,N_12495,N_12787);
nor U13116 (N_13116,N_12325,N_12861);
nor U13117 (N_13117,N_12547,N_12586);
or U13118 (N_13118,N_12597,N_12795);
nor U13119 (N_13119,N_12811,N_12929);
nand U13120 (N_13120,N_12789,N_12414);
nor U13121 (N_13121,N_12277,N_12567);
nor U13122 (N_13122,N_12346,N_12800);
nand U13123 (N_13123,N_12360,N_12455);
and U13124 (N_13124,N_12240,N_12178);
and U13125 (N_13125,N_12351,N_12809);
nor U13126 (N_13126,N_12968,N_12101);
and U13127 (N_13127,N_12055,N_12482);
or U13128 (N_13128,N_12303,N_12710);
nand U13129 (N_13129,N_12971,N_12200);
nand U13130 (N_13130,N_12607,N_12140);
nand U13131 (N_13131,N_12755,N_12545);
and U13132 (N_13132,N_12042,N_12978);
xnor U13133 (N_13133,N_12714,N_12284);
and U13134 (N_13134,N_12054,N_12948);
nor U13135 (N_13135,N_12474,N_12229);
nand U13136 (N_13136,N_12829,N_12361);
and U13137 (N_13137,N_12736,N_12686);
nor U13138 (N_13138,N_12757,N_12529);
or U13139 (N_13139,N_12307,N_12011);
xnor U13140 (N_13140,N_12201,N_12581);
xnor U13141 (N_13141,N_12711,N_12770);
nor U13142 (N_13142,N_12903,N_12329);
nand U13143 (N_13143,N_12148,N_12394);
and U13144 (N_13144,N_12184,N_12996);
nand U13145 (N_13145,N_12777,N_12245);
and U13146 (N_13146,N_12343,N_12693);
or U13147 (N_13147,N_12558,N_12420);
xnor U13148 (N_13148,N_12730,N_12330);
nor U13149 (N_13149,N_12685,N_12658);
and U13150 (N_13150,N_12604,N_12510);
nand U13151 (N_13151,N_12635,N_12271);
or U13152 (N_13152,N_12931,N_12802);
nor U13153 (N_13153,N_12803,N_12152);
or U13154 (N_13154,N_12637,N_12483);
nand U13155 (N_13155,N_12223,N_12182);
nor U13156 (N_13156,N_12517,N_12623);
xor U13157 (N_13157,N_12264,N_12682);
nor U13158 (N_13158,N_12142,N_12203);
xnor U13159 (N_13159,N_12831,N_12328);
or U13160 (N_13160,N_12562,N_12130);
xnor U13161 (N_13161,N_12709,N_12911);
or U13162 (N_13162,N_12259,N_12632);
nor U13163 (N_13163,N_12422,N_12514);
nor U13164 (N_13164,N_12678,N_12594);
xor U13165 (N_13165,N_12843,N_12554);
nand U13166 (N_13166,N_12703,N_12429);
or U13167 (N_13167,N_12273,N_12666);
or U13168 (N_13168,N_12863,N_12832);
and U13169 (N_13169,N_12097,N_12712);
xnor U13170 (N_13170,N_12128,N_12085);
and U13171 (N_13171,N_12272,N_12267);
or U13172 (N_13172,N_12304,N_12502);
and U13173 (N_13173,N_12279,N_12884);
and U13174 (N_13174,N_12553,N_12254);
nand U13175 (N_13175,N_12889,N_12765);
and U13176 (N_13176,N_12888,N_12435);
or U13177 (N_13177,N_12879,N_12070);
and U13178 (N_13178,N_12909,N_12726);
or U13179 (N_13179,N_12600,N_12263);
xnor U13180 (N_13180,N_12068,N_12782);
nand U13181 (N_13181,N_12470,N_12585);
or U13182 (N_13182,N_12938,N_12989);
and U13183 (N_13183,N_12928,N_12518);
nor U13184 (N_13184,N_12052,N_12583);
or U13185 (N_13185,N_12749,N_12501);
and U13186 (N_13186,N_12106,N_12023);
or U13187 (N_13187,N_12519,N_12926);
and U13188 (N_13188,N_12785,N_12135);
or U13189 (N_13189,N_12187,N_12352);
xor U13190 (N_13190,N_12662,N_12389);
nand U13191 (N_13191,N_12882,N_12258);
nand U13192 (N_13192,N_12890,N_12063);
or U13193 (N_13193,N_12366,N_12958);
or U13194 (N_13194,N_12655,N_12924);
and U13195 (N_13195,N_12664,N_12920);
and U13196 (N_13196,N_12370,N_12463);
xnor U13197 (N_13197,N_12243,N_12823);
nand U13198 (N_13198,N_12118,N_12117);
xnor U13199 (N_13199,N_12762,N_12488);
xor U13200 (N_13200,N_12235,N_12348);
or U13201 (N_13201,N_12575,N_12188);
or U13202 (N_13202,N_12812,N_12688);
and U13203 (N_13203,N_12166,N_12145);
nor U13204 (N_13204,N_12919,N_12029);
or U13205 (N_13205,N_12410,N_12419);
or U13206 (N_13206,N_12530,N_12649);
or U13207 (N_13207,N_12899,N_12602);
nand U13208 (N_13208,N_12119,N_12199);
or U13209 (N_13209,N_12239,N_12999);
xnor U13210 (N_13210,N_12098,N_12126);
or U13211 (N_13211,N_12698,N_12233);
nor U13212 (N_13212,N_12991,N_12080);
and U13213 (N_13213,N_12053,N_12760);
or U13214 (N_13214,N_12425,N_12563);
and U13215 (N_13215,N_12746,N_12480);
nor U13216 (N_13216,N_12696,N_12565);
nand U13217 (N_13217,N_12471,N_12516);
nand U13218 (N_13218,N_12695,N_12735);
and U13219 (N_13219,N_12476,N_12596);
or U13220 (N_13220,N_12992,N_12076);
nand U13221 (N_13221,N_12786,N_12675);
or U13222 (N_13222,N_12537,N_12621);
nor U13223 (N_13223,N_12398,N_12535);
nor U13224 (N_13224,N_12985,N_12741);
or U13225 (N_13225,N_12963,N_12496);
and U13226 (N_13226,N_12960,N_12845);
nand U13227 (N_13227,N_12852,N_12552);
and U13228 (N_13228,N_12967,N_12012);
or U13229 (N_13229,N_12167,N_12336);
and U13230 (N_13230,N_12608,N_12388);
and U13231 (N_13231,N_12643,N_12798);
nor U13232 (N_13232,N_12487,N_12190);
nor U13233 (N_13233,N_12384,N_12224);
and U13234 (N_13234,N_12393,N_12408);
nor U13235 (N_13235,N_12653,N_12704);
or U13236 (N_13236,N_12472,N_12661);
nand U13237 (N_13237,N_12137,N_12227);
nor U13238 (N_13238,N_12460,N_12149);
or U13239 (N_13239,N_12113,N_12975);
xnor U13240 (N_13240,N_12350,N_12952);
and U13241 (N_13241,N_12783,N_12622);
or U13242 (N_13242,N_12270,N_12708);
nor U13243 (N_13243,N_12940,N_12002);
and U13244 (N_13244,N_12478,N_12815);
xnor U13245 (N_13245,N_12446,N_12107);
or U13246 (N_13246,N_12297,N_12083);
nand U13247 (N_13247,N_12718,N_12773);
nand U13248 (N_13248,N_12673,N_12431);
or U13249 (N_13249,N_12788,N_12132);
or U13250 (N_13250,N_12739,N_12072);
and U13251 (N_13251,N_12218,N_12808);
nor U13252 (N_13252,N_12292,N_12957);
xor U13253 (N_13253,N_12423,N_12758);
nor U13254 (N_13254,N_12409,N_12354);
and U13255 (N_13255,N_12493,N_12225);
nor U13256 (N_13256,N_12833,N_12910);
and U13257 (N_13257,N_12372,N_12776);
nor U13258 (N_13258,N_12761,N_12536);
or U13259 (N_13259,N_12074,N_12862);
and U13260 (N_13260,N_12383,N_12794);
or U13261 (N_13261,N_12732,N_12867);
nand U13262 (N_13262,N_12274,N_12447);
or U13263 (N_13263,N_12615,N_12544);
and U13264 (N_13264,N_12075,N_12656);
or U13265 (N_13265,N_12921,N_12657);
nand U13266 (N_13266,N_12205,N_12209);
or U13267 (N_13267,N_12251,N_12896);
nand U13268 (N_13268,N_12720,N_12646);
nand U13269 (N_13269,N_12944,N_12707);
nor U13270 (N_13270,N_12143,N_12287);
and U13271 (N_13271,N_12174,N_12134);
nand U13272 (N_13272,N_12433,N_12018);
nand U13273 (N_13273,N_12935,N_12371);
and U13274 (N_13274,N_12573,N_12278);
and U13275 (N_13275,N_12421,N_12824);
and U13276 (N_13276,N_12231,N_12754);
nor U13277 (N_13277,N_12477,N_12731);
or U13278 (N_13278,N_12289,N_12387);
xor U13279 (N_13279,N_12830,N_12157);
nor U13280 (N_13280,N_12222,N_12663);
or U13281 (N_13281,N_12821,N_12778);
nand U13282 (N_13282,N_12990,N_12977);
xor U13283 (N_13283,N_12319,N_12533);
nand U13284 (N_13284,N_12525,N_12559);
nand U13285 (N_13285,N_12415,N_12660);
or U13286 (N_13286,N_12873,N_12907);
nand U13287 (N_13287,N_12959,N_12112);
nor U13288 (N_13288,N_12504,N_12327);
nand U13289 (N_13289,N_12219,N_12268);
nor U13290 (N_13290,N_12792,N_12840);
xnor U13291 (N_13291,N_12441,N_12939);
xor U13292 (N_13292,N_12013,N_12066);
and U13293 (N_13293,N_12043,N_12344);
or U13294 (N_13294,N_12887,N_12207);
nand U13295 (N_13295,N_12855,N_12671);
nand U13296 (N_13296,N_12473,N_12185);
nand U13297 (N_13297,N_12956,N_12291);
or U13298 (N_13298,N_12633,N_12230);
xor U13299 (N_13299,N_12069,N_12532);
nand U13300 (N_13300,N_12027,N_12522);
nor U13301 (N_13301,N_12362,N_12417);
or U13302 (N_13302,N_12456,N_12193);
nor U13303 (N_13303,N_12625,N_12858);
nand U13304 (N_13304,N_12093,N_12599);
and U13305 (N_13305,N_12309,N_12937);
or U13306 (N_13306,N_12440,N_12214);
and U13307 (N_13307,N_12902,N_12988);
nand U13308 (N_13308,N_12022,N_12674);
xnor U13309 (N_13309,N_12339,N_12490);
or U13310 (N_13310,N_12636,N_12047);
nor U13311 (N_13311,N_12974,N_12670);
and U13312 (N_13312,N_12550,N_12624);
or U13313 (N_13313,N_12111,N_12771);
nor U13314 (N_13314,N_12151,N_12058);
and U13315 (N_13315,N_12717,N_12403);
or U13316 (N_13316,N_12038,N_12453);
nand U13317 (N_13317,N_12298,N_12057);
nor U13318 (N_13318,N_12860,N_12121);
nand U13319 (N_13319,N_12381,N_12001);
nand U13320 (N_13320,N_12095,N_12310);
xor U13321 (N_13321,N_12246,N_12030);
nand U13322 (N_13322,N_12818,N_12173);
or U13323 (N_13323,N_12462,N_12822);
nor U13324 (N_13324,N_12236,N_12202);
nand U13325 (N_13325,N_12017,N_12192);
nand U13326 (N_13326,N_12528,N_12543);
or U13327 (N_13327,N_12768,N_12280);
and U13328 (N_13328,N_12073,N_12437);
nand U13329 (N_13329,N_12377,N_12349);
nand U13330 (N_13330,N_12834,N_12972);
nand U13331 (N_13331,N_12828,N_12560);
or U13332 (N_13332,N_12032,N_12503);
nor U13333 (N_13333,N_12131,N_12936);
and U13334 (N_13334,N_12198,N_12750);
or U13335 (N_13335,N_12449,N_12481);
nor U13336 (N_13336,N_12715,N_12020);
nand U13337 (N_13337,N_12308,N_12725);
nor U13338 (N_13338,N_12631,N_12242);
or U13339 (N_13339,N_12359,N_12466);
nor U13340 (N_13340,N_12723,N_12634);
or U13341 (N_13341,N_12687,N_12136);
xnor U13342 (N_13342,N_12606,N_12846);
nor U13343 (N_13343,N_12962,N_12286);
nor U13344 (N_13344,N_12090,N_12540);
nand U13345 (N_13345,N_12598,N_12314);
nand U13346 (N_13346,N_12133,N_12716);
nor U13347 (N_13347,N_12479,N_12028);
and U13348 (N_13348,N_12511,N_12241);
or U13349 (N_13349,N_12171,N_12973);
nand U13350 (N_13350,N_12041,N_12555);
nor U13351 (N_13351,N_12849,N_12549);
nor U13352 (N_13352,N_12091,N_12626);
nor U13353 (N_13353,N_12262,N_12994);
nor U13354 (N_13354,N_12611,N_12639);
nor U13355 (N_13355,N_12697,N_12141);
and U13356 (N_13356,N_12592,N_12342);
nor U13357 (N_13357,N_12508,N_12740);
and U13358 (N_13358,N_12317,N_12912);
nand U13359 (N_13359,N_12443,N_12061);
nand U13360 (N_13360,N_12868,N_12220);
nand U13361 (N_13361,N_12837,N_12261);
nand U13362 (N_13362,N_12587,N_12908);
nand U13363 (N_13363,N_12376,N_12541);
or U13364 (N_13364,N_12539,N_12426);
nand U13365 (N_13365,N_12257,N_12021);
nor U13366 (N_13366,N_12527,N_12835);
nor U13367 (N_13367,N_12087,N_12326);
nor U13368 (N_13368,N_12008,N_12589);
and U13369 (N_13369,N_12512,N_12071);
xor U13370 (N_13370,N_12299,N_12681);
or U13371 (N_13371,N_12363,N_12332);
nor U13372 (N_13372,N_12392,N_12743);
xor U13373 (N_13373,N_12520,N_12893);
nor U13374 (N_13374,N_12826,N_12556);
or U13375 (N_13375,N_12856,N_12159);
nor U13376 (N_13376,N_12432,N_12876);
or U13377 (N_13377,N_12497,N_12630);
and U13378 (N_13378,N_12146,N_12857);
or U13379 (N_13379,N_12062,N_12772);
or U13380 (N_13380,N_12124,N_12838);
nand U13381 (N_13381,N_12980,N_12290);
nor U13382 (N_13382,N_12814,N_12964);
nor U13383 (N_13383,N_12109,N_12791);
nor U13384 (N_13384,N_12927,N_12177);
nand U13385 (N_13385,N_12115,N_12048);
or U13386 (N_13386,N_12904,N_12515);
nor U13387 (N_13387,N_12337,N_12722);
or U13388 (N_13388,N_12294,N_12574);
nor U13389 (N_13389,N_12469,N_12064);
or U13390 (N_13390,N_12542,N_12179);
or U13391 (N_13391,N_12448,N_12642);
nand U13392 (N_13392,N_12538,N_12721);
nor U13393 (N_13393,N_12335,N_12486);
nor U13394 (N_13394,N_12025,N_12576);
xnor U13395 (N_13395,N_12950,N_12102);
and U13396 (N_13396,N_12614,N_12766);
nand U13397 (N_13397,N_12699,N_12641);
nand U13398 (N_13398,N_12374,N_12172);
or U13399 (N_13399,N_12943,N_12946);
or U13400 (N_13400,N_12970,N_12120);
nor U13401 (N_13401,N_12913,N_12734);
nor U13402 (N_13402,N_12505,N_12869);
nor U13403 (N_13403,N_12004,N_12756);
or U13404 (N_13404,N_12872,N_12499);
or U13405 (N_13405,N_12579,N_12084);
or U13406 (N_13406,N_12753,N_12806);
nor U13407 (N_13407,N_12684,N_12406);
nor U13408 (N_13408,N_12981,N_12513);
or U13409 (N_13409,N_12461,N_12181);
or U13410 (N_13410,N_12213,N_12859);
and U13411 (N_13411,N_12570,N_12250);
or U13412 (N_13412,N_12799,N_12728);
or U13413 (N_13413,N_12640,N_12580);
nor U13414 (N_13414,N_12413,N_12922);
and U13415 (N_13415,N_12331,N_12933);
and U13416 (N_13416,N_12380,N_12886);
nand U13417 (N_13417,N_12454,N_12680);
and U13418 (N_13418,N_12993,N_12211);
nor U13419 (N_13419,N_12340,N_12253);
and U13420 (N_13420,N_12060,N_12039);
and U13421 (N_13421,N_12683,N_12966);
or U13422 (N_13422,N_12491,N_12154);
nor U13423 (N_13423,N_12186,N_12260);
nor U13424 (N_13424,N_12668,N_12883);
and U13425 (N_13425,N_12445,N_12056);
or U13426 (N_13426,N_12232,N_12571);
nor U13427 (N_13427,N_12700,N_12727);
nand U13428 (N_13428,N_12713,N_12949);
and U13429 (N_13429,N_12217,N_12305);
or U13430 (N_13430,N_12165,N_12494);
nor U13431 (N_13431,N_12839,N_12796);
nand U13432 (N_13432,N_12302,N_12296);
nand U13433 (N_13433,N_12982,N_12100);
nor U13434 (N_13434,N_12900,N_12817);
nand U13435 (N_13435,N_12138,N_12742);
or U13436 (N_13436,N_12942,N_12313);
or U13437 (N_13437,N_12647,N_12997);
xor U13438 (N_13438,N_12813,N_12316);
or U13439 (N_13439,N_12015,N_12283);
xor U13440 (N_13440,N_12442,N_12969);
or U13441 (N_13441,N_12864,N_12105);
nor U13442 (N_13442,N_12875,N_12669);
or U13443 (N_13443,N_12457,N_12116);
nor U13444 (N_13444,N_12006,N_12007);
xnor U13445 (N_13445,N_12338,N_12411);
or U13446 (N_13446,N_12901,N_12096);
or U13447 (N_13447,N_12804,N_12551);
and U13448 (N_13448,N_12894,N_12191);
or U13449 (N_13449,N_12467,N_12092);
and U13450 (N_13450,N_12139,N_12577);
or U13451 (N_13451,N_12874,N_12582);
and U13452 (N_13452,N_12104,N_12498);
xor U13453 (N_13453,N_12797,N_12841);
or U13454 (N_13454,N_12905,N_12612);
or U13455 (N_13455,N_12451,N_12238);
nor U13456 (N_13456,N_12438,N_12781);
and U13457 (N_13457,N_12851,N_12378);
xor U13458 (N_13458,N_12780,N_12613);
nand U13459 (N_13459,N_12475,N_12401);
and U13460 (N_13460,N_12925,N_12333);
or U13461 (N_13461,N_12569,N_12848);
nor U13462 (N_13462,N_12256,N_12854);
nor U13463 (N_13463,N_12065,N_12405);
xor U13464 (N_13464,N_12871,N_12000);
or U13465 (N_13465,N_12255,N_12009);
and U13466 (N_13466,N_12395,N_12521);
or U13467 (N_13467,N_12593,N_12650);
and U13468 (N_13468,N_12609,N_12160);
and U13469 (N_13469,N_12285,N_12040);
nor U13470 (N_13470,N_12588,N_12769);
nor U13471 (N_13471,N_12168,N_12659);
and U13472 (N_13472,N_12169,N_12667);
nand U13473 (N_13473,N_12252,N_12546);
nand U13474 (N_13474,N_12318,N_12459);
and U13475 (N_13475,N_12983,N_12293);
and U13476 (N_13476,N_12037,N_12790);
nor U13477 (N_13477,N_12385,N_12334);
nor U13478 (N_13478,N_12610,N_12954);
nand U13479 (N_13479,N_12677,N_12428);
or U13480 (N_13480,N_12986,N_12998);
and U13481 (N_13481,N_12059,N_12898);
or U13482 (N_13482,N_12775,N_12619);
and U13483 (N_13483,N_12033,N_12237);
and U13484 (N_13484,N_12914,N_12844);
nor U13485 (N_13485,N_12391,N_12369);
or U13486 (N_13486,N_12282,N_12163);
and U13487 (N_13487,N_12356,N_12601);
or U13488 (N_13488,N_12906,N_12400);
nand U13489 (N_13489,N_12221,N_12249);
or U13490 (N_13490,N_12489,N_12368);
or U13491 (N_13491,N_12468,N_12465);
or U13492 (N_13492,N_12584,N_12424);
or U13493 (N_13493,N_12386,N_12492);
or U13494 (N_13494,N_12930,N_12005);
and U13495 (N_13495,N_12987,N_12692);
nor U13496 (N_13496,N_12046,N_12764);
xor U13497 (N_13497,N_12081,N_12158);
nand U13498 (N_13498,N_12628,N_12524);
xnor U13499 (N_13499,N_12676,N_12345);
or U13500 (N_13500,N_12197,N_12022);
and U13501 (N_13501,N_12239,N_12131);
xnor U13502 (N_13502,N_12549,N_12697);
and U13503 (N_13503,N_12447,N_12111);
nand U13504 (N_13504,N_12634,N_12682);
xnor U13505 (N_13505,N_12080,N_12204);
or U13506 (N_13506,N_12800,N_12375);
or U13507 (N_13507,N_12068,N_12950);
nand U13508 (N_13508,N_12975,N_12452);
nor U13509 (N_13509,N_12599,N_12701);
and U13510 (N_13510,N_12296,N_12649);
and U13511 (N_13511,N_12975,N_12362);
nor U13512 (N_13512,N_12746,N_12798);
xor U13513 (N_13513,N_12136,N_12801);
nand U13514 (N_13514,N_12137,N_12898);
nor U13515 (N_13515,N_12725,N_12301);
nand U13516 (N_13516,N_12490,N_12709);
nor U13517 (N_13517,N_12467,N_12601);
or U13518 (N_13518,N_12886,N_12645);
and U13519 (N_13519,N_12655,N_12327);
nand U13520 (N_13520,N_12442,N_12753);
nand U13521 (N_13521,N_12920,N_12253);
nand U13522 (N_13522,N_12723,N_12999);
nor U13523 (N_13523,N_12374,N_12539);
nor U13524 (N_13524,N_12905,N_12639);
or U13525 (N_13525,N_12486,N_12059);
nor U13526 (N_13526,N_12069,N_12928);
or U13527 (N_13527,N_12703,N_12754);
and U13528 (N_13528,N_12721,N_12971);
nor U13529 (N_13529,N_12991,N_12335);
nor U13530 (N_13530,N_12108,N_12125);
and U13531 (N_13531,N_12231,N_12098);
nand U13532 (N_13532,N_12569,N_12505);
or U13533 (N_13533,N_12336,N_12913);
nor U13534 (N_13534,N_12743,N_12430);
or U13535 (N_13535,N_12734,N_12648);
nand U13536 (N_13536,N_12961,N_12083);
and U13537 (N_13537,N_12448,N_12805);
or U13538 (N_13538,N_12363,N_12923);
nand U13539 (N_13539,N_12489,N_12564);
xor U13540 (N_13540,N_12728,N_12551);
and U13541 (N_13541,N_12678,N_12239);
xnor U13542 (N_13542,N_12034,N_12215);
and U13543 (N_13543,N_12318,N_12599);
and U13544 (N_13544,N_12530,N_12461);
nor U13545 (N_13545,N_12782,N_12764);
xnor U13546 (N_13546,N_12094,N_12495);
nor U13547 (N_13547,N_12969,N_12983);
and U13548 (N_13548,N_12818,N_12185);
nand U13549 (N_13549,N_12378,N_12521);
nor U13550 (N_13550,N_12141,N_12218);
and U13551 (N_13551,N_12175,N_12728);
and U13552 (N_13552,N_12071,N_12622);
xnor U13553 (N_13553,N_12337,N_12533);
nor U13554 (N_13554,N_12142,N_12049);
nor U13555 (N_13555,N_12377,N_12253);
nor U13556 (N_13556,N_12200,N_12482);
nor U13557 (N_13557,N_12038,N_12521);
nor U13558 (N_13558,N_12778,N_12446);
xnor U13559 (N_13559,N_12010,N_12159);
nor U13560 (N_13560,N_12340,N_12789);
xor U13561 (N_13561,N_12665,N_12335);
nand U13562 (N_13562,N_12626,N_12094);
or U13563 (N_13563,N_12834,N_12203);
or U13564 (N_13564,N_12981,N_12308);
nor U13565 (N_13565,N_12444,N_12387);
nand U13566 (N_13566,N_12371,N_12803);
nand U13567 (N_13567,N_12198,N_12577);
and U13568 (N_13568,N_12036,N_12503);
nor U13569 (N_13569,N_12330,N_12442);
and U13570 (N_13570,N_12870,N_12151);
xnor U13571 (N_13571,N_12648,N_12940);
nor U13572 (N_13572,N_12446,N_12361);
xor U13573 (N_13573,N_12073,N_12679);
or U13574 (N_13574,N_12327,N_12221);
nand U13575 (N_13575,N_12142,N_12827);
xor U13576 (N_13576,N_12031,N_12511);
and U13577 (N_13577,N_12640,N_12307);
or U13578 (N_13578,N_12105,N_12284);
and U13579 (N_13579,N_12664,N_12320);
and U13580 (N_13580,N_12253,N_12598);
nand U13581 (N_13581,N_12213,N_12432);
and U13582 (N_13582,N_12414,N_12080);
nand U13583 (N_13583,N_12448,N_12739);
nor U13584 (N_13584,N_12087,N_12649);
nor U13585 (N_13585,N_12598,N_12414);
and U13586 (N_13586,N_12490,N_12193);
and U13587 (N_13587,N_12664,N_12606);
nand U13588 (N_13588,N_12687,N_12935);
and U13589 (N_13589,N_12712,N_12735);
and U13590 (N_13590,N_12275,N_12733);
and U13591 (N_13591,N_12305,N_12572);
or U13592 (N_13592,N_12630,N_12735);
nand U13593 (N_13593,N_12200,N_12000);
nor U13594 (N_13594,N_12017,N_12805);
xnor U13595 (N_13595,N_12819,N_12073);
nand U13596 (N_13596,N_12035,N_12084);
and U13597 (N_13597,N_12234,N_12408);
or U13598 (N_13598,N_12532,N_12270);
nor U13599 (N_13599,N_12430,N_12032);
or U13600 (N_13600,N_12529,N_12977);
and U13601 (N_13601,N_12311,N_12166);
nor U13602 (N_13602,N_12701,N_12846);
nor U13603 (N_13603,N_12184,N_12083);
xnor U13604 (N_13604,N_12620,N_12166);
nor U13605 (N_13605,N_12452,N_12556);
xor U13606 (N_13606,N_12351,N_12715);
xor U13607 (N_13607,N_12723,N_12018);
nand U13608 (N_13608,N_12680,N_12215);
nor U13609 (N_13609,N_12797,N_12729);
nor U13610 (N_13610,N_12101,N_12483);
or U13611 (N_13611,N_12335,N_12121);
and U13612 (N_13612,N_12286,N_12444);
or U13613 (N_13613,N_12297,N_12054);
or U13614 (N_13614,N_12267,N_12778);
nor U13615 (N_13615,N_12678,N_12718);
nor U13616 (N_13616,N_12806,N_12023);
nor U13617 (N_13617,N_12199,N_12227);
or U13618 (N_13618,N_12277,N_12730);
nand U13619 (N_13619,N_12639,N_12616);
nand U13620 (N_13620,N_12802,N_12692);
or U13621 (N_13621,N_12621,N_12510);
or U13622 (N_13622,N_12716,N_12471);
nor U13623 (N_13623,N_12641,N_12451);
and U13624 (N_13624,N_12927,N_12002);
nand U13625 (N_13625,N_12885,N_12628);
nor U13626 (N_13626,N_12419,N_12141);
xor U13627 (N_13627,N_12092,N_12773);
or U13628 (N_13628,N_12754,N_12887);
nand U13629 (N_13629,N_12812,N_12718);
xnor U13630 (N_13630,N_12145,N_12372);
or U13631 (N_13631,N_12334,N_12748);
nand U13632 (N_13632,N_12333,N_12690);
nand U13633 (N_13633,N_12260,N_12171);
nor U13634 (N_13634,N_12169,N_12635);
nand U13635 (N_13635,N_12881,N_12407);
xnor U13636 (N_13636,N_12620,N_12524);
and U13637 (N_13637,N_12988,N_12534);
nand U13638 (N_13638,N_12354,N_12132);
nor U13639 (N_13639,N_12676,N_12583);
nor U13640 (N_13640,N_12386,N_12625);
xor U13641 (N_13641,N_12396,N_12578);
xnor U13642 (N_13642,N_12019,N_12477);
nor U13643 (N_13643,N_12122,N_12175);
and U13644 (N_13644,N_12101,N_12117);
nand U13645 (N_13645,N_12718,N_12287);
nand U13646 (N_13646,N_12663,N_12796);
xnor U13647 (N_13647,N_12791,N_12073);
nand U13648 (N_13648,N_12661,N_12200);
xnor U13649 (N_13649,N_12024,N_12135);
nor U13650 (N_13650,N_12808,N_12819);
or U13651 (N_13651,N_12997,N_12968);
xor U13652 (N_13652,N_12885,N_12878);
and U13653 (N_13653,N_12826,N_12681);
nand U13654 (N_13654,N_12899,N_12763);
or U13655 (N_13655,N_12705,N_12607);
or U13656 (N_13656,N_12799,N_12278);
and U13657 (N_13657,N_12033,N_12898);
nor U13658 (N_13658,N_12718,N_12712);
nor U13659 (N_13659,N_12873,N_12804);
nor U13660 (N_13660,N_12880,N_12792);
or U13661 (N_13661,N_12850,N_12112);
nor U13662 (N_13662,N_12072,N_12243);
nand U13663 (N_13663,N_12741,N_12380);
nor U13664 (N_13664,N_12706,N_12405);
nor U13665 (N_13665,N_12557,N_12813);
or U13666 (N_13666,N_12131,N_12758);
nor U13667 (N_13667,N_12697,N_12741);
nand U13668 (N_13668,N_12819,N_12246);
and U13669 (N_13669,N_12855,N_12422);
nor U13670 (N_13670,N_12102,N_12803);
nor U13671 (N_13671,N_12784,N_12494);
or U13672 (N_13672,N_12845,N_12106);
nor U13673 (N_13673,N_12168,N_12062);
or U13674 (N_13674,N_12648,N_12089);
or U13675 (N_13675,N_12581,N_12099);
or U13676 (N_13676,N_12170,N_12813);
or U13677 (N_13677,N_12102,N_12314);
nor U13678 (N_13678,N_12393,N_12499);
and U13679 (N_13679,N_12481,N_12179);
nand U13680 (N_13680,N_12417,N_12825);
or U13681 (N_13681,N_12264,N_12148);
and U13682 (N_13682,N_12066,N_12335);
nor U13683 (N_13683,N_12802,N_12789);
nor U13684 (N_13684,N_12809,N_12188);
and U13685 (N_13685,N_12488,N_12176);
and U13686 (N_13686,N_12868,N_12941);
nor U13687 (N_13687,N_12509,N_12799);
or U13688 (N_13688,N_12620,N_12156);
nor U13689 (N_13689,N_12158,N_12348);
xor U13690 (N_13690,N_12854,N_12585);
xor U13691 (N_13691,N_12978,N_12209);
or U13692 (N_13692,N_12413,N_12453);
nor U13693 (N_13693,N_12674,N_12525);
nand U13694 (N_13694,N_12368,N_12715);
nor U13695 (N_13695,N_12129,N_12471);
or U13696 (N_13696,N_12481,N_12035);
or U13697 (N_13697,N_12488,N_12611);
or U13698 (N_13698,N_12278,N_12127);
nor U13699 (N_13699,N_12230,N_12617);
and U13700 (N_13700,N_12900,N_12916);
nor U13701 (N_13701,N_12327,N_12975);
xnor U13702 (N_13702,N_12386,N_12320);
xnor U13703 (N_13703,N_12159,N_12897);
nor U13704 (N_13704,N_12562,N_12880);
nand U13705 (N_13705,N_12796,N_12505);
nand U13706 (N_13706,N_12872,N_12833);
nand U13707 (N_13707,N_12327,N_12690);
or U13708 (N_13708,N_12024,N_12349);
nor U13709 (N_13709,N_12990,N_12936);
and U13710 (N_13710,N_12730,N_12072);
xnor U13711 (N_13711,N_12193,N_12589);
nor U13712 (N_13712,N_12624,N_12451);
nor U13713 (N_13713,N_12143,N_12572);
xor U13714 (N_13714,N_12353,N_12313);
nand U13715 (N_13715,N_12875,N_12786);
nor U13716 (N_13716,N_12618,N_12461);
nor U13717 (N_13717,N_12743,N_12961);
nor U13718 (N_13718,N_12068,N_12186);
nand U13719 (N_13719,N_12560,N_12080);
nand U13720 (N_13720,N_12848,N_12912);
and U13721 (N_13721,N_12044,N_12804);
and U13722 (N_13722,N_12591,N_12291);
and U13723 (N_13723,N_12905,N_12960);
and U13724 (N_13724,N_12192,N_12883);
nand U13725 (N_13725,N_12276,N_12491);
and U13726 (N_13726,N_12016,N_12495);
nor U13727 (N_13727,N_12002,N_12562);
or U13728 (N_13728,N_12326,N_12562);
and U13729 (N_13729,N_12006,N_12936);
nand U13730 (N_13730,N_12737,N_12492);
nand U13731 (N_13731,N_12971,N_12717);
xnor U13732 (N_13732,N_12285,N_12614);
xor U13733 (N_13733,N_12376,N_12945);
nor U13734 (N_13734,N_12509,N_12939);
xnor U13735 (N_13735,N_12316,N_12267);
nor U13736 (N_13736,N_12212,N_12526);
or U13737 (N_13737,N_12406,N_12457);
nand U13738 (N_13738,N_12393,N_12480);
or U13739 (N_13739,N_12674,N_12703);
xor U13740 (N_13740,N_12557,N_12756);
and U13741 (N_13741,N_12246,N_12635);
or U13742 (N_13742,N_12181,N_12518);
nand U13743 (N_13743,N_12351,N_12286);
and U13744 (N_13744,N_12083,N_12865);
nor U13745 (N_13745,N_12882,N_12163);
and U13746 (N_13746,N_12696,N_12167);
and U13747 (N_13747,N_12216,N_12011);
nand U13748 (N_13748,N_12864,N_12103);
nand U13749 (N_13749,N_12371,N_12219);
and U13750 (N_13750,N_12023,N_12419);
or U13751 (N_13751,N_12944,N_12325);
or U13752 (N_13752,N_12809,N_12208);
or U13753 (N_13753,N_12890,N_12294);
nor U13754 (N_13754,N_12776,N_12246);
nor U13755 (N_13755,N_12026,N_12509);
xnor U13756 (N_13756,N_12646,N_12817);
or U13757 (N_13757,N_12104,N_12370);
nor U13758 (N_13758,N_12893,N_12968);
and U13759 (N_13759,N_12555,N_12687);
or U13760 (N_13760,N_12329,N_12662);
and U13761 (N_13761,N_12465,N_12743);
and U13762 (N_13762,N_12731,N_12552);
and U13763 (N_13763,N_12071,N_12716);
nand U13764 (N_13764,N_12223,N_12740);
and U13765 (N_13765,N_12524,N_12687);
and U13766 (N_13766,N_12377,N_12142);
nor U13767 (N_13767,N_12354,N_12047);
and U13768 (N_13768,N_12550,N_12035);
or U13769 (N_13769,N_12609,N_12934);
and U13770 (N_13770,N_12747,N_12440);
or U13771 (N_13771,N_12264,N_12477);
and U13772 (N_13772,N_12293,N_12840);
xnor U13773 (N_13773,N_12106,N_12707);
and U13774 (N_13774,N_12763,N_12295);
or U13775 (N_13775,N_12947,N_12387);
or U13776 (N_13776,N_12275,N_12473);
or U13777 (N_13777,N_12546,N_12068);
and U13778 (N_13778,N_12287,N_12944);
nand U13779 (N_13779,N_12315,N_12364);
nand U13780 (N_13780,N_12195,N_12160);
or U13781 (N_13781,N_12687,N_12451);
or U13782 (N_13782,N_12994,N_12604);
nand U13783 (N_13783,N_12988,N_12123);
and U13784 (N_13784,N_12382,N_12001);
or U13785 (N_13785,N_12528,N_12941);
nor U13786 (N_13786,N_12831,N_12792);
nor U13787 (N_13787,N_12012,N_12688);
nor U13788 (N_13788,N_12667,N_12611);
nand U13789 (N_13789,N_12497,N_12225);
xnor U13790 (N_13790,N_12402,N_12034);
xor U13791 (N_13791,N_12165,N_12320);
or U13792 (N_13792,N_12246,N_12003);
or U13793 (N_13793,N_12970,N_12452);
or U13794 (N_13794,N_12327,N_12247);
nand U13795 (N_13795,N_12594,N_12441);
or U13796 (N_13796,N_12259,N_12805);
nand U13797 (N_13797,N_12341,N_12364);
nand U13798 (N_13798,N_12955,N_12519);
nand U13799 (N_13799,N_12169,N_12482);
and U13800 (N_13800,N_12023,N_12021);
and U13801 (N_13801,N_12042,N_12326);
and U13802 (N_13802,N_12804,N_12026);
nor U13803 (N_13803,N_12759,N_12972);
or U13804 (N_13804,N_12141,N_12324);
or U13805 (N_13805,N_12796,N_12966);
nand U13806 (N_13806,N_12164,N_12114);
nor U13807 (N_13807,N_12212,N_12294);
nand U13808 (N_13808,N_12987,N_12521);
and U13809 (N_13809,N_12823,N_12349);
xor U13810 (N_13810,N_12549,N_12178);
or U13811 (N_13811,N_12590,N_12375);
or U13812 (N_13812,N_12511,N_12750);
and U13813 (N_13813,N_12032,N_12952);
nand U13814 (N_13814,N_12602,N_12875);
or U13815 (N_13815,N_12120,N_12702);
or U13816 (N_13816,N_12302,N_12575);
and U13817 (N_13817,N_12143,N_12786);
nand U13818 (N_13818,N_12621,N_12900);
or U13819 (N_13819,N_12325,N_12298);
or U13820 (N_13820,N_12237,N_12876);
nor U13821 (N_13821,N_12296,N_12465);
xnor U13822 (N_13822,N_12644,N_12983);
nand U13823 (N_13823,N_12153,N_12067);
or U13824 (N_13824,N_12682,N_12020);
xnor U13825 (N_13825,N_12163,N_12325);
or U13826 (N_13826,N_12701,N_12442);
and U13827 (N_13827,N_12962,N_12128);
nand U13828 (N_13828,N_12558,N_12414);
nor U13829 (N_13829,N_12394,N_12356);
nand U13830 (N_13830,N_12435,N_12073);
or U13831 (N_13831,N_12101,N_12121);
and U13832 (N_13832,N_12199,N_12379);
nor U13833 (N_13833,N_12036,N_12994);
nor U13834 (N_13834,N_12817,N_12848);
xor U13835 (N_13835,N_12721,N_12097);
nor U13836 (N_13836,N_12468,N_12779);
nor U13837 (N_13837,N_12923,N_12937);
xnor U13838 (N_13838,N_12556,N_12747);
or U13839 (N_13839,N_12242,N_12071);
or U13840 (N_13840,N_12815,N_12428);
and U13841 (N_13841,N_12688,N_12069);
nand U13842 (N_13842,N_12238,N_12780);
and U13843 (N_13843,N_12168,N_12760);
or U13844 (N_13844,N_12396,N_12049);
nand U13845 (N_13845,N_12938,N_12221);
or U13846 (N_13846,N_12565,N_12204);
or U13847 (N_13847,N_12381,N_12817);
xor U13848 (N_13848,N_12706,N_12012);
xnor U13849 (N_13849,N_12153,N_12468);
nand U13850 (N_13850,N_12685,N_12872);
xnor U13851 (N_13851,N_12718,N_12478);
and U13852 (N_13852,N_12387,N_12496);
or U13853 (N_13853,N_12597,N_12346);
and U13854 (N_13854,N_12716,N_12384);
or U13855 (N_13855,N_12905,N_12779);
and U13856 (N_13856,N_12394,N_12110);
nor U13857 (N_13857,N_12066,N_12248);
xnor U13858 (N_13858,N_12703,N_12710);
or U13859 (N_13859,N_12374,N_12418);
or U13860 (N_13860,N_12521,N_12659);
nand U13861 (N_13861,N_12716,N_12321);
or U13862 (N_13862,N_12618,N_12538);
or U13863 (N_13863,N_12923,N_12255);
nand U13864 (N_13864,N_12492,N_12277);
or U13865 (N_13865,N_12715,N_12644);
or U13866 (N_13866,N_12617,N_12285);
nand U13867 (N_13867,N_12105,N_12429);
or U13868 (N_13868,N_12093,N_12762);
or U13869 (N_13869,N_12049,N_12756);
nor U13870 (N_13870,N_12676,N_12436);
nand U13871 (N_13871,N_12992,N_12528);
nand U13872 (N_13872,N_12448,N_12506);
nand U13873 (N_13873,N_12036,N_12244);
xnor U13874 (N_13874,N_12214,N_12637);
and U13875 (N_13875,N_12859,N_12989);
nor U13876 (N_13876,N_12058,N_12209);
nand U13877 (N_13877,N_12218,N_12212);
and U13878 (N_13878,N_12069,N_12796);
nor U13879 (N_13879,N_12022,N_12977);
xnor U13880 (N_13880,N_12791,N_12661);
nor U13881 (N_13881,N_12963,N_12902);
nor U13882 (N_13882,N_12821,N_12856);
nor U13883 (N_13883,N_12789,N_12140);
nand U13884 (N_13884,N_12864,N_12286);
nor U13885 (N_13885,N_12738,N_12271);
and U13886 (N_13886,N_12357,N_12047);
nor U13887 (N_13887,N_12826,N_12469);
and U13888 (N_13888,N_12551,N_12459);
and U13889 (N_13889,N_12021,N_12851);
nor U13890 (N_13890,N_12836,N_12124);
or U13891 (N_13891,N_12901,N_12022);
nand U13892 (N_13892,N_12000,N_12691);
or U13893 (N_13893,N_12121,N_12192);
nand U13894 (N_13894,N_12601,N_12955);
nand U13895 (N_13895,N_12414,N_12588);
nor U13896 (N_13896,N_12381,N_12539);
or U13897 (N_13897,N_12766,N_12985);
or U13898 (N_13898,N_12807,N_12851);
and U13899 (N_13899,N_12149,N_12795);
or U13900 (N_13900,N_12031,N_12196);
nor U13901 (N_13901,N_12055,N_12636);
xor U13902 (N_13902,N_12986,N_12388);
nand U13903 (N_13903,N_12403,N_12809);
or U13904 (N_13904,N_12042,N_12685);
nand U13905 (N_13905,N_12588,N_12624);
nand U13906 (N_13906,N_12736,N_12319);
nand U13907 (N_13907,N_12192,N_12686);
and U13908 (N_13908,N_12764,N_12585);
nand U13909 (N_13909,N_12409,N_12086);
and U13910 (N_13910,N_12236,N_12265);
and U13911 (N_13911,N_12520,N_12313);
and U13912 (N_13912,N_12680,N_12244);
xor U13913 (N_13913,N_12356,N_12674);
or U13914 (N_13914,N_12139,N_12419);
nand U13915 (N_13915,N_12602,N_12250);
or U13916 (N_13916,N_12253,N_12409);
or U13917 (N_13917,N_12308,N_12157);
xor U13918 (N_13918,N_12925,N_12188);
nand U13919 (N_13919,N_12563,N_12876);
nand U13920 (N_13920,N_12922,N_12004);
and U13921 (N_13921,N_12085,N_12388);
nor U13922 (N_13922,N_12490,N_12792);
and U13923 (N_13923,N_12058,N_12080);
or U13924 (N_13924,N_12779,N_12382);
and U13925 (N_13925,N_12159,N_12228);
and U13926 (N_13926,N_12691,N_12265);
and U13927 (N_13927,N_12184,N_12312);
nor U13928 (N_13928,N_12558,N_12953);
nand U13929 (N_13929,N_12004,N_12562);
nand U13930 (N_13930,N_12748,N_12771);
xor U13931 (N_13931,N_12516,N_12598);
xnor U13932 (N_13932,N_12618,N_12583);
and U13933 (N_13933,N_12450,N_12420);
nand U13934 (N_13934,N_12990,N_12163);
and U13935 (N_13935,N_12578,N_12468);
nor U13936 (N_13936,N_12442,N_12370);
or U13937 (N_13937,N_12739,N_12785);
and U13938 (N_13938,N_12258,N_12338);
or U13939 (N_13939,N_12402,N_12433);
xor U13940 (N_13940,N_12406,N_12281);
and U13941 (N_13941,N_12705,N_12270);
nor U13942 (N_13942,N_12570,N_12852);
and U13943 (N_13943,N_12820,N_12485);
nand U13944 (N_13944,N_12023,N_12155);
nand U13945 (N_13945,N_12829,N_12176);
nor U13946 (N_13946,N_12312,N_12279);
nor U13947 (N_13947,N_12732,N_12547);
and U13948 (N_13948,N_12277,N_12631);
and U13949 (N_13949,N_12972,N_12664);
nor U13950 (N_13950,N_12709,N_12015);
nor U13951 (N_13951,N_12562,N_12569);
nor U13952 (N_13952,N_12490,N_12747);
nand U13953 (N_13953,N_12203,N_12811);
nor U13954 (N_13954,N_12863,N_12758);
or U13955 (N_13955,N_12262,N_12230);
or U13956 (N_13956,N_12914,N_12189);
xnor U13957 (N_13957,N_12287,N_12775);
xnor U13958 (N_13958,N_12680,N_12540);
nand U13959 (N_13959,N_12146,N_12990);
nand U13960 (N_13960,N_12508,N_12454);
or U13961 (N_13961,N_12877,N_12563);
and U13962 (N_13962,N_12159,N_12094);
nor U13963 (N_13963,N_12955,N_12734);
or U13964 (N_13964,N_12620,N_12492);
nor U13965 (N_13965,N_12264,N_12072);
or U13966 (N_13966,N_12242,N_12994);
or U13967 (N_13967,N_12196,N_12772);
nor U13968 (N_13968,N_12204,N_12231);
and U13969 (N_13969,N_12888,N_12719);
or U13970 (N_13970,N_12576,N_12150);
or U13971 (N_13971,N_12685,N_12618);
nor U13972 (N_13972,N_12038,N_12014);
xnor U13973 (N_13973,N_12143,N_12763);
or U13974 (N_13974,N_12251,N_12980);
and U13975 (N_13975,N_12664,N_12844);
and U13976 (N_13976,N_12781,N_12052);
nand U13977 (N_13977,N_12424,N_12261);
and U13978 (N_13978,N_12636,N_12170);
or U13979 (N_13979,N_12148,N_12190);
and U13980 (N_13980,N_12715,N_12010);
nand U13981 (N_13981,N_12754,N_12444);
or U13982 (N_13982,N_12204,N_12968);
and U13983 (N_13983,N_12553,N_12996);
nand U13984 (N_13984,N_12124,N_12940);
and U13985 (N_13985,N_12233,N_12015);
or U13986 (N_13986,N_12119,N_12690);
or U13987 (N_13987,N_12047,N_12534);
or U13988 (N_13988,N_12283,N_12960);
or U13989 (N_13989,N_12360,N_12451);
or U13990 (N_13990,N_12522,N_12222);
nor U13991 (N_13991,N_12537,N_12831);
nor U13992 (N_13992,N_12540,N_12427);
or U13993 (N_13993,N_12361,N_12833);
and U13994 (N_13994,N_12027,N_12945);
or U13995 (N_13995,N_12026,N_12776);
nand U13996 (N_13996,N_12637,N_12517);
or U13997 (N_13997,N_12825,N_12757);
nor U13998 (N_13998,N_12829,N_12420);
nor U13999 (N_13999,N_12743,N_12163);
nand U14000 (N_14000,N_13969,N_13616);
nand U14001 (N_14001,N_13805,N_13997);
and U14002 (N_14002,N_13188,N_13135);
nand U14003 (N_14003,N_13625,N_13473);
nand U14004 (N_14004,N_13324,N_13964);
and U14005 (N_14005,N_13892,N_13825);
or U14006 (N_14006,N_13962,N_13054);
and U14007 (N_14007,N_13191,N_13986);
xnor U14008 (N_14008,N_13077,N_13586);
and U14009 (N_14009,N_13666,N_13701);
nor U14010 (N_14010,N_13945,N_13430);
or U14011 (N_14011,N_13059,N_13799);
or U14012 (N_14012,N_13012,N_13201);
or U14013 (N_14013,N_13459,N_13779);
nand U14014 (N_14014,N_13500,N_13877);
nor U14015 (N_14015,N_13605,N_13461);
nor U14016 (N_14016,N_13309,N_13338);
nand U14017 (N_14017,N_13818,N_13774);
nor U14018 (N_14018,N_13631,N_13656);
nand U14019 (N_14019,N_13470,N_13770);
nand U14020 (N_14020,N_13662,N_13103);
and U14021 (N_14021,N_13957,N_13238);
nor U14022 (N_14022,N_13776,N_13959);
and U14023 (N_14023,N_13953,N_13780);
nand U14024 (N_14024,N_13136,N_13541);
and U14025 (N_14025,N_13761,N_13041);
nand U14026 (N_14026,N_13366,N_13325);
and U14027 (N_14027,N_13177,N_13222);
xnor U14028 (N_14028,N_13013,N_13767);
and U14029 (N_14029,N_13383,N_13963);
nor U14030 (N_14030,N_13123,N_13358);
nand U14031 (N_14031,N_13941,N_13693);
nand U14032 (N_14032,N_13518,N_13420);
nand U14033 (N_14033,N_13965,N_13539);
xnor U14034 (N_14034,N_13442,N_13471);
nand U14035 (N_14035,N_13574,N_13389);
and U14036 (N_14036,N_13249,N_13478);
and U14037 (N_14037,N_13529,N_13487);
nor U14038 (N_14038,N_13072,N_13122);
nor U14039 (N_14039,N_13764,N_13398);
and U14040 (N_14040,N_13102,N_13579);
or U14041 (N_14041,N_13460,N_13657);
or U14042 (N_14042,N_13166,N_13113);
or U14043 (N_14043,N_13956,N_13450);
nor U14044 (N_14044,N_13536,N_13567);
and U14045 (N_14045,N_13152,N_13340);
or U14046 (N_14046,N_13226,N_13407);
or U14047 (N_14047,N_13590,N_13243);
xor U14048 (N_14048,N_13221,N_13623);
or U14049 (N_14049,N_13516,N_13708);
nor U14050 (N_14050,N_13934,N_13068);
nand U14051 (N_14051,N_13772,N_13961);
or U14052 (N_14052,N_13350,N_13568);
xnor U14053 (N_14053,N_13663,N_13045);
xnor U14054 (N_14054,N_13233,N_13985);
and U14055 (N_14055,N_13486,N_13224);
nand U14056 (N_14056,N_13523,N_13749);
and U14057 (N_14057,N_13667,N_13786);
or U14058 (N_14058,N_13798,N_13317);
or U14059 (N_14059,N_13261,N_13995);
or U14060 (N_14060,N_13272,N_13328);
or U14061 (N_14061,N_13648,N_13791);
or U14062 (N_14062,N_13190,N_13276);
nor U14063 (N_14063,N_13722,N_13641);
nand U14064 (N_14064,N_13534,N_13411);
nor U14065 (N_14065,N_13427,N_13385);
nand U14066 (N_14066,N_13680,N_13329);
or U14067 (N_14067,N_13967,N_13946);
nand U14068 (N_14068,N_13333,N_13158);
xor U14069 (N_14069,N_13312,N_13092);
nand U14070 (N_14070,N_13245,N_13704);
xnor U14071 (N_14071,N_13668,N_13371);
nor U14072 (N_14072,N_13075,N_13337);
nand U14073 (N_14073,N_13843,N_13356);
or U14074 (N_14074,N_13007,N_13467);
xnor U14075 (N_14075,N_13160,N_13918);
xor U14076 (N_14076,N_13931,N_13869);
nor U14077 (N_14077,N_13828,N_13597);
and U14078 (N_14078,N_13495,N_13219);
nor U14079 (N_14079,N_13928,N_13409);
nor U14080 (N_14080,N_13562,N_13800);
or U14081 (N_14081,N_13748,N_13380);
or U14082 (N_14082,N_13996,N_13431);
and U14083 (N_14083,N_13204,N_13556);
or U14084 (N_14084,N_13862,N_13355);
nand U14085 (N_14085,N_13729,N_13530);
nand U14086 (N_14086,N_13917,N_13189);
and U14087 (N_14087,N_13766,N_13129);
or U14088 (N_14088,N_13935,N_13565);
or U14089 (N_14089,N_13638,N_13699);
nor U14090 (N_14090,N_13304,N_13402);
and U14091 (N_14091,N_13692,N_13857);
nor U14092 (N_14092,N_13308,N_13073);
and U14093 (N_14093,N_13794,N_13617);
or U14094 (N_14094,N_13876,N_13469);
nor U14095 (N_14095,N_13528,N_13033);
and U14096 (N_14096,N_13148,N_13532);
or U14097 (N_14097,N_13452,N_13681);
nand U14098 (N_14098,N_13480,N_13105);
and U14099 (N_14099,N_13697,N_13119);
nand U14100 (N_14100,N_13318,N_13739);
nor U14101 (N_14101,N_13115,N_13374);
xnor U14102 (N_14102,N_13895,N_13923);
nor U14103 (N_14103,N_13353,N_13365);
nand U14104 (N_14104,N_13335,N_13417);
xnor U14105 (N_14105,N_13030,N_13503);
or U14106 (N_14106,N_13808,N_13378);
and U14107 (N_14107,N_13582,N_13206);
nand U14108 (N_14108,N_13234,N_13302);
nor U14109 (N_14109,N_13730,N_13367);
or U14110 (N_14110,N_13140,N_13838);
and U14111 (N_14111,N_13978,N_13440);
xnor U14112 (N_14112,N_13698,N_13652);
and U14113 (N_14113,N_13179,N_13051);
nor U14114 (N_14114,N_13546,N_13632);
xor U14115 (N_14115,N_13745,N_13482);
and U14116 (N_14116,N_13720,N_13743);
xor U14117 (N_14117,N_13907,N_13133);
xor U14118 (N_14118,N_13071,N_13542);
nor U14119 (N_14119,N_13010,N_13989);
or U14120 (N_14120,N_13384,N_13575);
or U14121 (N_14121,N_13437,N_13540);
or U14122 (N_14122,N_13062,N_13581);
nor U14123 (N_14123,N_13472,N_13058);
nand U14124 (N_14124,N_13817,N_13639);
nand U14125 (N_14125,N_13858,N_13239);
and U14126 (N_14126,N_13228,N_13866);
and U14127 (N_14127,N_13036,N_13732);
nand U14128 (N_14128,N_13836,N_13802);
nand U14129 (N_14129,N_13479,N_13065);
or U14130 (N_14130,N_13282,N_13047);
or U14131 (N_14131,N_13455,N_13307);
nand U14132 (N_14132,N_13173,N_13576);
nand U14133 (N_14133,N_13476,N_13814);
or U14134 (N_14134,N_13438,N_13882);
and U14135 (N_14135,N_13138,N_13775);
xnor U14136 (N_14136,N_13100,N_13305);
nor U14137 (N_14137,N_13607,N_13481);
and U14138 (N_14138,N_13275,N_13126);
xor U14139 (N_14139,N_13551,N_13603);
or U14140 (N_14140,N_13872,N_13564);
and U14141 (N_14141,N_13181,N_13379);
and U14142 (N_14142,N_13019,N_13526);
or U14143 (N_14143,N_13214,N_13762);
and U14144 (N_14144,N_13194,N_13024);
xor U14145 (N_14145,N_13155,N_13841);
nor U14146 (N_14146,N_13008,N_13583);
nor U14147 (N_14147,N_13125,N_13313);
or U14148 (N_14148,N_13410,N_13104);
nand U14149 (N_14149,N_13273,N_13061);
or U14150 (N_14150,N_13971,N_13608);
or U14151 (N_14151,N_13498,N_13844);
or U14152 (N_14152,N_13533,N_13205);
nand U14153 (N_14153,N_13180,N_13053);
nand U14154 (N_14154,N_13506,N_13364);
and U14155 (N_14155,N_13975,N_13773);
and U14156 (N_14156,N_13376,N_13485);
and U14157 (N_14157,N_13684,N_13213);
nor U14158 (N_14158,N_13032,N_13695);
or U14159 (N_14159,N_13675,N_13419);
xor U14160 (N_14160,N_13390,N_13852);
nor U14161 (N_14161,N_13904,N_13588);
xnor U14162 (N_14162,N_13421,N_13099);
nand U14163 (N_14163,N_13199,N_13001);
nand U14164 (N_14164,N_13132,N_13203);
nand U14165 (N_14165,N_13970,N_13332);
and U14166 (N_14166,N_13973,N_13756);
xnor U14167 (N_14167,N_13446,N_13785);
nand U14168 (N_14168,N_13274,N_13991);
nand U14169 (N_14169,N_13783,N_13363);
and U14170 (N_14170,N_13422,N_13829);
nand U14171 (N_14171,N_13078,N_13393);
xnor U14172 (N_14172,N_13112,N_13792);
xnor U14173 (N_14173,N_13035,N_13845);
nor U14174 (N_14174,N_13170,N_13911);
nand U14175 (N_14175,N_13821,N_13354);
and U14176 (N_14176,N_13323,N_13369);
and U14177 (N_14177,N_13299,N_13893);
nand U14178 (N_14178,N_13050,N_13039);
xnor U14179 (N_14179,N_13968,N_13236);
or U14180 (N_14180,N_13504,N_13755);
nand U14181 (N_14181,N_13510,N_13860);
and U14182 (N_14182,N_13406,N_13824);
xor U14183 (N_14183,N_13057,N_13240);
nand U14184 (N_14184,N_13705,N_13741);
nand U14185 (N_14185,N_13003,N_13587);
nor U14186 (N_14186,N_13381,N_13670);
or U14187 (N_14187,N_13146,N_13781);
or U14188 (N_14188,N_13707,N_13508);
or U14189 (N_14189,N_13382,N_13489);
nand U14190 (N_14190,N_13981,N_13445);
nor U14191 (N_14191,N_13782,N_13207);
or U14192 (N_14192,N_13492,N_13833);
and U14193 (N_14193,N_13509,N_13933);
nand U14194 (N_14194,N_13700,N_13831);
and U14195 (N_14195,N_13908,N_13232);
nor U14196 (N_14196,N_13804,N_13801);
xor U14197 (N_14197,N_13880,N_13763);
or U14198 (N_14198,N_13477,N_13106);
or U14199 (N_14199,N_13111,N_13691);
nor U14200 (N_14200,N_13223,N_13859);
and U14201 (N_14201,N_13255,N_13633);
and U14202 (N_14202,N_13026,N_13496);
and U14203 (N_14203,N_13426,N_13063);
or U14204 (N_14204,N_13458,N_13905);
xor U14205 (N_14205,N_13490,N_13352);
nand U14206 (N_14206,N_13884,N_13271);
and U14207 (N_14207,N_13982,N_13595);
nor U14208 (N_14208,N_13294,N_13674);
or U14209 (N_14209,N_13640,N_13341);
nor U14210 (N_14210,N_13644,N_13686);
nor U14211 (N_14211,N_13230,N_13578);
xor U14212 (N_14212,N_13916,N_13277);
and U14213 (N_14213,N_13002,N_13871);
xor U14214 (N_14214,N_13344,N_13447);
or U14215 (N_14215,N_13217,N_13519);
nand U14216 (N_14216,N_13387,N_13643);
xor U14217 (N_14217,N_13734,N_13083);
nand U14218 (N_14218,N_13149,N_13628);
or U14219 (N_14219,N_13462,N_13719);
or U14220 (N_14220,N_13827,N_13789);
nand U14221 (N_14221,N_13919,N_13555);
nor U14222 (N_14222,N_13987,N_13598);
nand U14223 (N_14223,N_13940,N_13930);
and U14224 (N_14224,N_13044,N_13316);
nand U14225 (N_14225,N_13349,N_13690);
xor U14226 (N_14226,N_13851,N_13795);
nand U14227 (N_14227,N_13883,N_13184);
nand U14228 (N_14228,N_13327,N_13863);
nand U14229 (N_14229,N_13938,N_13793);
nor U14230 (N_14230,N_13563,N_13416);
xor U14231 (N_14231,N_13171,N_13837);
nand U14232 (N_14232,N_13830,N_13310);
or U14233 (N_14233,N_13647,N_13216);
and U14234 (N_14234,N_13635,N_13400);
nor U14235 (N_14235,N_13881,N_13257);
nor U14236 (N_14236,N_13006,N_13513);
or U14237 (N_14237,N_13321,N_13098);
nand U14238 (N_14238,N_13183,N_13157);
and U14239 (N_14239,N_13910,N_13254);
or U14240 (N_14240,N_13040,N_13022);
xor U14241 (N_14241,N_13293,N_13517);
nor U14242 (N_14242,N_13742,N_13569);
or U14243 (N_14243,N_13314,N_13235);
and U14244 (N_14244,N_13463,N_13088);
nand U14245 (N_14245,N_13089,N_13056);
and U14246 (N_14246,N_13456,N_13591);
and U14247 (N_14247,N_13849,N_13676);
nor U14248 (N_14248,N_13167,N_13303);
nor U14249 (N_14249,N_13637,N_13009);
and U14250 (N_14250,N_13535,N_13561);
nand U14251 (N_14251,N_13163,N_13491);
or U14252 (N_14252,N_13550,N_13602);
nor U14253 (N_14253,N_13464,N_13237);
nand U14254 (N_14254,N_13977,N_13156);
xnor U14255 (N_14255,N_13746,N_13474);
nand U14256 (N_14256,N_13218,N_13976);
and U14257 (N_14257,N_13178,N_13262);
or U14258 (N_14258,N_13453,N_13645);
or U14259 (N_14259,N_13658,N_13891);
or U14260 (N_14260,N_13401,N_13248);
nor U14261 (N_14261,N_13424,N_13418);
nand U14262 (N_14262,N_13027,N_13966);
xor U14263 (N_14263,N_13664,N_13028);
xnor U14264 (N_14264,N_13483,N_13428);
xnor U14265 (N_14265,N_13220,N_13484);
nor U14266 (N_14266,N_13765,N_13980);
or U14267 (N_14267,N_13673,N_13448);
and U14268 (N_14268,N_13209,N_13468);
xnor U14269 (N_14269,N_13840,N_13124);
nand U14270 (N_14270,N_13524,N_13894);
nand U14271 (N_14271,N_13947,N_13090);
nor U14272 (N_14272,N_13441,N_13853);
and U14273 (N_14273,N_13614,N_13839);
nor U14274 (N_14274,N_13343,N_13286);
xor U14275 (N_14275,N_13992,N_13005);
xor U14276 (N_14276,N_13711,N_13466);
nand U14277 (N_14277,N_13143,N_13733);
or U14278 (N_14278,N_13750,N_13377);
and U14279 (N_14279,N_13580,N_13787);
xnor U14280 (N_14280,N_13788,N_13423);
nor U14281 (N_14281,N_13291,N_13298);
nor U14282 (N_14282,N_13899,N_13703);
nand U14283 (N_14283,N_13758,N_13187);
nand U14284 (N_14284,N_13267,N_13898);
or U14285 (N_14285,N_13988,N_13347);
xnor U14286 (N_14286,N_13622,N_13856);
nand U14287 (N_14287,N_13936,N_13326);
nand U14288 (N_14288,N_13901,N_13599);
and U14289 (N_14289,N_13131,N_13646);
xnor U14290 (N_14290,N_13714,N_13672);
nand U14291 (N_14291,N_13016,N_13682);
xor U14292 (N_14292,N_13688,N_13724);
and U14293 (N_14293,N_13436,N_13300);
or U14294 (N_14294,N_13151,N_13162);
nand U14295 (N_14295,N_13070,N_13937);
and U14296 (N_14296,N_13336,N_13589);
nand U14297 (N_14297,N_13412,N_13769);
or U14298 (N_14298,N_13642,N_13475);
nor U14299 (N_14299,N_13896,N_13502);
nor U14300 (N_14300,N_13816,N_13429);
or U14301 (N_14301,N_13263,N_13879);
nand U14302 (N_14302,N_13999,N_13258);
nor U14303 (N_14303,N_13164,N_13796);
xor U14304 (N_14304,N_13678,N_13921);
nor U14305 (N_14305,N_13247,N_13117);
or U14306 (N_14306,N_13665,N_13159);
nand U14307 (N_14307,N_13979,N_13386);
nor U14308 (N_14308,N_13186,N_13694);
nor U14309 (N_14309,N_13611,N_13284);
and U14310 (N_14310,N_13949,N_13819);
or U14311 (N_14311,N_13515,N_13153);
nand U14312 (N_14312,N_13878,N_13958);
and U14313 (N_14313,N_13669,N_13096);
xnor U14314 (N_14314,N_13029,N_13037);
nand U14315 (N_14315,N_13403,N_13955);
or U14316 (N_14316,N_13835,N_13943);
nand U14317 (N_14317,N_13130,N_13554);
nor U14318 (N_14318,N_13270,N_13727);
nand U14319 (N_14319,N_13659,N_13052);
and U14320 (N_14320,N_13553,N_13134);
or U14321 (N_14321,N_13195,N_13738);
nor U14322 (N_14322,N_13259,N_13740);
xor U14323 (N_14323,N_13850,N_13241);
nor U14324 (N_14324,N_13289,N_13373);
or U14325 (N_14325,N_13048,N_13197);
nor U14326 (N_14326,N_13361,N_13998);
or U14327 (N_14327,N_13109,N_13505);
xnor U14328 (N_14328,N_13444,N_13736);
or U14329 (N_14329,N_13120,N_13025);
or U14330 (N_14330,N_13185,N_13281);
nand U14331 (N_14331,N_13944,N_13660);
or U14332 (N_14332,N_13621,N_13725);
or U14333 (N_14333,N_13139,N_13060);
or U14334 (N_14334,N_13443,N_13726);
or U14335 (N_14335,N_13889,N_13292);
xnor U14336 (N_14336,N_13903,N_13751);
and U14337 (N_14337,N_13709,N_13875);
or U14338 (N_14338,N_13950,N_13046);
and U14339 (N_14339,N_13368,N_13537);
nand U14340 (N_14340,N_13601,N_13334);
nand U14341 (N_14341,N_13687,N_13408);
or U14342 (N_14342,N_13522,N_13279);
or U14343 (N_14343,N_13269,N_13296);
and U14344 (N_14344,N_13544,N_13362);
and U14345 (N_14345,N_13777,N_13514);
nand U14346 (N_14346,N_13552,N_13434);
nor U14347 (N_14347,N_13834,N_13391);
or U14348 (N_14348,N_13121,N_13784);
or U14349 (N_14349,N_13549,N_13210);
nor U14350 (N_14350,N_13432,N_13168);
or U14351 (N_14351,N_13454,N_13813);
nor U14352 (N_14352,N_13229,N_13520);
nor U14353 (N_14353,N_13790,N_13538);
nand U14354 (N_14354,N_13759,N_13922);
nor U14355 (N_14355,N_13627,N_13572);
nor U14356 (N_14356,N_13926,N_13706);
and U14357 (N_14357,N_13842,N_13266);
nand U14358 (N_14358,N_13348,N_13671);
and U14359 (N_14359,N_13994,N_13810);
or U14360 (N_14360,N_13415,N_13952);
nor U14361 (N_14361,N_13942,N_13076);
nand U14362 (N_14362,N_13465,N_13066);
nand U14363 (N_14363,N_13080,N_13260);
nand U14364 (N_14364,N_13182,N_13141);
xnor U14365 (N_14365,N_13435,N_13372);
nand U14366 (N_14366,N_13984,N_13208);
and U14367 (N_14367,N_13874,N_13250);
and U14368 (N_14368,N_13165,N_13653);
xnor U14369 (N_14369,N_13118,N_13902);
and U14370 (N_14370,N_13330,N_13650);
xor U14371 (N_14371,N_13778,N_13754);
nor U14372 (N_14372,N_13085,N_13757);
or U14373 (N_14373,N_13624,N_13196);
or U14374 (N_14374,N_13457,N_13927);
or U14375 (N_14375,N_13861,N_13264);
or U14376 (N_14376,N_13735,N_13511);
xor U14377 (N_14377,N_13543,N_13512);
or U14378 (N_14378,N_13873,N_13888);
and U14379 (N_14379,N_13823,N_13499);
and U14380 (N_14380,N_13322,N_13848);
nor U14381 (N_14381,N_13507,N_13854);
nor U14382 (N_14382,N_13655,N_13696);
nand U14383 (N_14383,N_13906,N_13034);
and U14384 (N_14384,N_13974,N_13809);
or U14385 (N_14385,N_13909,N_13346);
and U14386 (N_14386,N_13357,N_13127);
nand U14387 (N_14387,N_13397,N_13501);
or U14388 (N_14388,N_13760,N_13174);
and U14389 (N_14389,N_13017,N_13375);
and U14390 (N_14390,N_13610,N_13449);
or U14391 (N_14391,N_13172,N_13094);
or U14392 (N_14392,N_13771,N_13244);
nand U14393 (N_14393,N_13287,N_13055);
or U14394 (N_14394,N_13744,N_13439);
nor U14395 (N_14395,N_13320,N_13116);
xor U14396 (N_14396,N_13600,N_13527);
and U14397 (N_14397,N_13951,N_13081);
or U14398 (N_14398,N_13095,N_13252);
nand U14399 (N_14399,N_13865,N_13086);
xnor U14400 (N_14400,N_13728,N_13731);
and U14401 (N_14401,N_13768,N_13620);
or U14402 (N_14402,N_13723,N_13815);
nand U14403 (N_14403,N_13084,N_13425);
or U14404 (N_14404,N_13451,N_13493);
or U14405 (N_14405,N_13613,N_13626);
nand U14406 (N_14406,N_13433,N_13392);
or U14407 (N_14407,N_13651,N_13630);
or U14408 (N_14408,N_13288,N_13594);
xor U14409 (N_14409,N_13079,N_13747);
xor U14410 (N_14410,N_13145,N_13091);
or U14411 (N_14411,N_13593,N_13192);
nand U14412 (N_14412,N_13606,N_13710);
nor U14413 (N_14413,N_13559,N_13913);
and U14414 (N_14414,N_13948,N_13887);
and U14415 (N_14415,N_13812,N_13634);
nand U14416 (N_14416,N_13198,N_13394);
nand U14417 (N_14417,N_13932,N_13011);
nand U14418 (N_14418,N_13864,N_13531);
or U14419 (N_14419,N_13547,N_13253);
nor U14420 (N_14420,N_13870,N_13885);
nand U14421 (N_14421,N_13717,N_13215);
or U14422 (N_14422,N_13737,N_13020);
nand U14423 (N_14423,N_13886,N_13242);
nor U14424 (N_14424,N_13311,N_13558);
nor U14425 (N_14425,N_13573,N_13150);
nand U14426 (N_14426,N_13114,N_13752);
nor U14427 (N_14427,N_13822,N_13405);
nand U14428 (N_14428,N_13175,N_13169);
nor U14429 (N_14429,N_13404,N_13097);
nand U14430 (N_14430,N_13212,N_13649);
nand U14431 (N_14431,N_13954,N_13021);
or U14432 (N_14432,N_13577,N_13176);
or U14433 (N_14433,N_13716,N_13345);
or U14434 (N_14434,N_13370,N_13718);
and U14435 (N_14435,N_13897,N_13211);
and U14436 (N_14436,N_13557,N_13414);
nor U14437 (N_14437,N_13712,N_13868);
and U14438 (N_14438,N_13990,N_13042);
nor U14439 (N_14439,N_13014,N_13049);
xnor U14440 (N_14440,N_13315,N_13604);
xnor U14441 (N_14441,N_13753,N_13101);
or U14442 (N_14442,N_13677,N_13082);
and U14443 (N_14443,N_13811,N_13912);
or U14444 (N_14444,N_13560,N_13280);
xor U14445 (N_14445,N_13797,N_13018);
or U14446 (N_14446,N_13297,N_13592);
and U14447 (N_14447,N_13915,N_13290);
nand U14448 (N_14448,N_13067,N_13846);
and U14449 (N_14449,N_13107,N_13108);
nand U14450 (N_14450,N_13144,N_13256);
nand U14451 (N_14451,N_13715,N_13295);
nor U14452 (N_14452,N_13683,N_13494);
xor U14453 (N_14453,N_13069,N_13685);
nor U14454 (N_14454,N_13301,N_13890);
and U14455 (N_14455,N_13571,N_13636);
and U14456 (N_14456,N_13993,N_13154);
or U14457 (N_14457,N_13200,N_13826);
nor U14458 (N_14458,N_13596,N_13359);
or U14459 (N_14459,N_13147,N_13832);
and U14460 (N_14460,N_13545,N_13615);
or U14461 (N_14461,N_13225,N_13806);
nand U14462 (N_14462,N_13820,N_13570);
nor U14463 (N_14463,N_13618,N_13629);
xnor U14464 (N_14464,N_13654,N_13251);
xnor U14465 (N_14465,N_13193,N_13721);
and U14466 (N_14466,N_13713,N_13142);
or U14467 (N_14467,N_13023,N_13087);
nor U14468 (N_14468,N_13137,N_13847);
and U14469 (N_14469,N_13278,N_13702);
nor U14470 (N_14470,N_13566,N_13548);
nand U14471 (N_14471,N_13585,N_13619);
nand U14472 (N_14472,N_13331,N_13043);
or U14473 (N_14473,N_13497,N_13285);
or U14474 (N_14474,N_13319,N_13351);
or U14475 (N_14475,N_13031,N_13925);
xor U14476 (N_14476,N_13972,N_13004);
nand U14477 (N_14477,N_13268,N_13488);
xor U14478 (N_14478,N_13227,N_13399);
nor U14479 (N_14479,N_13306,N_13900);
or U14480 (N_14480,N_13093,N_13807);
nor U14481 (N_14481,N_13342,N_13339);
and U14482 (N_14482,N_13939,N_13609);
and U14483 (N_14483,N_13525,N_13803);
nor U14484 (N_14484,N_13920,N_13360);
nor U14485 (N_14485,N_13246,N_13689);
and U14486 (N_14486,N_13960,N_13914);
and U14487 (N_14487,N_13231,N_13283);
xnor U14488 (N_14488,N_13521,N_13388);
or U14489 (N_14489,N_13929,N_13661);
nand U14490 (N_14490,N_13161,N_13038);
nor U14491 (N_14491,N_13413,N_13265);
nor U14492 (N_14492,N_13584,N_13202);
nand U14493 (N_14493,N_13015,N_13074);
nand U14494 (N_14494,N_13679,N_13396);
nand U14495 (N_14495,N_13110,N_13395);
nand U14496 (N_14496,N_13855,N_13000);
nor U14497 (N_14497,N_13128,N_13064);
nand U14498 (N_14498,N_13867,N_13612);
nand U14499 (N_14499,N_13924,N_13983);
xnor U14500 (N_14500,N_13208,N_13766);
nor U14501 (N_14501,N_13453,N_13267);
or U14502 (N_14502,N_13275,N_13866);
xor U14503 (N_14503,N_13806,N_13538);
xor U14504 (N_14504,N_13986,N_13539);
nand U14505 (N_14505,N_13961,N_13336);
nor U14506 (N_14506,N_13302,N_13908);
and U14507 (N_14507,N_13399,N_13949);
or U14508 (N_14508,N_13577,N_13535);
or U14509 (N_14509,N_13793,N_13505);
xor U14510 (N_14510,N_13611,N_13772);
nand U14511 (N_14511,N_13004,N_13541);
and U14512 (N_14512,N_13227,N_13162);
and U14513 (N_14513,N_13569,N_13898);
and U14514 (N_14514,N_13262,N_13252);
and U14515 (N_14515,N_13501,N_13417);
nor U14516 (N_14516,N_13338,N_13183);
or U14517 (N_14517,N_13782,N_13267);
or U14518 (N_14518,N_13476,N_13215);
or U14519 (N_14519,N_13025,N_13534);
nor U14520 (N_14520,N_13729,N_13187);
xnor U14521 (N_14521,N_13564,N_13579);
nand U14522 (N_14522,N_13620,N_13722);
xor U14523 (N_14523,N_13665,N_13842);
nor U14524 (N_14524,N_13305,N_13978);
and U14525 (N_14525,N_13060,N_13600);
and U14526 (N_14526,N_13930,N_13102);
nand U14527 (N_14527,N_13751,N_13457);
and U14528 (N_14528,N_13987,N_13037);
and U14529 (N_14529,N_13572,N_13426);
nand U14530 (N_14530,N_13503,N_13279);
nand U14531 (N_14531,N_13267,N_13389);
nand U14532 (N_14532,N_13606,N_13456);
and U14533 (N_14533,N_13107,N_13113);
nor U14534 (N_14534,N_13577,N_13326);
xnor U14535 (N_14535,N_13199,N_13841);
and U14536 (N_14536,N_13825,N_13354);
and U14537 (N_14537,N_13382,N_13284);
nor U14538 (N_14538,N_13730,N_13435);
or U14539 (N_14539,N_13602,N_13259);
and U14540 (N_14540,N_13452,N_13202);
nor U14541 (N_14541,N_13384,N_13822);
nor U14542 (N_14542,N_13756,N_13877);
nand U14543 (N_14543,N_13887,N_13858);
nand U14544 (N_14544,N_13645,N_13924);
nand U14545 (N_14545,N_13927,N_13746);
nor U14546 (N_14546,N_13999,N_13231);
nand U14547 (N_14547,N_13120,N_13419);
nor U14548 (N_14548,N_13300,N_13311);
and U14549 (N_14549,N_13974,N_13595);
nor U14550 (N_14550,N_13354,N_13174);
nor U14551 (N_14551,N_13578,N_13010);
nor U14552 (N_14552,N_13610,N_13006);
or U14553 (N_14553,N_13849,N_13396);
nor U14554 (N_14554,N_13561,N_13811);
xnor U14555 (N_14555,N_13460,N_13590);
nand U14556 (N_14556,N_13776,N_13232);
or U14557 (N_14557,N_13572,N_13093);
nor U14558 (N_14558,N_13337,N_13242);
xor U14559 (N_14559,N_13878,N_13391);
nor U14560 (N_14560,N_13358,N_13415);
nand U14561 (N_14561,N_13221,N_13897);
xnor U14562 (N_14562,N_13377,N_13837);
nand U14563 (N_14563,N_13979,N_13596);
and U14564 (N_14564,N_13970,N_13322);
nand U14565 (N_14565,N_13016,N_13101);
or U14566 (N_14566,N_13967,N_13424);
and U14567 (N_14567,N_13340,N_13201);
or U14568 (N_14568,N_13728,N_13862);
nand U14569 (N_14569,N_13951,N_13334);
nor U14570 (N_14570,N_13383,N_13547);
and U14571 (N_14571,N_13358,N_13396);
and U14572 (N_14572,N_13709,N_13935);
and U14573 (N_14573,N_13921,N_13109);
nand U14574 (N_14574,N_13067,N_13028);
xor U14575 (N_14575,N_13060,N_13870);
nand U14576 (N_14576,N_13927,N_13600);
or U14577 (N_14577,N_13621,N_13957);
nor U14578 (N_14578,N_13574,N_13192);
or U14579 (N_14579,N_13160,N_13249);
nand U14580 (N_14580,N_13355,N_13860);
nand U14581 (N_14581,N_13842,N_13896);
nand U14582 (N_14582,N_13546,N_13788);
and U14583 (N_14583,N_13083,N_13632);
nor U14584 (N_14584,N_13299,N_13900);
and U14585 (N_14585,N_13890,N_13400);
and U14586 (N_14586,N_13506,N_13534);
nor U14587 (N_14587,N_13694,N_13796);
and U14588 (N_14588,N_13967,N_13723);
nor U14589 (N_14589,N_13321,N_13016);
and U14590 (N_14590,N_13052,N_13703);
xor U14591 (N_14591,N_13009,N_13851);
nand U14592 (N_14592,N_13370,N_13616);
nor U14593 (N_14593,N_13114,N_13492);
nand U14594 (N_14594,N_13142,N_13831);
nand U14595 (N_14595,N_13091,N_13096);
nor U14596 (N_14596,N_13144,N_13435);
or U14597 (N_14597,N_13785,N_13965);
nand U14598 (N_14598,N_13828,N_13744);
and U14599 (N_14599,N_13495,N_13112);
nand U14600 (N_14600,N_13925,N_13811);
or U14601 (N_14601,N_13338,N_13875);
and U14602 (N_14602,N_13066,N_13897);
or U14603 (N_14603,N_13847,N_13396);
xnor U14604 (N_14604,N_13856,N_13880);
nor U14605 (N_14605,N_13809,N_13382);
and U14606 (N_14606,N_13302,N_13744);
nor U14607 (N_14607,N_13710,N_13498);
nand U14608 (N_14608,N_13113,N_13592);
nand U14609 (N_14609,N_13282,N_13493);
nor U14610 (N_14610,N_13826,N_13255);
nor U14611 (N_14611,N_13854,N_13262);
nand U14612 (N_14612,N_13459,N_13308);
xor U14613 (N_14613,N_13576,N_13350);
or U14614 (N_14614,N_13302,N_13415);
and U14615 (N_14615,N_13573,N_13474);
or U14616 (N_14616,N_13056,N_13893);
and U14617 (N_14617,N_13678,N_13474);
nand U14618 (N_14618,N_13369,N_13467);
and U14619 (N_14619,N_13092,N_13961);
nor U14620 (N_14620,N_13721,N_13940);
nand U14621 (N_14621,N_13262,N_13954);
or U14622 (N_14622,N_13762,N_13003);
nand U14623 (N_14623,N_13786,N_13397);
nand U14624 (N_14624,N_13016,N_13561);
nand U14625 (N_14625,N_13405,N_13185);
and U14626 (N_14626,N_13497,N_13042);
nand U14627 (N_14627,N_13173,N_13061);
or U14628 (N_14628,N_13176,N_13118);
nor U14629 (N_14629,N_13413,N_13631);
nor U14630 (N_14630,N_13718,N_13198);
nor U14631 (N_14631,N_13902,N_13437);
nand U14632 (N_14632,N_13036,N_13069);
and U14633 (N_14633,N_13333,N_13019);
nor U14634 (N_14634,N_13125,N_13065);
or U14635 (N_14635,N_13275,N_13407);
nor U14636 (N_14636,N_13858,N_13376);
and U14637 (N_14637,N_13659,N_13012);
nor U14638 (N_14638,N_13812,N_13407);
and U14639 (N_14639,N_13757,N_13061);
nor U14640 (N_14640,N_13220,N_13891);
nor U14641 (N_14641,N_13819,N_13774);
nor U14642 (N_14642,N_13029,N_13595);
and U14643 (N_14643,N_13608,N_13001);
or U14644 (N_14644,N_13286,N_13805);
or U14645 (N_14645,N_13615,N_13756);
and U14646 (N_14646,N_13212,N_13500);
or U14647 (N_14647,N_13766,N_13184);
xnor U14648 (N_14648,N_13710,N_13131);
nand U14649 (N_14649,N_13972,N_13897);
or U14650 (N_14650,N_13678,N_13844);
nand U14651 (N_14651,N_13101,N_13500);
and U14652 (N_14652,N_13643,N_13617);
xnor U14653 (N_14653,N_13049,N_13971);
or U14654 (N_14654,N_13242,N_13530);
nand U14655 (N_14655,N_13304,N_13648);
nor U14656 (N_14656,N_13858,N_13628);
nand U14657 (N_14657,N_13588,N_13603);
and U14658 (N_14658,N_13735,N_13039);
or U14659 (N_14659,N_13356,N_13218);
or U14660 (N_14660,N_13452,N_13305);
and U14661 (N_14661,N_13781,N_13046);
nand U14662 (N_14662,N_13596,N_13463);
nor U14663 (N_14663,N_13830,N_13407);
nand U14664 (N_14664,N_13524,N_13646);
and U14665 (N_14665,N_13134,N_13130);
or U14666 (N_14666,N_13123,N_13087);
and U14667 (N_14667,N_13397,N_13537);
nand U14668 (N_14668,N_13688,N_13969);
or U14669 (N_14669,N_13010,N_13811);
and U14670 (N_14670,N_13019,N_13746);
nor U14671 (N_14671,N_13512,N_13748);
nand U14672 (N_14672,N_13462,N_13126);
nand U14673 (N_14673,N_13842,N_13595);
nand U14674 (N_14674,N_13578,N_13782);
and U14675 (N_14675,N_13177,N_13211);
nor U14676 (N_14676,N_13479,N_13012);
and U14677 (N_14677,N_13438,N_13792);
and U14678 (N_14678,N_13010,N_13655);
nand U14679 (N_14679,N_13808,N_13417);
nand U14680 (N_14680,N_13653,N_13361);
or U14681 (N_14681,N_13328,N_13714);
or U14682 (N_14682,N_13420,N_13564);
and U14683 (N_14683,N_13157,N_13618);
nor U14684 (N_14684,N_13942,N_13124);
or U14685 (N_14685,N_13588,N_13411);
or U14686 (N_14686,N_13090,N_13392);
and U14687 (N_14687,N_13671,N_13833);
nor U14688 (N_14688,N_13125,N_13355);
nand U14689 (N_14689,N_13755,N_13910);
or U14690 (N_14690,N_13217,N_13298);
and U14691 (N_14691,N_13534,N_13829);
or U14692 (N_14692,N_13129,N_13044);
nor U14693 (N_14693,N_13238,N_13912);
and U14694 (N_14694,N_13554,N_13858);
or U14695 (N_14695,N_13909,N_13577);
nand U14696 (N_14696,N_13357,N_13598);
nor U14697 (N_14697,N_13782,N_13550);
nor U14698 (N_14698,N_13965,N_13841);
or U14699 (N_14699,N_13115,N_13560);
or U14700 (N_14700,N_13641,N_13420);
nand U14701 (N_14701,N_13459,N_13010);
and U14702 (N_14702,N_13429,N_13238);
or U14703 (N_14703,N_13995,N_13887);
nand U14704 (N_14704,N_13560,N_13427);
xor U14705 (N_14705,N_13168,N_13099);
or U14706 (N_14706,N_13174,N_13318);
or U14707 (N_14707,N_13821,N_13516);
nand U14708 (N_14708,N_13488,N_13312);
nor U14709 (N_14709,N_13127,N_13593);
or U14710 (N_14710,N_13602,N_13873);
nor U14711 (N_14711,N_13739,N_13427);
nor U14712 (N_14712,N_13350,N_13393);
or U14713 (N_14713,N_13753,N_13656);
nand U14714 (N_14714,N_13731,N_13921);
nand U14715 (N_14715,N_13544,N_13117);
and U14716 (N_14716,N_13301,N_13810);
nor U14717 (N_14717,N_13049,N_13482);
and U14718 (N_14718,N_13571,N_13397);
xor U14719 (N_14719,N_13618,N_13159);
nand U14720 (N_14720,N_13956,N_13027);
nor U14721 (N_14721,N_13982,N_13285);
nand U14722 (N_14722,N_13621,N_13293);
or U14723 (N_14723,N_13459,N_13073);
nor U14724 (N_14724,N_13691,N_13005);
nand U14725 (N_14725,N_13695,N_13317);
nand U14726 (N_14726,N_13289,N_13217);
nor U14727 (N_14727,N_13006,N_13578);
and U14728 (N_14728,N_13420,N_13740);
xnor U14729 (N_14729,N_13328,N_13162);
or U14730 (N_14730,N_13686,N_13563);
nand U14731 (N_14731,N_13809,N_13264);
nand U14732 (N_14732,N_13831,N_13736);
xor U14733 (N_14733,N_13966,N_13950);
nor U14734 (N_14734,N_13201,N_13944);
nand U14735 (N_14735,N_13985,N_13802);
or U14736 (N_14736,N_13851,N_13828);
xnor U14737 (N_14737,N_13393,N_13905);
nor U14738 (N_14738,N_13288,N_13743);
nor U14739 (N_14739,N_13706,N_13666);
and U14740 (N_14740,N_13019,N_13126);
and U14741 (N_14741,N_13158,N_13798);
and U14742 (N_14742,N_13188,N_13919);
or U14743 (N_14743,N_13010,N_13314);
nor U14744 (N_14744,N_13869,N_13902);
nand U14745 (N_14745,N_13177,N_13587);
or U14746 (N_14746,N_13815,N_13282);
or U14747 (N_14747,N_13287,N_13298);
and U14748 (N_14748,N_13937,N_13910);
nand U14749 (N_14749,N_13114,N_13429);
nand U14750 (N_14750,N_13434,N_13439);
or U14751 (N_14751,N_13758,N_13701);
or U14752 (N_14752,N_13950,N_13829);
nor U14753 (N_14753,N_13774,N_13238);
nand U14754 (N_14754,N_13732,N_13904);
nand U14755 (N_14755,N_13198,N_13471);
and U14756 (N_14756,N_13664,N_13711);
and U14757 (N_14757,N_13551,N_13124);
nor U14758 (N_14758,N_13384,N_13438);
or U14759 (N_14759,N_13326,N_13295);
nand U14760 (N_14760,N_13853,N_13030);
or U14761 (N_14761,N_13824,N_13621);
and U14762 (N_14762,N_13733,N_13364);
nand U14763 (N_14763,N_13273,N_13461);
or U14764 (N_14764,N_13415,N_13323);
or U14765 (N_14765,N_13951,N_13146);
and U14766 (N_14766,N_13257,N_13073);
and U14767 (N_14767,N_13530,N_13164);
and U14768 (N_14768,N_13240,N_13882);
or U14769 (N_14769,N_13277,N_13135);
nand U14770 (N_14770,N_13613,N_13955);
or U14771 (N_14771,N_13540,N_13778);
nor U14772 (N_14772,N_13818,N_13197);
and U14773 (N_14773,N_13336,N_13325);
xor U14774 (N_14774,N_13467,N_13205);
nand U14775 (N_14775,N_13326,N_13461);
nor U14776 (N_14776,N_13025,N_13702);
nand U14777 (N_14777,N_13468,N_13108);
and U14778 (N_14778,N_13307,N_13454);
xnor U14779 (N_14779,N_13032,N_13413);
and U14780 (N_14780,N_13249,N_13539);
nor U14781 (N_14781,N_13596,N_13483);
nand U14782 (N_14782,N_13588,N_13824);
nor U14783 (N_14783,N_13008,N_13447);
nor U14784 (N_14784,N_13075,N_13817);
nand U14785 (N_14785,N_13510,N_13946);
nand U14786 (N_14786,N_13412,N_13556);
and U14787 (N_14787,N_13523,N_13253);
and U14788 (N_14788,N_13265,N_13951);
and U14789 (N_14789,N_13157,N_13870);
and U14790 (N_14790,N_13102,N_13356);
nor U14791 (N_14791,N_13564,N_13266);
xor U14792 (N_14792,N_13863,N_13526);
xnor U14793 (N_14793,N_13329,N_13550);
xnor U14794 (N_14794,N_13678,N_13620);
or U14795 (N_14795,N_13491,N_13649);
and U14796 (N_14796,N_13974,N_13462);
and U14797 (N_14797,N_13699,N_13273);
or U14798 (N_14798,N_13365,N_13142);
nor U14799 (N_14799,N_13526,N_13176);
or U14800 (N_14800,N_13766,N_13348);
nor U14801 (N_14801,N_13276,N_13422);
nor U14802 (N_14802,N_13268,N_13583);
nand U14803 (N_14803,N_13828,N_13677);
and U14804 (N_14804,N_13589,N_13288);
xor U14805 (N_14805,N_13971,N_13259);
or U14806 (N_14806,N_13488,N_13964);
nor U14807 (N_14807,N_13172,N_13282);
and U14808 (N_14808,N_13010,N_13775);
nand U14809 (N_14809,N_13325,N_13278);
or U14810 (N_14810,N_13560,N_13100);
and U14811 (N_14811,N_13398,N_13943);
and U14812 (N_14812,N_13162,N_13819);
and U14813 (N_14813,N_13590,N_13300);
and U14814 (N_14814,N_13874,N_13263);
nand U14815 (N_14815,N_13973,N_13382);
or U14816 (N_14816,N_13918,N_13399);
nor U14817 (N_14817,N_13201,N_13874);
and U14818 (N_14818,N_13584,N_13750);
nand U14819 (N_14819,N_13722,N_13579);
and U14820 (N_14820,N_13343,N_13295);
nand U14821 (N_14821,N_13067,N_13850);
nor U14822 (N_14822,N_13303,N_13243);
or U14823 (N_14823,N_13335,N_13962);
and U14824 (N_14824,N_13037,N_13481);
xnor U14825 (N_14825,N_13500,N_13710);
nand U14826 (N_14826,N_13739,N_13212);
and U14827 (N_14827,N_13897,N_13317);
or U14828 (N_14828,N_13449,N_13678);
nand U14829 (N_14829,N_13532,N_13650);
nand U14830 (N_14830,N_13305,N_13630);
nand U14831 (N_14831,N_13876,N_13604);
and U14832 (N_14832,N_13884,N_13313);
and U14833 (N_14833,N_13645,N_13289);
nand U14834 (N_14834,N_13831,N_13694);
nor U14835 (N_14835,N_13713,N_13705);
or U14836 (N_14836,N_13431,N_13421);
nor U14837 (N_14837,N_13595,N_13158);
nand U14838 (N_14838,N_13961,N_13881);
nand U14839 (N_14839,N_13277,N_13088);
nor U14840 (N_14840,N_13704,N_13218);
nand U14841 (N_14841,N_13167,N_13785);
xnor U14842 (N_14842,N_13373,N_13588);
or U14843 (N_14843,N_13485,N_13904);
or U14844 (N_14844,N_13301,N_13892);
nand U14845 (N_14845,N_13589,N_13187);
xnor U14846 (N_14846,N_13943,N_13711);
xor U14847 (N_14847,N_13545,N_13071);
and U14848 (N_14848,N_13619,N_13499);
nor U14849 (N_14849,N_13738,N_13847);
nand U14850 (N_14850,N_13874,N_13483);
nand U14851 (N_14851,N_13482,N_13112);
or U14852 (N_14852,N_13459,N_13346);
nor U14853 (N_14853,N_13776,N_13589);
nor U14854 (N_14854,N_13350,N_13672);
nand U14855 (N_14855,N_13382,N_13636);
or U14856 (N_14856,N_13568,N_13531);
xor U14857 (N_14857,N_13362,N_13120);
and U14858 (N_14858,N_13670,N_13520);
nor U14859 (N_14859,N_13925,N_13104);
or U14860 (N_14860,N_13207,N_13430);
nor U14861 (N_14861,N_13606,N_13414);
nor U14862 (N_14862,N_13536,N_13792);
and U14863 (N_14863,N_13734,N_13422);
nor U14864 (N_14864,N_13941,N_13274);
nor U14865 (N_14865,N_13112,N_13955);
or U14866 (N_14866,N_13884,N_13995);
xnor U14867 (N_14867,N_13374,N_13525);
and U14868 (N_14868,N_13320,N_13865);
or U14869 (N_14869,N_13119,N_13454);
nor U14870 (N_14870,N_13654,N_13971);
or U14871 (N_14871,N_13742,N_13410);
or U14872 (N_14872,N_13710,N_13646);
nand U14873 (N_14873,N_13138,N_13634);
xor U14874 (N_14874,N_13592,N_13295);
or U14875 (N_14875,N_13719,N_13207);
and U14876 (N_14876,N_13378,N_13696);
or U14877 (N_14877,N_13732,N_13647);
nor U14878 (N_14878,N_13078,N_13147);
or U14879 (N_14879,N_13329,N_13758);
nor U14880 (N_14880,N_13703,N_13777);
nand U14881 (N_14881,N_13334,N_13992);
and U14882 (N_14882,N_13264,N_13156);
or U14883 (N_14883,N_13057,N_13316);
nand U14884 (N_14884,N_13395,N_13837);
or U14885 (N_14885,N_13031,N_13261);
and U14886 (N_14886,N_13482,N_13686);
and U14887 (N_14887,N_13060,N_13692);
nand U14888 (N_14888,N_13353,N_13355);
nor U14889 (N_14889,N_13929,N_13321);
nand U14890 (N_14890,N_13198,N_13637);
or U14891 (N_14891,N_13238,N_13946);
and U14892 (N_14892,N_13901,N_13435);
nor U14893 (N_14893,N_13097,N_13494);
nand U14894 (N_14894,N_13330,N_13889);
nand U14895 (N_14895,N_13390,N_13002);
and U14896 (N_14896,N_13916,N_13400);
or U14897 (N_14897,N_13451,N_13568);
or U14898 (N_14898,N_13584,N_13662);
and U14899 (N_14899,N_13018,N_13469);
or U14900 (N_14900,N_13498,N_13784);
nand U14901 (N_14901,N_13232,N_13029);
and U14902 (N_14902,N_13830,N_13760);
nand U14903 (N_14903,N_13727,N_13125);
or U14904 (N_14904,N_13958,N_13662);
nor U14905 (N_14905,N_13122,N_13569);
or U14906 (N_14906,N_13107,N_13011);
nor U14907 (N_14907,N_13329,N_13827);
nor U14908 (N_14908,N_13981,N_13036);
nor U14909 (N_14909,N_13331,N_13838);
and U14910 (N_14910,N_13225,N_13088);
or U14911 (N_14911,N_13957,N_13762);
and U14912 (N_14912,N_13898,N_13945);
or U14913 (N_14913,N_13401,N_13139);
and U14914 (N_14914,N_13809,N_13419);
nand U14915 (N_14915,N_13251,N_13124);
nand U14916 (N_14916,N_13656,N_13901);
and U14917 (N_14917,N_13350,N_13761);
nor U14918 (N_14918,N_13610,N_13014);
or U14919 (N_14919,N_13969,N_13475);
nand U14920 (N_14920,N_13051,N_13577);
or U14921 (N_14921,N_13677,N_13478);
nor U14922 (N_14922,N_13819,N_13990);
or U14923 (N_14923,N_13265,N_13203);
and U14924 (N_14924,N_13142,N_13289);
nor U14925 (N_14925,N_13440,N_13146);
nor U14926 (N_14926,N_13035,N_13127);
nor U14927 (N_14927,N_13804,N_13716);
nor U14928 (N_14928,N_13797,N_13923);
xnor U14929 (N_14929,N_13004,N_13167);
xnor U14930 (N_14930,N_13698,N_13097);
and U14931 (N_14931,N_13019,N_13723);
nor U14932 (N_14932,N_13771,N_13816);
and U14933 (N_14933,N_13410,N_13717);
or U14934 (N_14934,N_13613,N_13846);
nand U14935 (N_14935,N_13362,N_13366);
or U14936 (N_14936,N_13556,N_13434);
nor U14937 (N_14937,N_13917,N_13912);
and U14938 (N_14938,N_13870,N_13392);
nand U14939 (N_14939,N_13564,N_13719);
or U14940 (N_14940,N_13831,N_13155);
nand U14941 (N_14941,N_13212,N_13277);
or U14942 (N_14942,N_13561,N_13349);
or U14943 (N_14943,N_13240,N_13368);
nor U14944 (N_14944,N_13548,N_13147);
and U14945 (N_14945,N_13676,N_13832);
nand U14946 (N_14946,N_13803,N_13344);
and U14947 (N_14947,N_13781,N_13496);
and U14948 (N_14948,N_13176,N_13949);
nand U14949 (N_14949,N_13359,N_13360);
and U14950 (N_14950,N_13119,N_13477);
and U14951 (N_14951,N_13548,N_13987);
or U14952 (N_14952,N_13387,N_13629);
nand U14953 (N_14953,N_13240,N_13409);
and U14954 (N_14954,N_13561,N_13502);
nor U14955 (N_14955,N_13656,N_13984);
nand U14956 (N_14956,N_13179,N_13980);
or U14957 (N_14957,N_13948,N_13411);
or U14958 (N_14958,N_13328,N_13903);
xor U14959 (N_14959,N_13865,N_13404);
nand U14960 (N_14960,N_13451,N_13346);
nor U14961 (N_14961,N_13935,N_13677);
and U14962 (N_14962,N_13372,N_13733);
and U14963 (N_14963,N_13952,N_13991);
nand U14964 (N_14964,N_13724,N_13251);
nand U14965 (N_14965,N_13011,N_13094);
nor U14966 (N_14966,N_13174,N_13925);
nor U14967 (N_14967,N_13863,N_13481);
or U14968 (N_14968,N_13190,N_13129);
or U14969 (N_14969,N_13268,N_13698);
nor U14970 (N_14970,N_13480,N_13769);
nand U14971 (N_14971,N_13260,N_13831);
nor U14972 (N_14972,N_13904,N_13104);
or U14973 (N_14973,N_13756,N_13474);
and U14974 (N_14974,N_13451,N_13183);
and U14975 (N_14975,N_13924,N_13926);
nand U14976 (N_14976,N_13056,N_13841);
and U14977 (N_14977,N_13404,N_13103);
nor U14978 (N_14978,N_13355,N_13099);
or U14979 (N_14979,N_13064,N_13797);
nor U14980 (N_14980,N_13517,N_13867);
and U14981 (N_14981,N_13243,N_13020);
nor U14982 (N_14982,N_13243,N_13439);
or U14983 (N_14983,N_13412,N_13244);
xor U14984 (N_14984,N_13172,N_13653);
or U14985 (N_14985,N_13416,N_13216);
and U14986 (N_14986,N_13446,N_13718);
or U14987 (N_14987,N_13870,N_13330);
nor U14988 (N_14988,N_13575,N_13032);
nor U14989 (N_14989,N_13917,N_13864);
and U14990 (N_14990,N_13113,N_13233);
nor U14991 (N_14991,N_13603,N_13084);
and U14992 (N_14992,N_13929,N_13608);
and U14993 (N_14993,N_13738,N_13890);
or U14994 (N_14994,N_13036,N_13168);
xor U14995 (N_14995,N_13357,N_13592);
xnor U14996 (N_14996,N_13627,N_13140);
nand U14997 (N_14997,N_13687,N_13698);
xnor U14998 (N_14998,N_13047,N_13481);
or U14999 (N_14999,N_13214,N_13466);
nor UO_0 (O_0,N_14700,N_14927);
or UO_1 (O_1,N_14229,N_14337);
or UO_2 (O_2,N_14260,N_14887);
and UO_3 (O_3,N_14093,N_14864);
nor UO_4 (O_4,N_14424,N_14790);
nor UO_5 (O_5,N_14170,N_14781);
nor UO_6 (O_6,N_14101,N_14068);
and UO_7 (O_7,N_14282,N_14676);
and UO_8 (O_8,N_14694,N_14180);
or UO_9 (O_9,N_14262,N_14638);
and UO_10 (O_10,N_14690,N_14840);
or UO_11 (O_11,N_14920,N_14992);
or UO_12 (O_12,N_14867,N_14426);
and UO_13 (O_13,N_14963,N_14911);
nand UO_14 (O_14,N_14151,N_14332);
nand UO_15 (O_15,N_14258,N_14044);
or UO_16 (O_16,N_14739,N_14066);
nand UO_17 (O_17,N_14311,N_14361);
nand UO_18 (O_18,N_14748,N_14368);
and UO_19 (O_19,N_14327,N_14298);
nand UO_20 (O_20,N_14671,N_14320);
or UO_21 (O_21,N_14221,N_14344);
xor UO_22 (O_22,N_14423,N_14384);
or UO_23 (O_23,N_14073,N_14001);
or UO_24 (O_24,N_14412,N_14737);
nor UO_25 (O_25,N_14492,N_14787);
nor UO_26 (O_26,N_14405,N_14546);
nand UO_27 (O_27,N_14235,N_14427);
nor UO_28 (O_28,N_14554,N_14070);
xnor UO_29 (O_29,N_14286,N_14239);
and UO_30 (O_30,N_14242,N_14989);
nand UO_31 (O_31,N_14421,N_14633);
nand UO_32 (O_32,N_14226,N_14984);
nor UO_33 (O_33,N_14853,N_14662);
nor UO_34 (O_34,N_14884,N_14125);
or UO_35 (O_35,N_14827,N_14904);
and UO_36 (O_36,N_14977,N_14960);
nand UO_37 (O_37,N_14255,N_14205);
nor UO_38 (O_38,N_14744,N_14860);
xor UO_39 (O_39,N_14254,N_14461);
and UO_40 (O_40,N_14120,N_14331);
nand UO_41 (O_41,N_14196,N_14925);
nor UO_42 (O_42,N_14980,N_14348);
and UO_43 (O_43,N_14155,N_14617);
nand UO_44 (O_44,N_14576,N_14224);
nor UO_45 (O_45,N_14527,N_14306);
xor UO_46 (O_46,N_14782,N_14951);
nor UO_47 (O_47,N_14726,N_14789);
or UO_48 (O_48,N_14863,N_14571);
nand UO_49 (O_49,N_14000,N_14954);
nor UO_50 (O_50,N_14402,N_14702);
nor UO_51 (O_51,N_14483,N_14947);
or UO_52 (O_52,N_14683,N_14313);
nand UO_53 (O_53,N_14281,N_14914);
nand UO_54 (O_54,N_14241,N_14054);
or UO_55 (O_55,N_14187,N_14022);
and UO_56 (O_56,N_14006,N_14303);
or UO_57 (O_57,N_14552,N_14613);
and UO_58 (O_58,N_14708,N_14333);
xor UO_59 (O_59,N_14417,N_14654);
and UO_60 (O_60,N_14908,N_14463);
nor UO_61 (O_61,N_14341,N_14821);
or UO_62 (O_62,N_14641,N_14764);
and UO_63 (O_63,N_14563,N_14579);
nor UO_64 (O_64,N_14048,N_14682);
and UO_65 (O_65,N_14291,N_14635);
nor UO_66 (O_66,N_14026,N_14407);
or UO_67 (O_67,N_14362,N_14251);
and UO_68 (O_68,N_14450,N_14263);
or UO_69 (O_69,N_14288,N_14323);
or UO_70 (O_70,N_14144,N_14039);
and UO_71 (O_71,N_14050,N_14177);
or UO_72 (O_72,N_14439,N_14364);
and UO_73 (O_73,N_14592,N_14418);
nor UO_74 (O_74,N_14922,N_14406);
or UO_75 (O_75,N_14316,N_14334);
nand UO_76 (O_76,N_14266,N_14946);
nand UO_77 (O_77,N_14560,N_14043);
and UO_78 (O_78,N_14161,N_14674);
nor UO_79 (O_79,N_14959,N_14456);
nor UO_80 (O_80,N_14997,N_14668);
xnor UO_81 (O_81,N_14098,N_14888);
xnor UO_82 (O_82,N_14040,N_14141);
and UO_83 (O_83,N_14607,N_14097);
xnor UO_84 (O_84,N_14531,N_14422);
or UO_85 (O_85,N_14115,N_14698);
or UO_86 (O_86,N_14958,N_14970);
xnor UO_87 (O_87,N_14494,N_14627);
and UO_88 (O_88,N_14156,N_14113);
nor UO_89 (O_89,N_14523,N_14359);
nor UO_90 (O_90,N_14881,N_14695);
and UO_91 (O_91,N_14847,N_14755);
nor UO_92 (O_92,N_14515,N_14408);
nand UO_93 (O_93,N_14926,N_14498);
and UO_94 (O_94,N_14124,N_14248);
and UO_95 (O_95,N_14459,N_14064);
xnor UO_96 (O_96,N_14961,N_14176);
nor UO_97 (O_97,N_14645,N_14481);
and UO_98 (O_98,N_14893,N_14211);
nand UO_99 (O_99,N_14236,N_14256);
and UO_100 (O_100,N_14591,N_14479);
or UO_101 (O_101,N_14181,N_14317);
or UO_102 (O_102,N_14400,N_14559);
nor UO_103 (O_103,N_14716,N_14570);
xnor UO_104 (O_104,N_14106,N_14051);
or UO_105 (O_105,N_14091,N_14952);
nand UO_106 (O_106,N_14890,N_14660);
or UO_107 (O_107,N_14967,N_14469);
nor UO_108 (O_108,N_14019,N_14131);
or UO_109 (O_109,N_14257,N_14612);
nor UO_110 (O_110,N_14350,N_14185);
nand UO_111 (O_111,N_14453,N_14905);
nand UO_112 (O_112,N_14793,N_14939);
nand UO_113 (O_113,N_14058,N_14214);
nand UO_114 (O_114,N_14729,N_14856);
xor UO_115 (O_115,N_14548,N_14240);
nor UO_116 (O_116,N_14356,N_14688);
nor UO_117 (O_117,N_14514,N_14593);
or UO_118 (O_118,N_14347,N_14861);
and UO_119 (O_119,N_14501,N_14586);
xnor UO_120 (O_120,N_14604,N_14305);
nor UO_121 (O_121,N_14122,N_14495);
nor UO_122 (O_122,N_14965,N_14985);
nor UO_123 (O_123,N_14642,N_14990);
xor UO_124 (O_124,N_14105,N_14470);
nor UO_125 (O_125,N_14529,N_14711);
and UO_126 (O_126,N_14371,N_14778);
or UO_127 (O_127,N_14780,N_14833);
or UO_128 (O_128,N_14773,N_14705);
nor UO_129 (O_129,N_14901,N_14476);
or UO_130 (O_130,N_14249,N_14758);
or UO_131 (O_131,N_14072,N_14534);
and UO_132 (O_132,N_14330,N_14615);
xnor UO_133 (O_133,N_14455,N_14028);
and UO_134 (O_134,N_14216,N_14420);
nor UO_135 (O_135,N_14849,N_14810);
or UO_136 (O_136,N_14206,N_14493);
nor UO_137 (O_137,N_14971,N_14452);
xor UO_138 (O_138,N_14982,N_14981);
nor UO_139 (O_139,N_14968,N_14264);
or UO_140 (O_140,N_14973,N_14747);
nand UO_141 (O_141,N_14153,N_14460);
nor UO_142 (O_142,N_14880,N_14147);
and UO_143 (O_143,N_14616,N_14611);
nand UO_144 (O_144,N_14443,N_14500);
or UO_145 (O_145,N_14088,N_14843);
nand UO_146 (O_146,N_14274,N_14589);
or UO_147 (O_147,N_14474,N_14590);
nand UO_148 (O_148,N_14816,N_14772);
nand UO_149 (O_149,N_14724,N_14566);
nor UO_150 (O_150,N_14774,N_14133);
nor UO_151 (O_151,N_14065,N_14850);
and UO_152 (O_152,N_14142,N_14457);
or UO_153 (O_153,N_14536,N_14550);
nand UO_154 (O_154,N_14053,N_14511);
nor UO_155 (O_155,N_14677,N_14999);
and UO_156 (O_156,N_14983,N_14219);
and UO_157 (O_157,N_14626,N_14537);
or UO_158 (O_158,N_14857,N_14366);
nor UO_159 (O_159,N_14932,N_14987);
or UO_160 (O_160,N_14173,N_14814);
or UO_161 (O_161,N_14335,N_14369);
nand UO_162 (O_162,N_14631,N_14622);
and UO_163 (O_163,N_14841,N_14834);
nand UO_164 (O_164,N_14938,N_14375);
nand UO_165 (O_165,N_14329,N_14763);
nand UO_166 (O_166,N_14732,N_14564);
nand UO_167 (O_167,N_14004,N_14127);
nor UO_168 (O_168,N_14130,N_14381);
xnor UO_169 (O_169,N_14411,N_14409);
nand UO_170 (O_170,N_14831,N_14388);
or UO_171 (O_171,N_14447,N_14326);
and UO_172 (O_172,N_14033,N_14071);
nand UO_173 (O_173,N_14806,N_14906);
nand UO_174 (O_174,N_14038,N_14628);
and UO_175 (O_175,N_14035,N_14152);
or UO_176 (O_176,N_14165,N_14160);
or UO_177 (O_177,N_14619,N_14699);
or UO_178 (O_178,N_14049,N_14157);
and UO_179 (O_179,N_14745,N_14896);
or UO_180 (O_180,N_14618,N_14964);
nand UO_181 (O_181,N_14178,N_14055);
and UO_182 (O_182,N_14391,N_14753);
nor UO_183 (O_183,N_14605,N_14533);
nor UO_184 (O_184,N_14247,N_14458);
nand UO_185 (O_185,N_14302,N_14121);
and UO_186 (O_186,N_14136,N_14648);
nand UO_187 (O_187,N_14021,N_14786);
nor UO_188 (O_188,N_14697,N_14568);
or UO_189 (O_189,N_14309,N_14714);
or UO_190 (O_190,N_14653,N_14937);
and UO_191 (O_191,N_14410,N_14340);
nand UO_192 (O_192,N_14193,N_14034);
nor UO_193 (O_193,N_14791,N_14269);
nand UO_194 (O_194,N_14357,N_14355);
and UO_195 (O_195,N_14685,N_14974);
and UO_196 (O_196,N_14643,N_14110);
nand UO_197 (O_197,N_14882,N_14373);
nor UO_198 (O_198,N_14770,N_14942);
nand UO_199 (O_199,N_14567,N_14740);
nor UO_200 (O_200,N_14953,N_14525);
xor UO_201 (O_201,N_14112,N_14594);
or UO_202 (O_202,N_14454,N_14924);
xor UO_203 (O_203,N_14278,N_14299);
and UO_204 (O_204,N_14244,N_14132);
nor UO_205 (O_205,N_14077,N_14270);
xnor UO_206 (O_206,N_14923,N_14415);
or UO_207 (O_207,N_14885,N_14319);
nor UO_208 (O_208,N_14528,N_14602);
nor UO_209 (O_209,N_14150,N_14620);
and UO_210 (O_210,N_14217,N_14228);
nand UO_211 (O_211,N_14067,N_14488);
nand UO_212 (O_212,N_14203,N_14894);
or UO_213 (O_213,N_14099,N_14921);
xor UO_214 (O_214,N_14480,N_14765);
nor UO_215 (O_215,N_14489,N_14865);
or UO_216 (O_216,N_14762,N_14756);
or UO_217 (O_217,N_14032,N_14010);
nor UO_218 (O_218,N_14210,N_14741);
or UO_219 (O_219,N_14595,N_14749);
nor UO_220 (O_220,N_14596,N_14289);
or UO_221 (O_221,N_14015,N_14271);
nor UO_222 (O_222,N_14670,N_14587);
or UO_223 (O_223,N_14140,N_14213);
nand UO_224 (O_224,N_14875,N_14658);
nand UO_225 (O_225,N_14075,N_14636);
xnor UO_226 (O_226,N_14846,N_14553);
nor UO_227 (O_227,N_14541,N_14539);
xor UO_228 (O_228,N_14207,N_14730);
xor UO_229 (O_229,N_14295,N_14574);
and UO_230 (O_230,N_14601,N_14829);
nor UO_231 (O_231,N_14215,N_14855);
and UO_232 (O_232,N_14767,N_14222);
or UO_233 (O_233,N_14955,N_14374);
nand UO_234 (O_234,N_14832,N_14517);
or UO_235 (O_235,N_14376,N_14859);
and UO_236 (O_236,N_14159,N_14431);
and UO_237 (O_237,N_14813,N_14918);
nand UO_238 (O_238,N_14390,N_14315);
nor UO_239 (O_239,N_14365,N_14017);
and UO_240 (O_240,N_14530,N_14862);
or UO_241 (O_241,N_14839,N_14549);
nand UO_242 (O_242,N_14703,N_14046);
nor UO_243 (O_243,N_14118,N_14208);
and UO_244 (O_244,N_14647,N_14707);
or UO_245 (O_245,N_14759,N_14189);
nor UO_246 (O_246,N_14339,N_14569);
nand UO_247 (O_247,N_14891,N_14902);
and UO_248 (O_248,N_14092,N_14804);
nand UO_249 (O_249,N_14811,N_14148);
or UO_250 (O_250,N_14027,N_14524);
nor UO_251 (O_251,N_14975,N_14812);
nor UO_252 (O_252,N_14023,N_14087);
nor UO_253 (O_253,N_14752,N_14102);
and UO_254 (O_254,N_14499,N_14957);
or UO_255 (O_255,N_14830,N_14192);
and UO_256 (O_256,N_14950,N_14045);
nor UO_257 (O_257,N_14393,N_14387);
and UO_258 (O_258,N_14300,N_14598);
or UO_259 (O_259,N_14338,N_14792);
or UO_260 (O_260,N_14689,N_14684);
nor UO_261 (O_261,N_14581,N_14059);
nor UO_262 (O_262,N_14195,N_14910);
nor UO_263 (O_263,N_14292,N_14917);
or UO_264 (O_264,N_14029,N_14929);
or UO_265 (O_265,N_14675,N_14230);
nand UO_266 (O_266,N_14667,N_14915);
nor UO_267 (O_267,N_14279,N_14731);
xor UO_268 (O_268,N_14310,N_14808);
or UO_269 (O_269,N_14649,N_14284);
and UO_270 (O_270,N_14873,N_14652);
xor UO_271 (O_271,N_14232,N_14993);
nand UO_272 (O_272,N_14253,N_14526);
and UO_273 (O_273,N_14351,N_14487);
nand UO_274 (O_274,N_14809,N_14468);
nor UO_275 (O_275,N_14555,N_14686);
or UO_276 (O_276,N_14795,N_14640);
or UO_277 (O_277,N_14293,N_14512);
nand UO_278 (O_278,N_14135,N_14717);
or UO_279 (O_279,N_14720,N_14414);
and UO_280 (O_280,N_14265,N_14978);
xnor UO_281 (O_281,N_14532,N_14600);
and UO_282 (O_282,N_14430,N_14535);
nor UO_283 (O_283,N_14202,N_14883);
nor UO_284 (O_284,N_14389,N_14644);
or UO_285 (O_285,N_14183,N_14996);
and UO_286 (O_286,N_14014,N_14962);
or UO_287 (O_287,N_14941,N_14522);
nor UO_288 (O_288,N_14625,N_14261);
and UO_289 (O_289,N_14949,N_14324);
or UO_290 (O_290,N_14020,N_14785);
nor UO_291 (O_291,N_14584,N_14164);
and UO_292 (O_292,N_14505,N_14798);
xor UO_293 (O_293,N_14871,N_14743);
nand UO_294 (O_294,N_14346,N_14757);
nor UO_295 (O_295,N_14802,N_14507);
nor UO_296 (O_296,N_14353,N_14934);
or UO_297 (O_297,N_14047,N_14042);
nor UO_298 (O_298,N_14166,N_14945);
and UO_299 (O_299,N_14998,N_14462);
nand UO_300 (O_300,N_14307,N_14094);
and UO_301 (O_301,N_14428,N_14188);
and UO_302 (O_302,N_14002,N_14723);
xnor UO_303 (O_303,N_14931,N_14837);
or UO_304 (O_304,N_14234,N_14464);
and UO_305 (O_305,N_14624,N_14354);
nor UO_306 (O_306,N_14578,N_14966);
nand UO_307 (O_307,N_14396,N_14986);
nand UO_308 (O_308,N_14433,N_14725);
or UO_309 (O_309,N_14472,N_14370);
nand UO_310 (O_310,N_14486,N_14259);
nand UO_311 (O_311,N_14940,N_14991);
or UO_312 (O_312,N_14521,N_14637);
nor UO_313 (O_313,N_14672,N_14104);
or UO_314 (O_314,N_14083,N_14736);
or UO_315 (O_315,N_14441,N_14490);
and UO_316 (O_316,N_14403,N_14943);
and UO_317 (O_317,N_14687,N_14669);
nand UO_318 (O_318,N_14379,N_14169);
and UO_319 (O_319,N_14562,N_14444);
xnor UO_320 (O_320,N_14116,N_14972);
and UO_321 (O_321,N_14076,N_14588);
and UO_322 (O_322,N_14238,N_14416);
and UO_323 (O_323,N_14100,N_14976);
nand UO_324 (O_324,N_14434,N_14220);
nand UO_325 (O_325,N_14706,N_14162);
nand UO_326 (O_326,N_14886,N_14796);
or UO_327 (O_327,N_14629,N_14807);
nor UO_328 (O_328,N_14398,N_14079);
or UO_329 (O_329,N_14935,N_14466);
nand UO_330 (O_330,N_14143,N_14543);
nor UO_331 (O_331,N_14632,N_14138);
and UO_332 (O_332,N_14565,N_14691);
or UO_333 (O_333,N_14036,N_14769);
or UO_334 (O_334,N_14639,N_14056);
or UO_335 (O_335,N_14360,N_14727);
nor UO_336 (O_336,N_14037,N_14018);
and UO_337 (O_337,N_14614,N_14090);
xor UO_338 (O_338,N_14069,N_14382);
and UO_339 (O_339,N_14760,N_14776);
nand UO_340 (O_340,N_14503,N_14815);
nand UO_341 (O_341,N_14225,N_14820);
and UO_342 (O_342,N_14201,N_14465);
and UO_343 (O_343,N_14866,N_14606);
or UO_344 (O_344,N_14826,N_14003);
nand UO_345 (O_345,N_14710,N_14979);
or UO_346 (O_346,N_14089,N_14016);
nand UO_347 (O_347,N_14907,N_14673);
and UO_348 (O_348,N_14657,N_14750);
nor UO_349 (O_349,N_14779,N_14502);
and UO_350 (O_350,N_14007,N_14738);
nand UO_351 (O_351,N_14651,N_14399);
nand UO_352 (O_352,N_14928,N_14318);
nand UO_353 (O_353,N_14030,N_14312);
nand UO_354 (O_354,N_14878,N_14542);
and UO_355 (O_355,N_14805,N_14437);
and UO_356 (O_356,N_14060,N_14243);
or UO_357 (O_357,N_14558,N_14146);
or UO_358 (O_358,N_14095,N_14969);
xnor UO_359 (O_359,N_14848,N_14746);
or UO_360 (O_360,N_14074,N_14383);
or UO_361 (O_361,N_14715,N_14297);
and UO_362 (O_362,N_14062,N_14852);
nand UO_363 (O_363,N_14392,N_14103);
and UO_364 (O_364,N_14575,N_14218);
nand UO_365 (O_365,N_14585,N_14656);
or UO_366 (O_366,N_14547,N_14119);
nor UO_367 (O_367,N_14367,N_14704);
or UO_368 (O_368,N_14473,N_14761);
or UO_369 (O_369,N_14154,N_14342);
or UO_370 (O_370,N_14438,N_14446);
or UO_371 (O_371,N_14372,N_14948);
nand UO_372 (O_372,N_14024,N_14572);
nor UO_373 (O_373,N_14491,N_14285);
nand UO_374 (O_374,N_14768,N_14109);
nand UO_375 (O_375,N_14696,N_14081);
xnor UO_376 (O_376,N_14823,N_14478);
and UO_377 (O_377,N_14429,N_14471);
nor UO_378 (O_378,N_14322,N_14349);
and UO_379 (O_379,N_14204,N_14835);
xor UO_380 (O_380,N_14128,N_14419);
and UO_381 (O_381,N_14851,N_14801);
nand UO_382 (O_382,N_14892,N_14519);
nand UO_383 (O_383,N_14011,N_14573);
and UO_384 (O_384,N_14692,N_14250);
or UO_385 (O_385,N_14485,N_14449);
xor UO_386 (O_386,N_14874,N_14510);
nor UO_387 (O_387,N_14903,N_14276);
nand UO_388 (O_388,N_14538,N_14513);
nor UO_389 (O_389,N_14722,N_14008);
nor UO_390 (O_390,N_14520,N_14909);
or UO_391 (O_391,N_14191,N_14824);
or UO_392 (O_392,N_14267,N_14858);
or UO_393 (O_393,N_14919,N_14482);
nand UO_394 (O_394,N_14139,N_14484);
or UO_395 (O_395,N_14085,N_14377);
xor UO_396 (O_396,N_14080,N_14425);
and UO_397 (O_397,N_14868,N_14822);
nand UO_398 (O_398,N_14184,N_14123);
nor UO_399 (O_399,N_14819,N_14158);
nand UO_400 (O_400,N_14869,N_14845);
xnor UO_401 (O_401,N_14580,N_14363);
or UO_402 (O_402,N_14012,N_14448);
xor UO_403 (O_403,N_14742,N_14734);
nor UO_404 (O_404,N_14275,N_14944);
and UO_405 (O_405,N_14134,N_14872);
or UO_406 (O_406,N_14718,N_14397);
xnor UO_407 (O_407,N_14114,N_14630);
nand UO_408 (O_408,N_14895,N_14149);
or UO_409 (O_409,N_14111,N_14182);
xnor UO_410 (O_410,N_14916,N_14082);
or UO_411 (O_411,N_14728,N_14936);
nor UO_412 (O_412,N_14540,N_14386);
nand UO_413 (O_413,N_14233,N_14661);
nand UO_414 (O_414,N_14818,N_14296);
or UO_415 (O_415,N_14245,N_14129);
xor UO_416 (O_416,N_14401,N_14475);
or UO_417 (O_417,N_14561,N_14179);
and UO_418 (O_418,N_14031,N_14078);
or UO_419 (O_419,N_14988,N_14817);
nand UO_420 (O_420,N_14912,N_14799);
nor UO_421 (O_421,N_14506,N_14664);
or UO_422 (O_422,N_14190,N_14283);
and UO_423 (O_423,N_14496,N_14336);
or UO_424 (O_424,N_14783,N_14900);
and UO_425 (O_425,N_14380,N_14655);
or UO_426 (O_426,N_14681,N_14041);
nor UO_427 (O_427,N_14451,N_14693);
nor UO_428 (O_428,N_14343,N_14328);
nor UO_429 (O_429,N_14013,N_14440);
or UO_430 (O_430,N_14777,N_14325);
or UO_431 (O_431,N_14854,N_14803);
nand UO_432 (O_432,N_14784,N_14200);
or UO_433 (O_433,N_14287,N_14557);
and UO_434 (O_434,N_14582,N_14145);
nor UO_435 (O_435,N_14842,N_14057);
nand UO_436 (O_436,N_14733,N_14052);
and UO_437 (O_437,N_14663,N_14825);
and UO_438 (O_438,N_14436,N_14930);
and UO_439 (O_439,N_14198,N_14477);
or UO_440 (O_440,N_14603,N_14794);
and UO_441 (O_441,N_14701,N_14171);
xnor UO_442 (O_442,N_14117,N_14385);
nor UO_443 (O_443,N_14277,N_14137);
or UO_444 (O_444,N_14107,N_14504);
nor UO_445 (O_445,N_14308,N_14084);
and UO_446 (O_446,N_14913,N_14273);
or UO_447 (O_447,N_14665,N_14680);
nor UO_448 (O_448,N_14609,N_14771);
and UO_449 (O_449,N_14404,N_14800);
nand UO_450 (O_450,N_14174,N_14879);
or UO_451 (O_451,N_14435,N_14199);
nor UO_452 (O_452,N_14358,N_14646);
and UO_453 (O_453,N_14518,N_14623);
nor UO_454 (O_454,N_14227,N_14994);
and UO_455 (O_455,N_14844,N_14395);
or UO_456 (O_456,N_14709,N_14956);
nor UO_457 (O_457,N_14467,N_14754);
and UO_458 (O_458,N_14897,N_14197);
nor UO_459 (O_459,N_14209,N_14544);
nor UO_460 (O_460,N_14610,N_14678);
xor UO_461 (O_461,N_14005,N_14186);
or UO_462 (O_462,N_14650,N_14231);
xnor UO_463 (O_463,N_14378,N_14445);
or UO_464 (O_464,N_14025,N_14766);
nor UO_465 (O_465,N_14167,N_14108);
nor UO_466 (O_466,N_14516,N_14608);
xor UO_467 (O_467,N_14788,N_14352);
nor UO_468 (O_468,N_14294,N_14995);
or UO_469 (O_469,N_14194,N_14621);
xnor UO_470 (O_470,N_14096,N_14413);
nor UO_471 (O_471,N_14899,N_14345);
nor UO_472 (O_472,N_14838,N_14212);
nor UO_473 (O_473,N_14304,N_14394);
nor UO_474 (O_474,N_14237,N_14301);
or UO_475 (O_475,N_14712,N_14061);
nor UO_476 (O_476,N_14290,N_14545);
nand UO_477 (O_477,N_14551,N_14775);
and UO_478 (O_478,N_14442,N_14735);
nor UO_479 (O_479,N_14599,N_14009);
or UO_480 (O_480,N_14597,N_14634);
or UO_481 (O_481,N_14828,N_14321);
or UO_482 (O_482,N_14659,N_14898);
xor UO_483 (O_483,N_14168,N_14223);
nand UO_484 (O_484,N_14836,N_14508);
nor UO_485 (O_485,N_14889,N_14870);
and UO_486 (O_486,N_14126,N_14933);
nor UO_487 (O_487,N_14063,N_14751);
nand UO_488 (O_488,N_14246,N_14280);
or UO_489 (O_489,N_14172,N_14252);
or UO_490 (O_490,N_14666,N_14577);
xnor UO_491 (O_491,N_14497,N_14086);
nand UO_492 (O_492,N_14721,N_14583);
nand UO_493 (O_493,N_14797,N_14175);
nand UO_494 (O_494,N_14272,N_14314);
nand UO_495 (O_495,N_14877,N_14268);
and UO_496 (O_496,N_14876,N_14679);
and UO_497 (O_497,N_14432,N_14163);
or UO_498 (O_498,N_14719,N_14556);
and UO_499 (O_499,N_14509,N_14713);
or UO_500 (O_500,N_14137,N_14902);
and UO_501 (O_501,N_14950,N_14088);
or UO_502 (O_502,N_14246,N_14047);
or UO_503 (O_503,N_14252,N_14861);
and UO_504 (O_504,N_14304,N_14465);
nand UO_505 (O_505,N_14109,N_14667);
nor UO_506 (O_506,N_14623,N_14905);
xnor UO_507 (O_507,N_14810,N_14285);
nor UO_508 (O_508,N_14934,N_14328);
or UO_509 (O_509,N_14297,N_14205);
nand UO_510 (O_510,N_14222,N_14710);
nand UO_511 (O_511,N_14304,N_14168);
nand UO_512 (O_512,N_14648,N_14976);
xnor UO_513 (O_513,N_14686,N_14293);
and UO_514 (O_514,N_14870,N_14789);
xnor UO_515 (O_515,N_14942,N_14940);
and UO_516 (O_516,N_14543,N_14031);
and UO_517 (O_517,N_14141,N_14158);
and UO_518 (O_518,N_14088,N_14035);
and UO_519 (O_519,N_14131,N_14230);
nor UO_520 (O_520,N_14061,N_14865);
nor UO_521 (O_521,N_14585,N_14631);
and UO_522 (O_522,N_14410,N_14164);
nor UO_523 (O_523,N_14785,N_14232);
nand UO_524 (O_524,N_14737,N_14775);
or UO_525 (O_525,N_14250,N_14670);
xor UO_526 (O_526,N_14741,N_14735);
or UO_527 (O_527,N_14217,N_14625);
nor UO_528 (O_528,N_14555,N_14886);
or UO_529 (O_529,N_14448,N_14462);
nand UO_530 (O_530,N_14794,N_14361);
or UO_531 (O_531,N_14694,N_14616);
xor UO_532 (O_532,N_14279,N_14435);
or UO_533 (O_533,N_14399,N_14756);
nor UO_534 (O_534,N_14658,N_14361);
nand UO_535 (O_535,N_14810,N_14468);
nor UO_536 (O_536,N_14335,N_14990);
or UO_537 (O_537,N_14207,N_14887);
nor UO_538 (O_538,N_14767,N_14057);
or UO_539 (O_539,N_14421,N_14437);
nor UO_540 (O_540,N_14832,N_14116);
and UO_541 (O_541,N_14369,N_14577);
or UO_542 (O_542,N_14823,N_14175);
nand UO_543 (O_543,N_14370,N_14630);
nand UO_544 (O_544,N_14195,N_14270);
nand UO_545 (O_545,N_14421,N_14124);
and UO_546 (O_546,N_14304,N_14760);
or UO_547 (O_547,N_14964,N_14992);
nor UO_548 (O_548,N_14985,N_14473);
and UO_549 (O_549,N_14875,N_14343);
and UO_550 (O_550,N_14779,N_14374);
and UO_551 (O_551,N_14070,N_14111);
nand UO_552 (O_552,N_14949,N_14107);
and UO_553 (O_553,N_14272,N_14240);
and UO_554 (O_554,N_14900,N_14838);
or UO_555 (O_555,N_14338,N_14079);
nor UO_556 (O_556,N_14373,N_14834);
or UO_557 (O_557,N_14969,N_14026);
or UO_558 (O_558,N_14583,N_14547);
nand UO_559 (O_559,N_14694,N_14167);
nor UO_560 (O_560,N_14425,N_14812);
xor UO_561 (O_561,N_14045,N_14357);
xnor UO_562 (O_562,N_14485,N_14475);
xor UO_563 (O_563,N_14988,N_14037);
nand UO_564 (O_564,N_14585,N_14590);
nand UO_565 (O_565,N_14624,N_14392);
and UO_566 (O_566,N_14925,N_14073);
xnor UO_567 (O_567,N_14511,N_14326);
xnor UO_568 (O_568,N_14367,N_14736);
and UO_569 (O_569,N_14679,N_14535);
and UO_570 (O_570,N_14854,N_14809);
or UO_571 (O_571,N_14907,N_14512);
and UO_572 (O_572,N_14747,N_14279);
nand UO_573 (O_573,N_14988,N_14193);
nor UO_574 (O_574,N_14927,N_14461);
and UO_575 (O_575,N_14052,N_14476);
nor UO_576 (O_576,N_14486,N_14589);
nor UO_577 (O_577,N_14284,N_14179);
nor UO_578 (O_578,N_14087,N_14586);
nor UO_579 (O_579,N_14081,N_14390);
nand UO_580 (O_580,N_14954,N_14697);
and UO_581 (O_581,N_14435,N_14844);
and UO_582 (O_582,N_14038,N_14439);
or UO_583 (O_583,N_14066,N_14636);
nor UO_584 (O_584,N_14688,N_14121);
or UO_585 (O_585,N_14791,N_14240);
nor UO_586 (O_586,N_14896,N_14500);
and UO_587 (O_587,N_14738,N_14269);
nor UO_588 (O_588,N_14296,N_14513);
or UO_589 (O_589,N_14576,N_14474);
and UO_590 (O_590,N_14022,N_14019);
nand UO_591 (O_591,N_14700,N_14144);
and UO_592 (O_592,N_14362,N_14312);
or UO_593 (O_593,N_14657,N_14292);
and UO_594 (O_594,N_14640,N_14170);
nand UO_595 (O_595,N_14965,N_14633);
nor UO_596 (O_596,N_14588,N_14135);
or UO_597 (O_597,N_14673,N_14342);
nand UO_598 (O_598,N_14915,N_14541);
xnor UO_599 (O_599,N_14780,N_14297);
and UO_600 (O_600,N_14115,N_14099);
nor UO_601 (O_601,N_14465,N_14922);
nor UO_602 (O_602,N_14057,N_14108);
and UO_603 (O_603,N_14200,N_14998);
nand UO_604 (O_604,N_14713,N_14579);
or UO_605 (O_605,N_14879,N_14905);
nand UO_606 (O_606,N_14069,N_14605);
nor UO_607 (O_607,N_14686,N_14662);
or UO_608 (O_608,N_14167,N_14857);
nor UO_609 (O_609,N_14724,N_14755);
or UO_610 (O_610,N_14934,N_14930);
or UO_611 (O_611,N_14371,N_14840);
nor UO_612 (O_612,N_14389,N_14916);
or UO_613 (O_613,N_14628,N_14268);
nand UO_614 (O_614,N_14874,N_14743);
nor UO_615 (O_615,N_14720,N_14033);
and UO_616 (O_616,N_14433,N_14331);
xnor UO_617 (O_617,N_14806,N_14625);
nand UO_618 (O_618,N_14188,N_14374);
nor UO_619 (O_619,N_14096,N_14116);
or UO_620 (O_620,N_14518,N_14125);
and UO_621 (O_621,N_14866,N_14947);
and UO_622 (O_622,N_14688,N_14462);
nor UO_623 (O_623,N_14627,N_14340);
nor UO_624 (O_624,N_14105,N_14297);
nand UO_625 (O_625,N_14651,N_14925);
xnor UO_626 (O_626,N_14684,N_14531);
nor UO_627 (O_627,N_14374,N_14095);
and UO_628 (O_628,N_14585,N_14008);
nor UO_629 (O_629,N_14757,N_14192);
and UO_630 (O_630,N_14786,N_14153);
nor UO_631 (O_631,N_14511,N_14280);
nand UO_632 (O_632,N_14752,N_14606);
nor UO_633 (O_633,N_14573,N_14434);
and UO_634 (O_634,N_14582,N_14829);
nor UO_635 (O_635,N_14916,N_14990);
nand UO_636 (O_636,N_14481,N_14853);
and UO_637 (O_637,N_14682,N_14622);
nand UO_638 (O_638,N_14089,N_14391);
nand UO_639 (O_639,N_14141,N_14249);
or UO_640 (O_640,N_14548,N_14825);
or UO_641 (O_641,N_14742,N_14334);
nor UO_642 (O_642,N_14738,N_14463);
and UO_643 (O_643,N_14738,N_14217);
and UO_644 (O_644,N_14449,N_14889);
nor UO_645 (O_645,N_14792,N_14261);
and UO_646 (O_646,N_14373,N_14501);
nor UO_647 (O_647,N_14725,N_14301);
xnor UO_648 (O_648,N_14923,N_14800);
nand UO_649 (O_649,N_14704,N_14247);
nor UO_650 (O_650,N_14949,N_14936);
nor UO_651 (O_651,N_14765,N_14210);
nand UO_652 (O_652,N_14226,N_14463);
nand UO_653 (O_653,N_14035,N_14626);
nand UO_654 (O_654,N_14605,N_14380);
and UO_655 (O_655,N_14306,N_14645);
nor UO_656 (O_656,N_14939,N_14085);
nand UO_657 (O_657,N_14916,N_14759);
nand UO_658 (O_658,N_14242,N_14224);
nand UO_659 (O_659,N_14782,N_14282);
or UO_660 (O_660,N_14847,N_14209);
nand UO_661 (O_661,N_14920,N_14237);
nand UO_662 (O_662,N_14424,N_14030);
xnor UO_663 (O_663,N_14817,N_14929);
nor UO_664 (O_664,N_14584,N_14191);
and UO_665 (O_665,N_14251,N_14295);
xor UO_666 (O_666,N_14136,N_14708);
nand UO_667 (O_667,N_14964,N_14633);
or UO_668 (O_668,N_14325,N_14973);
nor UO_669 (O_669,N_14731,N_14828);
or UO_670 (O_670,N_14526,N_14880);
and UO_671 (O_671,N_14964,N_14156);
nor UO_672 (O_672,N_14796,N_14482);
xnor UO_673 (O_673,N_14191,N_14684);
nor UO_674 (O_674,N_14825,N_14564);
xnor UO_675 (O_675,N_14934,N_14182);
and UO_676 (O_676,N_14195,N_14894);
nand UO_677 (O_677,N_14861,N_14977);
nor UO_678 (O_678,N_14126,N_14068);
or UO_679 (O_679,N_14551,N_14969);
or UO_680 (O_680,N_14657,N_14439);
or UO_681 (O_681,N_14450,N_14025);
or UO_682 (O_682,N_14254,N_14061);
nand UO_683 (O_683,N_14479,N_14318);
xnor UO_684 (O_684,N_14368,N_14173);
and UO_685 (O_685,N_14322,N_14051);
or UO_686 (O_686,N_14814,N_14899);
and UO_687 (O_687,N_14927,N_14025);
and UO_688 (O_688,N_14068,N_14392);
and UO_689 (O_689,N_14753,N_14888);
nand UO_690 (O_690,N_14706,N_14518);
nor UO_691 (O_691,N_14246,N_14373);
or UO_692 (O_692,N_14555,N_14992);
nor UO_693 (O_693,N_14098,N_14903);
and UO_694 (O_694,N_14292,N_14164);
nand UO_695 (O_695,N_14944,N_14006);
or UO_696 (O_696,N_14362,N_14388);
nor UO_697 (O_697,N_14662,N_14524);
or UO_698 (O_698,N_14329,N_14117);
and UO_699 (O_699,N_14987,N_14081);
or UO_700 (O_700,N_14783,N_14151);
and UO_701 (O_701,N_14675,N_14507);
nor UO_702 (O_702,N_14404,N_14077);
xor UO_703 (O_703,N_14838,N_14615);
nor UO_704 (O_704,N_14277,N_14205);
nor UO_705 (O_705,N_14524,N_14217);
nand UO_706 (O_706,N_14497,N_14496);
nor UO_707 (O_707,N_14521,N_14805);
nor UO_708 (O_708,N_14969,N_14228);
and UO_709 (O_709,N_14118,N_14117);
or UO_710 (O_710,N_14198,N_14243);
xor UO_711 (O_711,N_14705,N_14526);
nand UO_712 (O_712,N_14683,N_14364);
nand UO_713 (O_713,N_14578,N_14636);
nor UO_714 (O_714,N_14423,N_14775);
or UO_715 (O_715,N_14298,N_14506);
nand UO_716 (O_716,N_14991,N_14978);
or UO_717 (O_717,N_14037,N_14172);
and UO_718 (O_718,N_14772,N_14383);
and UO_719 (O_719,N_14910,N_14199);
nor UO_720 (O_720,N_14892,N_14481);
or UO_721 (O_721,N_14725,N_14062);
and UO_722 (O_722,N_14060,N_14667);
nor UO_723 (O_723,N_14082,N_14700);
or UO_724 (O_724,N_14200,N_14737);
nor UO_725 (O_725,N_14617,N_14482);
and UO_726 (O_726,N_14056,N_14165);
or UO_727 (O_727,N_14114,N_14154);
or UO_728 (O_728,N_14469,N_14956);
nor UO_729 (O_729,N_14221,N_14075);
nor UO_730 (O_730,N_14736,N_14979);
nand UO_731 (O_731,N_14710,N_14262);
or UO_732 (O_732,N_14146,N_14369);
nor UO_733 (O_733,N_14432,N_14450);
nor UO_734 (O_734,N_14348,N_14076);
nand UO_735 (O_735,N_14704,N_14483);
xnor UO_736 (O_736,N_14260,N_14352);
nor UO_737 (O_737,N_14746,N_14532);
and UO_738 (O_738,N_14280,N_14965);
and UO_739 (O_739,N_14849,N_14181);
nor UO_740 (O_740,N_14066,N_14859);
nand UO_741 (O_741,N_14722,N_14492);
or UO_742 (O_742,N_14533,N_14055);
and UO_743 (O_743,N_14350,N_14233);
nand UO_744 (O_744,N_14857,N_14126);
or UO_745 (O_745,N_14596,N_14664);
and UO_746 (O_746,N_14755,N_14557);
or UO_747 (O_747,N_14913,N_14739);
nor UO_748 (O_748,N_14046,N_14196);
nand UO_749 (O_749,N_14678,N_14068);
xor UO_750 (O_750,N_14592,N_14395);
and UO_751 (O_751,N_14207,N_14075);
xor UO_752 (O_752,N_14248,N_14967);
or UO_753 (O_753,N_14924,N_14733);
nand UO_754 (O_754,N_14133,N_14066);
or UO_755 (O_755,N_14017,N_14161);
and UO_756 (O_756,N_14950,N_14394);
or UO_757 (O_757,N_14872,N_14039);
nor UO_758 (O_758,N_14679,N_14578);
nand UO_759 (O_759,N_14599,N_14034);
nand UO_760 (O_760,N_14018,N_14416);
nand UO_761 (O_761,N_14944,N_14060);
nand UO_762 (O_762,N_14856,N_14228);
nand UO_763 (O_763,N_14155,N_14616);
or UO_764 (O_764,N_14039,N_14497);
and UO_765 (O_765,N_14129,N_14468);
or UO_766 (O_766,N_14742,N_14748);
or UO_767 (O_767,N_14160,N_14825);
nand UO_768 (O_768,N_14187,N_14100);
nor UO_769 (O_769,N_14768,N_14694);
xor UO_770 (O_770,N_14665,N_14617);
nor UO_771 (O_771,N_14737,N_14129);
and UO_772 (O_772,N_14070,N_14215);
xor UO_773 (O_773,N_14121,N_14060);
or UO_774 (O_774,N_14987,N_14212);
nor UO_775 (O_775,N_14646,N_14373);
nor UO_776 (O_776,N_14787,N_14187);
xor UO_777 (O_777,N_14447,N_14550);
and UO_778 (O_778,N_14193,N_14517);
nor UO_779 (O_779,N_14500,N_14392);
nor UO_780 (O_780,N_14934,N_14500);
nand UO_781 (O_781,N_14663,N_14205);
or UO_782 (O_782,N_14892,N_14028);
and UO_783 (O_783,N_14735,N_14682);
or UO_784 (O_784,N_14762,N_14364);
nor UO_785 (O_785,N_14413,N_14145);
nand UO_786 (O_786,N_14240,N_14110);
nand UO_787 (O_787,N_14788,N_14180);
xor UO_788 (O_788,N_14493,N_14391);
or UO_789 (O_789,N_14210,N_14301);
or UO_790 (O_790,N_14907,N_14417);
nand UO_791 (O_791,N_14923,N_14943);
or UO_792 (O_792,N_14277,N_14518);
and UO_793 (O_793,N_14022,N_14625);
or UO_794 (O_794,N_14911,N_14897);
xnor UO_795 (O_795,N_14779,N_14063);
nor UO_796 (O_796,N_14496,N_14087);
nor UO_797 (O_797,N_14698,N_14073);
or UO_798 (O_798,N_14235,N_14625);
nand UO_799 (O_799,N_14185,N_14356);
nand UO_800 (O_800,N_14033,N_14886);
nor UO_801 (O_801,N_14766,N_14362);
and UO_802 (O_802,N_14743,N_14584);
or UO_803 (O_803,N_14403,N_14476);
nor UO_804 (O_804,N_14767,N_14710);
or UO_805 (O_805,N_14293,N_14273);
and UO_806 (O_806,N_14913,N_14305);
nand UO_807 (O_807,N_14165,N_14684);
nand UO_808 (O_808,N_14052,N_14452);
nor UO_809 (O_809,N_14408,N_14557);
or UO_810 (O_810,N_14436,N_14777);
nand UO_811 (O_811,N_14493,N_14270);
nand UO_812 (O_812,N_14497,N_14043);
and UO_813 (O_813,N_14825,N_14634);
and UO_814 (O_814,N_14588,N_14848);
and UO_815 (O_815,N_14088,N_14553);
and UO_816 (O_816,N_14058,N_14306);
xnor UO_817 (O_817,N_14056,N_14582);
or UO_818 (O_818,N_14157,N_14647);
nor UO_819 (O_819,N_14506,N_14415);
or UO_820 (O_820,N_14299,N_14351);
nor UO_821 (O_821,N_14632,N_14690);
or UO_822 (O_822,N_14366,N_14495);
or UO_823 (O_823,N_14843,N_14873);
xnor UO_824 (O_824,N_14074,N_14995);
nand UO_825 (O_825,N_14286,N_14226);
or UO_826 (O_826,N_14814,N_14110);
and UO_827 (O_827,N_14954,N_14456);
nor UO_828 (O_828,N_14198,N_14779);
nand UO_829 (O_829,N_14335,N_14345);
or UO_830 (O_830,N_14270,N_14022);
nor UO_831 (O_831,N_14968,N_14807);
and UO_832 (O_832,N_14920,N_14804);
nor UO_833 (O_833,N_14714,N_14348);
and UO_834 (O_834,N_14985,N_14982);
nand UO_835 (O_835,N_14152,N_14732);
and UO_836 (O_836,N_14787,N_14036);
or UO_837 (O_837,N_14507,N_14305);
nand UO_838 (O_838,N_14581,N_14289);
nor UO_839 (O_839,N_14122,N_14018);
and UO_840 (O_840,N_14597,N_14859);
nor UO_841 (O_841,N_14778,N_14913);
and UO_842 (O_842,N_14285,N_14124);
and UO_843 (O_843,N_14146,N_14149);
and UO_844 (O_844,N_14341,N_14779);
nand UO_845 (O_845,N_14816,N_14545);
or UO_846 (O_846,N_14711,N_14723);
nor UO_847 (O_847,N_14927,N_14241);
or UO_848 (O_848,N_14184,N_14508);
and UO_849 (O_849,N_14130,N_14648);
nand UO_850 (O_850,N_14746,N_14886);
xor UO_851 (O_851,N_14775,N_14473);
or UO_852 (O_852,N_14914,N_14242);
xor UO_853 (O_853,N_14420,N_14208);
xor UO_854 (O_854,N_14602,N_14299);
nor UO_855 (O_855,N_14347,N_14355);
and UO_856 (O_856,N_14824,N_14303);
or UO_857 (O_857,N_14324,N_14934);
or UO_858 (O_858,N_14510,N_14239);
xor UO_859 (O_859,N_14851,N_14092);
and UO_860 (O_860,N_14942,N_14250);
nor UO_861 (O_861,N_14744,N_14559);
nor UO_862 (O_862,N_14430,N_14866);
and UO_863 (O_863,N_14917,N_14729);
and UO_864 (O_864,N_14720,N_14566);
xnor UO_865 (O_865,N_14217,N_14853);
and UO_866 (O_866,N_14566,N_14176);
nand UO_867 (O_867,N_14189,N_14971);
or UO_868 (O_868,N_14735,N_14878);
nor UO_869 (O_869,N_14612,N_14318);
nor UO_870 (O_870,N_14019,N_14304);
nor UO_871 (O_871,N_14824,N_14898);
nor UO_872 (O_872,N_14684,N_14421);
or UO_873 (O_873,N_14406,N_14682);
xnor UO_874 (O_874,N_14456,N_14703);
xnor UO_875 (O_875,N_14117,N_14930);
nand UO_876 (O_876,N_14470,N_14216);
and UO_877 (O_877,N_14569,N_14113);
nor UO_878 (O_878,N_14067,N_14779);
and UO_879 (O_879,N_14582,N_14908);
and UO_880 (O_880,N_14910,N_14632);
and UO_881 (O_881,N_14035,N_14361);
nand UO_882 (O_882,N_14596,N_14629);
nor UO_883 (O_883,N_14529,N_14045);
or UO_884 (O_884,N_14039,N_14243);
and UO_885 (O_885,N_14538,N_14124);
and UO_886 (O_886,N_14924,N_14415);
and UO_887 (O_887,N_14973,N_14126);
or UO_888 (O_888,N_14554,N_14865);
and UO_889 (O_889,N_14349,N_14626);
or UO_890 (O_890,N_14352,N_14730);
nor UO_891 (O_891,N_14530,N_14382);
or UO_892 (O_892,N_14135,N_14879);
and UO_893 (O_893,N_14086,N_14711);
or UO_894 (O_894,N_14785,N_14362);
and UO_895 (O_895,N_14592,N_14121);
or UO_896 (O_896,N_14187,N_14684);
or UO_897 (O_897,N_14833,N_14768);
nor UO_898 (O_898,N_14010,N_14452);
nor UO_899 (O_899,N_14952,N_14254);
and UO_900 (O_900,N_14420,N_14047);
nor UO_901 (O_901,N_14436,N_14688);
and UO_902 (O_902,N_14545,N_14507);
nor UO_903 (O_903,N_14148,N_14629);
nand UO_904 (O_904,N_14582,N_14418);
nand UO_905 (O_905,N_14325,N_14617);
or UO_906 (O_906,N_14601,N_14695);
xor UO_907 (O_907,N_14538,N_14232);
xnor UO_908 (O_908,N_14798,N_14718);
or UO_909 (O_909,N_14901,N_14620);
nor UO_910 (O_910,N_14571,N_14713);
or UO_911 (O_911,N_14141,N_14104);
and UO_912 (O_912,N_14765,N_14379);
nand UO_913 (O_913,N_14476,N_14027);
or UO_914 (O_914,N_14794,N_14212);
nand UO_915 (O_915,N_14928,N_14311);
nor UO_916 (O_916,N_14995,N_14695);
or UO_917 (O_917,N_14133,N_14353);
and UO_918 (O_918,N_14609,N_14850);
and UO_919 (O_919,N_14465,N_14462);
and UO_920 (O_920,N_14437,N_14449);
or UO_921 (O_921,N_14676,N_14527);
and UO_922 (O_922,N_14614,N_14832);
nand UO_923 (O_923,N_14161,N_14019);
or UO_924 (O_924,N_14126,N_14297);
nor UO_925 (O_925,N_14478,N_14196);
nand UO_926 (O_926,N_14657,N_14650);
nand UO_927 (O_927,N_14973,N_14940);
nor UO_928 (O_928,N_14890,N_14961);
or UO_929 (O_929,N_14345,N_14963);
and UO_930 (O_930,N_14837,N_14965);
nor UO_931 (O_931,N_14069,N_14815);
and UO_932 (O_932,N_14139,N_14536);
nor UO_933 (O_933,N_14041,N_14590);
and UO_934 (O_934,N_14197,N_14689);
and UO_935 (O_935,N_14189,N_14686);
nand UO_936 (O_936,N_14070,N_14397);
xor UO_937 (O_937,N_14540,N_14621);
xnor UO_938 (O_938,N_14490,N_14736);
or UO_939 (O_939,N_14048,N_14265);
nor UO_940 (O_940,N_14335,N_14287);
nor UO_941 (O_941,N_14472,N_14418);
nand UO_942 (O_942,N_14212,N_14517);
nand UO_943 (O_943,N_14771,N_14097);
nor UO_944 (O_944,N_14466,N_14442);
nand UO_945 (O_945,N_14300,N_14157);
and UO_946 (O_946,N_14354,N_14295);
xnor UO_947 (O_947,N_14521,N_14849);
nor UO_948 (O_948,N_14157,N_14691);
nor UO_949 (O_949,N_14082,N_14539);
nor UO_950 (O_950,N_14089,N_14996);
nor UO_951 (O_951,N_14955,N_14354);
nor UO_952 (O_952,N_14135,N_14883);
nor UO_953 (O_953,N_14239,N_14892);
and UO_954 (O_954,N_14881,N_14619);
or UO_955 (O_955,N_14909,N_14583);
nor UO_956 (O_956,N_14318,N_14509);
and UO_957 (O_957,N_14833,N_14301);
nand UO_958 (O_958,N_14574,N_14736);
nor UO_959 (O_959,N_14539,N_14324);
nand UO_960 (O_960,N_14588,N_14416);
or UO_961 (O_961,N_14768,N_14737);
and UO_962 (O_962,N_14348,N_14618);
and UO_963 (O_963,N_14157,N_14154);
nand UO_964 (O_964,N_14866,N_14976);
nand UO_965 (O_965,N_14349,N_14088);
nand UO_966 (O_966,N_14564,N_14541);
and UO_967 (O_967,N_14605,N_14526);
xor UO_968 (O_968,N_14284,N_14205);
or UO_969 (O_969,N_14734,N_14891);
or UO_970 (O_970,N_14960,N_14947);
nor UO_971 (O_971,N_14933,N_14786);
and UO_972 (O_972,N_14841,N_14173);
and UO_973 (O_973,N_14325,N_14563);
nand UO_974 (O_974,N_14660,N_14483);
and UO_975 (O_975,N_14518,N_14028);
nand UO_976 (O_976,N_14804,N_14565);
nor UO_977 (O_977,N_14078,N_14648);
nand UO_978 (O_978,N_14498,N_14025);
or UO_979 (O_979,N_14549,N_14965);
or UO_980 (O_980,N_14373,N_14536);
and UO_981 (O_981,N_14621,N_14752);
xor UO_982 (O_982,N_14753,N_14591);
and UO_983 (O_983,N_14721,N_14940);
or UO_984 (O_984,N_14336,N_14964);
nand UO_985 (O_985,N_14808,N_14840);
nor UO_986 (O_986,N_14937,N_14993);
nand UO_987 (O_987,N_14026,N_14828);
nand UO_988 (O_988,N_14288,N_14738);
or UO_989 (O_989,N_14200,N_14168);
nand UO_990 (O_990,N_14602,N_14890);
xnor UO_991 (O_991,N_14247,N_14051);
and UO_992 (O_992,N_14028,N_14250);
xnor UO_993 (O_993,N_14758,N_14365);
nand UO_994 (O_994,N_14446,N_14125);
nor UO_995 (O_995,N_14866,N_14121);
and UO_996 (O_996,N_14228,N_14930);
nor UO_997 (O_997,N_14229,N_14932);
nor UO_998 (O_998,N_14696,N_14260);
nor UO_999 (O_999,N_14223,N_14577);
nand UO_1000 (O_1000,N_14046,N_14034);
nand UO_1001 (O_1001,N_14101,N_14676);
and UO_1002 (O_1002,N_14939,N_14632);
and UO_1003 (O_1003,N_14085,N_14115);
xnor UO_1004 (O_1004,N_14567,N_14283);
xnor UO_1005 (O_1005,N_14615,N_14837);
nand UO_1006 (O_1006,N_14752,N_14713);
xnor UO_1007 (O_1007,N_14651,N_14789);
nor UO_1008 (O_1008,N_14748,N_14749);
and UO_1009 (O_1009,N_14412,N_14188);
or UO_1010 (O_1010,N_14506,N_14935);
nand UO_1011 (O_1011,N_14651,N_14611);
xor UO_1012 (O_1012,N_14804,N_14581);
and UO_1013 (O_1013,N_14743,N_14435);
xor UO_1014 (O_1014,N_14261,N_14910);
nand UO_1015 (O_1015,N_14243,N_14751);
and UO_1016 (O_1016,N_14555,N_14279);
and UO_1017 (O_1017,N_14985,N_14640);
nand UO_1018 (O_1018,N_14108,N_14678);
or UO_1019 (O_1019,N_14085,N_14550);
nor UO_1020 (O_1020,N_14310,N_14938);
nor UO_1021 (O_1021,N_14176,N_14038);
or UO_1022 (O_1022,N_14277,N_14630);
or UO_1023 (O_1023,N_14987,N_14022);
nand UO_1024 (O_1024,N_14660,N_14616);
and UO_1025 (O_1025,N_14195,N_14690);
and UO_1026 (O_1026,N_14604,N_14685);
nand UO_1027 (O_1027,N_14998,N_14297);
nand UO_1028 (O_1028,N_14017,N_14392);
or UO_1029 (O_1029,N_14362,N_14979);
and UO_1030 (O_1030,N_14527,N_14483);
nand UO_1031 (O_1031,N_14631,N_14569);
nand UO_1032 (O_1032,N_14075,N_14128);
nand UO_1033 (O_1033,N_14860,N_14672);
xnor UO_1034 (O_1034,N_14844,N_14375);
and UO_1035 (O_1035,N_14168,N_14372);
nor UO_1036 (O_1036,N_14765,N_14625);
nor UO_1037 (O_1037,N_14144,N_14179);
nand UO_1038 (O_1038,N_14888,N_14206);
nor UO_1039 (O_1039,N_14109,N_14746);
or UO_1040 (O_1040,N_14362,N_14090);
or UO_1041 (O_1041,N_14516,N_14788);
or UO_1042 (O_1042,N_14202,N_14554);
and UO_1043 (O_1043,N_14454,N_14423);
xnor UO_1044 (O_1044,N_14292,N_14373);
or UO_1045 (O_1045,N_14337,N_14636);
and UO_1046 (O_1046,N_14703,N_14955);
or UO_1047 (O_1047,N_14949,N_14922);
and UO_1048 (O_1048,N_14499,N_14392);
and UO_1049 (O_1049,N_14978,N_14364);
nand UO_1050 (O_1050,N_14982,N_14500);
or UO_1051 (O_1051,N_14590,N_14271);
nor UO_1052 (O_1052,N_14036,N_14596);
nor UO_1053 (O_1053,N_14396,N_14414);
or UO_1054 (O_1054,N_14939,N_14420);
nand UO_1055 (O_1055,N_14573,N_14753);
and UO_1056 (O_1056,N_14738,N_14839);
or UO_1057 (O_1057,N_14287,N_14902);
or UO_1058 (O_1058,N_14074,N_14848);
nand UO_1059 (O_1059,N_14046,N_14251);
or UO_1060 (O_1060,N_14262,N_14317);
or UO_1061 (O_1061,N_14815,N_14542);
nand UO_1062 (O_1062,N_14558,N_14543);
nor UO_1063 (O_1063,N_14553,N_14522);
xor UO_1064 (O_1064,N_14327,N_14680);
and UO_1065 (O_1065,N_14107,N_14014);
nor UO_1066 (O_1066,N_14780,N_14821);
nand UO_1067 (O_1067,N_14431,N_14093);
or UO_1068 (O_1068,N_14656,N_14910);
nand UO_1069 (O_1069,N_14891,N_14555);
nor UO_1070 (O_1070,N_14584,N_14368);
or UO_1071 (O_1071,N_14459,N_14569);
or UO_1072 (O_1072,N_14962,N_14323);
nor UO_1073 (O_1073,N_14303,N_14189);
or UO_1074 (O_1074,N_14123,N_14316);
nor UO_1075 (O_1075,N_14131,N_14850);
xnor UO_1076 (O_1076,N_14640,N_14551);
or UO_1077 (O_1077,N_14407,N_14308);
or UO_1078 (O_1078,N_14821,N_14496);
nor UO_1079 (O_1079,N_14199,N_14434);
and UO_1080 (O_1080,N_14074,N_14878);
nand UO_1081 (O_1081,N_14562,N_14376);
and UO_1082 (O_1082,N_14130,N_14807);
nand UO_1083 (O_1083,N_14579,N_14369);
and UO_1084 (O_1084,N_14551,N_14809);
or UO_1085 (O_1085,N_14442,N_14094);
and UO_1086 (O_1086,N_14879,N_14464);
nand UO_1087 (O_1087,N_14500,N_14182);
nand UO_1088 (O_1088,N_14152,N_14106);
or UO_1089 (O_1089,N_14535,N_14652);
nor UO_1090 (O_1090,N_14499,N_14047);
nand UO_1091 (O_1091,N_14651,N_14073);
or UO_1092 (O_1092,N_14639,N_14761);
or UO_1093 (O_1093,N_14186,N_14347);
xor UO_1094 (O_1094,N_14907,N_14463);
and UO_1095 (O_1095,N_14132,N_14538);
and UO_1096 (O_1096,N_14240,N_14448);
or UO_1097 (O_1097,N_14657,N_14700);
or UO_1098 (O_1098,N_14344,N_14266);
or UO_1099 (O_1099,N_14348,N_14591);
or UO_1100 (O_1100,N_14638,N_14209);
or UO_1101 (O_1101,N_14648,N_14259);
and UO_1102 (O_1102,N_14144,N_14461);
and UO_1103 (O_1103,N_14721,N_14208);
or UO_1104 (O_1104,N_14207,N_14039);
nor UO_1105 (O_1105,N_14670,N_14475);
and UO_1106 (O_1106,N_14637,N_14110);
and UO_1107 (O_1107,N_14413,N_14425);
or UO_1108 (O_1108,N_14208,N_14143);
nand UO_1109 (O_1109,N_14741,N_14241);
or UO_1110 (O_1110,N_14771,N_14674);
nand UO_1111 (O_1111,N_14790,N_14390);
and UO_1112 (O_1112,N_14442,N_14645);
nand UO_1113 (O_1113,N_14420,N_14767);
or UO_1114 (O_1114,N_14713,N_14490);
and UO_1115 (O_1115,N_14012,N_14079);
and UO_1116 (O_1116,N_14357,N_14732);
nor UO_1117 (O_1117,N_14103,N_14985);
and UO_1118 (O_1118,N_14691,N_14821);
nand UO_1119 (O_1119,N_14799,N_14217);
xnor UO_1120 (O_1120,N_14910,N_14156);
or UO_1121 (O_1121,N_14953,N_14784);
nor UO_1122 (O_1122,N_14127,N_14728);
nor UO_1123 (O_1123,N_14866,N_14922);
nor UO_1124 (O_1124,N_14360,N_14317);
xnor UO_1125 (O_1125,N_14513,N_14323);
and UO_1126 (O_1126,N_14760,N_14525);
nand UO_1127 (O_1127,N_14531,N_14894);
nor UO_1128 (O_1128,N_14503,N_14422);
or UO_1129 (O_1129,N_14941,N_14326);
nand UO_1130 (O_1130,N_14213,N_14380);
or UO_1131 (O_1131,N_14984,N_14073);
xnor UO_1132 (O_1132,N_14945,N_14781);
or UO_1133 (O_1133,N_14322,N_14053);
nor UO_1134 (O_1134,N_14127,N_14068);
nand UO_1135 (O_1135,N_14981,N_14459);
and UO_1136 (O_1136,N_14960,N_14337);
nor UO_1137 (O_1137,N_14378,N_14480);
or UO_1138 (O_1138,N_14230,N_14227);
nand UO_1139 (O_1139,N_14277,N_14417);
nor UO_1140 (O_1140,N_14078,N_14349);
or UO_1141 (O_1141,N_14122,N_14370);
nand UO_1142 (O_1142,N_14970,N_14032);
and UO_1143 (O_1143,N_14751,N_14757);
nand UO_1144 (O_1144,N_14390,N_14277);
nand UO_1145 (O_1145,N_14082,N_14748);
xnor UO_1146 (O_1146,N_14063,N_14511);
nand UO_1147 (O_1147,N_14637,N_14977);
nand UO_1148 (O_1148,N_14930,N_14111);
nor UO_1149 (O_1149,N_14793,N_14486);
nor UO_1150 (O_1150,N_14125,N_14993);
nor UO_1151 (O_1151,N_14265,N_14271);
nor UO_1152 (O_1152,N_14514,N_14127);
nor UO_1153 (O_1153,N_14377,N_14364);
nand UO_1154 (O_1154,N_14395,N_14916);
nor UO_1155 (O_1155,N_14031,N_14690);
nand UO_1156 (O_1156,N_14096,N_14565);
and UO_1157 (O_1157,N_14354,N_14833);
xnor UO_1158 (O_1158,N_14439,N_14905);
nor UO_1159 (O_1159,N_14897,N_14903);
nor UO_1160 (O_1160,N_14535,N_14675);
or UO_1161 (O_1161,N_14410,N_14798);
nand UO_1162 (O_1162,N_14016,N_14050);
and UO_1163 (O_1163,N_14449,N_14619);
xnor UO_1164 (O_1164,N_14507,N_14310);
and UO_1165 (O_1165,N_14301,N_14197);
nand UO_1166 (O_1166,N_14159,N_14182);
and UO_1167 (O_1167,N_14225,N_14948);
nor UO_1168 (O_1168,N_14549,N_14176);
nand UO_1169 (O_1169,N_14853,N_14328);
or UO_1170 (O_1170,N_14453,N_14491);
nor UO_1171 (O_1171,N_14403,N_14769);
xnor UO_1172 (O_1172,N_14195,N_14661);
or UO_1173 (O_1173,N_14563,N_14378);
nand UO_1174 (O_1174,N_14380,N_14372);
nand UO_1175 (O_1175,N_14857,N_14173);
or UO_1176 (O_1176,N_14834,N_14605);
or UO_1177 (O_1177,N_14293,N_14216);
nand UO_1178 (O_1178,N_14102,N_14890);
xor UO_1179 (O_1179,N_14077,N_14721);
or UO_1180 (O_1180,N_14676,N_14903);
nor UO_1181 (O_1181,N_14553,N_14653);
or UO_1182 (O_1182,N_14853,N_14937);
and UO_1183 (O_1183,N_14446,N_14588);
xnor UO_1184 (O_1184,N_14566,N_14694);
or UO_1185 (O_1185,N_14168,N_14465);
nor UO_1186 (O_1186,N_14766,N_14960);
nand UO_1187 (O_1187,N_14954,N_14479);
xnor UO_1188 (O_1188,N_14648,N_14969);
and UO_1189 (O_1189,N_14599,N_14164);
nand UO_1190 (O_1190,N_14722,N_14129);
nand UO_1191 (O_1191,N_14238,N_14638);
and UO_1192 (O_1192,N_14493,N_14735);
nor UO_1193 (O_1193,N_14880,N_14572);
or UO_1194 (O_1194,N_14753,N_14725);
nand UO_1195 (O_1195,N_14429,N_14426);
nand UO_1196 (O_1196,N_14848,N_14260);
nor UO_1197 (O_1197,N_14779,N_14003);
nand UO_1198 (O_1198,N_14672,N_14793);
or UO_1199 (O_1199,N_14559,N_14326);
nor UO_1200 (O_1200,N_14548,N_14227);
or UO_1201 (O_1201,N_14751,N_14968);
xnor UO_1202 (O_1202,N_14282,N_14566);
nand UO_1203 (O_1203,N_14855,N_14816);
nor UO_1204 (O_1204,N_14537,N_14826);
nor UO_1205 (O_1205,N_14697,N_14366);
and UO_1206 (O_1206,N_14982,N_14668);
and UO_1207 (O_1207,N_14837,N_14355);
and UO_1208 (O_1208,N_14382,N_14323);
and UO_1209 (O_1209,N_14689,N_14710);
and UO_1210 (O_1210,N_14976,N_14678);
and UO_1211 (O_1211,N_14241,N_14322);
xnor UO_1212 (O_1212,N_14621,N_14628);
nor UO_1213 (O_1213,N_14419,N_14869);
nand UO_1214 (O_1214,N_14994,N_14597);
or UO_1215 (O_1215,N_14993,N_14111);
nand UO_1216 (O_1216,N_14776,N_14179);
and UO_1217 (O_1217,N_14700,N_14773);
nand UO_1218 (O_1218,N_14080,N_14190);
or UO_1219 (O_1219,N_14429,N_14201);
nand UO_1220 (O_1220,N_14722,N_14098);
nor UO_1221 (O_1221,N_14567,N_14144);
and UO_1222 (O_1222,N_14046,N_14534);
and UO_1223 (O_1223,N_14724,N_14707);
and UO_1224 (O_1224,N_14679,N_14001);
xor UO_1225 (O_1225,N_14585,N_14206);
nor UO_1226 (O_1226,N_14047,N_14833);
nor UO_1227 (O_1227,N_14602,N_14540);
nor UO_1228 (O_1228,N_14216,N_14714);
xor UO_1229 (O_1229,N_14730,N_14514);
nand UO_1230 (O_1230,N_14908,N_14322);
nor UO_1231 (O_1231,N_14934,N_14523);
nor UO_1232 (O_1232,N_14791,N_14324);
and UO_1233 (O_1233,N_14565,N_14827);
and UO_1234 (O_1234,N_14709,N_14380);
or UO_1235 (O_1235,N_14623,N_14736);
nor UO_1236 (O_1236,N_14655,N_14836);
or UO_1237 (O_1237,N_14062,N_14129);
nand UO_1238 (O_1238,N_14546,N_14296);
nand UO_1239 (O_1239,N_14805,N_14225);
or UO_1240 (O_1240,N_14602,N_14967);
nand UO_1241 (O_1241,N_14545,N_14869);
xnor UO_1242 (O_1242,N_14265,N_14196);
nand UO_1243 (O_1243,N_14957,N_14917);
or UO_1244 (O_1244,N_14595,N_14999);
nand UO_1245 (O_1245,N_14554,N_14084);
and UO_1246 (O_1246,N_14159,N_14376);
and UO_1247 (O_1247,N_14633,N_14897);
nand UO_1248 (O_1248,N_14418,N_14329);
nand UO_1249 (O_1249,N_14028,N_14391);
nand UO_1250 (O_1250,N_14285,N_14793);
nor UO_1251 (O_1251,N_14389,N_14183);
or UO_1252 (O_1252,N_14028,N_14837);
xnor UO_1253 (O_1253,N_14192,N_14954);
and UO_1254 (O_1254,N_14392,N_14220);
nand UO_1255 (O_1255,N_14509,N_14854);
nor UO_1256 (O_1256,N_14070,N_14645);
or UO_1257 (O_1257,N_14033,N_14991);
and UO_1258 (O_1258,N_14841,N_14239);
nor UO_1259 (O_1259,N_14064,N_14276);
nor UO_1260 (O_1260,N_14968,N_14983);
nand UO_1261 (O_1261,N_14940,N_14982);
nand UO_1262 (O_1262,N_14596,N_14147);
nor UO_1263 (O_1263,N_14839,N_14489);
or UO_1264 (O_1264,N_14640,N_14311);
or UO_1265 (O_1265,N_14357,N_14639);
and UO_1266 (O_1266,N_14001,N_14753);
or UO_1267 (O_1267,N_14975,N_14486);
nor UO_1268 (O_1268,N_14109,N_14580);
or UO_1269 (O_1269,N_14865,N_14464);
nand UO_1270 (O_1270,N_14499,N_14906);
or UO_1271 (O_1271,N_14745,N_14820);
nor UO_1272 (O_1272,N_14581,N_14227);
or UO_1273 (O_1273,N_14733,N_14952);
nand UO_1274 (O_1274,N_14152,N_14486);
or UO_1275 (O_1275,N_14270,N_14152);
nand UO_1276 (O_1276,N_14781,N_14915);
or UO_1277 (O_1277,N_14532,N_14650);
or UO_1278 (O_1278,N_14679,N_14644);
or UO_1279 (O_1279,N_14460,N_14222);
or UO_1280 (O_1280,N_14847,N_14623);
or UO_1281 (O_1281,N_14808,N_14060);
nand UO_1282 (O_1282,N_14263,N_14262);
xor UO_1283 (O_1283,N_14865,N_14834);
and UO_1284 (O_1284,N_14587,N_14254);
nor UO_1285 (O_1285,N_14776,N_14120);
xor UO_1286 (O_1286,N_14937,N_14623);
or UO_1287 (O_1287,N_14499,N_14427);
nand UO_1288 (O_1288,N_14946,N_14725);
nand UO_1289 (O_1289,N_14015,N_14299);
xnor UO_1290 (O_1290,N_14192,N_14064);
and UO_1291 (O_1291,N_14552,N_14393);
and UO_1292 (O_1292,N_14385,N_14230);
and UO_1293 (O_1293,N_14900,N_14249);
and UO_1294 (O_1294,N_14412,N_14971);
or UO_1295 (O_1295,N_14368,N_14649);
nand UO_1296 (O_1296,N_14859,N_14908);
nor UO_1297 (O_1297,N_14758,N_14698);
or UO_1298 (O_1298,N_14561,N_14476);
and UO_1299 (O_1299,N_14126,N_14927);
and UO_1300 (O_1300,N_14743,N_14610);
nor UO_1301 (O_1301,N_14295,N_14528);
or UO_1302 (O_1302,N_14296,N_14310);
nand UO_1303 (O_1303,N_14442,N_14892);
and UO_1304 (O_1304,N_14283,N_14548);
nand UO_1305 (O_1305,N_14869,N_14569);
nor UO_1306 (O_1306,N_14356,N_14595);
nand UO_1307 (O_1307,N_14127,N_14095);
and UO_1308 (O_1308,N_14440,N_14795);
and UO_1309 (O_1309,N_14011,N_14448);
xor UO_1310 (O_1310,N_14679,N_14598);
and UO_1311 (O_1311,N_14284,N_14856);
nor UO_1312 (O_1312,N_14818,N_14311);
and UO_1313 (O_1313,N_14648,N_14258);
nand UO_1314 (O_1314,N_14418,N_14535);
nor UO_1315 (O_1315,N_14634,N_14168);
nand UO_1316 (O_1316,N_14089,N_14266);
or UO_1317 (O_1317,N_14229,N_14384);
or UO_1318 (O_1318,N_14535,N_14006);
nand UO_1319 (O_1319,N_14187,N_14580);
xnor UO_1320 (O_1320,N_14286,N_14719);
and UO_1321 (O_1321,N_14916,N_14213);
nand UO_1322 (O_1322,N_14412,N_14732);
xor UO_1323 (O_1323,N_14915,N_14357);
xor UO_1324 (O_1324,N_14212,N_14900);
and UO_1325 (O_1325,N_14412,N_14060);
or UO_1326 (O_1326,N_14130,N_14267);
and UO_1327 (O_1327,N_14809,N_14857);
xor UO_1328 (O_1328,N_14068,N_14121);
or UO_1329 (O_1329,N_14498,N_14007);
and UO_1330 (O_1330,N_14938,N_14324);
nand UO_1331 (O_1331,N_14651,N_14755);
or UO_1332 (O_1332,N_14435,N_14652);
nor UO_1333 (O_1333,N_14631,N_14073);
nor UO_1334 (O_1334,N_14849,N_14727);
or UO_1335 (O_1335,N_14598,N_14560);
and UO_1336 (O_1336,N_14630,N_14117);
and UO_1337 (O_1337,N_14389,N_14029);
or UO_1338 (O_1338,N_14648,N_14213);
nor UO_1339 (O_1339,N_14174,N_14211);
nor UO_1340 (O_1340,N_14833,N_14424);
nand UO_1341 (O_1341,N_14441,N_14081);
and UO_1342 (O_1342,N_14541,N_14018);
or UO_1343 (O_1343,N_14589,N_14041);
nand UO_1344 (O_1344,N_14786,N_14580);
nor UO_1345 (O_1345,N_14748,N_14369);
or UO_1346 (O_1346,N_14512,N_14938);
or UO_1347 (O_1347,N_14489,N_14869);
nand UO_1348 (O_1348,N_14553,N_14365);
and UO_1349 (O_1349,N_14688,N_14156);
and UO_1350 (O_1350,N_14875,N_14767);
or UO_1351 (O_1351,N_14132,N_14433);
or UO_1352 (O_1352,N_14769,N_14445);
nand UO_1353 (O_1353,N_14981,N_14835);
and UO_1354 (O_1354,N_14255,N_14461);
and UO_1355 (O_1355,N_14722,N_14150);
or UO_1356 (O_1356,N_14548,N_14040);
and UO_1357 (O_1357,N_14765,N_14123);
nor UO_1358 (O_1358,N_14559,N_14199);
and UO_1359 (O_1359,N_14063,N_14877);
nor UO_1360 (O_1360,N_14962,N_14936);
nor UO_1361 (O_1361,N_14355,N_14700);
and UO_1362 (O_1362,N_14729,N_14293);
nand UO_1363 (O_1363,N_14792,N_14993);
or UO_1364 (O_1364,N_14581,N_14930);
and UO_1365 (O_1365,N_14867,N_14527);
and UO_1366 (O_1366,N_14742,N_14178);
nand UO_1367 (O_1367,N_14311,N_14126);
nand UO_1368 (O_1368,N_14600,N_14251);
xor UO_1369 (O_1369,N_14886,N_14775);
and UO_1370 (O_1370,N_14111,N_14355);
or UO_1371 (O_1371,N_14814,N_14416);
xnor UO_1372 (O_1372,N_14045,N_14287);
nand UO_1373 (O_1373,N_14508,N_14349);
nand UO_1374 (O_1374,N_14180,N_14440);
nor UO_1375 (O_1375,N_14198,N_14195);
nand UO_1376 (O_1376,N_14162,N_14699);
or UO_1377 (O_1377,N_14994,N_14078);
or UO_1378 (O_1378,N_14217,N_14952);
and UO_1379 (O_1379,N_14300,N_14192);
or UO_1380 (O_1380,N_14028,N_14812);
and UO_1381 (O_1381,N_14608,N_14272);
nand UO_1382 (O_1382,N_14594,N_14592);
nand UO_1383 (O_1383,N_14148,N_14567);
and UO_1384 (O_1384,N_14805,N_14364);
xor UO_1385 (O_1385,N_14789,N_14105);
nor UO_1386 (O_1386,N_14248,N_14739);
and UO_1387 (O_1387,N_14628,N_14977);
or UO_1388 (O_1388,N_14245,N_14787);
nand UO_1389 (O_1389,N_14668,N_14776);
xor UO_1390 (O_1390,N_14546,N_14683);
nor UO_1391 (O_1391,N_14734,N_14263);
nand UO_1392 (O_1392,N_14210,N_14638);
nor UO_1393 (O_1393,N_14457,N_14628);
nand UO_1394 (O_1394,N_14561,N_14360);
nor UO_1395 (O_1395,N_14778,N_14845);
nor UO_1396 (O_1396,N_14445,N_14602);
nand UO_1397 (O_1397,N_14367,N_14475);
nor UO_1398 (O_1398,N_14026,N_14793);
nor UO_1399 (O_1399,N_14487,N_14397);
nand UO_1400 (O_1400,N_14875,N_14773);
nor UO_1401 (O_1401,N_14202,N_14033);
or UO_1402 (O_1402,N_14842,N_14032);
nor UO_1403 (O_1403,N_14446,N_14516);
nor UO_1404 (O_1404,N_14705,N_14102);
nor UO_1405 (O_1405,N_14239,N_14833);
nand UO_1406 (O_1406,N_14291,N_14581);
and UO_1407 (O_1407,N_14679,N_14939);
or UO_1408 (O_1408,N_14168,N_14235);
or UO_1409 (O_1409,N_14772,N_14034);
xor UO_1410 (O_1410,N_14052,N_14198);
and UO_1411 (O_1411,N_14254,N_14894);
nand UO_1412 (O_1412,N_14281,N_14788);
nand UO_1413 (O_1413,N_14460,N_14549);
or UO_1414 (O_1414,N_14986,N_14199);
nor UO_1415 (O_1415,N_14163,N_14248);
nor UO_1416 (O_1416,N_14446,N_14805);
or UO_1417 (O_1417,N_14597,N_14059);
nand UO_1418 (O_1418,N_14126,N_14175);
or UO_1419 (O_1419,N_14416,N_14665);
and UO_1420 (O_1420,N_14921,N_14117);
nor UO_1421 (O_1421,N_14627,N_14702);
or UO_1422 (O_1422,N_14145,N_14271);
and UO_1423 (O_1423,N_14101,N_14146);
nand UO_1424 (O_1424,N_14672,N_14419);
nor UO_1425 (O_1425,N_14425,N_14053);
nor UO_1426 (O_1426,N_14015,N_14578);
nand UO_1427 (O_1427,N_14384,N_14620);
nor UO_1428 (O_1428,N_14142,N_14794);
and UO_1429 (O_1429,N_14890,N_14214);
nor UO_1430 (O_1430,N_14477,N_14687);
or UO_1431 (O_1431,N_14972,N_14706);
nand UO_1432 (O_1432,N_14068,N_14569);
nor UO_1433 (O_1433,N_14194,N_14387);
nand UO_1434 (O_1434,N_14811,N_14891);
xor UO_1435 (O_1435,N_14269,N_14776);
or UO_1436 (O_1436,N_14771,N_14973);
or UO_1437 (O_1437,N_14141,N_14623);
nand UO_1438 (O_1438,N_14786,N_14476);
nand UO_1439 (O_1439,N_14045,N_14066);
and UO_1440 (O_1440,N_14513,N_14244);
and UO_1441 (O_1441,N_14862,N_14618);
nand UO_1442 (O_1442,N_14940,N_14558);
nand UO_1443 (O_1443,N_14751,N_14786);
nand UO_1444 (O_1444,N_14015,N_14538);
or UO_1445 (O_1445,N_14863,N_14825);
nand UO_1446 (O_1446,N_14737,N_14780);
nor UO_1447 (O_1447,N_14213,N_14874);
and UO_1448 (O_1448,N_14228,N_14592);
and UO_1449 (O_1449,N_14062,N_14951);
nand UO_1450 (O_1450,N_14344,N_14589);
or UO_1451 (O_1451,N_14717,N_14381);
nor UO_1452 (O_1452,N_14095,N_14213);
or UO_1453 (O_1453,N_14226,N_14680);
or UO_1454 (O_1454,N_14904,N_14891);
or UO_1455 (O_1455,N_14913,N_14662);
and UO_1456 (O_1456,N_14884,N_14626);
and UO_1457 (O_1457,N_14366,N_14284);
or UO_1458 (O_1458,N_14699,N_14608);
nor UO_1459 (O_1459,N_14555,N_14262);
nor UO_1460 (O_1460,N_14005,N_14407);
nand UO_1461 (O_1461,N_14387,N_14854);
or UO_1462 (O_1462,N_14965,N_14873);
nand UO_1463 (O_1463,N_14096,N_14739);
nand UO_1464 (O_1464,N_14984,N_14731);
nand UO_1465 (O_1465,N_14992,N_14521);
and UO_1466 (O_1466,N_14305,N_14340);
nand UO_1467 (O_1467,N_14499,N_14785);
nor UO_1468 (O_1468,N_14193,N_14986);
nor UO_1469 (O_1469,N_14090,N_14006);
nor UO_1470 (O_1470,N_14125,N_14837);
nor UO_1471 (O_1471,N_14997,N_14721);
or UO_1472 (O_1472,N_14359,N_14362);
and UO_1473 (O_1473,N_14896,N_14076);
or UO_1474 (O_1474,N_14736,N_14205);
nand UO_1475 (O_1475,N_14517,N_14059);
xor UO_1476 (O_1476,N_14768,N_14853);
or UO_1477 (O_1477,N_14161,N_14080);
nor UO_1478 (O_1478,N_14949,N_14563);
and UO_1479 (O_1479,N_14273,N_14864);
xor UO_1480 (O_1480,N_14910,N_14006);
or UO_1481 (O_1481,N_14810,N_14266);
and UO_1482 (O_1482,N_14439,N_14929);
or UO_1483 (O_1483,N_14865,N_14594);
and UO_1484 (O_1484,N_14015,N_14071);
nand UO_1485 (O_1485,N_14266,N_14590);
or UO_1486 (O_1486,N_14089,N_14275);
nor UO_1487 (O_1487,N_14416,N_14672);
or UO_1488 (O_1488,N_14723,N_14808);
or UO_1489 (O_1489,N_14073,N_14391);
nand UO_1490 (O_1490,N_14372,N_14164);
nand UO_1491 (O_1491,N_14019,N_14828);
nor UO_1492 (O_1492,N_14226,N_14256);
or UO_1493 (O_1493,N_14680,N_14208);
or UO_1494 (O_1494,N_14049,N_14959);
nor UO_1495 (O_1495,N_14483,N_14884);
nor UO_1496 (O_1496,N_14984,N_14436);
and UO_1497 (O_1497,N_14654,N_14621);
or UO_1498 (O_1498,N_14176,N_14567);
nand UO_1499 (O_1499,N_14661,N_14388);
nor UO_1500 (O_1500,N_14807,N_14204);
or UO_1501 (O_1501,N_14373,N_14944);
or UO_1502 (O_1502,N_14656,N_14230);
nor UO_1503 (O_1503,N_14911,N_14487);
or UO_1504 (O_1504,N_14195,N_14055);
or UO_1505 (O_1505,N_14180,N_14380);
nand UO_1506 (O_1506,N_14755,N_14803);
nand UO_1507 (O_1507,N_14429,N_14793);
nand UO_1508 (O_1508,N_14474,N_14704);
nor UO_1509 (O_1509,N_14046,N_14556);
nand UO_1510 (O_1510,N_14491,N_14291);
nand UO_1511 (O_1511,N_14277,N_14949);
or UO_1512 (O_1512,N_14173,N_14654);
nor UO_1513 (O_1513,N_14622,N_14194);
nor UO_1514 (O_1514,N_14898,N_14006);
nor UO_1515 (O_1515,N_14854,N_14089);
nor UO_1516 (O_1516,N_14545,N_14917);
xor UO_1517 (O_1517,N_14952,N_14209);
or UO_1518 (O_1518,N_14804,N_14593);
or UO_1519 (O_1519,N_14716,N_14417);
nor UO_1520 (O_1520,N_14034,N_14119);
nor UO_1521 (O_1521,N_14218,N_14801);
or UO_1522 (O_1522,N_14736,N_14371);
nand UO_1523 (O_1523,N_14166,N_14558);
nand UO_1524 (O_1524,N_14512,N_14996);
or UO_1525 (O_1525,N_14343,N_14594);
xnor UO_1526 (O_1526,N_14590,N_14757);
nor UO_1527 (O_1527,N_14606,N_14410);
xnor UO_1528 (O_1528,N_14265,N_14463);
nand UO_1529 (O_1529,N_14793,N_14044);
nor UO_1530 (O_1530,N_14993,N_14164);
nor UO_1531 (O_1531,N_14581,N_14077);
nor UO_1532 (O_1532,N_14083,N_14387);
xor UO_1533 (O_1533,N_14267,N_14440);
nand UO_1534 (O_1534,N_14271,N_14696);
or UO_1535 (O_1535,N_14557,N_14599);
or UO_1536 (O_1536,N_14723,N_14222);
xor UO_1537 (O_1537,N_14634,N_14263);
nor UO_1538 (O_1538,N_14643,N_14662);
or UO_1539 (O_1539,N_14649,N_14875);
and UO_1540 (O_1540,N_14015,N_14052);
and UO_1541 (O_1541,N_14404,N_14722);
nand UO_1542 (O_1542,N_14385,N_14112);
or UO_1543 (O_1543,N_14483,N_14890);
and UO_1544 (O_1544,N_14151,N_14597);
xnor UO_1545 (O_1545,N_14703,N_14320);
xor UO_1546 (O_1546,N_14221,N_14109);
nor UO_1547 (O_1547,N_14814,N_14567);
and UO_1548 (O_1548,N_14370,N_14095);
nand UO_1549 (O_1549,N_14813,N_14858);
nor UO_1550 (O_1550,N_14416,N_14864);
nand UO_1551 (O_1551,N_14676,N_14587);
nor UO_1552 (O_1552,N_14088,N_14592);
nand UO_1553 (O_1553,N_14478,N_14803);
and UO_1554 (O_1554,N_14780,N_14413);
xor UO_1555 (O_1555,N_14792,N_14216);
or UO_1556 (O_1556,N_14763,N_14192);
and UO_1557 (O_1557,N_14558,N_14039);
and UO_1558 (O_1558,N_14169,N_14862);
and UO_1559 (O_1559,N_14664,N_14625);
nor UO_1560 (O_1560,N_14485,N_14446);
or UO_1561 (O_1561,N_14189,N_14635);
xor UO_1562 (O_1562,N_14415,N_14244);
nand UO_1563 (O_1563,N_14361,N_14043);
nand UO_1564 (O_1564,N_14236,N_14771);
xor UO_1565 (O_1565,N_14944,N_14517);
nand UO_1566 (O_1566,N_14582,N_14061);
nor UO_1567 (O_1567,N_14529,N_14009);
or UO_1568 (O_1568,N_14204,N_14078);
nand UO_1569 (O_1569,N_14292,N_14186);
xnor UO_1570 (O_1570,N_14861,N_14283);
or UO_1571 (O_1571,N_14970,N_14368);
nand UO_1572 (O_1572,N_14416,N_14537);
nor UO_1573 (O_1573,N_14563,N_14287);
nor UO_1574 (O_1574,N_14819,N_14448);
nor UO_1575 (O_1575,N_14977,N_14566);
or UO_1576 (O_1576,N_14786,N_14816);
nor UO_1577 (O_1577,N_14712,N_14636);
nor UO_1578 (O_1578,N_14520,N_14601);
or UO_1579 (O_1579,N_14969,N_14654);
xor UO_1580 (O_1580,N_14055,N_14480);
xnor UO_1581 (O_1581,N_14173,N_14505);
nor UO_1582 (O_1582,N_14600,N_14968);
nand UO_1583 (O_1583,N_14162,N_14343);
and UO_1584 (O_1584,N_14317,N_14997);
or UO_1585 (O_1585,N_14964,N_14927);
nand UO_1586 (O_1586,N_14330,N_14840);
nor UO_1587 (O_1587,N_14228,N_14295);
and UO_1588 (O_1588,N_14668,N_14876);
xor UO_1589 (O_1589,N_14881,N_14303);
or UO_1590 (O_1590,N_14432,N_14387);
or UO_1591 (O_1591,N_14027,N_14053);
xor UO_1592 (O_1592,N_14330,N_14088);
or UO_1593 (O_1593,N_14263,N_14033);
nor UO_1594 (O_1594,N_14566,N_14480);
or UO_1595 (O_1595,N_14271,N_14377);
nor UO_1596 (O_1596,N_14927,N_14239);
or UO_1597 (O_1597,N_14806,N_14192);
nor UO_1598 (O_1598,N_14328,N_14628);
or UO_1599 (O_1599,N_14213,N_14280);
nand UO_1600 (O_1600,N_14181,N_14350);
and UO_1601 (O_1601,N_14880,N_14740);
nor UO_1602 (O_1602,N_14543,N_14916);
or UO_1603 (O_1603,N_14078,N_14556);
nand UO_1604 (O_1604,N_14117,N_14073);
nor UO_1605 (O_1605,N_14745,N_14651);
and UO_1606 (O_1606,N_14036,N_14088);
nor UO_1607 (O_1607,N_14593,N_14408);
or UO_1608 (O_1608,N_14177,N_14515);
nand UO_1609 (O_1609,N_14177,N_14002);
nor UO_1610 (O_1610,N_14524,N_14242);
nand UO_1611 (O_1611,N_14170,N_14013);
or UO_1612 (O_1612,N_14023,N_14078);
xnor UO_1613 (O_1613,N_14133,N_14580);
nor UO_1614 (O_1614,N_14534,N_14025);
nor UO_1615 (O_1615,N_14910,N_14979);
nand UO_1616 (O_1616,N_14677,N_14752);
or UO_1617 (O_1617,N_14508,N_14671);
and UO_1618 (O_1618,N_14262,N_14836);
and UO_1619 (O_1619,N_14085,N_14450);
or UO_1620 (O_1620,N_14554,N_14994);
xor UO_1621 (O_1621,N_14551,N_14537);
nand UO_1622 (O_1622,N_14895,N_14566);
or UO_1623 (O_1623,N_14741,N_14107);
nor UO_1624 (O_1624,N_14175,N_14939);
nor UO_1625 (O_1625,N_14814,N_14932);
nand UO_1626 (O_1626,N_14769,N_14823);
and UO_1627 (O_1627,N_14689,N_14874);
nor UO_1628 (O_1628,N_14388,N_14427);
nor UO_1629 (O_1629,N_14539,N_14212);
nor UO_1630 (O_1630,N_14774,N_14400);
and UO_1631 (O_1631,N_14396,N_14742);
or UO_1632 (O_1632,N_14042,N_14055);
nor UO_1633 (O_1633,N_14932,N_14307);
and UO_1634 (O_1634,N_14869,N_14003);
or UO_1635 (O_1635,N_14068,N_14073);
nor UO_1636 (O_1636,N_14030,N_14470);
nor UO_1637 (O_1637,N_14782,N_14030);
or UO_1638 (O_1638,N_14485,N_14816);
and UO_1639 (O_1639,N_14993,N_14648);
nor UO_1640 (O_1640,N_14240,N_14615);
or UO_1641 (O_1641,N_14884,N_14768);
nor UO_1642 (O_1642,N_14556,N_14860);
xnor UO_1643 (O_1643,N_14957,N_14000);
nand UO_1644 (O_1644,N_14837,N_14060);
xor UO_1645 (O_1645,N_14078,N_14541);
xor UO_1646 (O_1646,N_14625,N_14873);
nand UO_1647 (O_1647,N_14485,N_14569);
and UO_1648 (O_1648,N_14233,N_14081);
xnor UO_1649 (O_1649,N_14215,N_14997);
nor UO_1650 (O_1650,N_14441,N_14975);
and UO_1651 (O_1651,N_14130,N_14427);
xnor UO_1652 (O_1652,N_14952,N_14863);
and UO_1653 (O_1653,N_14856,N_14225);
xor UO_1654 (O_1654,N_14613,N_14305);
nand UO_1655 (O_1655,N_14153,N_14241);
nor UO_1656 (O_1656,N_14081,N_14878);
or UO_1657 (O_1657,N_14505,N_14199);
or UO_1658 (O_1658,N_14202,N_14214);
xor UO_1659 (O_1659,N_14262,N_14231);
nand UO_1660 (O_1660,N_14103,N_14846);
and UO_1661 (O_1661,N_14540,N_14213);
nand UO_1662 (O_1662,N_14706,N_14758);
xor UO_1663 (O_1663,N_14876,N_14407);
xor UO_1664 (O_1664,N_14281,N_14852);
nor UO_1665 (O_1665,N_14869,N_14540);
xor UO_1666 (O_1666,N_14243,N_14920);
nor UO_1667 (O_1667,N_14502,N_14445);
nor UO_1668 (O_1668,N_14940,N_14805);
nand UO_1669 (O_1669,N_14397,N_14845);
or UO_1670 (O_1670,N_14009,N_14034);
nor UO_1671 (O_1671,N_14309,N_14117);
nor UO_1672 (O_1672,N_14632,N_14478);
nor UO_1673 (O_1673,N_14755,N_14620);
nor UO_1674 (O_1674,N_14151,N_14703);
nor UO_1675 (O_1675,N_14897,N_14821);
nor UO_1676 (O_1676,N_14074,N_14880);
and UO_1677 (O_1677,N_14805,N_14970);
and UO_1678 (O_1678,N_14725,N_14157);
and UO_1679 (O_1679,N_14234,N_14627);
and UO_1680 (O_1680,N_14812,N_14644);
nor UO_1681 (O_1681,N_14471,N_14703);
or UO_1682 (O_1682,N_14876,N_14448);
and UO_1683 (O_1683,N_14897,N_14581);
nand UO_1684 (O_1684,N_14824,N_14875);
or UO_1685 (O_1685,N_14545,N_14891);
or UO_1686 (O_1686,N_14229,N_14239);
and UO_1687 (O_1687,N_14215,N_14084);
and UO_1688 (O_1688,N_14241,N_14021);
or UO_1689 (O_1689,N_14753,N_14322);
and UO_1690 (O_1690,N_14353,N_14273);
or UO_1691 (O_1691,N_14670,N_14686);
nor UO_1692 (O_1692,N_14996,N_14746);
nor UO_1693 (O_1693,N_14956,N_14775);
and UO_1694 (O_1694,N_14932,N_14022);
xor UO_1695 (O_1695,N_14812,N_14420);
nor UO_1696 (O_1696,N_14617,N_14545);
nand UO_1697 (O_1697,N_14908,N_14074);
or UO_1698 (O_1698,N_14813,N_14359);
nand UO_1699 (O_1699,N_14019,N_14591);
or UO_1700 (O_1700,N_14964,N_14344);
and UO_1701 (O_1701,N_14168,N_14478);
nor UO_1702 (O_1702,N_14442,N_14803);
and UO_1703 (O_1703,N_14948,N_14317);
nand UO_1704 (O_1704,N_14393,N_14764);
and UO_1705 (O_1705,N_14902,N_14227);
nor UO_1706 (O_1706,N_14588,N_14374);
nand UO_1707 (O_1707,N_14966,N_14317);
nand UO_1708 (O_1708,N_14631,N_14003);
and UO_1709 (O_1709,N_14363,N_14091);
or UO_1710 (O_1710,N_14705,N_14505);
nor UO_1711 (O_1711,N_14986,N_14819);
nor UO_1712 (O_1712,N_14693,N_14295);
nor UO_1713 (O_1713,N_14632,N_14011);
nand UO_1714 (O_1714,N_14472,N_14189);
or UO_1715 (O_1715,N_14255,N_14377);
and UO_1716 (O_1716,N_14083,N_14317);
or UO_1717 (O_1717,N_14001,N_14371);
or UO_1718 (O_1718,N_14911,N_14379);
and UO_1719 (O_1719,N_14911,N_14815);
nand UO_1720 (O_1720,N_14855,N_14913);
or UO_1721 (O_1721,N_14363,N_14381);
or UO_1722 (O_1722,N_14293,N_14944);
nand UO_1723 (O_1723,N_14239,N_14083);
or UO_1724 (O_1724,N_14833,N_14735);
nand UO_1725 (O_1725,N_14837,N_14249);
nor UO_1726 (O_1726,N_14149,N_14507);
nor UO_1727 (O_1727,N_14758,N_14294);
and UO_1728 (O_1728,N_14753,N_14878);
and UO_1729 (O_1729,N_14587,N_14756);
nor UO_1730 (O_1730,N_14584,N_14336);
nand UO_1731 (O_1731,N_14863,N_14709);
and UO_1732 (O_1732,N_14157,N_14067);
xor UO_1733 (O_1733,N_14162,N_14886);
and UO_1734 (O_1734,N_14382,N_14317);
and UO_1735 (O_1735,N_14820,N_14873);
and UO_1736 (O_1736,N_14911,N_14448);
and UO_1737 (O_1737,N_14234,N_14738);
nor UO_1738 (O_1738,N_14628,N_14827);
nand UO_1739 (O_1739,N_14849,N_14458);
xor UO_1740 (O_1740,N_14218,N_14724);
xor UO_1741 (O_1741,N_14684,N_14217);
nand UO_1742 (O_1742,N_14844,N_14641);
nand UO_1743 (O_1743,N_14644,N_14363);
nand UO_1744 (O_1744,N_14113,N_14389);
xnor UO_1745 (O_1745,N_14108,N_14025);
xor UO_1746 (O_1746,N_14928,N_14387);
nor UO_1747 (O_1747,N_14011,N_14356);
nor UO_1748 (O_1748,N_14039,N_14146);
and UO_1749 (O_1749,N_14153,N_14946);
xor UO_1750 (O_1750,N_14325,N_14352);
nor UO_1751 (O_1751,N_14594,N_14640);
nor UO_1752 (O_1752,N_14364,N_14695);
nand UO_1753 (O_1753,N_14912,N_14430);
or UO_1754 (O_1754,N_14218,N_14944);
or UO_1755 (O_1755,N_14973,N_14057);
or UO_1756 (O_1756,N_14115,N_14152);
nor UO_1757 (O_1757,N_14925,N_14813);
xnor UO_1758 (O_1758,N_14202,N_14024);
or UO_1759 (O_1759,N_14420,N_14902);
nand UO_1760 (O_1760,N_14025,N_14208);
and UO_1761 (O_1761,N_14018,N_14296);
and UO_1762 (O_1762,N_14677,N_14998);
and UO_1763 (O_1763,N_14743,N_14009);
and UO_1764 (O_1764,N_14388,N_14818);
and UO_1765 (O_1765,N_14062,N_14749);
xor UO_1766 (O_1766,N_14766,N_14210);
nand UO_1767 (O_1767,N_14573,N_14978);
nor UO_1768 (O_1768,N_14637,N_14010);
and UO_1769 (O_1769,N_14397,N_14019);
nand UO_1770 (O_1770,N_14649,N_14638);
or UO_1771 (O_1771,N_14805,N_14550);
nor UO_1772 (O_1772,N_14172,N_14331);
nand UO_1773 (O_1773,N_14965,N_14579);
or UO_1774 (O_1774,N_14951,N_14537);
xor UO_1775 (O_1775,N_14479,N_14607);
nand UO_1776 (O_1776,N_14086,N_14873);
xnor UO_1777 (O_1777,N_14872,N_14136);
or UO_1778 (O_1778,N_14562,N_14526);
xnor UO_1779 (O_1779,N_14533,N_14477);
nor UO_1780 (O_1780,N_14525,N_14948);
or UO_1781 (O_1781,N_14210,N_14499);
nand UO_1782 (O_1782,N_14376,N_14526);
nor UO_1783 (O_1783,N_14955,N_14422);
and UO_1784 (O_1784,N_14959,N_14685);
or UO_1785 (O_1785,N_14495,N_14126);
and UO_1786 (O_1786,N_14259,N_14744);
nand UO_1787 (O_1787,N_14278,N_14558);
or UO_1788 (O_1788,N_14058,N_14003);
nand UO_1789 (O_1789,N_14698,N_14982);
or UO_1790 (O_1790,N_14599,N_14655);
and UO_1791 (O_1791,N_14703,N_14987);
xor UO_1792 (O_1792,N_14251,N_14073);
or UO_1793 (O_1793,N_14039,N_14680);
nand UO_1794 (O_1794,N_14926,N_14196);
nand UO_1795 (O_1795,N_14349,N_14099);
nor UO_1796 (O_1796,N_14303,N_14187);
and UO_1797 (O_1797,N_14469,N_14303);
nor UO_1798 (O_1798,N_14886,N_14460);
and UO_1799 (O_1799,N_14737,N_14886);
nor UO_1800 (O_1800,N_14365,N_14675);
nand UO_1801 (O_1801,N_14459,N_14226);
nor UO_1802 (O_1802,N_14707,N_14379);
nand UO_1803 (O_1803,N_14515,N_14815);
nor UO_1804 (O_1804,N_14979,N_14321);
or UO_1805 (O_1805,N_14371,N_14954);
nand UO_1806 (O_1806,N_14932,N_14521);
nor UO_1807 (O_1807,N_14993,N_14229);
nand UO_1808 (O_1808,N_14965,N_14440);
nor UO_1809 (O_1809,N_14986,N_14127);
nand UO_1810 (O_1810,N_14260,N_14060);
and UO_1811 (O_1811,N_14132,N_14591);
and UO_1812 (O_1812,N_14075,N_14931);
nor UO_1813 (O_1813,N_14215,N_14244);
or UO_1814 (O_1814,N_14608,N_14211);
nand UO_1815 (O_1815,N_14430,N_14199);
nor UO_1816 (O_1816,N_14497,N_14892);
and UO_1817 (O_1817,N_14514,N_14370);
nand UO_1818 (O_1818,N_14347,N_14278);
xnor UO_1819 (O_1819,N_14870,N_14453);
nor UO_1820 (O_1820,N_14023,N_14249);
and UO_1821 (O_1821,N_14968,N_14268);
nor UO_1822 (O_1822,N_14819,N_14080);
xor UO_1823 (O_1823,N_14760,N_14235);
or UO_1824 (O_1824,N_14094,N_14407);
and UO_1825 (O_1825,N_14645,N_14726);
nor UO_1826 (O_1826,N_14086,N_14322);
or UO_1827 (O_1827,N_14065,N_14780);
nand UO_1828 (O_1828,N_14656,N_14485);
nand UO_1829 (O_1829,N_14213,N_14023);
nand UO_1830 (O_1830,N_14553,N_14126);
nand UO_1831 (O_1831,N_14231,N_14342);
nand UO_1832 (O_1832,N_14856,N_14534);
nand UO_1833 (O_1833,N_14468,N_14861);
nor UO_1834 (O_1834,N_14337,N_14257);
nand UO_1835 (O_1835,N_14009,N_14883);
xnor UO_1836 (O_1836,N_14396,N_14925);
nor UO_1837 (O_1837,N_14942,N_14578);
or UO_1838 (O_1838,N_14809,N_14512);
nand UO_1839 (O_1839,N_14114,N_14452);
nor UO_1840 (O_1840,N_14822,N_14271);
and UO_1841 (O_1841,N_14221,N_14604);
xor UO_1842 (O_1842,N_14185,N_14172);
xor UO_1843 (O_1843,N_14303,N_14780);
nand UO_1844 (O_1844,N_14395,N_14451);
or UO_1845 (O_1845,N_14628,N_14045);
or UO_1846 (O_1846,N_14668,N_14758);
nor UO_1847 (O_1847,N_14240,N_14457);
and UO_1848 (O_1848,N_14701,N_14977);
or UO_1849 (O_1849,N_14416,N_14629);
or UO_1850 (O_1850,N_14751,N_14620);
nand UO_1851 (O_1851,N_14330,N_14393);
and UO_1852 (O_1852,N_14064,N_14564);
nor UO_1853 (O_1853,N_14233,N_14901);
or UO_1854 (O_1854,N_14788,N_14170);
xor UO_1855 (O_1855,N_14465,N_14964);
nand UO_1856 (O_1856,N_14695,N_14825);
nand UO_1857 (O_1857,N_14187,N_14506);
or UO_1858 (O_1858,N_14532,N_14311);
and UO_1859 (O_1859,N_14296,N_14370);
or UO_1860 (O_1860,N_14074,N_14920);
and UO_1861 (O_1861,N_14903,N_14642);
nand UO_1862 (O_1862,N_14379,N_14249);
nand UO_1863 (O_1863,N_14659,N_14237);
or UO_1864 (O_1864,N_14946,N_14461);
and UO_1865 (O_1865,N_14860,N_14966);
nor UO_1866 (O_1866,N_14140,N_14529);
xor UO_1867 (O_1867,N_14898,N_14192);
nor UO_1868 (O_1868,N_14162,N_14709);
nor UO_1869 (O_1869,N_14282,N_14904);
xnor UO_1870 (O_1870,N_14459,N_14969);
or UO_1871 (O_1871,N_14390,N_14402);
and UO_1872 (O_1872,N_14842,N_14695);
nand UO_1873 (O_1873,N_14118,N_14302);
xnor UO_1874 (O_1874,N_14939,N_14673);
or UO_1875 (O_1875,N_14604,N_14211);
and UO_1876 (O_1876,N_14700,N_14947);
nor UO_1877 (O_1877,N_14888,N_14019);
and UO_1878 (O_1878,N_14198,N_14296);
nor UO_1879 (O_1879,N_14721,N_14353);
and UO_1880 (O_1880,N_14100,N_14189);
or UO_1881 (O_1881,N_14965,N_14812);
nand UO_1882 (O_1882,N_14377,N_14055);
or UO_1883 (O_1883,N_14543,N_14777);
or UO_1884 (O_1884,N_14749,N_14653);
or UO_1885 (O_1885,N_14206,N_14852);
and UO_1886 (O_1886,N_14083,N_14004);
nor UO_1887 (O_1887,N_14682,N_14852);
nor UO_1888 (O_1888,N_14545,N_14005);
nor UO_1889 (O_1889,N_14898,N_14656);
nand UO_1890 (O_1890,N_14396,N_14595);
or UO_1891 (O_1891,N_14745,N_14940);
nor UO_1892 (O_1892,N_14875,N_14130);
or UO_1893 (O_1893,N_14920,N_14145);
or UO_1894 (O_1894,N_14824,N_14786);
or UO_1895 (O_1895,N_14337,N_14158);
or UO_1896 (O_1896,N_14637,N_14678);
and UO_1897 (O_1897,N_14252,N_14886);
xor UO_1898 (O_1898,N_14176,N_14020);
and UO_1899 (O_1899,N_14374,N_14542);
and UO_1900 (O_1900,N_14133,N_14454);
or UO_1901 (O_1901,N_14037,N_14400);
and UO_1902 (O_1902,N_14210,N_14083);
or UO_1903 (O_1903,N_14072,N_14848);
or UO_1904 (O_1904,N_14973,N_14381);
or UO_1905 (O_1905,N_14064,N_14743);
nand UO_1906 (O_1906,N_14826,N_14207);
nand UO_1907 (O_1907,N_14432,N_14506);
or UO_1908 (O_1908,N_14385,N_14039);
nor UO_1909 (O_1909,N_14165,N_14920);
nand UO_1910 (O_1910,N_14611,N_14598);
or UO_1911 (O_1911,N_14859,N_14314);
nor UO_1912 (O_1912,N_14749,N_14365);
and UO_1913 (O_1913,N_14901,N_14563);
nor UO_1914 (O_1914,N_14452,N_14211);
nand UO_1915 (O_1915,N_14633,N_14778);
nand UO_1916 (O_1916,N_14236,N_14036);
nand UO_1917 (O_1917,N_14623,N_14073);
and UO_1918 (O_1918,N_14763,N_14233);
and UO_1919 (O_1919,N_14963,N_14972);
nand UO_1920 (O_1920,N_14154,N_14125);
nor UO_1921 (O_1921,N_14646,N_14327);
and UO_1922 (O_1922,N_14030,N_14025);
or UO_1923 (O_1923,N_14352,N_14342);
xor UO_1924 (O_1924,N_14347,N_14718);
or UO_1925 (O_1925,N_14480,N_14860);
or UO_1926 (O_1926,N_14910,N_14715);
nand UO_1927 (O_1927,N_14236,N_14843);
nand UO_1928 (O_1928,N_14401,N_14441);
and UO_1929 (O_1929,N_14445,N_14537);
or UO_1930 (O_1930,N_14840,N_14894);
nor UO_1931 (O_1931,N_14158,N_14041);
or UO_1932 (O_1932,N_14077,N_14936);
nand UO_1933 (O_1933,N_14655,N_14700);
nand UO_1934 (O_1934,N_14836,N_14878);
nor UO_1935 (O_1935,N_14790,N_14844);
or UO_1936 (O_1936,N_14293,N_14548);
nor UO_1937 (O_1937,N_14122,N_14938);
and UO_1938 (O_1938,N_14493,N_14132);
and UO_1939 (O_1939,N_14633,N_14802);
and UO_1940 (O_1940,N_14317,N_14349);
and UO_1941 (O_1941,N_14721,N_14259);
xor UO_1942 (O_1942,N_14883,N_14381);
and UO_1943 (O_1943,N_14495,N_14771);
and UO_1944 (O_1944,N_14944,N_14643);
nor UO_1945 (O_1945,N_14228,N_14829);
or UO_1946 (O_1946,N_14490,N_14913);
or UO_1947 (O_1947,N_14043,N_14666);
nand UO_1948 (O_1948,N_14740,N_14264);
nor UO_1949 (O_1949,N_14459,N_14944);
nor UO_1950 (O_1950,N_14536,N_14606);
and UO_1951 (O_1951,N_14525,N_14900);
or UO_1952 (O_1952,N_14829,N_14463);
nor UO_1953 (O_1953,N_14732,N_14655);
nor UO_1954 (O_1954,N_14690,N_14447);
nor UO_1955 (O_1955,N_14512,N_14773);
nor UO_1956 (O_1956,N_14036,N_14188);
or UO_1957 (O_1957,N_14698,N_14079);
nor UO_1958 (O_1958,N_14957,N_14417);
or UO_1959 (O_1959,N_14641,N_14697);
nor UO_1960 (O_1960,N_14992,N_14432);
nor UO_1961 (O_1961,N_14566,N_14284);
or UO_1962 (O_1962,N_14367,N_14022);
xnor UO_1963 (O_1963,N_14454,N_14098);
nor UO_1964 (O_1964,N_14774,N_14763);
nor UO_1965 (O_1965,N_14988,N_14005);
xnor UO_1966 (O_1966,N_14501,N_14241);
nor UO_1967 (O_1967,N_14774,N_14102);
nor UO_1968 (O_1968,N_14684,N_14467);
nor UO_1969 (O_1969,N_14579,N_14785);
and UO_1970 (O_1970,N_14416,N_14127);
nor UO_1971 (O_1971,N_14761,N_14516);
nor UO_1972 (O_1972,N_14878,N_14958);
nand UO_1973 (O_1973,N_14758,N_14757);
nor UO_1974 (O_1974,N_14222,N_14747);
nor UO_1975 (O_1975,N_14225,N_14080);
and UO_1976 (O_1976,N_14460,N_14161);
nor UO_1977 (O_1977,N_14110,N_14477);
and UO_1978 (O_1978,N_14849,N_14700);
or UO_1979 (O_1979,N_14056,N_14428);
nand UO_1980 (O_1980,N_14066,N_14132);
and UO_1981 (O_1981,N_14452,N_14016);
nor UO_1982 (O_1982,N_14965,N_14102);
xor UO_1983 (O_1983,N_14656,N_14276);
nand UO_1984 (O_1984,N_14566,N_14792);
nand UO_1985 (O_1985,N_14659,N_14243);
nor UO_1986 (O_1986,N_14461,N_14072);
or UO_1987 (O_1987,N_14635,N_14610);
nor UO_1988 (O_1988,N_14609,N_14483);
and UO_1989 (O_1989,N_14792,N_14930);
xnor UO_1990 (O_1990,N_14711,N_14280);
nand UO_1991 (O_1991,N_14171,N_14151);
and UO_1992 (O_1992,N_14866,N_14369);
nor UO_1993 (O_1993,N_14801,N_14180);
nor UO_1994 (O_1994,N_14781,N_14523);
nand UO_1995 (O_1995,N_14929,N_14189);
nand UO_1996 (O_1996,N_14586,N_14780);
xor UO_1997 (O_1997,N_14789,N_14228);
nand UO_1998 (O_1998,N_14614,N_14606);
and UO_1999 (O_1999,N_14209,N_14225);
endmodule