module basic_1000_10000_1500_5_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_833,In_199);
and U1 (N_1,In_696,In_248);
nor U2 (N_2,In_799,In_467);
and U3 (N_3,In_135,In_619);
and U4 (N_4,In_111,In_52);
nand U5 (N_5,In_536,In_98);
or U6 (N_6,In_877,In_126);
and U7 (N_7,In_582,In_965);
and U8 (N_8,In_943,In_798);
xor U9 (N_9,In_889,In_597);
and U10 (N_10,In_795,In_214);
or U11 (N_11,In_992,In_342);
nand U12 (N_12,In_923,In_263);
nand U13 (N_13,In_985,In_955);
nand U14 (N_14,In_269,In_870);
or U15 (N_15,In_846,In_80);
or U16 (N_16,In_181,In_821);
nor U17 (N_17,In_437,In_223);
nand U18 (N_18,In_625,In_447);
and U19 (N_19,In_499,In_91);
or U20 (N_20,In_986,In_410);
xnor U21 (N_21,In_497,In_634);
or U22 (N_22,In_903,In_577);
or U23 (N_23,In_152,In_188);
nor U24 (N_24,In_587,In_874);
xor U25 (N_25,In_86,In_501);
and U26 (N_26,In_537,In_106);
nand U27 (N_27,In_907,In_974);
nor U28 (N_28,In_809,In_288);
nor U29 (N_29,In_864,In_201);
nor U30 (N_30,In_995,In_443);
or U31 (N_31,In_975,In_706);
nand U32 (N_32,In_742,In_491);
and U33 (N_33,In_861,In_669);
or U34 (N_34,In_952,In_883);
nand U35 (N_35,In_891,In_145);
and U36 (N_36,In_568,In_811);
xor U37 (N_37,In_963,In_403);
and U38 (N_38,In_949,In_843);
nand U39 (N_39,In_748,In_487);
nand U40 (N_40,In_924,In_186);
nor U41 (N_41,In_946,In_378);
xnor U42 (N_42,In_740,In_412);
and U43 (N_43,In_588,In_901);
nand U44 (N_44,In_298,In_600);
or U45 (N_45,In_67,In_972);
xor U46 (N_46,In_656,In_520);
xnor U47 (N_47,In_761,In_739);
or U48 (N_48,In_319,In_234);
and U49 (N_49,In_778,In_277);
nor U50 (N_50,In_236,In_104);
xnor U51 (N_51,In_158,In_650);
nand U52 (N_52,In_708,In_76);
and U53 (N_53,In_21,In_917);
nand U54 (N_54,In_939,In_814);
nand U55 (N_55,In_123,In_139);
xor U56 (N_56,In_43,In_753);
or U57 (N_57,In_835,In_872);
nand U58 (N_58,In_215,In_289);
or U59 (N_59,In_959,In_449);
or U60 (N_60,In_562,In_482);
nand U61 (N_61,In_200,In_929);
or U62 (N_62,In_813,In_876);
and U63 (N_63,In_657,In_154);
or U64 (N_64,In_140,In_477);
nand U65 (N_65,In_39,In_859);
xnor U66 (N_66,In_405,In_324);
and U67 (N_67,In_572,In_341);
nor U68 (N_68,In_415,In_621);
nor U69 (N_69,In_167,In_693);
nor U70 (N_70,In_278,In_244);
or U71 (N_71,In_980,In_17);
xnor U72 (N_72,In_388,In_727);
and U73 (N_73,In_168,In_950);
nor U74 (N_74,In_579,In_287);
and U75 (N_75,In_810,In_559);
xnor U76 (N_76,In_141,In_225);
nor U77 (N_77,In_459,In_598);
nor U78 (N_78,In_113,In_496);
or U79 (N_79,In_430,In_383);
nand U80 (N_80,In_75,In_724);
or U81 (N_81,In_328,In_481);
nand U82 (N_82,In_348,In_681);
nand U83 (N_83,In_744,In_601);
xnor U84 (N_84,In_42,In_738);
nand U85 (N_85,In_33,In_602);
nor U86 (N_86,In_816,In_511);
and U87 (N_87,In_114,In_112);
nor U88 (N_88,In_60,In_984);
or U89 (N_89,In_30,In_393);
nor U90 (N_90,In_815,In_717);
and U91 (N_91,In_245,In_485);
nand U92 (N_92,In_309,In_591);
or U93 (N_93,In_573,In_228);
nand U94 (N_94,In_808,In_649);
and U95 (N_95,In_764,In_465);
nor U96 (N_96,In_732,In_221);
or U97 (N_97,In_541,In_590);
nor U98 (N_98,In_551,In_688);
and U99 (N_99,In_899,In_962);
and U100 (N_100,In_124,In_838);
or U101 (N_101,In_375,In_70);
nand U102 (N_102,In_564,In_19);
xnor U103 (N_103,In_531,In_928);
xor U104 (N_104,In_432,In_533);
or U105 (N_105,In_676,In_517);
xor U106 (N_106,In_323,In_61);
nor U107 (N_107,In_62,In_203);
or U108 (N_108,In_322,In_756);
xor U109 (N_109,In_989,In_902);
xor U110 (N_110,In_958,In_664);
or U111 (N_111,In_643,In_15);
and U112 (N_112,In_36,In_852);
or U113 (N_113,In_170,In_222);
nand U114 (N_114,In_295,In_208);
xor U115 (N_115,In_133,In_353);
nor U116 (N_116,In_519,In_930);
and U117 (N_117,In_697,In_489);
xor U118 (N_118,In_1,In_401);
and U119 (N_119,In_402,In_8);
nor U120 (N_120,In_291,In_824);
and U121 (N_121,In_646,In_9);
xnor U122 (N_122,In_906,In_580);
or U123 (N_123,In_720,In_78);
nand U124 (N_124,In_191,In_831);
or U125 (N_125,In_494,In_768);
or U126 (N_126,In_754,In_28);
xor U127 (N_127,In_911,In_49);
and U128 (N_128,In_174,In_888);
and U129 (N_129,In_645,In_913);
nand U130 (N_130,In_151,In_553);
nor U131 (N_131,In_421,In_780);
nor U132 (N_132,In_435,In_82);
xor U133 (N_133,In_468,In_612);
or U134 (N_134,In_63,In_853);
nand U135 (N_135,In_450,In_349);
and U136 (N_136,In_472,In_128);
or U137 (N_137,In_609,In_918);
and U138 (N_138,In_428,In_805);
xor U139 (N_139,In_436,In_411);
or U140 (N_140,In_414,In_318);
nand U141 (N_141,In_973,In_711);
or U142 (N_142,In_686,In_13);
and U143 (N_143,In_794,In_894);
nor U144 (N_144,In_534,In_565);
and U145 (N_145,In_781,In_555);
nand U146 (N_146,In_997,In_521);
or U147 (N_147,In_473,In_325);
nand U148 (N_148,In_292,In_95);
or U149 (N_149,In_599,In_674);
and U150 (N_150,In_272,In_660);
or U151 (N_151,In_77,In_760);
and U152 (N_152,In_26,In_108);
and U153 (N_153,In_610,In_212);
and U154 (N_154,In_66,In_624);
nor U155 (N_155,In_779,In_954);
nor U156 (N_156,In_953,In_823);
and U157 (N_157,In_125,In_187);
or U158 (N_158,In_440,In_211);
xor U159 (N_159,In_510,In_942);
xnor U160 (N_160,In_366,In_647);
xor U161 (N_161,In_528,In_190);
nand U162 (N_162,In_886,In_490);
and U163 (N_163,In_119,In_343);
and U164 (N_164,In_197,In_335);
and U165 (N_165,In_219,In_464);
and U166 (N_166,In_364,In_265);
and U167 (N_167,In_777,In_977);
xnor U168 (N_168,In_585,In_968);
and U169 (N_169,In_595,In_561);
nor U170 (N_170,In_249,In_458);
or U171 (N_171,In_546,In_293);
or U172 (N_172,In_849,In_189);
nor U173 (N_173,In_72,In_358);
and U174 (N_174,In_801,In_680);
xnor U175 (N_175,In_38,In_229);
xnor U176 (N_176,In_317,In_340);
and U177 (N_177,In_936,In_800);
and U178 (N_178,In_312,In_763);
nand U179 (N_179,In_790,In_539);
nand U180 (N_180,In_150,In_14);
nor U181 (N_181,In_793,In_850);
and U182 (N_182,In_661,In_429);
nor U183 (N_183,In_948,In_854);
or U184 (N_184,In_32,In_937);
nor U185 (N_185,In_932,In_178);
and U186 (N_186,In_180,In_50);
and U187 (N_187,In_981,In_444);
and U188 (N_188,In_31,In_784);
and U189 (N_189,In_767,In_788);
nand U190 (N_190,In_385,In_636);
xor U191 (N_191,In_479,In_507);
xnor U192 (N_192,In_659,In_177);
xnor U193 (N_193,In_502,In_392);
or U194 (N_194,In_716,In_702);
and U195 (N_195,In_550,In_842);
xor U196 (N_196,In_148,In_217);
nand U197 (N_197,In_185,In_545);
xor U198 (N_198,In_433,In_839);
or U199 (N_199,In_58,In_327);
nor U200 (N_200,In_99,In_857);
or U201 (N_201,In_6,In_136);
xor U202 (N_202,In_765,In_334);
or U203 (N_203,In_423,In_276);
xnor U204 (N_204,In_848,In_456);
xnor U205 (N_205,In_721,In_240);
or U206 (N_206,In_868,In_275);
or U207 (N_207,In_301,In_766);
nand U208 (N_208,In_500,In_408);
or U209 (N_209,In_184,In_605);
or U210 (N_210,In_284,In_990);
nor U211 (N_211,In_302,In_122);
and U212 (N_212,In_755,In_130);
xor U213 (N_213,In_653,In_161);
or U214 (N_214,In_804,In_478);
nor U215 (N_215,In_470,In_149);
and U216 (N_216,In_153,In_374);
and U217 (N_217,In_270,In_817);
or U218 (N_218,In_548,In_871);
and U219 (N_219,In_896,In_352);
and U220 (N_220,In_614,In_417);
or U221 (N_221,In_728,In_578);
and U222 (N_222,In_227,In_538);
or U223 (N_223,In_216,In_231);
or U224 (N_224,In_606,In_710);
xnor U225 (N_225,In_120,In_957);
and U226 (N_226,In_827,In_469);
xnor U227 (N_227,In_452,In_770);
nor U228 (N_228,In_569,In_925);
or U229 (N_229,In_747,In_514);
and U230 (N_230,In_723,In_685);
or U231 (N_231,In_271,In_55);
and U232 (N_232,In_68,In_644);
xnor U233 (N_233,In_395,In_836);
nand U234 (N_234,In_143,In_927);
nand U235 (N_235,In_785,In_27);
or U236 (N_236,In_282,In_549);
or U237 (N_237,In_407,In_841);
nand U238 (N_238,In_851,In_530);
nand U239 (N_239,In_819,In_751);
nor U240 (N_240,In_776,In_344);
nand U241 (N_241,In_97,In_2);
nor U242 (N_242,In_283,In_563);
nor U243 (N_243,In_757,In_107);
nor U244 (N_244,In_210,In_361);
xor U245 (N_245,In_329,In_247);
nor U246 (N_246,In_544,In_285);
and U247 (N_247,In_762,In_858);
xor U248 (N_248,In_637,In_183);
nor U249 (N_249,In_162,In_235);
or U250 (N_250,In_832,In_476);
or U251 (N_251,In_315,In_983);
or U252 (N_252,In_845,In_641);
nor U253 (N_253,In_782,In_442);
xor U254 (N_254,In_668,In_567);
nand U255 (N_255,In_867,In_424);
or U256 (N_256,In_892,In_23);
nand U257 (N_257,In_37,In_796);
nand U258 (N_258,In_369,In_338);
nand U259 (N_259,In_916,In_233);
and U260 (N_260,In_103,In_121);
xor U261 (N_261,In_455,In_310);
nand U262 (N_262,In_552,In_771);
nand U263 (N_263,In_791,In_812);
and U264 (N_264,In_583,In_689);
nand U265 (N_265,In_462,In_792);
nand U266 (N_266,In_956,In_991);
xnor U267 (N_267,In_475,In_743);
or U268 (N_268,In_193,In_694);
nand U269 (N_269,In_255,In_155);
xor U270 (N_270,In_759,In_999);
nand U271 (N_271,In_252,In_504);
nand U272 (N_272,In_752,In_44);
and U273 (N_273,In_856,In_53);
nand U274 (N_274,In_722,In_613);
and U275 (N_275,In_206,In_220);
nand U276 (N_276,In_59,In_797);
nand U277 (N_277,In_673,In_296);
nand U278 (N_278,In_806,In_390);
nand U279 (N_279,In_439,In_300);
nand U280 (N_280,In_243,In_789);
nand U281 (N_281,In_371,In_627);
and U282 (N_282,In_367,In_884);
or U283 (N_283,In_509,In_434);
and U284 (N_284,In_926,In_786);
nand U285 (N_285,In_41,In_346);
and U286 (N_286,In_608,In_313);
nor U287 (N_287,In_869,In_703);
and U288 (N_288,In_357,In_3);
and U289 (N_289,In_709,In_714);
or U290 (N_290,In_783,In_137);
and U291 (N_291,In_628,In_45);
nand U292 (N_292,In_74,In_273);
xor U293 (N_293,In_362,In_453);
nor U294 (N_294,In_438,In_527);
nand U295 (N_295,In_921,In_667);
nor U296 (N_296,In_640,In_182);
or U297 (N_297,In_994,In_626);
nand U298 (N_298,In_993,In_57);
nor U299 (N_299,In_830,In_264);
and U300 (N_300,In_967,In_20);
xor U301 (N_301,In_35,In_675);
and U302 (N_302,In_397,In_418);
or U303 (N_303,In_48,In_607);
and U304 (N_304,In_157,In_413);
nor U305 (N_305,In_242,In_132);
and U306 (N_306,In_844,In_982);
and U307 (N_307,In_314,In_718);
nand U308 (N_308,In_914,In_945);
nor U309 (N_309,In_18,In_204);
xnor U310 (N_310,In_46,In_701);
xnor U311 (N_311,In_198,In_679);
nand U312 (N_312,In_879,In_574);
or U313 (N_313,In_192,In_775);
nor U314 (N_314,In_90,In_279);
nand U315 (N_315,In_529,In_758);
xnor U316 (N_316,In_376,In_620);
or U317 (N_317,In_363,In_304);
and U318 (N_318,In_5,In_226);
or U319 (N_319,In_0,In_29);
nor U320 (N_320,In_540,In_426);
and U321 (N_321,In_508,In_652);
nor U322 (N_322,In_34,In_900);
nand U323 (N_323,In_735,In_678);
and U324 (N_324,In_7,In_360);
xor U325 (N_325,In_655,In_267);
nor U326 (N_326,In_73,In_332);
xor U327 (N_327,In_492,In_175);
xnor U328 (N_328,In_331,In_40);
or U329 (N_329,In_422,In_988);
or U330 (N_330,In_337,In_746);
and U331 (N_331,In_372,In_919);
nor U332 (N_332,In_505,In_268);
xor U333 (N_333,In_261,In_259);
nand U334 (N_334,In_750,In_594);
or U335 (N_335,In_909,In_825);
and U336 (N_336,In_399,In_966);
nand U337 (N_337,In_604,In_173);
and U338 (N_338,In_726,In_345);
nor U339 (N_339,In_166,In_241);
nand U340 (N_340,In_146,In_306);
nand U341 (N_341,In_622,In_257);
and U342 (N_342,In_557,In_651);
nand U343 (N_343,In_658,In_523);
and U344 (N_344,In_642,In_611);
or U345 (N_345,In_733,In_115);
and U346 (N_346,In_290,In_56);
xor U347 (N_347,In_951,In_513);
xnor U348 (N_348,In_774,In_488);
xor U349 (N_349,In_665,In_10);
xnor U350 (N_350,In_847,In_880);
xor U351 (N_351,In_142,In_575);
nand U352 (N_352,In_134,In_670);
nor U353 (N_353,In_230,In_617);
nor U354 (N_354,In_632,In_542);
or U355 (N_355,In_394,In_905);
nor U356 (N_356,In_976,In_165);
or U357 (N_357,In_51,In_725);
xor U358 (N_358,In_592,In_560);
nand U359 (N_359,In_71,In_89);
or U360 (N_360,In_695,In_603);
and U361 (N_361,In_730,In_885);
xnor U362 (N_362,In_878,In_589);
and U363 (N_363,In_209,In_355);
nand U364 (N_364,In_908,In_160);
xnor U365 (N_365,In_741,In_102);
or U366 (N_366,In_525,In_535);
xor U367 (N_367,In_895,In_159);
xor U368 (N_368,In_466,In_631);
and U369 (N_369,In_515,In_260);
and U370 (N_370,In_840,In_556);
nand U371 (N_371,In_281,In_196);
and U372 (N_372,In_558,In_630);
or U373 (N_373,In_941,In_299);
xnor U374 (N_374,In_969,In_205);
nand U375 (N_375,In_807,In_239);
or U376 (N_376,In_359,In_915);
and U377 (N_377,In_321,In_736);
xnor U378 (N_378,In_87,In_127);
xnor U379 (N_379,In_512,In_386);
or U380 (N_380,In_922,In_749);
nor U381 (N_381,In_910,In_84);
nor U382 (N_382,In_4,In_224);
xnor U383 (N_383,In_365,In_933);
nor U384 (N_384,In_368,In_65);
nand U385 (N_385,In_47,In_570);
nor U386 (N_386,In_860,In_409);
xnor U387 (N_387,In_446,In_866);
nor U388 (N_388,In_944,In_887);
xnor U389 (N_389,In_12,In_330);
and U390 (N_390,In_566,In_931);
nor U391 (N_391,In_493,In_109);
and U392 (N_392,In_638,In_96);
nor U393 (N_393,In_826,In_463);
nor U394 (N_394,In_22,In_863);
nor U395 (N_395,In_495,In_384);
and U396 (N_396,In_576,In_524);
and U397 (N_397,In_699,In_663);
nand U398 (N_398,In_404,In_169);
nand U399 (N_399,In_947,In_93);
xor U400 (N_400,In_54,In_94);
nor U401 (N_401,In_875,In_677);
nand U402 (N_402,In_461,In_581);
nand U403 (N_403,In_339,In_303);
nand U404 (N_404,In_266,In_246);
and U405 (N_405,In_380,In_391);
or U406 (N_406,In_769,In_882);
xnor U407 (N_407,In_996,In_498);
and U408 (N_408,In_970,In_897);
and U409 (N_409,In_305,In_172);
or U410 (N_410,In_81,In_406);
xor U411 (N_411,In_554,In_398);
xnor U412 (N_412,In_690,In_971);
xnor U413 (N_413,In_639,In_547);
xnor U414 (N_414,In_961,In_262);
nand U415 (N_415,In_862,In_336);
or U416 (N_416,In_448,In_129);
or U417 (N_417,In_987,In_828);
and U418 (N_418,In_593,In_297);
nand U419 (N_419,In_350,In_171);
nand U420 (N_420,In_818,In_280);
nor U421 (N_421,In_138,In_719);
xnor U422 (N_422,In_506,In_745);
and U423 (N_423,In_633,In_881);
or U424 (N_424,In_938,In_503);
and U425 (N_425,In_773,In_457);
nor U426 (N_426,In_935,In_347);
and U427 (N_427,In_890,In_253);
and U428 (N_428,In_416,In_731);
nand U429 (N_429,In_427,In_964);
xnor U430 (N_430,In_176,In_307);
nand U431 (N_431,In_802,In_734);
and U432 (N_432,In_195,In_131);
nand U433 (N_433,In_940,In_202);
nor U434 (N_434,In_682,In_381);
and U435 (N_435,In_483,In_311);
or U436 (N_436,In_379,In_420);
xor U437 (N_437,In_616,In_454);
or U438 (N_438,In_715,In_912);
or U439 (N_439,In_586,In_855);
and U440 (N_440,In_354,In_460);
or U441 (N_441,In_308,In_232);
or U442 (N_442,In_474,In_400);
xnor U443 (N_443,In_865,In_772);
and U444 (N_444,In_904,In_101);
nand U445 (N_445,In_213,In_571);
nand U446 (N_446,In_671,In_445);
xor U447 (N_447,In_672,In_687);
xnor U448 (N_448,In_700,In_834);
nand U449 (N_449,In_618,In_156);
or U450 (N_450,In_373,In_526);
nor U451 (N_451,In_584,In_286);
nor U452 (N_452,In_237,In_419);
nand U453 (N_453,In_707,In_666);
and U454 (N_454,In_387,In_471);
and U455 (N_455,In_635,In_820);
nor U456 (N_456,In_274,In_898);
nand U457 (N_457,In_88,In_164);
xor U458 (N_458,In_396,In_370);
nor U459 (N_459,In_79,In_333);
nand U460 (N_460,In_698,In_648);
xnor U461 (N_461,In_654,In_729);
xnor U462 (N_462,In_934,In_829);
nand U463 (N_463,In_147,In_662);
or U464 (N_464,In_486,In_451);
or U465 (N_465,In_979,In_684);
nor U466 (N_466,In_83,In_250);
xor U467 (N_467,In_144,In_16);
or U468 (N_468,In_377,In_431);
and U469 (N_469,In_24,In_105);
or U470 (N_470,In_320,In_532);
and U471 (N_471,In_683,In_629);
or U472 (N_472,In_692,In_382);
nand U473 (N_473,In_518,In_117);
nor U474 (N_474,In_998,In_163);
or U475 (N_475,In_207,In_251);
and U476 (N_476,In_596,In_11);
nor U477 (N_477,In_787,In_258);
and U478 (N_478,In_615,In_351);
or U479 (N_479,In_893,In_256);
nand U480 (N_480,In_704,In_118);
nand U481 (N_481,In_441,In_978);
xnor U482 (N_482,In_712,In_705);
nor U483 (N_483,In_194,In_356);
or U484 (N_484,In_64,In_920);
nand U485 (N_485,In_822,In_543);
nor U486 (N_486,In_179,In_737);
and U487 (N_487,In_837,In_92);
xor U488 (N_488,In_254,In_85);
nor U489 (N_489,In_218,In_326);
nor U490 (N_490,In_516,In_425);
xnor U491 (N_491,In_389,In_623);
nor U492 (N_492,In_522,In_803);
xor U493 (N_493,In_110,In_69);
nand U494 (N_494,In_713,In_691);
xnor U495 (N_495,In_116,In_316);
or U496 (N_496,In_25,In_480);
or U497 (N_497,In_873,In_238);
nor U498 (N_498,In_484,In_960);
and U499 (N_499,In_100,In_294);
nand U500 (N_500,In_68,In_522);
nand U501 (N_501,In_525,In_871);
and U502 (N_502,In_885,In_964);
xor U503 (N_503,In_29,In_923);
nor U504 (N_504,In_628,In_836);
xnor U505 (N_505,In_196,In_314);
or U506 (N_506,In_869,In_464);
xor U507 (N_507,In_279,In_954);
and U508 (N_508,In_425,In_751);
and U509 (N_509,In_18,In_696);
xnor U510 (N_510,In_372,In_758);
nor U511 (N_511,In_44,In_550);
xor U512 (N_512,In_34,In_114);
or U513 (N_513,In_290,In_190);
and U514 (N_514,In_174,In_426);
nand U515 (N_515,In_358,In_652);
nand U516 (N_516,In_188,In_983);
nor U517 (N_517,In_280,In_916);
or U518 (N_518,In_134,In_262);
nor U519 (N_519,In_632,In_596);
nand U520 (N_520,In_471,In_289);
xor U521 (N_521,In_254,In_436);
or U522 (N_522,In_798,In_132);
or U523 (N_523,In_633,In_812);
nand U524 (N_524,In_691,In_495);
and U525 (N_525,In_424,In_793);
and U526 (N_526,In_942,In_432);
xor U527 (N_527,In_602,In_774);
nor U528 (N_528,In_740,In_843);
and U529 (N_529,In_363,In_707);
nor U530 (N_530,In_646,In_992);
and U531 (N_531,In_319,In_395);
nor U532 (N_532,In_410,In_402);
or U533 (N_533,In_554,In_156);
nand U534 (N_534,In_704,In_500);
xnor U535 (N_535,In_306,In_645);
xor U536 (N_536,In_445,In_837);
or U537 (N_537,In_745,In_422);
and U538 (N_538,In_796,In_416);
and U539 (N_539,In_808,In_384);
or U540 (N_540,In_741,In_179);
or U541 (N_541,In_755,In_290);
nor U542 (N_542,In_972,In_589);
xnor U543 (N_543,In_8,In_348);
nand U544 (N_544,In_22,In_326);
nand U545 (N_545,In_994,In_533);
xnor U546 (N_546,In_96,In_804);
or U547 (N_547,In_677,In_941);
or U548 (N_548,In_390,In_807);
nand U549 (N_549,In_916,In_942);
and U550 (N_550,In_412,In_145);
or U551 (N_551,In_463,In_364);
nor U552 (N_552,In_96,In_294);
or U553 (N_553,In_339,In_495);
xnor U554 (N_554,In_453,In_128);
nand U555 (N_555,In_814,In_145);
or U556 (N_556,In_826,In_646);
nand U557 (N_557,In_625,In_823);
nor U558 (N_558,In_413,In_451);
nand U559 (N_559,In_417,In_295);
nor U560 (N_560,In_28,In_405);
or U561 (N_561,In_206,In_45);
nor U562 (N_562,In_628,In_272);
and U563 (N_563,In_292,In_368);
xnor U564 (N_564,In_486,In_318);
nor U565 (N_565,In_1,In_944);
nor U566 (N_566,In_660,In_334);
nand U567 (N_567,In_915,In_976);
xor U568 (N_568,In_277,In_353);
and U569 (N_569,In_834,In_221);
or U570 (N_570,In_511,In_989);
xor U571 (N_571,In_851,In_232);
and U572 (N_572,In_722,In_187);
or U573 (N_573,In_164,In_801);
nand U574 (N_574,In_30,In_853);
and U575 (N_575,In_513,In_114);
or U576 (N_576,In_809,In_947);
nor U577 (N_577,In_50,In_395);
and U578 (N_578,In_433,In_578);
xor U579 (N_579,In_989,In_72);
xnor U580 (N_580,In_982,In_551);
and U581 (N_581,In_829,In_538);
and U582 (N_582,In_685,In_486);
xnor U583 (N_583,In_621,In_858);
nor U584 (N_584,In_219,In_132);
xor U585 (N_585,In_851,In_926);
nand U586 (N_586,In_159,In_56);
xnor U587 (N_587,In_894,In_665);
xnor U588 (N_588,In_215,In_59);
xor U589 (N_589,In_724,In_398);
nor U590 (N_590,In_676,In_441);
or U591 (N_591,In_380,In_717);
nor U592 (N_592,In_533,In_443);
nor U593 (N_593,In_369,In_511);
and U594 (N_594,In_470,In_749);
or U595 (N_595,In_277,In_791);
and U596 (N_596,In_962,In_334);
or U597 (N_597,In_291,In_490);
xnor U598 (N_598,In_5,In_858);
nand U599 (N_599,In_108,In_46);
nor U600 (N_600,In_280,In_682);
and U601 (N_601,In_967,In_417);
and U602 (N_602,In_885,In_820);
or U603 (N_603,In_803,In_319);
and U604 (N_604,In_113,In_102);
xnor U605 (N_605,In_274,In_523);
nor U606 (N_606,In_526,In_630);
and U607 (N_607,In_603,In_77);
or U608 (N_608,In_68,In_505);
xor U609 (N_609,In_657,In_442);
and U610 (N_610,In_97,In_460);
nor U611 (N_611,In_435,In_588);
and U612 (N_612,In_921,In_742);
nor U613 (N_613,In_21,In_864);
or U614 (N_614,In_899,In_684);
nor U615 (N_615,In_710,In_53);
xor U616 (N_616,In_579,In_751);
nor U617 (N_617,In_273,In_992);
nand U618 (N_618,In_729,In_10);
xnor U619 (N_619,In_201,In_477);
xor U620 (N_620,In_527,In_297);
or U621 (N_621,In_691,In_370);
nand U622 (N_622,In_14,In_1);
xnor U623 (N_623,In_3,In_735);
and U624 (N_624,In_842,In_587);
xor U625 (N_625,In_536,In_978);
and U626 (N_626,In_255,In_201);
nand U627 (N_627,In_443,In_426);
nand U628 (N_628,In_583,In_740);
nor U629 (N_629,In_12,In_357);
nor U630 (N_630,In_926,In_718);
nand U631 (N_631,In_812,In_50);
or U632 (N_632,In_440,In_550);
xnor U633 (N_633,In_624,In_875);
or U634 (N_634,In_989,In_76);
and U635 (N_635,In_995,In_97);
nand U636 (N_636,In_326,In_241);
xor U637 (N_637,In_116,In_804);
nand U638 (N_638,In_108,In_772);
or U639 (N_639,In_758,In_332);
nor U640 (N_640,In_75,In_331);
xor U641 (N_641,In_200,In_865);
nand U642 (N_642,In_305,In_589);
nor U643 (N_643,In_809,In_311);
and U644 (N_644,In_192,In_129);
xor U645 (N_645,In_634,In_260);
and U646 (N_646,In_321,In_778);
nor U647 (N_647,In_283,In_848);
and U648 (N_648,In_59,In_55);
nand U649 (N_649,In_844,In_428);
or U650 (N_650,In_921,In_957);
or U651 (N_651,In_688,In_649);
nand U652 (N_652,In_739,In_589);
nand U653 (N_653,In_195,In_369);
xor U654 (N_654,In_956,In_356);
xor U655 (N_655,In_365,In_416);
xnor U656 (N_656,In_302,In_895);
xnor U657 (N_657,In_133,In_998);
nand U658 (N_658,In_214,In_577);
xor U659 (N_659,In_193,In_716);
or U660 (N_660,In_853,In_100);
and U661 (N_661,In_132,In_899);
xor U662 (N_662,In_286,In_495);
xnor U663 (N_663,In_657,In_810);
or U664 (N_664,In_625,In_258);
xnor U665 (N_665,In_29,In_181);
nor U666 (N_666,In_548,In_857);
and U667 (N_667,In_301,In_176);
and U668 (N_668,In_793,In_299);
or U669 (N_669,In_364,In_425);
and U670 (N_670,In_633,In_486);
and U671 (N_671,In_926,In_50);
and U672 (N_672,In_45,In_215);
and U673 (N_673,In_286,In_837);
nor U674 (N_674,In_806,In_874);
xor U675 (N_675,In_83,In_814);
nor U676 (N_676,In_155,In_430);
or U677 (N_677,In_390,In_460);
or U678 (N_678,In_890,In_883);
xnor U679 (N_679,In_846,In_843);
nor U680 (N_680,In_104,In_736);
xnor U681 (N_681,In_481,In_586);
nor U682 (N_682,In_331,In_704);
xnor U683 (N_683,In_740,In_500);
and U684 (N_684,In_610,In_432);
xnor U685 (N_685,In_800,In_645);
nand U686 (N_686,In_416,In_968);
nand U687 (N_687,In_286,In_392);
xnor U688 (N_688,In_801,In_425);
xnor U689 (N_689,In_936,In_611);
and U690 (N_690,In_921,In_101);
nand U691 (N_691,In_892,In_990);
nor U692 (N_692,In_965,In_493);
nor U693 (N_693,In_93,In_606);
nor U694 (N_694,In_930,In_348);
or U695 (N_695,In_97,In_478);
xnor U696 (N_696,In_188,In_687);
or U697 (N_697,In_89,In_109);
or U698 (N_698,In_147,In_668);
and U699 (N_699,In_655,In_428);
xnor U700 (N_700,In_866,In_304);
nand U701 (N_701,In_619,In_208);
or U702 (N_702,In_832,In_155);
xor U703 (N_703,In_487,In_881);
nand U704 (N_704,In_94,In_601);
and U705 (N_705,In_938,In_767);
and U706 (N_706,In_372,In_819);
nand U707 (N_707,In_571,In_908);
xnor U708 (N_708,In_865,In_361);
and U709 (N_709,In_378,In_587);
and U710 (N_710,In_297,In_364);
nand U711 (N_711,In_61,In_706);
nand U712 (N_712,In_238,In_401);
or U713 (N_713,In_38,In_522);
nor U714 (N_714,In_11,In_514);
and U715 (N_715,In_731,In_720);
nand U716 (N_716,In_840,In_877);
nor U717 (N_717,In_681,In_743);
nor U718 (N_718,In_919,In_611);
nor U719 (N_719,In_685,In_421);
xor U720 (N_720,In_584,In_396);
and U721 (N_721,In_783,In_428);
nand U722 (N_722,In_424,In_812);
nor U723 (N_723,In_797,In_573);
or U724 (N_724,In_471,In_293);
and U725 (N_725,In_157,In_827);
xnor U726 (N_726,In_449,In_337);
or U727 (N_727,In_235,In_280);
nor U728 (N_728,In_430,In_443);
or U729 (N_729,In_28,In_988);
nand U730 (N_730,In_697,In_877);
and U731 (N_731,In_645,In_721);
and U732 (N_732,In_704,In_391);
and U733 (N_733,In_430,In_666);
and U734 (N_734,In_841,In_978);
nor U735 (N_735,In_384,In_786);
nor U736 (N_736,In_782,In_703);
nor U737 (N_737,In_973,In_250);
nor U738 (N_738,In_641,In_494);
or U739 (N_739,In_936,In_678);
and U740 (N_740,In_403,In_756);
and U741 (N_741,In_115,In_333);
or U742 (N_742,In_720,In_285);
xor U743 (N_743,In_643,In_129);
nor U744 (N_744,In_923,In_734);
nand U745 (N_745,In_66,In_794);
or U746 (N_746,In_290,In_642);
and U747 (N_747,In_66,In_557);
and U748 (N_748,In_467,In_780);
and U749 (N_749,In_429,In_921);
and U750 (N_750,In_337,In_187);
and U751 (N_751,In_230,In_319);
and U752 (N_752,In_735,In_22);
nor U753 (N_753,In_154,In_267);
nor U754 (N_754,In_573,In_555);
and U755 (N_755,In_797,In_865);
xor U756 (N_756,In_18,In_108);
or U757 (N_757,In_523,In_33);
nand U758 (N_758,In_281,In_908);
or U759 (N_759,In_298,In_978);
nor U760 (N_760,In_606,In_51);
and U761 (N_761,In_922,In_733);
nand U762 (N_762,In_528,In_874);
and U763 (N_763,In_989,In_265);
or U764 (N_764,In_217,In_70);
and U765 (N_765,In_419,In_631);
or U766 (N_766,In_230,In_852);
or U767 (N_767,In_309,In_529);
nor U768 (N_768,In_95,In_704);
nor U769 (N_769,In_55,In_663);
nor U770 (N_770,In_125,In_633);
xnor U771 (N_771,In_208,In_882);
or U772 (N_772,In_238,In_817);
xnor U773 (N_773,In_259,In_553);
or U774 (N_774,In_778,In_722);
and U775 (N_775,In_998,In_852);
and U776 (N_776,In_813,In_309);
and U777 (N_777,In_852,In_394);
or U778 (N_778,In_94,In_482);
xor U779 (N_779,In_950,In_642);
nor U780 (N_780,In_892,In_326);
nor U781 (N_781,In_394,In_91);
nor U782 (N_782,In_362,In_225);
xnor U783 (N_783,In_950,In_974);
nor U784 (N_784,In_618,In_319);
nand U785 (N_785,In_402,In_311);
and U786 (N_786,In_997,In_647);
xnor U787 (N_787,In_409,In_249);
nand U788 (N_788,In_259,In_117);
and U789 (N_789,In_888,In_864);
nor U790 (N_790,In_825,In_464);
nand U791 (N_791,In_160,In_528);
or U792 (N_792,In_394,In_296);
and U793 (N_793,In_646,In_236);
nand U794 (N_794,In_324,In_453);
and U795 (N_795,In_617,In_442);
or U796 (N_796,In_881,In_322);
nand U797 (N_797,In_252,In_944);
xnor U798 (N_798,In_777,In_125);
nor U799 (N_799,In_544,In_53);
xnor U800 (N_800,In_633,In_776);
nor U801 (N_801,In_667,In_628);
nor U802 (N_802,In_850,In_923);
nand U803 (N_803,In_691,In_796);
xnor U804 (N_804,In_239,In_977);
nor U805 (N_805,In_30,In_684);
nand U806 (N_806,In_325,In_506);
nor U807 (N_807,In_652,In_879);
xnor U808 (N_808,In_580,In_495);
and U809 (N_809,In_708,In_64);
and U810 (N_810,In_877,In_562);
xnor U811 (N_811,In_321,In_441);
xor U812 (N_812,In_769,In_579);
and U813 (N_813,In_86,In_685);
or U814 (N_814,In_920,In_957);
nor U815 (N_815,In_419,In_937);
nand U816 (N_816,In_197,In_56);
nor U817 (N_817,In_507,In_33);
xor U818 (N_818,In_578,In_820);
or U819 (N_819,In_958,In_312);
and U820 (N_820,In_475,In_965);
xor U821 (N_821,In_775,In_87);
xnor U822 (N_822,In_557,In_488);
xnor U823 (N_823,In_698,In_173);
or U824 (N_824,In_763,In_663);
or U825 (N_825,In_262,In_479);
xor U826 (N_826,In_256,In_706);
xor U827 (N_827,In_146,In_771);
xnor U828 (N_828,In_150,In_145);
or U829 (N_829,In_269,In_757);
xnor U830 (N_830,In_229,In_55);
nand U831 (N_831,In_362,In_149);
nand U832 (N_832,In_77,In_508);
and U833 (N_833,In_479,In_257);
and U834 (N_834,In_323,In_624);
nand U835 (N_835,In_118,In_76);
xnor U836 (N_836,In_282,In_703);
nor U837 (N_837,In_932,In_2);
xor U838 (N_838,In_855,In_465);
xor U839 (N_839,In_590,In_540);
or U840 (N_840,In_524,In_753);
nand U841 (N_841,In_600,In_348);
or U842 (N_842,In_87,In_588);
nor U843 (N_843,In_639,In_781);
xor U844 (N_844,In_875,In_20);
xor U845 (N_845,In_861,In_729);
nor U846 (N_846,In_226,In_607);
nand U847 (N_847,In_665,In_945);
xnor U848 (N_848,In_827,In_271);
xnor U849 (N_849,In_707,In_742);
nand U850 (N_850,In_276,In_692);
nor U851 (N_851,In_595,In_793);
nor U852 (N_852,In_460,In_620);
nor U853 (N_853,In_78,In_975);
and U854 (N_854,In_598,In_538);
nor U855 (N_855,In_357,In_190);
or U856 (N_856,In_427,In_530);
xnor U857 (N_857,In_795,In_21);
or U858 (N_858,In_850,In_144);
or U859 (N_859,In_2,In_429);
or U860 (N_860,In_189,In_526);
nor U861 (N_861,In_11,In_450);
xor U862 (N_862,In_167,In_272);
and U863 (N_863,In_957,In_324);
or U864 (N_864,In_640,In_451);
nand U865 (N_865,In_826,In_992);
or U866 (N_866,In_385,In_488);
nand U867 (N_867,In_339,In_955);
xnor U868 (N_868,In_141,In_206);
and U869 (N_869,In_804,In_86);
or U870 (N_870,In_867,In_902);
xor U871 (N_871,In_940,In_992);
nor U872 (N_872,In_41,In_914);
and U873 (N_873,In_864,In_566);
and U874 (N_874,In_36,In_371);
or U875 (N_875,In_676,In_819);
and U876 (N_876,In_834,In_691);
xor U877 (N_877,In_962,In_360);
nor U878 (N_878,In_394,In_231);
or U879 (N_879,In_306,In_178);
nand U880 (N_880,In_711,In_503);
xor U881 (N_881,In_361,In_551);
or U882 (N_882,In_573,In_818);
nand U883 (N_883,In_571,In_214);
nand U884 (N_884,In_247,In_406);
or U885 (N_885,In_410,In_690);
xor U886 (N_886,In_312,In_338);
or U887 (N_887,In_646,In_249);
and U888 (N_888,In_266,In_238);
and U889 (N_889,In_335,In_746);
or U890 (N_890,In_897,In_646);
and U891 (N_891,In_908,In_228);
nand U892 (N_892,In_383,In_722);
nor U893 (N_893,In_787,In_640);
xor U894 (N_894,In_452,In_905);
xor U895 (N_895,In_214,In_392);
nor U896 (N_896,In_586,In_777);
nand U897 (N_897,In_977,In_767);
or U898 (N_898,In_294,In_289);
nand U899 (N_899,In_527,In_890);
nand U900 (N_900,In_397,In_867);
or U901 (N_901,In_820,In_48);
and U902 (N_902,In_728,In_46);
xor U903 (N_903,In_692,In_917);
nor U904 (N_904,In_757,In_569);
and U905 (N_905,In_347,In_927);
nor U906 (N_906,In_628,In_551);
xor U907 (N_907,In_790,In_829);
nor U908 (N_908,In_317,In_914);
and U909 (N_909,In_907,In_437);
nand U910 (N_910,In_362,In_897);
or U911 (N_911,In_250,In_569);
or U912 (N_912,In_788,In_255);
nand U913 (N_913,In_335,In_804);
nor U914 (N_914,In_392,In_610);
nand U915 (N_915,In_996,In_516);
nor U916 (N_916,In_981,In_870);
xnor U917 (N_917,In_436,In_617);
xnor U918 (N_918,In_839,In_679);
nand U919 (N_919,In_642,In_560);
or U920 (N_920,In_340,In_655);
nor U921 (N_921,In_501,In_491);
xnor U922 (N_922,In_7,In_927);
or U923 (N_923,In_670,In_128);
xor U924 (N_924,In_685,In_463);
or U925 (N_925,In_452,In_563);
nand U926 (N_926,In_975,In_173);
or U927 (N_927,In_931,In_297);
or U928 (N_928,In_349,In_311);
nand U929 (N_929,In_302,In_351);
xnor U930 (N_930,In_871,In_273);
xnor U931 (N_931,In_975,In_634);
xor U932 (N_932,In_278,In_24);
and U933 (N_933,In_75,In_394);
and U934 (N_934,In_979,In_882);
and U935 (N_935,In_737,In_283);
and U936 (N_936,In_923,In_772);
and U937 (N_937,In_390,In_951);
and U938 (N_938,In_80,In_183);
nor U939 (N_939,In_978,In_252);
nor U940 (N_940,In_246,In_924);
xnor U941 (N_941,In_285,In_589);
xor U942 (N_942,In_920,In_926);
or U943 (N_943,In_15,In_138);
nor U944 (N_944,In_379,In_62);
nor U945 (N_945,In_974,In_298);
and U946 (N_946,In_56,In_715);
nand U947 (N_947,In_438,In_954);
or U948 (N_948,In_917,In_821);
or U949 (N_949,In_877,In_954);
or U950 (N_950,In_714,In_20);
nand U951 (N_951,In_858,In_890);
nor U952 (N_952,In_419,In_578);
xnor U953 (N_953,In_3,In_132);
nand U954 (N_954,In_715,In_292);
or U955 (N_955,In_450,In_124);
xnor U956 (N_956,In_577,In_720);
xor U957 (N_957,In_412,In_639);
or U958 (N_958,In_988,In_229);
or U959 (N_959,In_254,In_914);
or U960 (N_960,In_801,In_702);
and U961 (N_961,In_963,In_472);
xnor U962 (N_962,In_708,In_143);
nand U963 (N_963,In_389,In_828);
or U964 (N_964,In_758,In_614);
or U965 (N_965,In_820,In_399);
nor U966 (N_966,In_782,In_571);
nor U967 (N_967,In_975,In_130);
and U968 (N_968,In_13,In_957);
nand U969 (N_969,In_298,In_238);
xnor U970 (N_970,In_134,In_109);
nor U971 (N_971,In_778,In_121);
nand U972 (N_972,In_669,In_773);
nor U973 (N_973,In_269,In_952);
nand U974 (N_974,In_343,In_634);
nand U975 (N_975,In_648,In_497);
xnor U976 (N_976,In_103,In_854);
nor U977 (N_977,In_533,In_76);
nor U978 (N_978,In_235,In_502);
or U979 (N_979,In_135,In_5);
xnor U980 (N_980,In_367,In_401);
xor U981 (N_981,In_926,In_900);
and U982 (N_982,In_36,In_373);
and U983 (N_983,In_998,In_356);
nor U984 (N_984,In_350,In_924);
nor U985 (N_985,In_506,In_974);
or U986 (N_986,In_268,In_910);
and U987 (N_987,In_363,In_462);
nand U988 (N_988,In_224,In_228);
nand U989 (N_989,In_835,In_465);
xnor U990 (N_990,In_59,In_532);
or U991 (N_991,In_532,In_238);
xnor U992 (N_992,In_403,In_98);
or U993 (N_993,In_931,In_627);
and U994 (N_994,In_903,In_691);
or U995 (N_995,In_38,In_199);
xor U996 (N_996,In_878,In_842);
xor U997 (N_997,In_719,In_213);
xnor U998 (N_998,In_443,In_188);
nor U999 (N_999,In_722,In_33);
nor U1000 (N_1000,In_204,In_457);
and U1001 (N_1001,In_170,In_600);
or U1002 (N_1002,In_30,In_422);
xor U1003 (N_1003,In_641,In_135);
xor U1004 (N_1004,In_392,In_411);
nor U1005 (N_1005,In_345,In_618);
and U1006 (N_1006,In_687,In_926);
or U1007 (N_1007,In_572,In_57);
or U1008 (N_1008,In_414,In_894);
and U1009 (N_1009,In_739,In_374);
or U1010 (N_1010,In_146,In_840);
or U1011 (N_1011,In_428,In_400);
and U1012 (N_1012,In_704,In_648);
xnor U1013 (N_1013,In_911,In_63);
xnor U1014 (N_1014,In_31,In_832);
or U1015 (N_1015,In_193,In_751);
and U1016 (N_1016,In_528,In_759);
or U1017 (N_1017,In_71,In_817);
and U1018 (N_1018,In_5,In_988);
and U1019 (N_1019,In_839,In_250);
and U1020 (N_1020,In_641,In_59);
nor U1021 (N_1021,In_559,In_618);
nor U1022 (N_1022,In_217,In_433);
xnor U1023 (N_1023,In_79,In_269);
nand U1024 (N_1024,In_714,In_198);
nand U1025 (N_1025,In_472,In_911);
xnor U1026 (N_1026,In_378,In_437);
and U1027 (N_1027,In_199,In_829);
nor U1028 (N_1028,In_523,In_915);
or U1029 (N_1029,In_205,In_166);
and U1030 (N_1030,In_281,In_775);
nand U1031 (N_1031,In_868,In_825);
nand U1032 (N_1032,In_927,In_979);
or U1033 (N_1033,In_560,In_172);
nor U1034 (N_1034,In_115,In_491);
and U1035 (N_1035,In_809,In_617);
and U1036 (N_1036,In_240,In_907);
nor U1037 (N_1037,In_29,In_186);
or U1038 (N_1038,In_493,In_991);
or U1039 (N_1039,In_839,In_68);
nand U1040 (N_1040,In_949,In_672);
xor U1041 (N_1041,In_636,In_536);
xor U1042 (N_1042,In_116,In_782);
nand U1043 (N_1043,In_929,In_857);
nor U1044 (N_1044,In_858,In_270);
nand U1045 (N_1045,In_37,In_59);
and U1046 (N_1046,In_785,In_129);
or U1047 (N_1047,In_395,In_364);
nor U1048 (N_1048,In_623,In_261);
and U1049 (N_1049,In_46,In_471);
nor U1050 (N_1050,In_216,In_120);
or U1051 (N_1051,In_125,In_860);
nand U1052 (N_1052,In_197,In_351);
and U1053 (N_1053,In_791,In_831);
and U1054 (N_1054,In_804,In_538);
or U1055 (N_1055,In_825,In_290);
and U1056 (N_1056,In_532,In_729);
or U1057 (N_1057,In_701,In_308);
nor U1058 (N_1058,In_869,In_968);
and U1059 (N_1059,In_659,In_262);
nor U1060 (N_1060,In_743,In_187);
or U1061 (N_1061,In_348,In_160);
and U1062 (N_1062,In_800,In_426);
and U1063 (N_1063,In_851,In_702);
xnor U1064 (N_1064,In_356,In_135);
nand U1065 (N_1065,In_11,In_686);
nor U1066 (N_1066,In_512,In_607);
nand U1067 (N_1067,In_135,In_399);
xnor U1068 (N_1068,In_56,In_396);
and U1069 (N_1069,In_232,In_869);
xnor U1070 (N_1070,In_894,In_259);
xor U1071 (N_1071,In_404,In_104);
nor U1072 (N_1072,In_29,In_496);
xor U1073 (N_1073,In_602,In_911);
nand U1074 (N_1074,In_20,In_719);
nor U1075 (N_1075,In_929,In_12);
nand U1076 (N_1076,In_444,In_911);
nand U1077 (N_1077,In_710,In_368);
xnor U1078 (N_1078,In_747,In_496);
or U1079 (N_1079,In_640,In_526);
xor U1080 (N_1080,In_629,In_68);
nor U1081 (N_1081,In_757,In_994);
xor U1082 (N_1082,In_960,In_308);
xor U1083 (N_1083,In_893,In_656);
and U1084 (N_1084,In_578,In_814);
nor U1085 (N_1085,In_499,In_41);
xor U1086 (N_1086,In_490,In_63);
and U1087 (N_1087,In_321,In_493);
nand U1088 (N_1088,In_346,In_569);
or U1089 (N_1089,In_746,In_665);
xnor U1090 (N_1090,In_708,In_390);
nor U1091 (N_1091,In_774,In_351);
nor U1092 (N_1092,In_937,In_395);
and U1093 (N_1093,In_68,In_88);
or U1094 (N_1094,In_166,In_67);
xor U1095 (N_1095,In_175,In_185);
nand U1096 (N_1096,In_880,In_88);
xnor U1097 (N_1097,In_371,In_842);
nand U1098 (N_1098,In_987,In_684);
xor U1099 (N_1099,In_157,In_131);
or U1100 (N_1100,In_103,In_925);
nand U1101 (N_1101,In_365,In_571);
nand U1102 (N_1102,In_657,In_541);
and U1103 (N_1103,In_830,In_144);
xor U1104 (N_1104,In_549,In_121);
and U1105 (N_1105,In_181,In_616);
nor U1106 (N_1106,In_144,In_563);
nand U1107 (N_1107,In_671,In_356);
nor U1108 (N_1108,In_680,In_947);
xnor U1109 (N_1109,In_441,In_13);
xor U1110 (N_1110,In_262,In_540);
and U1111 (N_1111,In_975,In_217);
xor U1112 (N_1112,In_670,In_618);
nor U1113 (N_1113,In_513,In_183);
and U1114 (N_1114,In_56,In_839);
nor U1115 (N_1115,In_71,In_279);
nand U1116 (N_1116,In_704,In_531);
nand U1117 (N_1117,In_154,In_628);
nand U1118 (N_1118,In_948,In_546);
xnor U1119 (N_1119,In_504,In_520);
or U1120 (N_1120,In_943,In_201);
or U1121 (N_1121,In_391,In_654);
and U1122 (N_1122,In_653,In_376);
xor U1123 (N_1123,In_355,In_570);
xor U1124 (N_1124,In_591,In_361);
nand U1125 (N_1125,In_766,In_981);
and U1126 (N_1126,In_657,In_564);
and U1127 (N_1127,In_990,In_232);
xnor U1128 (N_1128,In_573,In_874);
nor U1129 (N_1129,In_20,In_122);
nand U1130 (N_1130,In_425,In_16);
xnor U1131 (N_1131,In_986,In_227);
nor U1132 (N_1132,In_826,In_487);
xor U1133 (N_1133,In_999,In_731);
or U1134 (N_1134,In_592,In_367);
nand U1135 (N_1135,In_169,In_160);
xor U1136 (N_1136,In_360,In_232);
and U1137 (N_1137,In_77,In_28);
or U1138 (N_1138,In_345,In_189);
and U1139 (N_1139,In_641,In_893);
nor U1140 (N_1140,In_341,In_289);
nand U1141 (N_1141,In_537,In_614);
or U1142 (N_1142,In_489,In_139);
and U1143 (N_1143,In_720,In_64);
and U1144 (N_1144,In_912,In_108);
and U1145 (N_1145,In_730,In_471);
nand U1146 (N_1146,In_44,In_259);
xnor U1147 (N_1147,In_163,In_60);
or U1148 (N_1148,In_284,In_571);
and U1149 (N_1149,In_788,In_445);
nand U1150 (N_1150,In_223,In_354);
or U1151 (N_1151,In_7,In_129);
xnor U1152 (N_1152,In_218,In_343);
nand U1153 (N_1153,In_147,In_493);
nand U1154 (N_1154,In_315,In_139);
and U1155 (N_1155,In_291,In_88);
xor U1156 (N_1156,In_788,In_784);
or U1157 (N_1157,In_239,In_573);
nor U1158 (N_1158,In_618,In_477);
nand U1159 (N_1159,In_594,In_22);
and U1160 (N_1160,In_81,In_569);
and U1161 (N_1161,In_141,In_81);
and U1162 (N_1162,In_573,In_569);
or U1163 (N_1163,In_284,In_429);
nand U1164 (N_1164,In_677,In_626);
nor U1165 (N_1165,In_515,In_429);
xnor U1166 (N_1166,In_963,In_925);
xnor U1167 (N_1167,In_651,In_437);
and U1168 (N_1168,In_722,In_556);
or U1169 (N_1169,In_647,In_199);
nand U1170 (N_1170,In_327,In_86);
nor U1171 (N_1171,In_591,In_327);
nor U1172 (N_1172,In_710,In_640);
and U1173 (N_1173,In_998,In_925);
or U1174 (N_1174,In_730,In_439);
xor U1175 (N_1175,In_569,In_829);
and U1176 (N_1176,In_941,In_617);
or U1177 (N_1177,In_809,In_185);
nand U1178 (N_1178,In_872,In_667);
nor U1179 (N_1179,In_909,In_248);
or U1180 (N_1180,In_68,In_367);
and U1181 (N_1181,In_844,In_531);
nor U1182 (N_1182,In_161,In_363);
xor U1183 (N_1183,In_810,In_951);
and U1184 (N_1184,In_667,In_803);
xnor U1185 (N_1185,In_627,In_586);
nor U1186 (N_1186,In_290,In_236);
xnor U1187 (N_1187,In_317,In_120);
or U1188 (N_1188,In_416,In_497);
or U1189 (N_1189,In_637,In_90);
nor U1190 (N_1190,In_881,In_143);
nand U1191 (N_1191,In_221,In_814);
nand U1192 (N_1192,In_937,In_885);
nand U1193 (N_1193,In_146,In_206);
xor U1194 (N_1194,In_815,In_316);
or U1195 (N_1195,In_51,In_726);
xnor U1196 (N_1196,In_75,In_368);
or U1197 (N_1197,In_283,In_43);
and U1198 (N_1198,In_442,In_823);
and U1199 (N_1199,In_536,In_282);
or U1200 (N_1200,In_122,In_676);
and U1201 (N_1201,In_433,In_49);
or U1202 (N_1202,In_355,In_192);
nand U1203 (N_1203,In_515,In_883);
nand U1204 (N_1204,In_787,In_851);
and U1205 (N_1205,In_428,In_408);
nand U1206 (N_1206,In_104,In_545);
nand U1207 (N_1207,In_654,In_780);
nand U1208 (N_1208,In_95,In_850);
xnor U1209 (N_1209,In_794,In_775);
nand U1210 (N_1210,In_195,In_859);
nor U1211 (N_1211,In_233,In_607);
or U1212 (N_1212,In_681,In_953);
or U1213 (N_1213,In_850,In_128);
and U1214 (N_1214,In_308,In_620);
xnor U1215 (N_1215,In_39,In_651);
and U1216 (N_1216,In_960,In_662);
nor U1217 (N_1217,In_636,In_931);
nor U1218 (N_1218,In_841,In_188);
and U1219 (N_1219,In_796,In_61);
and U1220 (N_1220,In_415,In_627);
or U1221 (N_1221,In_650,In_800);
nand U1222 (N_1222,In_340,In_979);
or U1223 (N_1223,In_894,In_86);
or U1224 (N_1224,In_779,In_419);
nand U1225 (N_1225,In_273,In_409);
or U1226 (N_1226,In_135,In_483);
nand U1227 (N_1227,In_741,In_155);
nand U1228 (N_1228,In_860,In_485);
nor U1229 (N_1229,In_888,In_853);
nor U1230 (N_1230,In_221,In_963);
nand U1231 (N_1231,In_360,In_914);
or U1232 (N_1232,In_34,In_685);
xnor U1233 (N_1233,In_505,In_337);
nand U1234 (N_1234,In_635,In_741);
and U1235 (N_1235,In_141,In_709);
nand U1236 (N_1236,In_50,In_970);
xnor U1237 (N_1237,In_671,In_157);
and U1238 (N_1238,In_964,In_620);
nor U1239 (N_1239,In_326,In_102);
xnor U1240 (N_1240,In_850,In_557);
and U1241 (N_1241,In_522,In_630);
nor U1242 (N_1242,In_959,In_475);
nor U1243 (N_1243,In_980,In_964);
nand U1244 (N_1244,In_912,In_153);
xnor U1245 (N_1245,In_995,In_251);
nor U1246 (N_1246,In_667,In_274);
nor U1247 (N_1247,In_32,In_211);
nor U1248 (N_1248,In_285,In_10);
or U1249 (N_1249,In_35,In_831);
xor U1250 (N_1250,In_895,In_524);
or U1251 (N_1251,In_56,In_326);
xnor U1252 (N_1252,In_794,In_71);
and U1253 (N_1253,In_595,In_447);
xnor U1254 (N_1254,In_835,In_485);
nand U1255 (N_1255,In_278,In_852);
xnor U1256 (N_1256,In_445,In_54);
xor U1257 (N_1257,In_931,In_328);
xor U1258 (N_1258,In_385,In_169);
xnor U1259 (N_1259,In_639,In_610);
nand U1260 (N_1260,In_847,In_545);
and U1261 (N_1261,In_107,In_597);
nor U1262 (N_1262,In_592,In_619);
or U1263 (N_1263,In_132,In_330);
xnor U1264 (N_1264,In_718,In_635);
nor U1265 (N_1265,In_136,In_376);
nor U1266 (N_1266,In_322,In_209);
and U1267 (N_1267,In_580,In_755);
xor U1268 (N_1268,In_139,In_192);
and U1269 (N_1269,In_347,In_165);
nor U1270 (N_1270,In_252,In_173);
xor U1271 (N_1271,In_223,In_412);
or U1272 (N_1272,In_794,In_294);
and U1273 (N_1273,In_592,In_756);
and U1274 (N_1274,In_39,In_594);
nand U1275 (N_1275,In_279,In_385);
and U1276 (N_1276,In_601,In_786);
xor U1277 (N_1277,In_950,In_733);
xor U1278 (N_1278,In_832,In_154);
nor U1279 (N_1279,In_577,In_741);
xnor U1280 (N_1280,In_654,In_581);
and U1281 (N_1281,In_130,In_822);
nand U1282 (N_1282,In_735,In_552);
and U1283 (N_1283,In_357,In_933);
nand U1284 (N_1284,In_325,In_274);
xnor U1285 (N_1285,In_193,In_219);
or U1286 (N_1286,In_511,In_365);
and U1287 (N_1287,In_885,In_386);
xor U1288 (N_1288,In_185,In_53);
nand U1289 (N_1289,In_421,In_288);
nand U1290 (N_1290,In_408,In_962);
nor U1291 (N_1291,In_578,In_624);
nand U1292 (N_1292,In_552,In_202);
xnor U1293 (N_1293,In_901,In_75);
xnor U1294 (N_1294,In_209,In_805);
nor U1295 (N_1295,In_354,In_812);
and U1296 (N_1296,In_418,In_757);
xnor U1297 (N_1297,In_767,In_530);
xor U1298 (N_1298,In_827,In_382);
nand U1299 (N_1299,In_355,In_26);
xor U1300 (N_1300,In_337,In_378);
nor U1301 (N_1301,In_513,In_459);
xnor U1302 (N_1302,In_889,In_25);
nor U1303 (N_1303,In_916,In_178);
xor U1304 (N_1304,In_424,In_69);
or U1305 (N_1305,In_692,In_329);
nand U1306 (N_1306,In_120,In_704);
or U1307 (N_1307,In_283,In_785);
nand U1308 (N_1308,In_527,In_673);
and U1309 (N_1309,In_250,In_670);
and U1310 (N_1310,In_866,In_263);
or U1311 (N_1311,In_615,In_541);
and U1312 (N_1312,In_908,In_242);
xnor U1313 (N_1313,In_735,In_490);
nor U1314 (N_1314,In_984,In_442);
xor U1315 (N_1315,In_22,In_957);
and U1316 (N_1316,In_876,In_319);
or U1317 (N_1317,In_38,In_234);
and U1318 (N_1318,In_857,In_752);
and U1319 (N_1319,In_453,In_7);
nand U1320 (N_1320,In_792,In_148);
nand U1321 (N_1321,In_673,In_39);
xnor U1322 (N_1322,In_25,In_397);
nor U1323 (N_1323,In_979,In_50);
nand U1324 (N_1324,In_334,In_225);
nor U1325 (N_1325,In_701,In_866);
and U1326 (N_1326,In_817,In_911);
nand U1327 (N_1327,In_89,In_36);
and U1328 (N_1328,In_283,In_570);
and U1329 (N_1329,In_16,In_195);
nor U1330 (N_1330,In_67,In_546);
nor U1331 (N_1331,In_363,In_65);
or U1332 (N_1332,In_324,In_478);
and U1333 (N_1333,In_983,In_598);
nand U1334 (N_1334,In_633,In_530);
and U1335 (N_1335,In_922,In_258);
or U1336 (N_1336,In_969,In_53);
xor U1337 (N_1337,In_111,In_593);
or U1338 (N_1338,In_845,In_21);
nand U1339 (N_1339,In_94,In_497);
and U1340 (N_1340,In_113,In_642);
nand U1341 (N_1341,In_736,In_213);
or U1342 (N_1342,In_921,In_814);
and U1343 (N_1343,In_738,In_661);
and U1344 (N_1344,In_387,In_50);
or U1345 (N_1345,In_205,In_139);
nand U1346 (N_1346,In_401,In_217);
nand U1347 (N_1347,In_673,In_915);
or U1348 (N_1348,In_80,In_954);
xor U1349 (N_1349,In_326,In_841);
or U1350 (N_1350,In_29,In_139);
nand U1351 (N_1351,In_167,In_188);
nor U1352 (N_1352,In_696,In_249);
nor U1353 (N_1353,In_706,In_377);
and U1354 (N_1354,In_6,In_5);
xor U1355 (N_1355,In_323,In_954);
or U1356 (N_1356,In_68,In_180);
xnor U1357 (N_1357,In_770,In_692);
nand U1358 (N_1358,In_599,In_638);
nand U1359 (N_1359,In_335,In_301);
xor U1360 (N_1360,In_776,In_125);
and U1361 (N_1361,In_50,In_336);
xnor U1362 (N_1362,In_678,In_286);
nand U1363 (N_1363,In_453,In_375);
and U1364 (N_1364,In_120,In_931);
nand U1365 (N_1365,In_474,In_670);
or U1366 (N_1366,In_802,In_632);
or U1367 (N_1367,In_917,In_586);
nand U1368 (N_1368,In_891,In_554);
and U1369 (N_1369,In_239,In_662);
and U1370 (N_1370,In_831,In_910);
and U1371 (N_1371,In_360,In_514);
or U1372 (N_1372,In_511,In_691);
and U1373 (N_1373,In_427,In_563);
and U1374 (N_1374,In_867,In_714);
xor U1375 (N_1375,In_74,In_801);
xor U1376 (N_1376,In_571,In_733);
nand U1377 (N_1377,In_38,In_636);
xnor U1378 (N_1378,In_167,In_675);
or U1379 (N_1379,In_206,In_5);
or U1380 (N_1380,In_798,In_745);
nor U1381 (N_1381,In_274,In_253);
xor U1382 (N_1382,In_581,In_267);
xnor U1383 (N_1383,In_150,In_963);
xor U1384 (N_1384,In_179,In_245);
nand U1385 (N_1385,In_196,In_974);
nand U1386 (N_1386,In_130,In_392);
or U1387 (N_1387,In_8,In_303);
nor U1388 (N_1388,In_576,In_556);
nand U1389 (N_1389,In_511,In_245);
nand U1390 (N_1390,In_890,In_126);
nor U1391 (N_1391,In_856,In_875);
and U1392 (N_1392,In_678,In_863);
xnor U1393 (N_1393,In_224,In_210);
and U1394 (N_1394,In_634,In_415);
and U1395 (N_1395,In_670,In_572);
and U1396 (N_1396,In_412,In_444);
and U1397 (N_1397,In_190,In_914);
or U1398 (N_1398,In_525,In_819);
or U1399 (N_1399,In_536,In_220);
xor U1400 (N_1400,In_435,In_759);
xor U1401 (N_1401,In_729,In_279);
nor U1402 (N_1402,In_995,In_160);
nand U1403 (N_1403,In_530,In_794);
xor U1404 (N_1404,In_110,In_583);
or U1405 (N_1405,In_532,In_606);
and U1406 (N_1406,In_685,In_89);
xnor U1407 (N_1407,In_894,In_97);
and U1408 (N_1408,In_316,In_938);
or U1409 (N_1409,In_383,In_975);
nand U1410 (N_1410,In_310,In_829);
and U1411 (N_1411,In_254,In_767);
and U1412 (N_1412,In_681,In_438);
xor U1413 (N_1413,In_484,In_715);
xnor U1414 (N_1414,In_463,In_756);
or U1415 (N_1415,In_492,In_331);
and U1416 (N_1416,In_428,In_120);
and U1417 (N_1417,In_449,In_833);
or U1418 (N_1418,In_243,In_225);
nor U1419 (N_1419,In_320,In_517);
or U1420 (N_1420,In_220,In_885);
nor U1421 (N_1421,In_96,In_172);
nor U1422 (N_1422,In_35,In_697);
xnor U1423 (N_1423,In_299,In_865);
or U1424 (N_1424,In_870,In_785);
and U1425 (N_1425,In_66,In_541);
and U1426 (N_1426,In_476,In_335);
xor U1427 (N_1427,In_707,In_940);
nand U1428 (N_1428,In_962,In_460);
nor U1429 (N_1429,In_349,In_903);
or U1430 (N_1430,In_814,In_64);
nand U1431 (N_1431,In_993,In_266);
and U1432 (N_1432,In_362,In_816);
xor U1433 (N_1433,In_641,In_289);
or U1434 (N_1434,In_775,In_910);
xor U1435 (N_1435,In_57,In_22);
and U1436 (N_1436,In_358,In_158);
or U1437 (N_1437,In_396,In_569);
nand U1438 (N_1438,In_343,In_175);
xnor U1439 (N_1439,In_456,In_936);
nor U1440 (N_1440,In_959,In_842);
nand U1441 (N_1441,In_833,In_584);
xnor U1442 (N_1442,In_480,In_98);
nor U1443 (N_1443,In_696,In_468);
nand U1444 (N_1444,In_609,In_651);
or U1445 (N_1445,In_887,In_708);
nand U1446 (N_1446,In_835,In_711);
and U1447 (N_1447,In_888,In_443);
or U1448 (N_1448,In_623,In_277);
or U1449 (N_1449,In_949,In_572);
nand U1450 (N_1450,In_285,In_528);
and U1451 (N_1451,In_474,In_568);
nand U1452 (N_1452,In_749,In_406);
xor U1453 (N_1453,In_464,In_189);
nand U1454 (N_1454,In_266,In_794);
or U1455 (N_1455,In_344,In_732);
nor U1456 (N_1456,In_796,In_195);
xnor U1457 (N_1457,In_980,In_413);
and U1458 (N_1458,In_891,In_621);
and U1459 (N_1459,In_652,In_708);
xnor U1460 (N_1460,In_589,In_872);
and U1461 (N_1461,In_809,In_500);
nand U1462 (N_1462,In_327,In_272);
and U1463 (N_1463,In_861,In_579);
nand U1464 (N_1464,In_510,In_144);
and U1465 (N_1465,In_204,In_929);
and U1466 (N_1466,In_927,In_781);
nor U1467 (N_1467,In_119,In_120);
nand U1468 (N_1468,In_62,In_64);
xnor U1469 (N_1469,In_400,In_765);
nor U1470 (N_1470,In_209,In_217);
xor U1471 (N_1471,In_581,In_0);
nand U1472 (N_1472,In_265,In_677);
nand U1473 (N_1473,In_451,In_517);
and U1474 (N_1474,In_40,In_626);
nand U1475 (N_1475,In_254,In_864);
xnor U1476 (N_1476,In_916,In_716);
nand U1477 (N_1477,In_984,In_651);
and U1478 (N_1478,In_136,In_965);
and U1479 (N_1479,In_611,In_530);
nand U1480 (N_1480,In_542,In_573);
nand U1481 (N_1481,In_704,In_714);
xnor U1482 (N_1482,In_238,In_656);
nand U1483 (N_1483,In_518,In_595);
and U1484 (N_1484,In_140,In_906);
nor U1485 (N_1485,In_552,In_654);
or U1486 (N_1486,In_538,In_644);
and U1487 (N_1487,In_853,In_376);
or U1488 (N_1488,In_830,In_636);
nor U1489 (N_1489,In_49,In_620);
xnor U1490 (N_1490,In_970,In_632);
and U1491 (N_1491,In_711,In_500);
or U1492 (N_1492,In_367,In_368);
nor U1493 (N_1493,In_145,In_718);
nand U1494 (N_1494,In_592,In_130);
nand U1495 (N_1495,In_345,In_809);
and U1496 (N_1496,In_602,In_313);
nand U1497 (N_1497,In_327,In_137);
and U1498 (N_1498,In_993,In_980);
and U1499 (N_1499,In_584,In_734);
nand U1500 (N_1500,In_695,In_750);
nand U1501 (N_1501,In_303,In_512);
and U1502 (N_1502,In_251,In_972);
and U1503 (N_1503,In_134,In_140);
or U1504 (N_1504,In_70,In_88);
xor U1505 (N_1505,In_782,In_70);
and U1506 (N_1506,In_618,In_654);
or U1507 (N_1507,In_98,In_990);
nor U1508 (N_1508,In_780,In_620);
and U1509 (N_1509,In_242,In_661);
and U1510 (N_1510,In_206,In_298);
or U1511 (N_1511,In_912,In_763);
xnor U1512 (N_1512,In_677,In_122);
nor U1513 (N_1513,In_80,In_977);
xor U1514 (N_1514,In_679,In_540);
xor U1515 (N_1515,In_509,In_392);
nor U1516 (N_1516,In_233,In_207);
nor U1517 (N_1517,In_891,In_355);
nor U1518 (N_1518,In_402,In_524);
or U1519 (N_1519,In_736,In_29);
xnor U1520 (N_1520,In_440,In_105);
nand U1521 (N_1521,In_753,In_371);
xor U1522 (N_1522,In_46,In_217);
nand U1523 (N_1523,In_567,In_685);
and U1524 (N_1524,In_850,In_966);
nand U1525 (N_1525,In_872,In_579);
or U1526 (N_1526,In_679,In_300);
xnor U1527 (N_1527,In_307,In_184);
or U1528 (N_1528,In_600,In_82);
and U1529 (N_1529,In_489,In_324);
nand U1530 (N_1530,In_11,In_231);
nand U1531 (N_1531,In_745,In_86);
xnor U1532 (N_1532,In_830,In_635);
and U1533 (N_1533,In_912,In_257);
or U1534 (N_1534,In_464,In_84);
or U1535 (N_1535,In_55,In_403);
and U1536 (N_1536,In_111,In_324);
or U1537 (N_1537,In_399,In_284);
nor U1538 (N_1538,In_752,In_236);
or U1539 (N_1539,In_531,In_635);
or U1540 (N_1540,In_100,In_672);
nor U1541 (N_1541,In_334,In_15);
and U1542 (N_1542,In_537,In_314);
nor U1543 (N_1543,In_635,In_244);
and U1544 (N_1544,In_356,In_458);
or U1545 (N_1545,In_324,In_600);
nand U1546 (N_1546,In_434,In_267);
and U1547 (N_1547,In_940,In_31);
nor U1548 (N_1548,In_420,In_601);
or U1549 (N_1549,In_747,In_321);
or U1550 (N_1550,In_958,In_297);
nor U1551 (N_1551,In_292,In_198);
or U1552 (N_1552,In_146,In_910);
nor U1553 (N_1553,In_632,In_150);
or U1554 (N_1554,In_553,In_972);
or U1555 (N_1555,In_248,In_782);
and U1556 (N_1556,In_927,In_276);
xor U1557 (N_1557,In_286,In_277);
nor U1558 (N_1558,In_871,In_136);
and U1559 (N_1559,In_774,In_960);
nor U1560 (N_1560,In_370,In_175);
xor U1561 (N_1561,In_506,In_496);
and U1562 (N_1562,In_321,In_204);
and U1563 (N_1563,In_383,In_210);
and U1564 (N_1564,In_165,In_110);
nor U1565 (N_1565,In_519,In_778);
or U1566 (N_1566,In_453,In_94);
and U1567 (N_1567,In_464,In_533);
or U1568 (N_1568,In_567,In_991);
nor U1569 (N_1569,In_549,In_516);
or U1570 (N_1570,In_685,In_951);
and U1571 (N_1571,In_172,In_411);
and U1572 (N_1572,In_772,In_596);
and U1573 (N_1573,In_153,In_128);
or U1574 (N_1574,In_615,In_256);
xor U1575 (N_1575,In_216,In_61);
or U1576 (N_1576,In_873,In_82);
nor U1577 (N_1577,In_550,In_580);
nor U1578 (N_1578,In_432,In_725);
nor U1579 (N_1579,In_954,In_505);
nand U1580 (N_1580,In_519,In_331);
nor U1581 (N_1581,In_333,In_924);
or U1582 (N_1582,In_969,In_508);
xnor U1583 (N_1583,In_675,In_129);
nor U1584 (N_1584,In_434,In_804);
and U1585 (N_1585,In_705,In_306);
nor U1586 (N_1586,In_697,In_10);
xor U1587 (N_1587,In_68,In_288);
or U1588 (N_1588,In_116,In_228);
xnor U1589 (N_1589,In_635,In_585);
xnor U1590 (N_1590,In_636,In_743);
and U1591 (N_1591,In_259,In_831);
xor U1592 (N_1592,In_202,In_776);
nand U1593 (N_1593,In_369,In_265);
nand U1594 (N_1594,In_217,In_151);
nand U1595 (N_1595,In_376,In_516);
or U1596 (N_1596,In_334,In_808);
nor U1597 (N_1597,In_438,In_89);
and U1598 (N_1598,In_609,In_901);
or U1599 (N_1599,In_220,In_97);
xor U1600 (N_1600,In_623,In_293);
nand U1601 (N_1601,In_593,In_353);
nand U1602 (N_1602,In_167,In_621);
nor U1603 (N_1603,In_569,In_962);
nor U1604 (N_1604,In_429,In_166);
nor U1605 (N_1605,In_16,In_722);
xor U1606 (N_1606,In_959,In_241);
and U1607 (N_1607,In_139,In_379);
nand U1608 (N_1608,In_862,In_672);
nor U1609 (N_1609,In_464,In_628);
or U1610 (N_1610,In_464,In_939);
and U1611 (N_1611,In_445,In_348);
or U1612 (N_1612,In_252,In_556);
xnor U1613 (N_1613,In_161,In_198);
nor U1614 (N_1614,In_430,In_652);
nor U1615 (N_1615,In_130,In_783);
xor U1616 (N_1616,In_631,In_613);
or U1617 (N_1617,In_313,In_99);
and U1618 (N_1618,In_794,In_469);
nor U1619 (N_1619,In_465,In_446);
and U1620 (N_1620,In_398,In_932);
nor U1621 (N_1621,In_591,In_406);
and U1622 (N_1622,In_944,In_324);
xor U1623 (N_1623,In_890,In_603);
nand U1624 (N_1624,In_300,In_844);
nand U1625 (N_1625,In_273,In_278);
nor U1626 (N_1626,In_304,In_399);
nand U1627 (N_1627,In_822,In_567);
or U1628 (N_1628,In_20,In_31);
and U1629 (N_1629,In_955,In_127);
nand U1630 (N_1630,In_144,In_570);
xor U1631 (N_1631,In_675,In_732);
or U1632 (N_1632,In_299,In_316);
nor U1633 (N_1633,In_288,In_214);
nor U1634 (N_1634,In_889,In_506);
or U1635 (N_1635,In_913,In_956);
xor U1636 (N_1636,In_469,In_649);
xor U1637 (N_1637,In_273,In_299);
xor U1638 (N_1638,In_456,In_208);
and U1639 (N_1639,In_456,In_234);
or U1640 (N_1640,In_23,In_924);
nand U1641 (N_1641,In_41,In_125);
nor U1642 (N_1642,In_986,In_374);
nand U1643 (N_1643,In_102,In_96);
nor U1644 (N_1644,In_975,In_972);
nand U1645 (N_1645,In_852,In_200);
xor U1646 (N_1646,In_552,In_724);
nand U1647 (N_1647,In_266,In_485);
nor U1648 (N_1648,In_95,In_176);
nor U1649 (N_1649,In_582,In_28);
nand U1650 (N_1650,In_724,In_986);
xor U1651 (N_1651,In_985,In_949);
xnor U1652 (N_1652,In_333,In_943);
xnor U1653 (N_1653,In_755,In_712);
xor U1654 (N_1654,In_779,In_851);
nor U1655 (N_1655,In_750,In_273);
and U1656 (N_1656,In_939,In_541);
xor U1657 (N_1657,In_722,In_785);
and U1658 (N_1658,In_847,In_649);
nor U1659 (N_1659,In_981,In_760);
nor U1660 (N_1660,In_906,In_55);
xor U1661 (N_1661,In_795,In_857);
xnor U1662 (N_1662,In_736,In_824);
nor U1663 (N_1663,In_283,In_814);
or U1664 (N_1664,In_174,In_674);
xnor U1665 (N_1665,In_6,In_580);
or U1666 (N_1666,In_697,In_844);
nor U1667 (N_1667,In_631,In_885);
and U1668 (N_1668,In_21,In_646);
nand U1669 (N_1669,In_753,In_233);
xor U1670 (N_1670,In_246,In_612);
xor U1671 (N_1671,In_943,In_927);
xnor U1672 (N_1672,In_7,In_245);
nand U1673 (N_1673,In_926,In_374);
and U1674 (N_1674,In_238,In_999);
nand U1675 (N_1675,In_399,In_445);
xor U1676 (N_1676,In_385,In_463);
xor U1677 (N_1677,In_975,In_564);
nand U1678 (N_1678,In_410,In_472);
nor U1679 (N_1679,In_180,In_250);
xor U1680 (N_1680,In_247,In_134);
nand U1681 (N_1681,In_360,In_223);
and U1682 (N_1682,In_171,In_365);
xor U1683 (N_1683,In_619,In_605);
and U1684 (N_1684,In_680,In_24);
xnor U1685 (N_1685,In_543,In_329);
xor U1686 (N_1686,In_965,In_620);
nand U1687 (N_1687,In_807,In_945);
nor U1688 (N_1688,In_144,In_531);
xor U1689 (N_1689,In_338,In_395);
nand U1690 (N_1690,In_170,In_660);
xnor U1691 (N_1691,In_551,In_760);
nor U1692 (N_1692,In_245,In_229);
xnor U1693 (N_1693,In_654,In_272);
xnor U1694 (N_1694,In_416,In_904);
and U1695 (N_1695,In_184,In_295);
or U1696 (N_1696,In_2,In_157);
nor U1697 (N_1697,In_916,In_821);
and U1698 (N_1698,In_382,In_937);
nand U1699 (N_1699,In_45,In_172);
nand U1700 (N_1700,In_590,In_327);
or U1701 (N_1701,In_806,In_140);
nand U1702 (N_1702,In_880,In_836);
xor U1703 (N_1703,In_347,In_670);
and U1704 (N_1704,In_921,In_897);
xor U1705 (N_1705,In_942,In_115);
and U1706 (N_1706,In_88,In_513);
or U1707 (N_1707,In_170,In_579);
nor U1708 (N_1708,In_120,In_153);
nor U1709 (N_1709,In_999,In_220);
nor U1710 (N_1710,In_776,In_735);
and U1711 (N_1711,In_900,In_36);
nor U1712 (N_1712,In_295,In_501);
nor U1713 (N_1713,In_194,In_752);
and U1714 (N_1714,In_69,In_332);
and U1715 (N_1715,In_320,In_153);
nand U1716 (N_1716,In_188,In_261);
nor U1717 (N_1717,In_132,In_823);
nor U1718 (N_1718,In_85,In_392);
and U1719 (N_1719,In_770,In_958);
and U1720 (N_1720,In_321,In_384);
nor U1721 (N_1721,In_453,In_144);
nor U1722 (N_1722,In_969,In_581);
or U1723 (N_1723,In_291,In_455);
nor U1724 (N_1724,In_152,In_421);
xnor U1725 (N_1725,In_699,In_683);
xnor U1726 (N_1726,In_666,In_685);
or U1727 (N_1727,In_803,In_445);
nor U1728 (N_1728,In_858,In_39);
nor U1729 (N_1729,In_918,In_695);
or U1730 (N_1730,In_240,In_744);
xnor U1731 (N_1731,In_726,In_54);
and U1732 (N_1732,In_207,In_395);
xnor U1733 (N_1733,In_635,In_703);
nand U1734 (N_1734,In_368,In_774);
and U1735 (N_1735,In_248,In_948);
xor U1736 (N_1736,In_756,In_73);
or U1737 (N_1737,In_117,In_585);
xnor U1738 (N_1738,In_613,In_304);
nand U1739 (N_1739,In_825,In_822);
nand U1740 (N_1740,In_112,In_201);
or U1741 (N_1741,In_891,In_565);
xnor U1742 (N_1742,In_951,In_284);
or U1743 (N_1743,In_565,In_558);
xnor U1744 (N_1744,In_775,In_440);
xnor U1745 (N_1745,In_290,In_665);
or U1746 (N_1746,In_425,In_594);
or U1747 (N_1747,In_731,In_203);
and U1748 (N_1748,In_861,In_722);
or U1749 (N_1749,In_833,In_527);
nand U1750 (N_1750,In_633,In_917);
xor U1751 (N_1751,In_265,In_964);
xor U1752 (N_1752,In_561,In_911);
xor U1753 (N_1753,In_395,In_927);
and U1754 (N_1754,In_380,In_421);
or U1755 (N_1755,In_533,In_346);
and U1756 (N_1756,In_97,In_325);
nor U1757 (N_1757,In_487,In_33);
or U1758 (N_1758,In_299,In_701);
nand U1759 (N_1759,In_327,In_283);
nand U1760 (N_1760,In_771,In_619);
nand U1761 (N_1761,In_394,In_776);
nor U1762 (N_1762,In_968,In_187);
xnor U1763 (N_1763,In_82,In_354);
or U1764 (N_1764,In_923,In_18);
or U1765 (N_1765,In_756,In_794);
xor U1766 (N_1766,In_813,In_992);
or U1767 (N_1767,In_861,In_831);
or U1768 (N_1768,In_24,In_299);
and U1769 (N_1769,In_125,In_806);
nand U1770 (N_1770,In_551,In_907);
nand U1771 (N_1771,In_657,In_628);
and U1772 (N_1772,In_69,In_448);
xnor U1773 (N_1773,In_823,In_857);
nor U1774 (N_1774,In_687,In_323);
nand U1775 (N_1775,In_396,In_594);
nor U1776 (N_1776,In_841,In_280);
nand U1777 (N_1777,In_356,In_338);
and U1778 (N_1778,In_131,In_879);
nor U1779 (N_1779,In_799,In_491);
or U1780 (N_1780,In_500,In_95);
nor U1781 (N_1781,In_904,In_24);
and U1782 (N_1782,In_989,In_481);
nor U1783 (N_1783,In_960,In_859);
or U1784 (N_1784,In_983,In_369);
nand U1785 (N_1785,In_382,In_392);
and U1786 (N_1786,In_637,In_392);
or U1787 (N_1787,In_952,In_820);
or U1788 (N_1788,In_203,In_124);
and U1789 (N_1789,In_420,In_585);
xor U1790 (N_1790,In_241,In_462);
xor U1791 (N_1791,In_387,In_335);
or U1792 (N_1792,In_834,In_910);
or U1793 (N_1793,In_825,In_431);
or U1794 (N_1794,In_332,In_167);
nor U1795 (N_1795,In_369,In_245);
nand U1796 (N_1796,In_231,In_746);
nor U1797 (N_1797,In_554,In_222);
or U1798 (N_1798,In_661,In_469);
nor U1799 (N_1799,In_936,In_657);
and U1800 (N_1800,In_625,In_840);
nor U1801 (N_1801,In_916,In_74);
or U1802 (N_1802,In_848,In_219);
nand U1803 (N_1803,In_944,In_829);
nor U1804 (N_1804,In_923,In_577);
or U1805 (N_1805,In_731,In_130);
nand U1806 (N_1806,In_112,In_939);
and U1807 (N_1807,In_539,In_823);
or U1808 (N_1808,In_804,In_656);
nand U1809 (N_1809,In_859,In_459);
or U1810 (N_1810,In_651,In_637);
and U1811 (N_1811,In_597,In_220);
nor U1812 (N_1812,In_527,In_925);
xor U1813 (N_1813,In_204,In_908);
nand U1814 (N_1814,In_466,In_762);
and U1815 (N_1815,In_799,In_548);
nand U1816 (N_1816,In_77,In_856);
nand U1817 (N_1817,In_105,In_586);
nor U1818 (N_1818,In_551,In_187);
nor U1819 (N_1819,In_602,In_909);
nor U1820 (N_1820,In_833,In_548);
or U1821 (N_1821,In_201,In_696);
nor U1822 (N_1822,In_707,In_593);
nor U1823 (N_1823,In_238,In_688);
and U1824 (N_1824,In_228,In_977);
nor U1825 (N_1825,In_417,In_102);
and U1826 (N_1826,In_386,In_936);
or U1827 (N_1827,In_760,In_505);
nor U1828 (N_1828,In_83,In_974);
and U1829 (N_1829,In_716,In_224);
or U1830 (N_1830,In_74,In_170);
or U1831 (N_1831,In_195,In_635);
nand U1832 (N_1832,In_293,In_692);
nand U1833 (N_1833,In_316,In_587);
nor U1834 (N_1834,In_695,In_698);
xor U1835 (N_1835,In_835,In_802);
nor U1836 (N_1836,In_663,In_952);
nor U1837 (N_1837,In_568,In_18);
xnor U1838 (N_1838,In_289,In_951);
nand U1839 (N_1839,In_203,In_730);
nor U1840 (N_1840,In_881,In_269);
nand U1841 (N_1841,In_516,In_716);
nor U1842 (N_1842,In_363,In_366);
and U1843 (N_1843,In_137,In_850);
nand U1844 (N_1844,In_921,In_262);
nand U1845 (N_1845,In_787,In_667);
and U1846 (N_1846,In_640,In_518);
nand U1847 (N_1847,In_525,In_907);
nor U1848 (N_1848,In_644,In_287);
nor U1849 (N_1849,In_259,In_329);
and U1850 (N_1850,In_962,In_103);
or U1851 (N_1851,In_401,In_325);
nand U1852 (N_1852,In_710,In_485);
or U1853 (N_1853,In_998,In_140);
and U1854 (N_1854,In_571,In_370);
xnor U1855 (N_1855,In_744,In_981);
or U1856 (N_1856,In_755,In_337);
xor U1857 (N_1857,In_685,In_277);
or U1858 (N_1858,In_446,In_573);
and U1859 (N_1859,In_832,In_873);
and U1860 (N_1860,In_652,In_227);
or U1861 (N_1861,In_26,In_847);
xnor U1862 (N_1862,In_53,In_374);
nor U1863 (N_1863,In_157,In_993);
or U1864 (N_1864,In_172,In_356);
xor U1865 (N_1865,In_657,In_949);
or U1866 (N_1866,In_213,In_565);
xor U1867 (N_1867,In_452,In_778);
and U1868 (N_1868,In_748,In_552);
nor U1869 (N_1869,In_192,In_71);
or U1870 (N_1870,In_867,In_370);
and U1871 (N_1871,In_51,In_64);
and U1872 (N_1872,In_542,In_409);
xor U1873 (N_1873,In_63,In_129);
nor U1874 (N_1874,In_116,In_331);
xor U1875 (N_1875,In_721,In_469);
xnor U1876 (N_1876,In_756,In_190);
nor U1877 (N_1877,In_208,In_25);
nand U1878 (N_1878,In_564,In_297);
nor U1879 (N_1879,In_907,In_856);
nor U1880 (N_1880,In_941,In_173);
xnor U1881 (N_1881,In_125,In_816);
and U1882 (N_1882,In_305,In_754);
or U1883 (N_1883,In_699,In_478);
nand U1884 (N_1884,In_201,In_534);
nand U1885 (N_1885,In_61,In_463);
and U1886 (N_1886,In_699,In_646);
nand U1887 (N_1887,In_586,In_475);
and U1888 (N_1888,In_181,In_992);
nor U1889 (N_1889,In_594,In_667);
nand U1890 (N_1890,In_398,In_916);
nor U1891 (N_1891,In_166,In_952);
nand U1892 (N_1892,In_612,In_372);
or U1893 (N_1893,In_810,In_564);
and U1894 (N_1894,In_917,In_337);
and U1895 (N_1895,In_712,In_626);
and U1896 (N_1896,In_382,In_648);
or U1897 (N_1897,In_700,In_945);
nor U1898 (N_1898,In_481,In_760);
nand U1899 (N_1899,In_392,In_80);
and U1900 (N_1900,In_723,In_22);
xnor U1901 (N_1901,In_625,In_988);
nand U1902 (N_1902,In_487,In_986);
and U1903 (N_1903,In_261,In_469);
nand U1904 (N_1904,In_315,In_990);
and U1905 (N_1905,In_458,In_786);
xnor U1906 (N_1906,In_805,In_504);
or U1907 (N_1907,In_131,In_259);
and U1908 (N_1908,In_904,In_108);
xnor U1909 (N_1909,In_395,In_320);
and U1910 (N_1910,In_69,In_896);
nor U1911 (N_1911,In_824,In_616);
xor U1912 (N_1912,In_143,In_576);
or U1913 (N_1913,In_218,In_707);
nor U1914 (N_1914,In_224,In_614);
or U1915 (N_1915,In_445,In_139);
and U1916 (N_1916,In_583,In_863);
and U1917 (N_1917,In_695,In_942);
and U1918 (N_1918,In_965,In_437);
and U1919 (N_1919,In_308,In_1);
nand U1920 (N_1920,In_848,In_150);
or U1921 (N_1921,In_435,In_262);
xnor U1922 (N_1922,In_472,In_565);
or U1923 (N_1923,In_599,In_280);
nand U1924 (N_1924,In_92,In_619);
nor U1925 (N_1925,In_544,In_293);
and U1926 (N_1926,In_922,In_367);
or U1927 (N_1927,In_273,In_248);
or U1928 (N_1928,In_980,In_723);
or U1929 (N_1929,In_215,In_252);
nor U1930 (N_1930,In_56,In_926);
nor U1931 (N_1931,In_776,In_129);
and U1932 (N_1932,In_271,In_849);
and U1933 (N_1933,In_571,In_735);
xor U1934 (N_1934,In_6,In_259);
and U1935 (N_1935,In_139,In_108);
xor U1936 (N_1936,In_16,In_616);
nand U1937 (N_1937,In_537,In_783);
xor U1938 (N_1938,In_321,In_813);
or U1939 (N_1939,In_379,In_333);
xor U1940 (N_1940,In_585,In_598);
nand U1941 (N_1941,In_119,In_176);
nand U1942 (N_1942,In_205,In_194);
or U1943 (N_1943,In_91,In_720);
and U1944 (N_1944,In_201,In_915);
xnor U1945 (N_1945,In_941,In_1);
xor U1946 (N_1946,In_290,In_495);
nand U1947 (N_1947,In_749,In_698);
nor U1948 (N_1948,In_281,In_78);
nand U1949 (N_1949,In_244,In_368);
xor U1950 (N_1950,In_2,In_244);
nor U1951 (N_1951,In_451,In_866);
xnor U1952 (N_1952,In_521,In_252);
nand U1953 (N_1953,In_840,In_45);
xor U1954 (N_1954,In_81,In_788);
nor U1955 (N_1955,In_289,In_944);
nand U1956 (N_1956,In_660,In_903);
xor U1957 (N_1957,In_360,In_496);
xnor U1958 (N_1958,In_907,In_660);
or U1959 (N_1959,In_9,In_597);
or U1960 (N_1960,In_320,In_496);
nand U1961 (N_1961,In_224,In_803);
xor U1962 (N_1962,In_161,In_525);
and U1963 (N_1963,In_992,In_43);
nand U1964 (N_1964,In_562,In_386);
nor U1965 (N_1965,In_611,In_730);
and U1966 (N_1966,In_444,In_793);
nand U1967 (N_1967,In_606,In_355);
or U1968 (N_1968,In_40,In_356);
nor U1969 (N_1969,In_766,In_323);
nor U1970 (N_1970,In_643,In_977);
and U1971 (N_1971,In_612,In_61);
xnor U1972 (N_1972,In_790,In_92);
nor U1973 (N_1973,In_514,In_141);
nor U1974 (N_1974,In_673,In_962);
nor U1975 (N_1975,In_945,In_568);
nor U1976 (N_1976,In_329,In_181);
and U1977 (N_1977,In_154,In_460);
nand U1978 (N_1978,In_748,In_785);
nand U1979 (N_1979,In_452,In_444);
and U1980 (N_1980,In_675,In_935);
or U1981 (N_1981,In_735,In_329);
xor U1982 (N_1982,In_90,In_6);
nand U1983 (N_1983,In_631,In_170);
xnor U1984 (N_1984,In_375,In_606);
nor U1985 (N_1985,In_848,In_660);
nand U1986 (N_1986,In_628,In_28);
or U1987 (N_1987,In_908,In_976);
and U1988 (N_1988,In_638,In_289);
or U1989 (N_1989,In_577,In_262);
and U1990 (N_1990,In_347,In_568);
or U1991 (N_1991,In_686,In_748);
nand U1992 (N_1992,In_548,In_732);
or U1993 (N_1993,In_66,In_270);
xnor U1994 (N_1994,In_759,In_490);
or U1995 (N_1995,In_374,In_280);
nor U1996 (N_1996,In_847,In_984);
and U1997 (N_1997,In_119,In_237);
or U1998 (N_1998,In_780,In_942);
xnor U1999 (N_1999,In_389,In_881);
or U2000 (N_2000,N_1540,N_486);
xnor U2001 (N_2001,N_1405,N_1102);
nor U2002 (N_2002,N_1712,N_1134);
nand U2003 (N_2003,N_223,N_130);
nand U2004 (N_2004,N_259,N_893);
and U2005 (N_2005,N_15,N_504);
nor U2006 (N_2006,N_334,N_1968);
nor U2007 (N_2007,N_1193,N_1688);
and U2008 (N_2008,N_1326,N_1575);
xor U2009 (N_2009,N_1289,N_704);
xnor U2010 (N_2010,N_733,N_613);
and U2011 (N_2011,N_1436,N_337);
or U2012 (N_2012,N_972,N_1789);
xnor U2013 (N_2013,N_1745,N_99);
xnor U2014 (N_2014,N_668,N_1814);
nor U2015 (N_2015,N_1450,N_12);
and U2016 (N_2016,N_1933,N_1681);
and U2017 (N_2017,N_1463,N_1374);
nor U2018 (N_2018,N_1828,N_29);
nand U2019 (N_2019,N_1981,N_392);
nand U2020 (N_2020,N_952,N_1578);
and U2021 (N_2021,N_522,N_597);
and U2022 (N_2022,N_479,N_147);
xor U2023 (N_2023,N_589,N_1003);
nand U2024 (N_2024,N_1258,N_938);
or U2025 (N_2025,N_1737,N_1880);
nor U2026 (N_2026,N_1181,N_163);
xnor U2027 (N_2027,N_903,N_1999);
and U2028 (N_2028,N_1888,N_34);
or U2029 (N_2029,N_1534,N_168);
xnor U2030 (N_2030,N_491,N_145);
and U2031 (N_2031,N_1332,N_1277);
and U2032 (N_2032,N_1039,N_1899);
nand U2033 (N_2033,N_1139,N_1455);
and U2034 (N_2034,N_739,N_712);
or U2035 (N_2035,N_1963,N_821);
or U2036 (N_2036,N_902,N_539);
nand U2037 (N_2037,N_289,N_1925);
xor U2038 (N_2038,N_1602,N_265);
xnor U2039 (N_2039,N_1654,N_1546);
nand U2040 (N_2040,N_1187,N_167);
or U2041 (N_2041,N_761,N_1089);
nor U2042 (N_2042,N_117,N_1379);
nor U2043 (N_2043,N_576,N_21);
nand U2044 (N_2044,N_806,N_1090);
nand U2045 (N_2045,N_1592,N_181);
and U2046 (N_2046,N_978,N_50);
and U2047 (N_2047,N_1641,N_325);
nor U2048 (N_2048,N_499,N_1419);
xor U2049 (N_2049,N_1320,N_976);
and U2050 (N_2050,N_907,N_1972);
nand U2051 (N_2051,N_305,N_1846);
xor U2052 (N_2052,N_1731,N_667);
or U2053 (N_2053,N_135,N_572);
nor U2054 (N_2054,N_1409,N_274);
or U2055 (N_2055,N_1708,N_1831);
nand U2056 (N_2056,N_1816,N_180);
xor U2057 (N_2057,N_1410,N_69);
and U2058 (N_2058,N_1829,N_1603);
xor U2059 (N_2059,N_1148,N_418);
xor U2060 (N_2060,N_1229,N_197);
or U2061 (N_2061,N_1759,N_1541);
or U2062 (N_2062,N_1156,N_549);
or U2063 (N_2063,N_644,N_681);
nor U2064 (N_2064,N_1357,N_1551);
and U2065 (N_2065,N_184,N_1497);
or U2066 (N_2066,N_204,N_533);
nor U2067 (N_2067,N_57,N_1883);
or U2068 (N_2068,N_927,N_1794);
and U2069 (N_2069,N_1553,N_1358);
nor U2070 (N_2070,N_1686,N_965);
nand U2071 (N_2071,N_309,N_1834);
nand U2072 (N_2072,N_900,N_788);
xor U2073 (N_2073,N_997,N_885);
and U2074 (N_2074,N_1446,N_1190);
nor U2075 (N_2075,N_1041,N_1426);
and U2076 (N_2076,N_472,N_27);
or U2077 (N_2077,N_0,N_396);
nand U2078 (N_2078,N_1360,N_627);
or U2079 (N_2079,N_1991,N_971);
or U2080 (N_2080,N_1161,N_105);
nand U2081 (N_2081,N_1848,N_1083);
nor U2082 (N_2082,N_556,N_370);
nand U2083 (N_2083,N_1271,N_1478);
and U2084 (N_2084,N_1319,N_308);
xnor U2085 (N_2085,N_581,N_1496);
or U2086 (N_2086,N_1854,N_579);
or U2087 (N_2087,N_1109,N_782);
nand U2088 (N_2088,N_45,N_544);
nor U2089 (N_2089,N_1792,N_870);
and U2090 (N_2090,N_1055,N_721);
nor U2091 (N_2091,N_769,N_1830);
xor U2092 (N_2092,N_201,N_666);
and U2093 (N_2093,N_1653,N_1480);
nor U2094 (N_2094,N_489,N_1199);
nand U2095 (N_2095,N_993,N_208);
and U2096 (N_2096,N_1559,N_567);
xnor U2097 (N_2097,N_1233,N_1870);
nand U2098 (N_2098,N_101,N_537);
nor U2099 (N_2099,N_632,N_359);
nor U2100 (N_2100,N_235,N_1778);
or U2101 (N_2101,N_1609,N_438);
and U2102 (N_2102,N_1869,N_925);
xor U2103 (N_2103,N_1965,N_1622);
xor U2104 (N_2104,N_1385,N_1254);
or U2105 (N_2105,N_58,N_257);
nor U2106 (N_2106,N_1097,N_1656);
or U2107 (N_2107,N_1605,N_1537);
nand U2108 (N_2108,N_879,N_715);
nor U2109 (N_2109,N_1475,N_1075);
and U2110 (N_2110,N_451,N_784);
nand U2111 (N_2111,N_1489,N_1866);
and U2112 (N_2112,N_1432,N_1433);
and U2113 (N_2113,N_642,N_1570);
or U2114 (N_2114,N_1844,N_1642);
nor U2115 (N_2115,N_153,N_894);
xnor U2116 (N_2116,N_1918,N_1563);
nand U2117 (N_2117,N_1110,N_1961);
xnor U2118 (N_2118,N_1797,N_1321);
or U2119 (N_2119,N_1547,N_409);
and U2120 (N_2120,N_1997,N_66);
nand U2121 (N_2121,N_1781,N_839);
or U2122 (N_2122,N_1153,N_1472);
and U2123 (N_2123,N_293,N_104);
xnor U2124 (N_2124,N_897,N_427);
and U2125 (N_2125,N_1847,N_550);
or U2126 (N_2126,N_497,N_960);
xnor U2127 (N_2127,N_146,N_633);
and U2128 (N_2128,N_2,N_1112);
nand U2129 (N_2129,N_570,N_215);
nand U2130 (N_2130,N_110,N_836);
nand U2131 (N_2131,N_79,N_395);
nand U2132 (N_2132,N_1214,N_1131);
or U2133 (N_2133,N_561,N_1516);
and U2134 (N_2134,N_1926,N_1152);
nand U2135 (N_2135,N_939,N_776);
xnor U2136 (N_2136,N_1328,N_1821);
nor U2137 (N_2137,N_516,N_920);
nor U2138 (N_2138,N_336,N_906);
xor U2139 (N_2139,N_781,N_1425);
xor U2140 (N_2140,N_413,N_690);
and U2141 (N_2141,N_1774,N_618);
nand U2142 (N_2142,N_1142,N_899);
or U2143 (N_2143,N_880,N_1221);
nor U2144 (N_2144,N_303,N_56);
xor U2145 (N_2145,N_1660,N_1389);
nand U2146 (N_2146,N_689,N_1191);
nor U2147 (N_2147,N_990,N_1140);
or U2148 (N_2148,N_1849,N_331);
and U2149 (N_2149,N_410,N_1135);
and U2150 (N_2150,N_1552,N_916);
nand U2151 (N_2151,N_1544,N_1339);
or U2152 (N_2152,N_908,N_703);
and U2153 (N_2153,N_801,N_492);
nor U2154 (N_2154,N_943,N_1411);
nor U2155 (N_2155,N_192,N_1186);
nand U2156 (N_2156,N_86,N_311);
or U2157 (N_2157,N_575,N_1293);
nor U2158 (N_2158,N_1598,N_89);
and U2159 (N_2159,N_1730,N_92);
xor U2160 (N_2160,N_1351,N_129);
or U2161 (N_2161,N_115,N_1263);
or U2162 (N_2162,N_940,N_394);
and U2163 (N_2163,N_1456,N_865);
and U2164 (N_2164,N_1823,N_1872);
nor U2165 (N_2165,N_1951,N_1716);
or U2166 (N_2166,N_455,N_573);
and U2167 (N_2167,N_1005,N_536);
xor U2168 (N_2168,N_217,N_1531);
or U2169 (N_2169,N_808,N_218);
nand U2170 (N_2170,N_95,N_76);
or U2171 (N_2171,N_1967,N_1414);
nand U2172 (N_2172,N_1735,N_481);
nor U2173 (N_2173,N_709,N_1066);
xnor U2174 (N_2174,N_1356,N_1045);
and U2175 (N_2175,N_1934,N_1723);
nor U2176 (N_2176,N_1255,N_652);
nand U2177 (N_2177,N_1770,N_1477);
nand U2178 (N_2178,N_1071,N_1533);
or U2179 (N_2179,N_1396,N_365);
or U2180 (N_2180,N_292,N_407);
and U2181 (N_2181,N_1920,N_827);
nor U2182 (N_2182,N_1348,N_634);
or U2183 (N_2183,N_719,N_324);
xnor U2184 (N_2184,N_1224,N_912);
nand U2185 (N_2185,N_1371,N_416);
nand U2186 (N_2186,N_493,N_598);
xor U2187 (N_2187,N_229,N_1912);
nor U2188 (N_2188,N_1068,N_249);
and U2189 (N_2189,N_1160,N_1207);
nor U2190 (N_2190,N_1772,N_1035);
or U2191 (N_2191,N_725,N_1744);
nor U2192 (N_2192,N_1395,N_1067);
or U2193 (N_2193,N_1373,N_250);
xor U2194 (N_2194,N_811,N_838);
nor U2195 (N_2195,N_1978,N_710);
xnor U2196 (N_2196,N_1070,N_1752);
nand U2197 (N_2197,N_1885,N_1994);
xnor U2198 (N_2198,N_1099,N_926);
nor U2199 (N_2199,N_1215,N_429);
xor U2200 (N_2200,N_1889,N_1932);
nand U2201 (N_2201,N_97,N_1345);
and U2202 (N_2202,N_1275,N_1825);
or U2203 (N_2203,N_844,N_1474);
nand U2204 (N_2204,N_807,N_1801);
and U2205 (N_2205,N_488,N_434);
and U2206 (N_2206,N_258,N_476);
xnor U2207 (N_2207,N_1467,N_1125);
nand U2208 (N_2208,N_1201,N_1564);
nor U2209 (N_2209,N_1343,N_840);
and U2210 (N_2210,N_1648,N_166);
and U2211 (N_2211,N_1817,N_1011);
and U2212 (N_2212,N_1136,N_1865);
nand U2213 (N_2213,N_774,N_1182);
or U2214 (N_2214,N_564,N_546);
xnor U2215 (N_2215,N_152,N_871);
and U2216 (N_2216,N_756,N_65);
or U2217 (N_2217,N_285,N_992);
nand U2218 (N_2218,N_998,N_1212);
nand U2219 (N_2219,N_953,N_1941);
nand U2220 (N_2220,N_186,N_850);
nand U2221 (N_2221,N_64,N_1490);
nand U2222 (N_2222,N_818,N_1945);
and U2223 (N_2223,N_852,N_1388);
nor U2224 (N_2224,N_553,N_881);
xnor U2225 (N_2225,N_722,N_1227);
and U2226 (N_2226,N_1582,N_1053);
nand U2227 (N_2227,N_172,N_1625);
and U2228 (N_2228,N_1047,N_1107);
and U2229 (N_2229,N_841,N_373);
or U2230 (N_2230,N_417,N_1760);
and U2231 (N_2231,N_272,N_213);
and U2232 (N_2232,N_1088,N_1128);
and U2233 (N_2233,N_699,N_1464);
xnor U2234 (N_2234,N_606,N_1699);
nor U2235 (N_2235,N_955,N_720);
nand U2236 (N_2236,N_755,N_1966);
xor U2237 (N_2237,N_819,N_1282);
nand U2238 (N_2238,N_787,N_357);
nand U2239 (N_2239,N_1040,N_1783);
nor U2240 (N_2240,N_674,N_1741);
or U2241 (N_2241,N_1307,N_1037);
and U2242 (N_2242,N_1593,N_237);
and U2243 (N_2243,N_1093,N_1556);
and U2244 (N_2244,N_1391,N_1691);
nand U2245 (N_2245,N_1150,N_1590);
xor U2246 (N_2246,N_886,N_1469);
xnor U2247 (N_2247,N_320,N_421);
nor U2248 (N_2248,N_347,N_1476);
and U2249 (N_2249,N_538,N_692);
xnor U2250 (N_2250,N_1437,N_1957);
nor U2251 (N_2251,N_1919,N_1317);
xor U2252 (N_2252,N_846,N_1813);
nand U2253 (N_2253,N_39,N_1521);
xnor U2254 (N_2254,N_49,N_251);
nor U2255 (N_2255,N_1165,N_946);
nand U2256 (N_2256,N_1508,N_1733);
xor U2257 (N_2257,N_1010,N_366);
or U2258 (N_2258,N_1687,N_1174);
nand U2259 (N_2259,N_1714,N_1836);
nor U2260 (N_2260,N_981,N_16);
nand U2261 (N_2261,N_1381,N_1674);
and U2262 (N_2262,N_1851,N_941);
nand U2263 (N_2263,N_1228,N_741);
nand U2264 (N_2264,N_1771,N_3);
nand U2265 (N_2265,N_1629,N_1495);
and U2266 (N_2266,N_603,N_1871);
xnor U2267 (N_2267,N_7,N_156);
xnor U2268 (N_2268,N_680,N_588);
xnor U2269 (N_2269,N_1627,N_1274);
nor U2270 (N_2270,N_1751,N_817);
nor U2271 (N_2271,N_1331,N_380);
or U2272 (N_2272,N_1014,N_1818);
xor U2273 (N_2273,N_348,N_1754);
nor U2274 (N_2274,N_1178,N_310);
and U2275 (N_2275,N_1639,N_369);
nand U2276 (N_2276,N_221,N_737);
and U2277 (N_2277,N_386,N_1689);
xnor U2278 (N_2278,N_517,N_512);
nor U2279 (N_2279,N_771,N_1030);
xnor U2280 (N_2280,N_495,N_53);
or U2281 (N_2281,N_1158,N_584);
nand U2282 (N_2282,N_684,N_638);
or U2283 (N_2283,N_748,N_47);
xnor U2284 (N_2284,N_1724,N_48);
nor U2285 (N_2285,N_649,N_502);
xnor U2286 (N_2286,N_1393,N_1557);
and U2287 (N_2287,N_1042,N_1790);
nand U2288 (N_2288,N_1705,N_1113);
or U2289 (N_2289,N_1623,N_768);
nand U2290 (N_2290,N_914,N_980);
and U2291 (N_2291,N_1278,N_595);
nand U2292 (N_2292,N_975,N_1747);
nand U2293 (N_2293,N_1591,N_171);
or U2294 (N_2294,N_374,N_1498);
nand U2295 (N_2295,N_1631,N_754);
xnor U2296 (N_2296,N_1764,N_1492);
nand U2297 (N_2297,N_295,N_1555);
nor U2298 (N_2298,N_1344,N_1742);
nand U2299 (N_2299,N_639,N_764);
nand U2300 (N_2300,N_1337,N_1329);
xnor U2301 (N_2301,N_483,N_1837);
nor U2302 (N_2302,N_261,N_1264);
or U2303 (N_2303,N_454,N_134);
nor U2304 (N_2304,N_713,N_1915);
nor U2305 (N_2305,N_1749,N_727);
xor U2306 (N_2306,N_645,N_343);
xor U2307 (N_2307,N_560,N_67);
nand U2308 (N_2308,N_738,N_133);
nand U2309 (N_2309,N_170,N_1361);
and U2310 (N_2310,N_1788,N_874);
nand U2311 (N_2311,N_1529,N_612);
nand U2312 (N_2312,N_519,N_1359);
nor U2313 (N_2313,N_1798,N_982);
nand U2314 (N_2314,N_542,N_1399);
or U2315 (N_2315,N_1197,N_1101);
or U2316 (N_2316,N_1860,N_1897);
nor U2317 (N_2317,N_1124,N_333);
nand U2318 (N_2318,N_1130,N_695);
nand U2319 (N_2319,N_1038,N_273);
and U2320 (N_2320,N_388,N_890);
xor U2321 (N_2321,N_450,N_1727);
and U2322 (N_2322,N_759,N_1440);
or U2323 (N_2323,N_1558,N_376);
or U2324 (N_2324,N_629,N_521);
xnor U2325 (N_2325,N_643,N_1511);
nor U2326 (N_2326,N_1937,N_1487);
or U2327 (N_2327,N_277,N_1952);
nor U2328 (N_2328,N_677,N_339);
nor U2329 (N_2329,N_1311,N_30);
xor U2330 (N_2330,N_414,N_1665);
and U2331 (N_2331,N_404,N_753);
xnor U2332 (N_2332,N_1990,N_484);
nor U2333 (N_2333,N_1262,N_1459);
xor U2334 (N_2334,N_963,N_387);
and U2335 (N_2335,N_207,N_669);
nor U2336 (N_2336,N_125,N_1884);
and U2337 (N_2337,N_1261,N_22);
nor U2338 (N_2338,N_321,N_1185);
nand U2339 (N_2339,N_1672,N_909);
and U2340 (N_2340,N_800,N_616);
nor U2341 (N_2341,N_1183,N_238);
xor U2342 (N_2342,N_335,N_1970);
nor U2343 (N_2343,N_25,N_1611);
xor U2344 (N_2344,N_480,N_358);
and U2345 (N_2345,N_1679,N_586);
or U2346 (N_2346,N_464,N_1921);
or U2347 (N_2347,N_1924,N_52);
or U2348 (N_2348,N_765,N_1554);
nor U2349 (N_2349,N_1898,N_1748);
nor U2350 (N_2350,N_1523,N_262);
nand U2351 (N_2351,N_1281,N_766);
xor U2352 (N_2352,N_158,N_1402);
xor U2353 (N_2353,N_405,N_1095);
nor U2354 (N_2354,N_508,N_1064);
and U2355 (N_2355,N_735,N_1765);
nand U2356 (N_2356,N_1256,N_475);
nor U2357 (N_2357,N_1857,N_114);
nor U2358 (N_2358,N_1021,N_1209);
nor U2359 (N_2359,N_160,N_1877);
nand U2360 (N_2360,N_301,N_1314);
nand U2361 (N_2361,N_1782,N_578);
and U2362 (N_2362,N_785,N_917);
xor U2363 (N_2363,N_1382,N_636);
xnor U2364 (N_2364,N_469,N_1930);
and U2365 (N_2365,N_1632,N_933);
xnor U2366 (N_2366,N_658,N_651);
or U2367 (N_2367,N_1795,N_1767);
or U2368 (N_2368,N_1572,N_82);
or U2369 (N_2369,N_611,N_1740);
or U2370 (N_2370,N_1892,N_142);
xnor U2371 (N_2371,N_922,N_468);
nor U2372 (N_2372,N_1059,N_1294);
or U2373 (N_2373,N_1408,N_1028);
and U2374 (N_2374,N_1719,N_592);
nor U2375 (N_2375,N_1586,N_127);
nor U2376 (N_2376,N_1766,N_1856);
and U2377 (N_2377,N_1988,N_28);
nor U2378 (N_2378,N_225,N_164);
and U2379 (N_2379,N_290,N_1842);
nand U2380 (N_2380,N_1194,N_1859);
or U2381 (N_2381,N_529,N_936);
and U2382 (N_2382,N_1601,N_747);
xor U2383 (N_2383,N_530,N_1188);
nand U2384 (N_2384,N_9,N_1400);
nor U2385 (N_2385,N_1483,N_1079);
nand U2386 (N_2386,N_956,N_1597);
xor U2387 (N_2387,N_367,N_883);
xor U2388 (N_2388,N_1939,N_1330);
or U2389 (N_2389,N_1969,N_1237);
nor U2390 (N_2390,N_541,N_1651);
or U2391 (N_2391,N_1875,N_1647);
xor U2392 (N_2392,N_1211,N_397);
nor U2393 (N_2393,N_1364,N_1973);
xnor U2394 (N_2394,N_884,N_1610);
and U2395 (N_2395,N_283,N_1273);
and U2396 (N_2396,N_1953,N_510);
nand U2397 (N_2397,N_691,N_625);
xnor U2398 (N_2398,N_1176,N_1671);
nand U2399 (N_2399,N_1678,N_1878);
xnor U2400 (N_2400,N_1300,N_196);
xor U2401 (N_2401,N_1001,N_1649);
nor U2402 (N_2402,N_1901,N_477);
and U2403 (N_2403,N_73,N_1707);
or U2404 (N_2404,N_1443,N_317);
or U2405 (N_2405,N_1811,N_26);
and U2406 (N_2406,N_379,N_1718);
nor U2407 (N_2407,N_1950,N_1468);
nor U2408 (N_2408,N_1205,N_702);
nor U2409 (N_2409,N_707,N_33);
and U2410 (N_2410,N_867,N_242);
nand U2411 (N_2411,N_126,N_887);
xor U2412 (N_2412,N_1236,N_1734);
nand U2413 (N_2413,N_1874,N_1151);
nand U2414 (N_2414,N_770,N_718);
nand U2415 (N_2415,N_1304,N_490);
and U2416 (N_2416,N_460,N_842);
nor U2417 (N_2417,N_222,N_985);
and U2418 (N_2418,N_1159,N_1670);
and U2419 (N_2419,N_1757,N_1138);
xor U2420 (N_2420,N_1202,N_1362);
nand U2421 (N_2421,N_847,N_281);
or U2422 (N_2422,N_128,N_1100);
xnor U2423 (N_2423,N_831,N_403);
and U2424 (N_2424,N_1333,N_270);
nor U2425 (N_2425,N_219,N_661);
nand U2426 (N_2426,N_1077,N_1635);
nand U2427 (N_2427,N_804,N_1535);
xnor U2428 (N_2428,N_1822,N_590);
and U2429 (N_2429,N_494,N_1279);
xnor U2430 (N_2430,N_1530,N_306);
and U2431 (N_2431,N_994,N_515);
and U2432 (N_2432,N_401,N_1646);
xor U2433 (N_2433,N_1094,N_1545);
or U2434 (N_2434,N_122,N_31);
or U2435 (N_2435,N_1980,N_772);
nand U2436 (N_2436,N_1074,N_154);
or U2437 (N_2437,N_1896,N_1164);
or U2438 (N_2438,N_1615,N_383);
and U2439 (N_2439,N_1887,N_140);
or U2440 (N_2440,N_845,N_299);
xor U2441 (N_2441,N_1004,N_1607);
nor U2442 (N_2442,N_1845,N_1522);
or U2443 (N_2443,N_799,N_1057);
nand U2444 (N_2444,N_314,N_1034);
or U2445 (N_2445,N_330,N_169);
nand U2446 (N_2446,N_1427,N_858);
and U2447 (N_2447,N_534,N_408);
xnor U2448 (N_2448,N_1470,N_121);
and U2449 (N_2449,N_1655,N_676);
or U2450 (N_2450,N_1481,N_1750);
nand U2451 (N_2451,N_473,N_577);
nand U2452 (N_2452,N_520,N_863);
xnor U2453 (N_2453,N_191,N_1108);
xnor U2454 (N_2454,N_1694,N_1786);
and U2455 (N_2455,N_706,N_513);
xor U2456 (N_2456,N_1827,N_1574);
nor U2457 (N_2457,N_202,N_1532);
xnor U2458 (N_2458,N_1213,N_199);
or U2459 (N_2459,N_1514,N_1485);
nor U2460 (N_2460,N_1179,N_829);
xnor U2461 (N_2461,N_1503,N_316);
and U2462 (N_2462,N_593,N_1111);
or U2463 (N_2463,N_518,N_1208);
or U2464 (N_2464,N_1420,N_605);
or U2465 (N_2465,N_580,N_1527);
nand U2466 (N_2466,N_243,N_447);
xnor U2467 (N_2467,N_463,N_1891);
xor U2468 (N_2468,N_596,N_437);
and U2469 (N_2469,N_816,N_123);
or U2470 (N_2470,N_433,N_1230);
xnor U2471 (N_2471,N_83,N_532);
and U2472 (N_2472,N_1473,N_1098);
nand U2473 (N_2473,N_332,N_607);
xor U2474 (N_2474,N_1423,N_1983);
xor U2475 (N_2475,N_1613,N_1886);
and U2476 (N_2476,N_1805,N_1335);
xnor U2477 (N_2477,N_120,N_974);
nor U2478 (N_2478,N_1882,N_59);
nor U2479 (N_2479,N_1895,N_449);
nor U2480 (N_2480,N_964,N_795);
and U2481 (N_2481,N_1421,N_1637);
nor U2482 (N_2482,N_752,N_1149);
nand U2483 (N_2483,N_815,N_1787);
nor U2484 (N_2484,N_1031,N_1367);
or U2485 (N_2485,N_319,N_1612);
and U2486 (N_2486,N_812,N_1738);
or U2487 (N_2487,N_231,N_796);
xor U2488 (N_2488,N_75,N_724);
and U2489 (N_2489,N_1796,N_1577);
nor U2490 (N_2490,N_535,N_393);
nand U2491 (N_2491,N_1043,N_1499);
xnor U2492 (N_2492,N_411,N_71);
or U2493 (N_2493,N_61,N_200);
xnor U2494 (N_2494,N_1200,N_182);
nand U2495 (N_2495,N_141,N_1447);
nor U2496 (N_2496,N_1491,N_620);
and U2497 (N_2497,N_1500,N_621);
and U2498 (N_2498,N_792,N_1962);
nand U2499 (N_2499,N_915,N_138);
nand U2500 (N_2500,N_877,N_1458);
nand U2501 (N_2501,N_425,N_23);
xor U2502 (N_2502,N_1561,N_1280);
and U2503 (N_2503,N_1044,N_1244);
nand U2504 (N_2504,N_1155,N_412);
or U2505 (N_2505,N_1196,N_1698);
or U2506 (N_2506,N_540,N_1616);
xnor U2507 (N_2507,N_835,N_948);
or U2508 (N_2508,N_400,N_989);
or U2509 (N_2509,N_1016,N_1413);
nor U2510 (N_2510,N_1287,N_300);
or U2511 (N_2511,N_1667,N_1784);
nor U2512 (N_2512,N_378,N_1163);
xor U2513 (N_2513,N_1982,N_708);
xor U2514 (N_2514,N_304,N_843);
nor U2515 (N_2515,N_951,N_1267);
nand U2516 (N_2516,N_657,N_1793);
and U2517 (N_2517,N_1501,N_1019);
xor U2518 (N_2518,N_1082,N_1729);
nand U2519 (N_2519,N_1448,N_1336);
or U2520 (N_2520,N_1407,N_857);
or U2521 (N_2521,N_635,N_1573);
nand U2522 (N_2522,N_780,N_783);
xor U2523 (N_2523,N_551,N_55);
nor U2524 (N_2524,N_1302,N_1020);
nand U2525 (N_2525,N_1905,N_1682);
or U2526 (N_2526,N_43,N_701);
xor U2527 (N_2527,N_967,N_174);
and U2528 (N_2528,N_749,N_626);
nand U2529 (N_2529,N_100,N_391);
xor U2530 (N_2530,N_1517,N_1022);
nor U2531 (N_2531,N_1,N_1630);
or U2532 (N_2532,N_986,N_209);
xor U2533 (N_2533,N_98,N_420);
nand U2534 (N_2534,N_382,N_1791);
nand U2535 (N_2535,N_1693,N_587);
xnor U2536 (N_2536,N_1218,N_470);
nor U2537 (N_2537,N_1231,N_1428);
xnor U2538 (N_2538,N_390,N_1415);
nor U2539 (N_2539,N_823,N_687);
nor U2540 (N_2540,N_1235,N_1567);
or U2541 (N_2541,N_1550,N_1668);
nand U2542 (N_2542,N_711,N_507);
xnor U2543 (N_2543,N_1217,N_583);
and U2544 (N_2544,N_1334,N_1652);
nand U2545 (N_2545,N_183,N_1758);
nand U2546 (N_2546,N_1942,N_445);
nand U2547 (N_2547,N_1755,N_1141);
nand U2548 (N_2548,N_1434,N_745);
or U2549 (N_2549,N_1662,N_1864);
nor U2550 (N_2550,N_1599,N_1835);
nand U2551 (N_2551,N_431,N_349);
or U2552 (N_2552,N_950,N_566);
nand U2553 (N_2553,N_1316,N_1513);
nand U2554 (N_2554,N_1494,N_288);
or U2555 (N_2555,N_1947,N_1313);
nand U2556 (N_2556,N_1638,N_525);
nor U2557 (N_2557,N_1608,N_1488);
nand U2558 (N_2558,N_1838,N_660);
nand U2559 (N_2559,N_1568,N_547);
or U2560 (N_2560,N_1614,N_1873);
and U2561 (N_2561,N_94,N_452);
or U2562 (N_2562,N_1132,N_1562);
xnor U2563 (N_2563,N_779,N_1223);
xnor U2564 (N_2564,N_679,N_1171);
nor U2565 (N_2565,N_928,N_1370);
xor U2566 (N_2566,N_653,N_214);
xnor U2567 (N_2567,N_91,N_143);
nand U2568 (N_2568,N_1269,N_1394);
nor U2569 (N_2569,N_1505,N_1833);
nor U2570 (N_2570,N_1826,N_506);
xor U2571 (N_2571,N_1078,N_1424);
xnor U2572 (N_2572,N_565,N_315);
nor U2573 (N_2573,N_1596,N_977);
nand U2574 (N_2574,N_1539,N_514);
and U2575 (N_2575,N_944,N_1525);
xnor U2576 (N_2576,N_1518,N_205);
nand U2577 (N_2577,N_723,N_1007);
and U2578 (N_2578,N_1266,N_20);
and U2579 (N_2579,N_381,N_1192);
xnor U2580 (N_2580,N_1913,N_1026);
nand U2581 (N_2581,N_1702,N_1995);
or U2582 (N_2582,N_1916,N_220);
nand U2583 (N_2583,N_1722,N_1986);
xnor U2584 (N_2584,N_509,N_675);
or U2585 (N_2585,N_1123,N_617);
and U2586 (N_2586,N_1536,N_1971);
or U2587 (N_2587,N_1117,N_1692);
and U2588 (N_2588,N_1820,N_1365);
xor U2589 (N_2589,N_945,N_988);
nand U2590 (N_2590,N_851,N_1115);
xor U2591 (N_2591,N_323,N_155);
nor U2592 (N_2592,N_1585,N_1310);
or U2593 (N_2593,N_1881,N_1085);
nand U2594 (N_2594,N_1144,N_1676);
nor U2595 (N_2595,N_1318,N_921);
or U2596 (N_2596,N_526,N_809);
xnor U2597 (N_2597,N_1084,N_678);
xnor U2598 (N_2598,N_124,N_1862);
and U2599 (N_2599,N_1769,N_1861);
and U2600 (N_2600,N_428,N_1018);
nand U2601 (N_2601,N_557,N_1312);
and U2602 (N_2602,N_1519,N_112);
and U2603 (N_2603,N_1566,N_424);
nand U2604 (N_2604,N_1528,N_1780);
xnor U2605 (N_2605,N_1048,N_1587);
nor U2606 (N_2606,N_1029,N_107);
and U2607 (N_2607,N_698,N_150);
or U2608 (N_2608,N_524,N_1452);
nor U2609 (N_2609,N_1170,N_81);
nand U2610 (N_2610,N_904,N_1025);
or U2611 (N_2611,N_608,N_1776);
nand U2612 (N_2612,N_1543,N_1069);
nand U2613 (N_2613,N_1372,N_810);
or U2614 (N_2614,N_1046,N_108);
xnor U2615 (N_2615,N_1060,N_959);
and U2616 (N_2616,N_1509,N_1584);
nor U2617 (N_2617,N_361,N_896);
xnor U2618 (N_2618,N_599,N_1173);
xnor U2619 (N_2619,N_1841,N_318);
and U2620 (N_2620,N_892,N_1697);
xor U2621 (N_2621,N_554,N_1929);
or U2622 (N_2622,N_1979,N_1852);
and U2623 (N_2623,N_1524,N_245);
nand U2624 (N_2624,N_987,N_930);
or U2625 (N_2625,N_1189,N_1506);
or U2626 (N_2626,N_1761,N_1058);
and U2627 (N_2627,N_1375,N_432);
and U2628 (N_2628,N_600,N_1376);
xor U2629 (N_2629,N_686,N_1938);
or U2630 (N_2630,N_834,N_1619);
nand U2631 (N_2631,N_1569,N_1147);
or U2632 (N_2632,N_1955,N_889);
and U2633 (N_2633,N_326,N_1210);
nand U2634 (N_2634,N_743,N_558);
and U2635 (N_2635,N_957,N_574);
and U2636 (N_2636,N_869,N_1232);
nand U2637 (N_2637,N_559,N_384);
nand U2638 (N_2638,N_5,N_18);
nand U2639 (N_2639,N_1618,N_352);
nor U2640 (N_2640,N_1404,N_1992);
nor U2641 (N_2641,N_1297,N_1133);
and U2642 (N_2642,N_531,N_630);
nand U2643 (N_2643,N_267,N_910);
xnor U2644 (N_2644,N_1907,N_271);
xnor U2645 (N_2645,N_1685,N_777);
and U2646 (N_2646,N_1549,N_1911);
or U2647 (N_2647,N_328,N_1479);
nor U2648 (N_2648,N_1216,N_1355);
nor U2649 (N_2649,N_824,N_457);
nand U2650 (N_2650,N_640,N_662);
or U2651 (N_2651,N_62,N_1119);
and U2652 (N_2652,N_1204,N_833);
or U2653 (N_2653,N_1268,N_179);
or U2654 (N_2654,N_1721,N_935);
nor U2655 (N_2655,N_602,N_268);
nor U2656 (N_2656,N_113,N_878);
nor U2657 (N_2657,N_1248,N_1808);
nor U2658 (N_2658,N_1943,N_1368);
nand U2659 (N_2659,N_1775,N_919);
xnor U2660 (N_2660,N_1664,N_338);
or U2661 (N_2661,N_1341,N_175);
xnor U2662 (N_2662,N_1036,N_1325);
xnor U2663 (N_2663,N_873,N_805);
nor U2664 (N_2664,N_1105,N_406);
xnor U2665 (N_2665,N_279,N_226);
nor U2666 (N_2666,N_991,N_312);
and U2667 (N_2667,N_1076,N_37);
nand U2668 (N_2668,N_1976,N_482);
and U2669 (N_2669,N_1520,N_1438);
nand U2670 (N_2670,N_1008,N_206);
xnor U2671 (N_2671,N_1683,N_498);
xor U2672 (N_2672,N_730,N_1800);
xor U2673 (N_2673,N_1143,N_227);
and U2674 (N_2674,N_1677,N_1482);
nand U2675 (N_2675,N_728,N_688);
nand U2676 (N_2676,N_1690,N_856);
nor U2677 (N_2677,N_423,N_1804);
xnor U2678 (N_2678,N_341,N_872);
nor U2679 (N_2679,N_1739,N_961);
nor U2680 (N_2680,N_610,N_911);
or U2681 (N_2681,N_1732,N_442);
nand U2682 (N_2682,N_364,N_322);
nor U2683 (N_2683,N_1065,N_426);
nand U2684 (N_2684,N_232,N_1439);
and U2685 (N_2685,N_732,N_898);
nor U2686 (N_2686,N_1720,N_203);
nand U2687 (N_2687,N_1129,N_1386);
nand U2688 (N_2688,N_276,N_462);
xnor U2689 (N_2689,N_446,N_1746);
xor U2690 (N_2690,N_233,N_1908);
and U2691 (N_2691,N_999,N_876);
nor U2692 (N_2692,N_790,N_1390);
or U2693 (N_2693,N_663,N_1219);
nand U2694 (N_2694,N_415,N_1931);
nor U2695 (N_2695,N_1948,N_329);
xnor U2696 (N_2696,N_195,N_736);
nor U2697 (N_2697,N_1696,N_1777);
xor U2698 (N_2698,N_1779,N_1015);
nor U2699 (N_2699,N_656,N_1996);
nand U2700 (N_2700,N_789,N_1091);
and U2701 (N_2701,N_1288,N_954);
xor U2702 (N_2702,N_646,N_773);
xor U2703 (N_2703,N_830,N_913);
and U2704 (N_2704,N_1451,N_511);
xnor U2705 (N_2705,N_327,N_1206);
nor U2706 (N_2706,N_545,N_1465);
or U2707 (N_2707,N_1960,N_1704);
and U2708 (N_2708,N_1000,N_569);
and U2709 (N_2709,N_1024,N_13);
and U2710 (N_2710,N_165,N_1422);
nor U2711 (N_2711,N_371,N_1137);
and U2712 (N_2712,N_1172,N_1241);
xnor U2713 (N_2713,N_1162,N_1560);
nor U2714 (N_2714,N_1377,N_80);
nand U2715 (N_2715,N_1291,N_848);
xor U2716 (N_2716,N_284,N_1709);
and U2717 (N_2717,N_1242,N_116);
xnor U2718 (N_2718,N_1643,N_444);
xnor U2719 (N_2719,N_1073,N_1579);
and U2720 (N_2720,N_193,N_813);
nor U2721 (N_2721,N_291,N_478);
and U2722 (N_2722,N_705,N_615);
xnor U2723 (N_2723,N_794,N_282);
and U2724 (N_2724,N_177,N_861);
or U2725 (N_2725,N_1773,N_1106);
and U2726 (N_2726,N_1595,N_659);
nor U2727 (N_2727,N_1958,N_1180);
nand U2728 (N_2728,N_1661,N_854);
nor U2729 (N_2729,N_767,N_778);
and U2730 (N_2730,N_694,N_1906);
or U2731 (N_2731,N_296,N_1087);
nand U2732 (N_2732,N_1051,N_825);
or U2733 (N_2733,N_923,N_1272);
and U2734 (N_2734,N_1762,N_106);
xor U2735 (N_2735,N_1753,N_1657);
xor U2736 (N_2736,N_1636,N_360);
or U2737 (N_2737,N_973,N_1324);
or U2738 (N_2738,N_673,N_1118);
nand U2739 (N_2739,N_543,N_467);
nand U2740 (N_2740,N_716,N_355);
xor U2741 (N_2741,N_868,N_1954);
nand U2742 (N_2742,N_1380,N_672);
or U2743 (N_2743,N_422,N_6);
and U2744 (N_2744,N_1713,N_1902);
and U2745 (N_2745,N_1167,N_372);
nand U2746 (N_2746,N_1581,N_1049);
nor U2747 (N_2747,N_1238,N_1736);
or U2748 (N_2748,N_1565,N_1675);
or U2749 (N_2749,N_1305,N_252);
or U2750 (N_2750,N_1819,N_1175);
or U2751 (N_2751,N_683,N_302);
nor U2752 (N_2752,N_527,N_1249);
nor U2753 (N_2753,N_1815,N_1168);
and U2754 (N_2754,N_1717,N_1270);
nor U2755 (N_2755,N_1645,N_1666);
nor U2756 (N_2756,N_24,N_1604);
and U2757 (N_2757,N_96,N_487);
nor U2758 (N_2758,N_1803,N_46);
nand U2759 (N_2759,N_609,N_647);
nand U2760 (N_2760,N_1418,N_1462);
or U2761 (N_2761,N_1012,N_820);
xor U2762 (N_2762,N_1542,N_563);
nand U2763 (N_2763,N_1284,N_131);
nor U2764 (N_2764,N_937,N_1429);
xor U2765 (N_2765,N_968,N_280);
xor U2766 (N_2766,N_623,N_1306);
nand U2767 (N_2767,N_1056,N_1589);
or U2768 (N_2768,N_1484,N_1234);
or U2769 (N_2769,N_1285,N_436);
xnor U2770 (N_2770,N_430,N_1121);
nand U2771 (N_2771,N_471,N_1383);
nor U2772 (N_2772,N_1526,N_1756);
and U2773 (N_2773,N_1435,N_1342);
or U2774 (N_2774,N_1894,N_1347);
nor U2775 (N_2775,N_375,N_1538);
xnor U2776 (N_2776,N_266,N_1703);
nand U2777 (N_2777,N_239,N_757);
xor U2778 (N_2778,N_655,N_562);
or U2779 (N_2779,N_1669,N_744);
nor U2780 (N_2780,N_1092,N_1853);
xor U2781 (N_2781,N_190,N_966);
or U2782 (N_2782,N_41,N_1726);
nor U2783 (N_2783,N_439,N_760);
nand U2784 (N_2784,N_255,N_552);
xnor U2785 (N_2785,N_1700,N_1812);
and U2786 (N_2786,N_11,N_1626);
or U2787 (N_2787,N_670,N_1922);
nor U2788 (N_2788,N_109,N_1169);
or U2789 (N_2789,N_614,N_503);
nor U2790 (N_2790,N_1363,N_758);
xor U2791 (N_2791,N_1009,N_1240);
nor U2792 (N_2792,N_54,N_236);
or U2793 (N_2793,N_70,N_1340);
xor U2794 (N_2794,N_354,N_700);
nand U2795 (N_2795,N_230,N_864);
nor U2796 (N_2796,N_1220,N_1617);
nor U2797 (N_2797,N_837,N_1504);
xor U2798 (N_2798,N_93,N_1588);
nand U2799 (N_2799,N_1292,N_176);
nand U2800 (N_2800,N_342,N_1430);
and U2801 (N_2801,N_505,N_1806);
nor U2802 (N_2802,N_1416,N_934);
nand U2803 (N_2803,N_763,N_294);
and U2804 (N_2804,N_1807,N_1283);
nand U2805 (N_2805,N_287,N_1122);
nand U2806 (N_2806,N_459,N_1928);
nor U2807 (N_2807,N_1239,N_1984);
and U2808 (N_2808,N_1855,N_1350);
xor U2809 (N_2809,N_346,N_178);
nor U2810 (N_2810,N_918,N_742);
or U2811 (N_2811,N_1352,N_241);
xnor U2812 (N_2812,N_173,N_1867);
or U2813 (N_2813,N_1936,N_194);
and U2814 (N_2814,N_1198,N_35);
nand U2815 (N_2815,N_798,N_895);
and U2816 (N_2816,N_1412,N_826);
nand U2817 (N_2817,N_1659,N_443);
or U2818 (N_2818,N_1259,N_1072);
and U2819 (N_2819,N_185,N_1397);
nor U2820 (N_2820,N_1050,N_762);
or U2821 (N_2821,N_85,N_924);
nand U2822 (N_2822,N_1449,N_1120);
nand U2823 (N_2823,N_1103,N_313);
xnor U2824 (N_2824,N_682,N_1052);
or U2825 (N_2825,N_1701,N_103);
or U2826 (N_2826,N_458,N_1145);
and U2827 (N_2827,N_1493,N_161);
nor U2828 (N_2828,N_19,N_1634);
or U2829 (N_2829,N_1964,N_151);
and U2830 (N_2830,N_38,N_1354);
and U2831 (N_2831,N_211,N_949);
nand U2832 (N_2832,N_1768,N_1850);
or U2833 (N_2833,N_1606,N_8);
nand U2834 (N_2834,N_1032,N_1650);
nor U2835 (N_2835,N_1054,N_501);
or U2836 (N_2836,N_162,N_1863);
and U2837 (N_2837,N_984,N_1431);
or U2838 (N_2838,N_803,N_1222);
nand U2839 (N_2839,N_1299,N_1904);
and U2840 (N_2840,N_42,N_1417);
xor U2841 (N_2841,N_717,N_351);
and U2842 (N_2842,N_1985,N_582);
and U2843 (N_2843,N_1127,N_1903);
and U2844 (N_2844,N_970,N_1166);
or U2845 (N_2845,N_641,N_1398);
xor U2846 (N_2846,N_119,N_224);
nand U2847 (N_2847,N_983,N_1763);
and U2848 (N_2848,N_68,N_601);
and U2849 (N_2849,N_594,N_419);
and U2850 (N_2850,N_90,N_159);
and U2851 (N_2851,N_1515,N_619);
or U2852 (N_2852,N_465,N_1658);
or U2853 (N_2853,N_1977,N_1308);
and U2854 (N_2854,N_385,N_1809);
and U2855 (N_2855,N_1154,N_866);
or U2856 (N_2856,N_1096,N_1917);
nor U2857 (N_2857,N_10,N_1944);
nor U2858 (N_2858,N_362,N_286);
and U2859 (N_2859,N_1548,N_1286);
xor U2860 (N_2860,N_246,N_1387);
or U2861 (N_2861,N_88,N_44);
and U2862 (N_2862,N_855,N_1301);
nand U2863 (N_2863,N_228,N_1033);
nor U2864 (N_2864,N_624,N_853);
xor U2865 (N_2865,N_995,N_253);
or U2866 (N_2866,N_132,N_740);
nor U2867 (N_2867,N_1909,N_1384);
xnor U2868 (N_2868,N_932,N_1710);
nand U2869 (N_2869,N_1728,N_157);
xor U2870 (N_2870,N_1116,N_1725);
nand U2871 (N_2871,N_1743,N_585);
xor U2872 (N_2872,N_1510,N_849);
nor U2873 (N_2873,N_1378,N_344);
xor U2874 (N_2874,N_40,N_118);
xnor U2875 (N_2875,N_1253,N_234);
and U2876 (N_2876,N_1366,N_216);
nor U2877 (N_2877,N_1927,N_1673);
and U2878 (N_2878,N_1843,N_1177);
nor U2879 (N_2879,N_356,N_244);
and U2880 (N_2880,N_60,N_1502);
nand U2881 (N_2881,N_1706,N_1923);
or U2882 (N_2882,N_648,N_1644);
or U2883 (N_2883,N_1628,N_1322);
and U2884 (N_2884,N_671,N_188);
and U2885 (N_2885,N_746,N_148);
nor U2886 (N_2886,N_1063,N_1309);
and U2887 (N_2887,N_1353,N_1369);
nand U2888 (N_2888,N_1684,N_654);
nand U2889 (N_2889,N_1195,N_363);
or U2890 (N_2890,N_189,N_1940);
nor U2891 (N_2891,N_875,N_797);
nand U2892 (N_2892,N_139,N_1401);
and U2893 (N_2893,N_17,N_345);
and U2894 (N_2894,N_51,N_210);
xnor U2895 (N_2895,N_693,N_1695);
nor U2896 (N_2896,N_622,N_212);
nor U2897 (N_2897,N_1315,N_1257);
nor U2898 (N_2898,N_1507,N_77);
nor U2899 (N_2899,N_1914,N_905);
xnor U2900 (N_2900,N_474,N_697);
xnor U2901 (N_2901,N_1081,N_637);
xnor U2902 (N_2902,N_1583,N_832);
nor U2903 (N_2903,N_1840,N_1017);
nor U2904 (N_2904,N_1454,N_1975);
nor U2905 (N_2905,N_1013,N_979);
nand U2906 (N_2906,N_1061,N_275);
nor U2907 (N_2907,N_389,N_1346);
or U2908 (N_2908,N_1246,N_1890);
xor U2909 (N_2909,N_729,N_377);
nand U2910 (N_2910,N_1868,N_72);
and U2911 (N_2911,N_1512,N_1260);
and U2912 (N_2912,N_1006,N_1879);
xnor U2913 (N_2913,N_1893,N_1949);
nand U2914 (N_2914,N_555,N_353);
nand U2915 (N_2915,N_1580,N_1876);
nand U2916 (N_2916,N_136,N_1900);
nor U2917 (N_2917,N_1276,N_1471);
xnor U2918 (N_2918,N_1989,N_448);
nor U2919 (N_2919,N_441,N_1680);
and U2920 (N_2920,N_1250,N_440);
nor U2921 (N_2921,N_1251,N_1600);
and U2922 (N_2922,N_1444,N_859);
nand U2923 (N_2923,N_568,N_1298);
xnor U2924 (N_2924,N_102,N_631);
and U2925 (N_2925,N_350,N_298);
xnor U2926 (N_2926,N_1303,N_1453);
and U2927 (N_2927,N_734,N_14);
nand U2928 (N_2928,N_1226,N_1946);
or U2929 (N_2929,N_340,N_1245);
or U2930 (N_2930,N_1247,N_1974);
and U2931 (N_2931,N_793,N_523);
nand U2932 (N_2932,N_254,N_882);
and U2933 (N_2933,N_1571,N_969);
nor U2934 (N_2934,N_1987,N_1441);
xor U2935 (N_2935,N_461,N_1290);
or U2936 (N_2936,N_862,N_1086);
nor U2937 (N_2937,N_901,N_1023);
nand U2938 (N_2938,N_1910,N_1327);
nand U2939 (N_2939,N_1338,N_1027);
nor U2940 (N_2940,N_775,N_962);
nand U2941 (N_2941,N_456,N_398);
nand U2942 (N_2942,N_1296,N_1621);
nor U2943 (N_2943,N_500,N_731);
xnor U2944 (N_2944,N_665,N_240);
xnor U2945 (N_2945,N_1594,N_1624);
or U2946 (N_2946,N_604,N_942);
nor U2947 (N_2947,N_4,N_63);
nor U2948 (N_2948,N_947,N_278);
xnor U2949 (N_2949,N_1252,N_1466);
xor U2950 (N_2950,N_1802,N_1002);
xor U2951 (N_2951,N_466,N_1146);
nor U2952 (N_2952,N_1403,N_929);
or U2953 (N_2953,N_1935,N_453);
or U2954 (N_2954,N_264,N_1858);
xor U2955 (N_2955,N_1998,N_1785);
and U2956 (N_2956,N_87,N_1062);
xor U2957 (N_2957,N_269,N_726);
nor U2958 (N_2958,N_368,N_78);
or U2959 (N_2959,N_1243,N_1126);
nand U2960 (N_2960,N_247,N_1799);
xor U2961 (N_2961,N_263,N_187);
nor U2962 (N_2962,N_1295,N_1832);
nor U2963 (N_2963,N_307,N_1993);
or U2964 (N_2964,N_548,N_1715);
xor U2965 (N_2965,N_260,N_802);
or U2966 (N_2966,N_84,N_32);
xnor U2967 (N_2967,N_485,N_1265);
and U2968 (N_2968,N_1442,N_996);
nor U2969 (N_2969,N_256,N_1620);
and U2970 (N_2970,N_1323,N_750);
nor U2971 (N_2971,N_1663,N_751);
nor U2972 (N_2972,N_931,N_814);
nor U2973 (N_2973,N_1486,N_1576);
or U2974 (N_2974,N_435,N_571);
xor U2975 (N_2975,N_1956,N_1711);
nand U2976 (N_2976,N_74,N_822);
xor U2977 (N_2977,N_1460,N_111);
xnor U2978 (N_2978,N_786,N_297);
nor U2979 (N_2979,N_1633,N_402);
nand U2980 (N_2980,N_1461,N_714);
nor U2981 (N_2981,N_36,N_591);
nand U2982 (N_2982,N_248,N_1959);
xnor U2983 (N_2983,N_1157,N_891);
nand U2984 (N_2984,N_696,N_1114);
and U2985 (N_2985,N_1104,N_198);
nor U2986 (N_2986,N_528,N_828);
or U2987 (N_2987,N_1839,N_650);
xnor U2988 (N_2988,N_1080,N_1824);
nor U2989 (N_2989,N_1184,N_1640);
nand U2990 (N_2990,N_860,N_1445);
or U2991 (N_2991,N_1457,N_958);
nor U2992 (N_2992,N_144,N_888);
and U2993 (N_2993,N_1406,N_791);
xnor U2994 (N_2994,N_399,N_1810);
and U2995 (N_2995,N_137,N_664);
xnor U2996 (N_2996,N_149,N_1203);
and U2997 (N_2997,N_685,N_1225);
or U2998 (N_2998,N_1349,N_628);
nand U2999 (N_2999,N_1392,N_496);
nand U3000 (N_3000,N_1375,N_1326);
nor U3001 (N_3001,N_2,N_1784);
xnor U3002 (N_3002,N_578,N_1742);
and U3003 (N_3003,N_1199,N_287);
and U3004 (N_3004,N_1197,N_365);
nand U3005 (N_3005,N_415,N_456);
or U3006 (N_3006,N_494,N_126);
or U3007 (N_3007,N_1050,N_1854);
nand U3008 (N_3008,N_1121,N_1227);
xor U3009 (N_3009,N_613,N_1461);
nor U3010 (N_3010,N_412,N_1240);
and U3011 (N_3011,N_410,N_889);
nand U3012 (N_3012,N_841,N_1284);
or U3013 (N_3013,N_38,N_1135);
and U3014 (N_3014,N_1710,N_1970);
nand U3015 (N_3015,N_1470,N_80);
and U3016 (N_3016,N_711,N_615);
nand U3017 (N_3017,N_874,N_1453);
nor U3018 (N_3018,N_1549,N_850);
and U3019 (N_3019,N_1899,N_1942);
and U3020 (N_3020,N_1168,N_1340);
or U3021 (N_3021,N_1508,N_1686);
xnor U3022 (N_3022,N_271,N_1281);
or U3023 (N_3023,N_270,N_160);
nor U3024 (N_3024,N_249,N_474);
and U3025 (N_3025,N_595,N_1486);
nand U3026 (N_3026,N_38,N_264);
and U3027 (N_3027,N_1529,N_24);
xnor U3028 (N_3028,N_222,N_1714);
nand U3029 (N_3029,N_390,N_572);
and U3030 (N_3030,N_15,N_646);
xor U3031 (N_3031,N_1328,N_1635);
or U3032 (N_3032,N_1182,N_104);
or U3033 (N_3033,N_1075,N_1386);
nand U3034 (N_3034,N_952,N_1527);
xor U3035 (N_3035,N_515,N_1203);
xnor U3036 (N_3036,N_478,N_1969);
or U3037 (N_3037,N_636,N_44);
and U3038 (N_3038,N_1242,N_1643);
or U3039 (N_3039,N_868,N_406);
or U3040 (N_3040,N_880,N_1745);
xnor U3041 (N_3041,N_1779,N_1746);
xor U3042 (N_3042,N_956,N_913);
and U3043 (N_3043,N_1139,N_153);
xnor U3044 (N_3044,N_1707,N_438);
and U3045 (N_3045,N_857,N_750);
nand U3046 (N_3046,N_1268,N_882);
and U3047 (N_3047,N_1129,N_418);
or U3048 (N_3048,N_823,N_265);
or U3049 (N_3049,N_666,N_1312);
and U3050 (N_3050,N_1992,N_463);
xnor U3051 (N_3051,N_450,N_615);
xnor U3052 (N_3052,N_940,N_1839);
or U3053 (N_3053,N_1435,N_413);
nand U3054 (N_3054,N_1796,N_398);
nor U3055 (N_3055,N_560,N_753);
nor U3056 (N_3056,N_692,N_1299);
nor U3057 (N_3057,N_1250,N_435);
nand U3058 (N_3058,N_159,N_1096);
xor U3059 (N_3059,N_857,N_1171);
nand U3060 (N_3060,N_371,N_1576);
or U3061 (N_3061,N_1976,N_1509);
and U3062 (N_3062,N_1215,N_299);
or U3063 (N_3063,N_833,N_1495);
or U3064 (N_3064,N_648,N_670);
nor U3065 (N_3065,N_1479,N_1860);
nand U3066 (N_3066,N_279,N_568);
nand U3067 (N_3067,N_383,N_1274);
and U3068 (N_3068,N_634,N_1137);
nor U3069 (N_3069,N_781,N_357);
nor U3070 (N_3070,N_1993,N_1812);
and U3071 (N_3071,N_328,N_1986);
and U3072 (N_3072,N_696,N_1330);
nor U3073 (N_3073,N_1280,N_971);
nand U3074 (N_3074,N_1348,N_55);
nor U3075 (N_3075,N_1192,N_422);
or U3076 (N_3076,N_969,N_871);
nand U3077 (N_3077,N_110,N_1118);
nand U3078 (N_3078,N_1996,N_1882);
and U3079 (N_3079,N_1785,N_517);
and U3080 (N_3080,N_812,N_793);
or U3081 (N_3081,N_101,N_26);
nor U3082 (N_3082,N_1532,N_845);
nor U3083 (N_3083,N_1541,N_78);
and U3084 (N_3084,N_1547,N_1337);
nand U3085 (N_3085,N_682,N_851);
nor U3086 (N_3086,N_1802,N_1383);
xor U3087 (N_3087,N_930,N_1002);
nor U3088 (N_3088,N_1023,N_1528);
nor U3089 (N_3089,N_996,N_985);
nor U3090 (N_3090,N_558,N_623);
nand U3091 (N_3091,N_254,N_1644);
nand U3092 (N_3092,N_523,N_1610);
and U3093 (N_3093,N_1777,N_1247);
nand U3094 (N_3094,N_736,N_713);
xnor U3095 (N_3095,N_1831,N_1862);
xor U3096 (N_3096,N_192,N_1333);
nor U3097 (N_3097,N_1258,N_1097);
and U3098 (N_3098,N_965,N_193);
nand U3099 (N_3099,N_8,N_1434);
nor U3100 (N_3100,N_819,N_1167);
nand U3101 (N_3101,N_274,N_1987);
xor U3102 (N_3102,N_744,N_1010);
nor U3103 (N_3103,N_1057,N_1070);
and U3104 (N_3104,N_998,N_1553);
nor U3105 (N_3105,N_664,N_133);
nand U3106 (N_3106,N_373,N_981);
or U3107 (N_3107,N_449,N_929);
xnor U3108 (N_3108,N_745,N_1565);
xor U3109 (N_3109,N_459,N_1646);
nor U3110 (N_3110,N_1076,N_220);
nand U3111 (N_3111,N_1732,N_1358);
and U3112 (N_3112,N_1412,N_1068);
or U3113 (N_3113,N_1857,N_1635);
and U3114 (N_3114,N_1238,N_885);
nor U3115 (N_3115,N_1161,N_547);
and U3116 (N_3116,N_1259,N_1021);
nand U3117 (N_3117,N_661,N_1546);
nor U3118 (N_3118,N_156,N_733);
or U3119 (N_3119,N_229,N_1842);
and U3120 (N_3120,N_1021,N_372);
xnor U3121 (N_3121,N_1878,N_684);
nand U3122 (N_3122,N_66,N_53);
or U3123 (N_3123,N_1831,N_106);
and U3124 (N_3124,N_25,N_1106);
or U3125 (N_3125,N_1604,N_546);
nand U3126 (N_3126,N_1896,N_1360);
and U3127 (N_3127,N_1029,N_1835);
nor U3128 (N_3128,N_470,N_1744);
nor U3129 (N_3129,N_459,N_1995);
xor U3130 (N_3130,N_1688,N_202);
and U3131 (N_3131,N_1381,N_1504);
or U3132 (N_3132,N_867,N_1787);
nor U3133 (N_3133,N_963,N_1275);
nor U3134 (N_3134,N_61,N_54);
xnor U3135 (N_3135,N_1236,N_378);
nand U3136 (N_3136,N_1744,N_574);
or U3137 (N_3137,N_1935,N_934);
and U3138 (N_3138,N_1337,N_704);
or U3139 (N_3139,N_1959,N_289);
and U3140 (N_3140,N_575,N_1592);
nand U3141 (N_3141,N_509,N_763);
nor U3142 (N_3142,N_176,N_1555);
xnor U3143 (N_3143,N_1137,N_1100);
nor U3144 (N_3144,N_536,N_544);
and U3145 (N_3145,N_1844,N_1513);
nor U3146 (N_3146,N_589,N_479);
xnor U3147 (N_3147,N_1548,N_1672);
nor U3148 (N_3148,N_442,N_1643);
nand U3149 (N_3149,N_1624,N_1321);
nand U3150 (N_3150,N_216,N_1244);
nor U3151 (N_3151,N_468,N_325);
xnor U3152 (N_3152,N_852,N_777);
nand U3153 (N_3153,N_1019,N_723);
or U3154 (N_3154,N_1567,N_1641);
nor U3155 (N_3155,N_184,N_690);
nand U3156 (N_3156,N_584,N_986);
nand U3157 (N_3157,N_648,N_998);
xor U3158 (N_3158,N_1652,N_790);
nor U3159 (N_3159,N_814,N_553);
nand U3160 (N_3160,N_122,N_1775);
xor U3161 (N_3161,N_1202,N_1521);
xnor U3162 (N_3162,N_1008,N_1210);
nor U3163 (N_3163,N_1159,N_1345);
nand U3164 (N_3164,N_1421,N_432);
and U3165 (N_3165,N_184,N_415);
and U3166 (N_3166,N_91,N_659);
nand U3167 (N_3167,N_1257,N_690);
nor U3168 (N_3168,N_891,N_342);
and U3169 (N_3169,N_704,N_1075);
xor U3170 (N_3170,N_472,N_466);
or U3171 (N_3171,N_738,N_1104);
and U3172 (N_3172,N_646,N_496);
or U3173 (N_3173,N_42,N_603);
nor U3174 (N_3174,N_1650,N_593);
nor U3175 (N_3175,N_1225,N_1717);
or U3176 (N_3176,N_1659,N_1277);
or U3177 (N_3177,N_1658,N_1664);
or U3178 (N_3178,N_562,N_1);
and U3179 (N_3179,N_1240,N_838);
nor U3180 (N_3180,N_1301,N_1749);
or U3181 (N_3181,N_1782,N_1812);
or U3182 (N_3182,N_1010,N_264);
nand U3183 (N_3183,N_779,N_738);
xor U3184 (N_3184,N_987,N_594);
nand U3185 (N_3185,N_857,N_1894);
nand U3186 (N_3186,N_400,N_1052);
nand U3187 (N_3187,N_1778,N_997);
nor U3188 (N_3188,N_394,N_1407);
and U3189 (N_3189,N_1842,N_1638);
or U3190 (N_3190,N_232,N_1780);
xnor U3191 (N_3191,N_1280,N_301);
xor U3192 (N_3192,N_258,N_1954);
and U3193 (N_3193,N_1191,N_625);
nor U3194 (N_3194,N_731,N_1353);
nor U3195 (N_3195,N_1083,N_1020);
or U3196 (N_3196,N_1878,N_664);
nand U3197 (N_3197,N_1398,N_782);
nand U3198 (N_3198,N_1263,N_1041);
nand U3199 (N_3199,N_811,N_1060);
xnor U3200 (N_3200,N_1767,N_1744);
or U3201 (N_3201,N_1295,N_1741);
xor U3202 (N_3202,N_1879,N_1108);
and U3203 (N_3203,N_767,N_1566);
nor U3204 (N_3204,N_1235,N_416);
xnor U3205 (N_3205,N_732,N_97);
nor U3206 (N_3206,N_718,N_1502);
nor U3207 (N_3207,N_866,N_1112);
nor U3208 (N_3208,N_91,N_1446);
nand U3209 (N_3209,N_616,N_987);
nor U3210 (N_3210,N_1419,N_1358);
xor U3211 (N_3211,N_1303,N_641);
nand U3212 (N_3212,N_1727,N_1387);
xor U3213 (N_3213,N_1437,N_1629);
xnor U3214 (N_3214,N_1662,N_1128);
nor U3215 (N_3215,N_431,N_52);
nor U3216 (N_3216,N_413,N_1235);
nor U3217 (N_3217,N_1260,N_1295);
or U3218 (N_3218,N_817,N_1114);
and U3219 (N_3219,N_1124,N_1156);
or U3220 (N_3220,N_471,N_552);
and U3221 (N_3221,N_764,N_28);
and U3222 (N_3222,N_460,N_107);
nand U3223 (N_3223,N_1789,N_31);
or U3224 (N_3224,N_218,N_1958);
nor U3225 (N_3225,N_1667,N_1636);
xor U3226 (N_3226,N_894,N_1426);
nor U3227 (N_3227,N_1906,N_1980);
and U3228 (N_3228,N_462,N_1067);
nor U3229 (N_3229,N_1659,N_814);
or U3230 (N_3230,N_1570,N_1561);
nor U3231 (N_3231,N_192,N_1135);
xor U3232 (N_3232,N_1607,N_795);
xnor U3233 (N_3233,N_1533,N_1011);
nor U3234 (N_3234,N_1301,N_1639);
xor U3235 (N_3235,N_1097,N_1583);
and U3236 (N_3236,N_1768,N_983);
xnor U3237 (N_3237,N_284,N_927);
nor U3238 (N_3238,N_1315,N_419);
and U3239 (N_3239,N_552,N_389);
and U3240 (N_3240,N_105,N_557);
nand U3241 (N_3241,N_1017,N_1952);
or U3242 (N_3242,N_621,N_627);
and U3243 (N_3243,N_64,N_1094);
xor U3244 (N_3244,N_1955,N_344);
xnor U3245 (N_3245,N_955,N_169);
xor U3246 (N_3246,N_197,N_268);
nand U3247 (N_3247,N_1982,N_766);
and U3248 (N_3248,N_58,N_787);
xnor U3249 (N_3249,N_1270,N_1046);
and U3250 (N_3250,N_693,N_173);
nor U3251 (N_3251,N_1784,N_1020);
or U3252 (N_3252,N_1615,N_585);
nand U3253 (N_3253,N_252,N_749);
nor U3254 (N_3254,N_415,N_716);
xor U3255 (N_3255,N_165,N_890);
nor U3256 (N_3256,N_194,N_1569);
nand U3257 (N_3257,N_186,N_991);
xor U3258 (N_3258,N_1739,N_863);
nor U3259 (N_3259,N_163,N_1742);
nor U3260 (N_3260,N_1665,N_601);
or U3261 (N_3261,N_1373,N_700);
nor U3262 (N_3262,N_876,N_663);
and U3263 (N_3263,N_1014,N_783);
and U3264 (N_3264,N_1747,N_941);
nor U3265 (N_3265,N_1999,N_395);
xor U3266 (N_3266,N_112,N_583);
xnor U3267 (N_3267,N_1646,N_952);
xnor U3268 (N_3268,N_1149,N_692);
or U3269 (N_3269,N_998,N_1841);
xor U3270 (N_3270,N_54,N_1876);
nand U3271 (N_3271,N_1183,N_1216);
and U3272 (N_3272,N_598,N_843);
and U3273 (N_3273,N_1758,N_1031);
nor U3274 (N_3274,N_1292,N_1897);
or U3275 (N_3275,N_914,N_1978);
and U3276 (N_3276,N_1563,N_727);
nor U3277 (N_3277,N_1341,N_255);
and U3278 (N_3278,N_1985,N_406);
nor U3279 (N_3279,N_1784,N_1869);
nor U3280 (N_3280,N_227,N_756);
xnor U3281 (N_3281,N_476,N_1887);
xor U3282 (N_3282,N_397,N_1909);
xnor U3283 (N_3283,N_1575,N_14);
nor U3284 (N_3284,N_792,N_23);
or U3285 (N_3285,N_1062,N_341);
and U3286 (N_3286,N_743,N_202);
nor U3287 (N_3287,N_1335,N_159);
xnor U3288 (N_3288,N_897,N_10);
xnor U3289 (N_3289,N_404,N_258);
nand U3290 (N_3290,N_1483,N_835);
and U3291 (N_3291,N_281,N_82);
xnor U3292 (N_3292,N_1461,N_1622);
or U3293 (N_3293,N_1632,N_1843);
and U3294 (N_3294,N_873,N_1110);
nor U3295 (N_3295,N_424,N_135);
and U3296 (N_3296,N_1678,N_1883);
or U3297 (N_3297,N_1375,N_959);
nor U3298 (N_3298,N_1562,N_13);
and U3299 (N_3299,N_1781,N_270);
or U3300 (N_3300,N_1161,N_487);
nand U3301 (N_3301,N_866,N_120);
nand U3302 (N_3302,N_978,N_1010);
or U3303 (N_3303,N_412,N_508);
xnor U3304 (N_3304,N_1009,N_942);
xnor U3305 (N_3305,N_411,N_961);
or U3306 (N_3306,N_749,N_196);
nand U3307 (N_3307,N_201,N_67);
xor U3308 (N_3308,N_1097,N_745);
and U3309 (N_3309,N_461,N_1282);
and U3310 (N_3310,N_508,N_1491);
nor U3311 (N_3311,N_1889,N_1024);
and U3312 (N_3312,N_1000,N_220);
or U3313 (N_3313,N_1282,N_1781);
nor U3314 (N_3314,N_342,N_194);
nand U3315 (N_3315,N_32,N_175);
nor U3316 (N_3316,N_1703,N_1182);
and U3317 (N_3317,N_1237,N_1150);
and U3318 (N_3318,N_870,N_188);
nor U3319 (N_3319,N_971,N_384);
and U3320 (N_3320,N_1322,N_1645);
nand U3321 (N_3321,N_873,N_138);
xor U3322 (N_3322,N_527,N_1379);
nand U3323 (N_3323,N_685,N_421);
nand U3324 (N_3324,N_757,N_889);
xor U3325 (N_3325,N_1125,N_1084);
and U3326 (N_3326,N_272,N_1979);
nor U3327 (N_3327,N_1562,N_560);
xor U3328 (N_3328,N_651,N_362);
xnor U3329 (N_3329,N_605,N_1676);
or U3330 (N_3330,N_265,N_1414);
nand U3331 (N_3331,N_1565,N_1901);
and U3332 (N_3332,N_171,N_778);
nand U3333 (N_3333,N_815,N_1227);
and U3334 (N_3334,N_1092,N_1862);
xor U3335 (N_3335,N_531,N_732);
nor U3336 (N_3336,N_1976,N_1743);
nor U3337 (N_3337,N_737,N_58);
or U3338 (N_3338,N_1110,N_981);
and U3339 (N_3339,N_1432,N_104);
nand U3340 (N_3340,N_264,N_98);
xor U3341 (N_3341,N_1259,N_1067);
or U3342 (N_3342,N_1942,N_579);
nor U3343 (N_3343,N_1427,N_101);
and U3344 (N_3344,N_1748,N_1897);
xor U3345 (N_3345,N_903,N_1164);
nand U3346 (N_3346,N_814,N_662);
or U3347 (N_3347,N_776,N_1163);
and U3348 (N_3348,N_1014,N_1350);
and U3349 (N_3349,N_1758,N_1144);
and U3350 (N_3350,N_1068,N_583);
nor U3351 (N_3351,N_714,N_821);
nand U3352 (N_3352,N_5,N_1973);
nor U3353 (N_3353,N_939,N_991);
or U3354 (N_3354,N_1412,N_1556);
and U3355 (N_3355,N_1144,N_603);
and U3356 (N_3356,N_1756,N_177);
or U3357 (N_3357,N_822,N_106);
and U3358 (N_3358,N_1892,N_447);
or U3359 (N_3359,N_1306,N_1736);
and U3360 (N_3360,N_1965,N_1449);
and U3361 (N_3361,N_41,N_1123);
nand U3362 (N_3362,N_873,N_550);
xnor U3363 (N_3363,N_1754,N_1907);
or U3364 (N_3364,N_1394,N_69);
and U3365 (N_3365,N_954,N_1524);
or U3366 (N_3366,N_1800,N_1204);
nand U3367 (N_3367,N_1286,N_1712);
nor U3368 (N_3368,N_1774,N_371);
nand U3369 (N_3369,N_1499,N_462);
nand U3370 (N_3370,N_238,N_435);
nand U3371 (N_3371,N_1632,N_1245);
xor U3372 (N_3372,N_1588,N_461);
or U3373 (N_3373,N_1847,N_1454);
or U3374 (N_3374,N_697,N_71);
xnor U3375 (N_3375,N_234,N_538);
nor U3376 (N_3376,N_1651,N_1504);
or U3377 (N_3377,N_615,N_1643);
and U3378 (N_3378,N_1114,N_1552);
nor U3379 (N_3379,N_155,N_165);
and U3380 (N_3380,N_1562,N_1883);
and U3381 (N_3381,N_1821,N_1201);
or U3382 (N_3382,N_851,N_81);
nor U3383 (N_3383,N_1191,N_191);
nor U3384 (N_3384,N_56,N_922);
and U3385 (N_3385,N_741,N_829);
and U3386 (N_3386,N_809,N_703);
xor U3387 (N_3387,N_1628,N_951);
nor U3388 (N_3388,N_99,N_290);
xnor U3389 (N_3389,N_193,N_1298);
nor U3390 (N_3390,N_721,N_1553);
or U3391 (N_3391,N_1152,N_1341);
nand U3392 (N_3392,N_994,N_843);
nand U3393 (N_3393,N_1915,N_1418);
or U3394 (N_3394,N_543,N_796);
and U3395 (N_3395,N_905,N_1938);
or U3396 (N_3396,N_1079,N_953);
and U3397 (N_3397,N_1333,N_188);
nand U3398 (N_3398,N_11,N_1564);
nand U3399 (N_3399,N_168,N_1123);
and U3400 (N_3400,N_155,N_41);
nor U3401 (N_3401,N_1836,N_1024);
xor U3402 (N_3402,N_1885,N_1082);
and U3403 (N_3403,N_1947,N_848);
xnor U3404 (N_3404,N_1591,N_1676);
or U3405 (N_3405,N_1784,N_251);
or U3406 (N_3406,N_1312,N_1664);
nand U3407 (N_3407,N_1563,N_1772);
nor U3408 (N_3408,N_1767,N_1178);
nand U3409 (N_3409,N_1913,N_36);
and U3410 (N_3410,N_1854,N_984);
nor U3411 (N_3411,N_1450,N_633);
nand U3412 (N_3412,N_1259,N_1964);
nor U3413 (N_3413,N_428,N_200);
nor U3414 (N_3414,N_1732,N_736);
nor U3415 (N_3415,N_1936,N_724);
or U3416 (N_3416,N_1062,N_656);
nand U3417 (N_3417,N_86,N_1028);
nand U3418 (N_3418,N_1802,N_1254);
and U3419 (N_3419,N_1033,N_363);
nand U3420 (N_3420,N_50,N_1664);
or U3421 (N_3421,N_1070,N_272);
xor U3422 (N_3422,N_1118,N_1106);
and U3423 (N_3423,N_1929,N_723);
xnor U3424 (N_3424,N_973,N_374);
nor U3425 (N_3425,N_707,N_598);
xnor U3426 (N_3426,N_239,N_1330);
nor U3427 (N_3427,N_380,N_1107);
nand U3428 (N_3428,N_51,N_294);
nor U3429 (N_3429,N_500,N_1494);
or U3430 (N_3430,N_804,N_1558);
nor U3431 (N_3431,N_852,N_356);
nand U3432 (N_3432,N_1078,N_1179);
xnor U3433 (N_3433,N_267,N_665);
nor U3434 (N_3434,N_1295,N_94);
nor U3435 (N_3435,N_1147,N_319);
nand U3436 (N_3436,N_1707,N_476);
nand U3437 (N_3437,N_1134,N_1532);
nor U3438 (N_3438,N_1865,N_680);
or U3439 (N_3439,N_1018,N_933);
xor U3440 (N_3440,N_1875,N_1385);
xor U3441 (N_3441,N_1678,N_641);
or U3442 (N_3442,N_1768,N_295);
nor U3443 (N_3443,N_998,N_43);
or U3444 (N_3444,N_629,N_156);
nor U3445 (N_3445,N_207,N_1080);
and U3446 (N_3446,N_714,N_502);
nand U3447 (N_3447,N_120,N_230);
and U3448 (N_3448,N_1759,N_850);
nand U3449 (N_3449,N_408,N_1779);
or U3450 (N_3450,N_1378,N_1396);
nor U3451 (N_3451,N_1332,N_1317);
nand U3452 (N_3452,N_363,N_245);
nor U3453 (N_3453,N_77,N_404);
and U3454 (N_3454,N_695,N_402);
or U3455 (N_3455,N_538,N_1025);
nand U3456 (N_3456,N_319,N_771);
and U3457 (N_3457,N_612,N_1170);
nor U3458 (N_3458,N_1927,N_1712);
xnor U3459 (N_3459,N_524,N_1739);
nor U3460 (N_3460,N_891,N_1278);
nand U3461 (N_3461,N_1392,N_867);
and U3462 (N_3462,N_734,N_1013);
nand U3463 (N_3463,N_244,N_494);
nand U3464 (N_3464,N_1566,N_282);
nor U3465 (N_3465,N_569,N_1750);
and U3466 (N_3466,N_1515,N_1934);
xor U3467 (N_3467,N_1935,N_216);
or U3468 (N_3468,N_567,N_729);
or U3469 (N_3469,N_519,N_1541);
nor U3470 (N_3470,N_266,N_902);
xor U3471 (N_3471,N_1360,N_181);
nor U3472 (N_3472,N_1913,N_1093);
or U3473 (N_3473,N_432,N_1056);
xor U3474 (N_3474,N_571,N_1475);
nor U3475 (N_3475,N_831,N_1515);
nor U3476 (N_3476,N_517,N_1709);
or U3477 (N_3477,N_1739,N_1037);
and U3478 (N_3478,N_580,N_1189);
nand U3479 (N_3479,N_836,N_1417);
and U3480 (N_3480,N_1672,N_1078);
xnor U3481 (N_3481,N_1520,N_1264);
nor U3482 (N_3482,N_881,N_1261);
nor U3483 (N_3483,N_1698,N_944);
xnor U3484 (N_3484,N_1280,N_1166);
nor U3485 (N_3485,N_1331,N_1908);
nor U3486 (N_3486,N_1048,N_1999);
nand U3487 (N_3487,N_1662,N_1346);
or U3488 (N_3488,N_1890,N_518);
nor U3489 (N_3489,N_1591,N_1558);
or U3490 (N_3490,N_14,N_834);
nand U3491 (N_3491,N_281,N_976);
and U3492 (N_3492,N_1955,N_805);
xor U3493 (N_3493,N_968,N_1846);
and U3494 (N_3494,N_1897,N_1399);
and U3495 (N_3495,N_1618,N_1573);
nor U3496 (N_3496,N_338,N_659);
xnor U3497 (N_3497,N_1827,N_1479);
nand U3498 (N_3498,N_1669,N_902);
or U3499 (N_3499,N_1587,N_385);
and U3500 (N_3500,N_1052,N_1732);
xor U3501 (N_3501,N_679,N_370);
and U3502 (N_3502,N_1723,N_1072);
nand U3503 (N_3503,N_1408,N_219);
nand U3504 (N_3504,N_505,N_975);
and U3505 (N_3505,N_434,N_1642);
or U3506 (N_3506,N_459,N_418);
and U3507 (N_3507,N_1893,N_117);
nor U3508 (N_3508,N_465,N_1214);
nand U3509 (N_3509,N_1427,N_1792);
nor U3510 (N_3510,N_1798,N_1365);
nand U3511 (N_3511,N_267,N_78);
or U3512 (N_3512,N_1568,N_1230);
or U3513 (N_3513,N_7,N_1707);
and U3514 (N_3514,N_1070,N_761);
nor U3515 (N_3515,N_292,N_1842);
or U3516 (N_3516,N_464,N_1486);
or U3517 (N_3517,N_1049,N_1449);
nor U3518 (N_3518,N_242,N_1957);
and U3519 (N_3519,N_1929,N_1521);
nor U3520 (N_3520,N_1314,N_433);
nor U3521 (N_3521,N_1742,N_1227);
and U3522 (N_3522,N_1232,N_1922);
nand U3523 (N_3523,N_1482,N_1131);
nor U3524 (N_3524,N_1998,N_423);
xor U3525 (N_3525,N_1058,N_1350);
xnor U3526 (N_3526,N_1192,N_1809);
and U3527 (N_3527,N_909,N_925);
nor U3528 (N_3528,N_203,N_1109);
nor U3529 (N_3529,N_157,N_1002);
nand U3530 (N_3530,N_1303,N_1671);
nand U3531 (N_3531,N_1282,N_100);
or U3532 (N_3532,N_1876,N_1009);
nor U3533 (N_3533,N_680,N_1133);
xor U3534 (N_3534,N_113,N_1554);
or U3535 (N_3535,N_977,N_989);
nand U3536 (N_3536,N_1146,N_954);
nand U3537 (N_3537,N_606,N_561);
nand U3538 (N_3538,N_370,N_378);
or U3539 (N_3539,N_676,N_436);
nand U3540 (N_3540,N_1387,N_1344);
xor U3541 (N_3541,N_1669,N_453);
nor U3542 (N_3542,N_1777,N_939);
and U3543 (N_3543,N_294,N_687);
nand U3544 (N_3544,N_903,N_208);
nand U3545 (N_3545,N_1873,N_1809);
or U3546 (N_3546,N_1447,N_91);
nand U3547 (N_3547,N_964,N_1630);
or U3548 (N_3548,N_1216,N_67);
xor U3549 (N_3549,N_821,N_961);
nand U3550 (N_3550,N_1661,N_1301);
and U3551 (N_3551,N_732,N_580);
nand U3552 (N_3552,N_297,N_500);
nor U3553 (N_3553,N_1633,N_336);
and U3554 (N_3554,N_261,N_1834);
and U3555 (N_3555,N_395,N_1536);
xnor U3556 (N_3556,N_1010,N_1991);
or U3557 (N_3557,N_1077,N_708);
nor U3558 (N_3558,N_458,N_1744);
nand U3559 (N_3559,N_1959,N_659);
nor U3560 (N_3560,N_381,N_1244);
nor U3561 (N_3561,N_1813,N_811);
nand U3562 (N_3562,N_1534,N_1217);
xor U3563 (N_3563,N_184,N_995);
nor U3564 (N_3564,N_576,N_1678);
xnor U3565 (N_3565,N_1642,N_695);
nor U3566 (N_3566,N_545,N_1690);
or U3567 (N_3567,N_1881,N_1771);
nor U3568 (N_3568,N_76,N_1383);
or U3569 (N_3569,N_1161,N_768);
nor U3570 (N_3570,N_970,N_1197);
or U3571 (N_3571,N_1231,N_985);
or U3572 (N_3572,N_1972,N_127);
nand U3573 (N_3573,N_1199,N_538);
and U3574 (N_3574,N_1918,N_130);
nand U3575 (N_3575,N_1550,N_946);
or U3576 (N_3576,N_1094,N_682);
or U3577 (N_3577,N_761,N_1703);
nand U3578 (N_3578,N_663,N_1791);
or U3579 (N_3579,N_417,N_552);
nor U3580 (N_3580,N_1256,N_241);
or U3581 (N_3581,N_264,N_998);
and U3582 (N_3582,N_1929,N_288);
or U3583 (N_3583,N_543,N_1904);
or U3584 (N_3584,N_1034,N_338);
nand U3585 (N_3585,N_1620,N_1608);
nand U3586 (N_3586,N_1577,N_1639);
nand U3587 (N_3587,N_495,N_1210);
and U3588 (N_3588,N_1761,N_1963);
xnor U3589 (N_3589,N_795,N_1570);
or U3590 (N_3590,N_521,N_417);
xor U3591 (N_3591,N_1870,N_889);
and U3592 (N_3592,N_1499,N_194);
nor U3593 (N_3593,N_1112,N_1240);
or U3594 (N_3594,N_608,N_746);
xor U3595 (N_3595,N_891,N_1858);
and U3596 (N_3596,N_239,N_1322);
nor U3597 (N_3597,N_420,N_240);
xor U3598 (N_3598,N_702,N_1884);
nand U3599 (N_3599,N_380,N_1633);
nand U3600 (N_3600,N_353,N_1580);
xor U3601 (N_3601,N_601,N_1296);
or U3602 (N_3602,N_596,N_1763);
nor U3603 (N_3603,N_80,N_696);
nor U3604 (N_3604,N_1970,N_550);
nor U3605 (N_3605,N_637,N_892);
or U3606 (N_3606,N_279,N_653);
nor U3607 (N_3607,N_424,N_26);
and U3608 (N_3608,N_1521,N_1599);
xnor U3609 (N_3609,N_305,N_34);
and U3610 (N_3610,N_118,N_613);
and U3611 (N_3611,N_404,N_1497);
nor U3612 (N_3612,N_366,N_793);
nand U3613 (N_3613,N_335,N_1374);
xor U3614 (N_3614,N_1932,N_1203);
and U3615 (N_3615,N_1689,N_627);
or U3616 (N_3616,N_183,N_672);
nand U3617 (N_3617,N_1665,N_1501);
or U3618 (N_3618,N_1127,N_1820);
nand U3619 (N_3619,N_721,N_1830);
xnor U3620 (N_3620,N_1241,N_1603);
and U3621 (N_3621,N_458,N_3);
nand U3622 (N_3622,N_28,N_1438);
nor U3623 (N_3623,N_1816,N_1703);
xnor U3624 (N_3624,N_1974,N_1869);
and U3625 (N_3625,N_843,N_292);
and U3626 (N_3626,N_1019,N_1781);
nor U3627 (N_3627,N_184,N_1597);
and U3628 (N_3628,N_434,N_1748);
nor U3629 (N_3629,N_1628,N_10);
nand U3630 (N_3630,N_680,N_125);
xor U3631 (N_3631,N_801,N_1241);
or U3632 (N_3632,N_840,N_492);
or U3633 (N_3633,N_516,N_1124);
or U3634 (N_3634,N_208,N_652);
nor U3635 (N_3635,N_1833,N_829);
and U3636 (N_3636,N_1583,N_1090);
nor U3637 (N_3637,N_674,N_1798);
or U3638 (N_3638,N_1288,N_1680);
or U3639 (N_3639,N_147,N_38);
nand U3640 (N_3640,N_480,N_1979);
and U3641 (N_3641,N_511,N_784);
xnor U3642 (N_3642,N_1849,N_260);
nand U3643 (N_3643,N_424,N_1707);
or U3644 (N_3644,N_1032,N_19);
xor U3645 (N_3645,N_848,N_1461);
or U3646 (N_3646,N_176,N_1009);
nand U3647 (N_3647,N_279,N_1845);
xor U3648 (N_3648,N_1156,N_1470);
xnor U3649 (N_3649,N_857,N_1401);
or U3650 (N_3650,N_1110,N_741);
or U3651 (N_3651,N_1038,N_998);
nand U3652 (N_3652,N_1901,N_1550);
xor U3653 (N_3653,N_726,N_1404);
and U3654 (N_3654,N_1925,N_756);
xor U3655 (N_3655,N_57,N_140);
xor U3656 (N_3656,N_1803,N_1364);
xnor U3657 (N_3657,N_1699,N_1071);
and U3658 (N_3658,N_225,N_970);
or U3659 (N_3659,N_913,N_1472);
or U3660 (N_3660,N_668,N_1339);
or U3661 (N_3661,N_1627,N_666);
nor U3662 (N_3662,N_1897,N_843);
nor U3663 (N_3663,N_1746,N_1028);
or U3664 (N_3664,N_1077,N_934);
nor U3665 (N_3665,N_797,N_1759);
nor U3666 (N_3666,N_1938,N_1403);
or U3667 (N_3667,N_750,N_845);
or U3668 (N_3668,N_1865,N_705);
or U3669 (N_3669,N_976,N_1812);
or U3670 (N_3670,N_746,N_1699);
and U3671 (N_3671,N_1810,N_142);
and U3672 (N_3672,N_129,N_1433);
nand U3673 (N_3673,N_491,N_222);
or U3674 (N_3674,N_1270,N_1532);
xor U3675 (N_3675,N_945,N_1471);
nor U3676 (N_3676,N_79,N_1462);
nand U3677 (N_3677,N_1718,N_1110);
nor U3678 (N_3678,N_1985,N_1395);
nand U3679 (N_3679,N_1326,N_344);
or U3680 (N_3680,N_339,N_1056);
nor U3681 (N_3681,N_627,N_1316);
nand U3682 (N_3682,N_1656,N_803);
or U3683 (N_3683,N_498,N_117);
and U3684 (N_3684,N_1542,N_1298);
xor U3685 (N_3685,N_242,N_156);
and U3686 (N_3686,N_711,N_203);
nand U3687 (N_3687,N_1124,N_144);
and U3688 (N_3688,N_543,N_730);
or U3689 (N_3689,N_909,N_572);
or U3690 (N_3690,N_1260,N_511);
and U3691 (N_3691,N_1239,N_791);
or U3692 (N_3692,N_650,N_1478);
xnor U3693 (N_3693,N_1271,N_854);
nor U3694 (N_3694,N_1024,N_1070);
and U3695 (N_3695,N_339,N_921);
and U3696 (N_3696,N_653,N_1044);
nand U3697 (N_3697,N_195,N_1960);
or U3698 (N_3698,N_384,N_59);
nor U3699 (N_3699,N_1194,N_1190);
or U3700 (N_3700,N_439,N_1240);
nand U3701 (N_3701,N_436,N_1170);
xor U3702 (N_3702,N_547,N_1213);
or U3703 (N_3703,N_1611,N_15);
and U3704 (N_3704,N_967,N_1854);
xor U3705 (N_3705,N_1144,N_682);
nand U3706 (N_3706,N_698,N_642);
xor U3707 (N_3707,N_456,N_706);
xor U3708 (N_3708,N_574,N_1133);
nand U3709 (N_3709,N_760,N_1751);
or U3710 (N_3710,N_1710,N_1684);
xor U3711 (N_3711,N_1719,N_848);
nor U3712 (N_3712,N_1448,N_506);
and U3713 (N_3713,N_1234,N_412);
or U3714 (N_3714,N_1115,N_792);
and U3715 (N_3715,N_1372,N_1972);
nor U3716 (N_3716,N_39,N_759);
or U3717 (N_3717,N_879,N_495);
or U3718 (N_3718,N_177,N_439);
or U3719 (N_3719,N_282,N_1831);
or U3720 (N_3720,N_1913,N_1375);
or U3721 (N_3721,N_136,N_1643);
xor U3722 (N_3722,N_193,N_388);
nor U3723 (N_3723,N_1278,N_1738);
or U3724 (N_3724,N_460,N_703);
or U3725 (N_3725,N_28,N_1909);
or U3726 (N_3726,N_996,N_1779);
or U3727 (N_3727,N_1824,N_1490);
and U3728 (N_3728,N_1495,N_1039);
nor U3729 (N_3729,N_224,N_780);
nand U3730 (N_3730,N_834,N_222);
nor U3731 (N_3731,N_1704,N_508);
xnor U3732 (N_3732,N_433,N_418);
and U3733 (N_3733,N_1112,N_1146);
or U3734 (N_3734,N_800,N_1125);
xor U3735 (N_3735,N_1083,N_90);
nor U3736 (N_3736,N_1686,N_17);
and U3737 (N_3737,N_843,N_1665);
nand U3738 (N_3738,N_1479,N_414);
xnor U3739 (N_3739,N_1790,N_11);
or U3740 (N_3740,N_916,N_927);
and U3741 (N_3741,N_584,N_418);
and U3742 (N_3742,N_1121,N_1965);
and U3743 (N_3743,N_1979,N_1448);
nor U3744 (N_3744,N_491,N_1357);
xnor U3745 (N_3745,N_273,N_1832);
nand U3746 (N_3746,N_599,N_649);
xnor U3747 (N_3747,N_1743,N_1465);
and U3748 (N_3748,N_1960,N_876);
nor U3749 (N_3749,N_448,N_1139);
nand U3750 (N_3750,N_1908,N_1191);
nor U3751 (N_3751,N_136,N_845);
and U3752 (N_3752,N_1592,N_212);
nand U3753 (N_3753,N_84,N_957);
nand U3754 (N_3754,N_320,N_471);
xnor U3755 (N_3755,N_671,N_1355);
nor U3756 (N_3756,N_440,N_1826);
xnor U3757 (N_3757,N_687,N_637);
nand U3758 (N_3758,N_1712,N_915);
or U3759 (N_3759,N_1339,N_1551);
or U3760 (N_3760,N_438,N_1520);
and U3761 (N_3761,N_554,N_889);
and U3762 (N_3762,N_1899,N_1208);
xnor U3763 (N_3763,N_751,N_804);
nand U3764 (N_3764,N_1550,N_1338);
nand U3765 (N_3765,N_1401,N_1854);
xnor U3766 (N_3766,N_1656,N_1688);
and U3767 (N_3767,N_42,N_1013);
and U3768 (N_3768,N_1668,N_861);
nand U3769 (N_3769,N_1386,N_1635);
or U3770 (N_3770,N_940,N_338);
nor U3771 (N_3771,N_1560,N_1723);
nor U3772 (N_3772,N_1007,N_972);
nand U3773 (N_3773,N_1519,N_140);
and U3774 (N_3774,N_468,N_214);
xnor U3775 (N_3775,N_880,N_1898);
or U3776 (N_3776,N_1945,N_1174);
and U3777 (N_3777,N_1583,N_1232);
or U3778 (N_3778,N_872,N_1186);
nand U3779 (N_3779,N_1736,N_1033);
or U3780 (N_3780,N_1534,N_1222);
xnor U3781 (N_3781,N_465,N_1653);
nor U3782 (N_3782,N_1623,N_309);
xor U3783 (N_3783,N_1160,N_961);
or U3784 (N_3784,N_941,N_722);
nand U3785 (N_3785,N_205,N_1719);
or U3786 (N_3786,N_669,N_1309);
and U3787 (N_3787,N_198,N_680);
nor U3788 (N_3788,N_1764,N_1938);
or U3789 (N_3789,N_992,N_723);
xnor U3790 (N_3790,N_136,N_740);
nor U3791 (N_3791,N_1536,N_501);
nand U3792 (N_3792,N_1232,N_408);
nand U3793 (N_3793,N_1158,N_405);
nand U3794 (N_3794,N_1832,N_1596);
nor U3795 (N_3795,N_590,N_1278);
and U3796 (N_3796,N_509,N_1236);
xor U3797 (N_3797,N_482,N_525);
nand U3798 (N_3798,N_664,N_1147);
or U3799 (N_3799,N_1856,N_1133);
xnor U3800 (N_3800,N_1539,N_1428);
xnor U3801 (N_3801,N_156,N_1945);
xor U3802 (N_3802,N_528,N_389);
nand U3803 (N_3803,N_378,N_972);
nand U3804 (N_3804,N_1450,N_580);
or U3805 (N_3805,N_494,N_125);
and U3806 (N_3806,N_791,N_1461);
nand U3807 (N_3807,N_311,N_1557);
nand U3808 (N_3808,N_1722,N_1960);
nand U3809 (N_3809,N_1203,N_359);
nor U3810 (N_3810,N_79,N_1272);
xor U3811 (N_3811,N_1098,N_648);
xnor U3812 (N_3812,N_695,N_1062);
nor U3813 (N_3813,N_1944,N_1922);
nor U3814 (N_3814,N_1881,N_1563);
nand U3815 (N_3815,N_138,N_1624);
nand U3816 (N_3816,N_722,N_1986);
or U3817 (N_3817,N_452,N_1799);
nor U3818 (N_3818,N_592,N_116);
nand U3819 (N_3819,N_184,N_1900);
xor U3820 (N_3820,N_1946,N_889);
and U3821 (N_3821,N_56,N_1311);
nor U3822 (N_3822,N_332,N_17);
xor U3823 (N_3823,N_590,N_1081);
nor U3824 (N_3824,N_1869,N_482);
or U3825 (N_3825,N_472,N_1504);
xnor U3826 (N_3826,N_698,N_803);
nor U3827 (N_3827,N_1738,N_1564);
and U3828 (N_3828,N_1261,N_278);
nor U3829 (N_3829,N_1245,N_31);
xnor U3830 (N_3830,N_1727,N_1236);
or U3831 (N_3831,N_1794,N_1835);
and U3832 (N_3832,N_488,N_308);
or U3833 (N_3833,N_1916,N_279);
xnor U3834 (N_3834,N_648,N_1965);
xnor U3835 (N_3835,N_1916,N_1173);
or U3836 (N_3836,N_185,N_955);
xnor U3837 (N_3837,N_1921,N_764);
and U3838 (N_3838,N_1196,N_707);
xnor U3839 (N_3839,N_850,N_685);
nand U3840 (N_3840,N_242,N_777);
and U3841 (N_3841,N_687,N_623);
nor U3842 (N_3842,N_1398,N_727);
or U3843 (N_3843,N_12,N_1223);
nor U3844 (N_3844,N_661,N_1536);
or U3845 (N_3845,N_1975,N_873);
xnor U3846 (N_3846,N_797,N_1702);
or U3847 (N_3847,N_1317,N_1012);
or U3848 (N_3848,N_1056,N_402);
nor U3849 (N_3849,N_266,N_1933);
xor U3850 (N_3850,N_614,N_1318);
nor U3851 (N_3851,N_202,N_681);
or U3852 (N_3852,N_1052,N_437);
and U3853 (N_3853,N_1879,N_176);
nand U3854 (N_3854,N_1160,N_1812);
and U3855 (N_3855,N_237,N_979);
xor U3856 (N_3856,N_1263,N_853);
and U3857 (N_3857,N_1955,N_204);
nand U3858 (N_3858,N_1032,N_768);
xor U3859 (N_3859,N_1943,N_1410);
and U3860 (N_3860,N_100,N_767);
nor U3861 (N_3861,N_113,N_1150);
and U3862 (N_3862,N_334,N_866);
xnor U3863 (N_3863,N_1397,N_990);
xor U3864 (N_3864,N_293,N_255);
xnor U3865 (N_3865,N_57,N_1063);
nand U3866 (N_3866,N_1740,N_319);
nand U3867 (N_3867,N_268,N_1395);
xnor U3868 (N_3868,N_441,N_587);
nand U3869 (N_3869,N_221,N_57);
nand U3870 (N_3870,N_1356,N_1284);
xor U3871 (N_3871,N_1121,N_781);
nand U3872 (N_3872,N_208,N_668);
nor U3873 (N_3873,N_1476,N_1024);
nand U3874 (N_3874,N_1571,N_351);
nand U3875 (N_3875,N_1875,N_350);
or U3876 (N_3876,N_597,N_1186);
and U3877 (N_3877,N_202,N_242);
xor U3878 (N_3878,N_359,N_293);
xnor U3879 (N_3879,N_108,N_1285);
or U3880 (N_3880,N_56,N_1684);
nor U3881 (N_3881,N_1850,N_78);
or U3882 (N_3882,N_931,N_1024);
nand U3883 (N_3883,N_923,N_1980);
nor U3884 (N_3884,N_36,N_811);
xnor U3885 (N_3885,N_134,N_1168);
nand U3886 (N_3886,N_556,N_1664);
and U3887 (N_3887,N_515,N_1069);
and U3888 (N_3888,N_437,N_694);
xor U3889 (N_3889,N_1902,N_847);
or U3890 (N_3890,N_1719,N_362);
and U3891 (N_3891,N_1677,N_1546);
or U3892 (N_3892,N_1069,N_203);
and U3893 (N_3893,N_1093,N_600);
nor U3894 (N_3894,N_820,N_1930);
xor U3895 (N_3895,N_1263,N_1190);
xnor U3896 (N_3896,N_461,N_1291);
nor U3897 (N_3897,N_926,N_866);
xnor U3898 (N_3898,N_643,N_1144);
nand U3899 (N_3899,N_138,N_1532);
xnor U3900 (N_3900,N_1391,N_1513);
or U3901 (N_3901,N_930,N_1765);
or U3902 (N_3902,N_417,N_1133);
xor U3903 (N_3903,N_764,N_78);
and U3904 (N_3904,N_886,N_1766);
or U3905 (N_3905,N_868,N_1457);
or U3906 (N_3906,N_1632,N_1298);
nor U3907 (N_3907,N_229,N_884);
nor U3908 (N_3908,N_667,N_1252);
nor U3909 (N_3909,N_225,N_1890);
and U3910 (N_3910,N_712,N_254);
xnor U3911 (N_3911,N_151,N_1439);
and U3912 (N_3912,N_765,N_729);
xnor U3913 (N_3913,N_1775,N_1464);
xnor U3914 (N_3914,N_239,N_1050);
or U3915 (N_3915,N_1887,N_1272);
nor U3916 (N_3916,N_496,N_1);
nand U3917 (N_3917,N_865,N_345);
nor U3918 (N_3918,N_769,N_1571);
and U3919 (N_3919,N_1091,N_613);
nand U3920 (N_3920,N_1448,N_898);
or U3921 (N_3921,N_1118,N_70);
nor U3922 (N_3922,N_988,N_638);
xnor U3923 (N_3923,N_621,N_958);
and U3924 (N_3924,N_1081,N_1579);
xor U3925 (N_3925,N_989,N_552);
xnor U3926 (N_3926,N_1903,N_15);
or U3927 (N_3927,N_356,N_1023);
nand U3928 (N_3928,N_84,N_237);
nor U3929 (N_3929,N_1259,N_1077);
nor U3930 (N_3930,N_525,N_1295);
and U3931 (N_3931,N_1328,N_1921);
or U3932 (N_3932,N_1442,N_1418);
xnor U3933 (N_3933,N_1775,N_388);
nand U3934 (N_3934,N_734,N_781);
nand U3935 (N_3935,N_1273,N_903);
nor U3936 (N_3936,N_315,N_787);
xor U3937 (N_3937,N_98,N_296);
nand U3938 (N_3938,N_1836,N_1236);
xor U3939 (N_3939,N_6,N_1143);
nand U3940 (N_3940,N_170,N_1655);
xnor U3941 (N_3941,N_319,N_1661);
xnor U3942 (N_3942,N_1072,N_496);
or U3943 (N_3943,N_1702,N_1682);
nand U3944 (N_3944,N_1928,N_821);
or U3945 (N_3945,N_1655,N_598);
or U3946 (N_3946,N_1316,N_1549);
or U3947 (N_3947,N_38,N_125);
nand U3948 (N_3948,N_1404,N_1255);
xnor U3949 (N_3949,N_872,N_1446);
nor U3950 (N_3950,N_119,N_1812);
nor U3951 (N_3951,N_1059,N_1862);
or U3952 (N_3952,N_1579,N_1490);
nor U3953 (N_3953,N_834,N_422);
and U3954 (N_3954,N_818,N_350);
nor U3955 (N_3955,N_1665,N_1659);
or U3956 (N_3956,N_771,N_309);
or U3957 (N_3957,N_1548,N_1001);
or U3958 (N_3958,N_1730,N_1192);
nand U3959 (N_3959,N_1612,N_943);
nand U3960 (N_3960,N_517,N_1252);
or U3961 (N_3961,N_1256,N_15);
nor U3962 (N_3962,N_943,N_1332);
nor U3963 (N_3963,N_570,N_1493);
nand U3964 (N_3964,N_1264,N_48);
nand U3965 (N_3965,N_1327,N_1388);
and U3966 (N_3966,N_382,N_981);
nand U3967 (N_3967,N_415,N_194);
nand U3968 (N_3968,N_1250,N_904);
nor U3969 (N_3969,N_698,N_450);
nand U3970 (N_3970,N_802,N_1401);
nor U3971 (N_3971,N_110,N_142);
or U3972 (N_3972,N_217,N_997);
and U3973 (N_3973,N_1448,N_1982);
or U3974 (N_3974,N_486,N_532);
and U3975 (N_3975,N_1604,N_1112);
or U3976 (N_3976,N_1205,N_1054);
and U3977 (N_3977,N_1784,N_1939);
or U3978 (N_3978,N_1221,N_1863);
or U3979 (N_3979,N_982,N_410);
nand U3980 (N_3980,N_241,N_295);
nand U3981 (N_3981,N_1615,N_396);
xnor U3982 (N_3982,N_434,N_1771);
xnor U3983 (N_3983,N_363,N_942);
nor U3984 (N_3984,N_171,N_1493);
nand U3985 (N_3985,N_1024,N_612);
or U3986 (N_3986,N_782,N_23);
and U3987 (N_3987,N_1928,N_174);
xor U3988 (N_3988,N_218,N_1765);
xor U3989 (N_3989,N_1014,N_982);
and U3990 (N_3990,N_509,N_5);
or U3991 (N_3991,N_1750,N_396);
or U3992 (N_3992,N_37,N_700);
or U3993 (N_3993,N_58,N_704);
xor U3994 (N_3994,N_758,N_655);
nor U3995 (N_3995,N_1094,N_503);
and U3996 (N_3996,N_1601,N_685);
or U3997 (N_3997,N_928,N_435);
or U3998 (N_3998,N_1780,N_1926);
xnor U3999 (N_3999,N_896,N_570);
nand U4000 (N_4000,N_3780,N_3201);
and U4001 (N_4001,N_2997,N_2785);
or U4002 (N_4002,N_3659,N_2898);
xnor U4003 (N_4003,N_3617,N_2244);
and U4004 (N_4004,N_2152,N_2350);
or U4005 (N_4005,N_3606,N_3031);
and U4006 (N_4006,N_3507,N_2086);
nand U4007 (N_4007,N_3670,N_2605);
or U4008 (N_4008,N_3210,N_3766);
or U4009 (N_4009,N_2031,N_2459);
xnor U4010 (N_4010,N_2636,N_3563);
and U4011 (N_4011,N_3550,N_2767);
or U4012 (N_4012,N_2932,N_2071);
nor U4013 (N_4013,N_2540,N_3239);
nand U4014 (N_4014,N_2133,N_3404);
and U4015 (N_4015,N_3386,N_3097);
xor U4016 (N_4016,N_3783,N_3789);
nand U4017 (N_4017,N_2589,N_3823);
xor U4018 (N_4018,N_2649,N_3166);
nor U4019 (N_4019,N_3523,N_3229);
xor U4020 (N_4020,N_2131,N_2922);
and U4021 (N_4021,N_2120,N_2562);
xnor U4022 (N_4022,N_3358,N_3080);
xnor U4023 (N_4023,N_3407,N_2948);
nand U4024 (N_4024,N_2382,N_2514);
nor U4025 (N_4025,N_3504,N_2571);
and U4026 (N_4026,N_3827,N_2205);
and U4027 (N_4027,N_2675,N_2563);
or U4028 (N_4028,N_3989,N_3534);
nand U4029 (N_4029,N_2447,N_2134);
and U4030 (N_4030,N_3213,N_2918);
xnor U4031 (N_4031,N_3866,N_2236);
and U4032 (N_4032,N_2537,N_2189);
nand U4033 (N_4033,N_3921,N_2822);
or U4034 (N_4034,N_3824,N_3944);
or U4035 (N_4035,N_3014,N_2465);
or U4036 (N_4036,N_3748,N_3499);
nand U4037 (N_4037,N_2479,N_3214);
nor U4038 (N_4038,N_2863,N_2288);
nor U4039 (N_4039,N_2983,N_3400);
xnor U4040 (N_4040,N_2678,N_3599);
and U4041 (N_4041,N_3368,N_3555);
and U4042 (N_4042,N_3657,N_2659);
or U4043 (N_4043,N_3806,N_2130);
nand U4044 (N_4044,N_3947,N_3770);
xor U4045 (N_4045,N_2566,N_2705);
nand U4046 (N_4046,N_2125,N_3942);
xnor U4047 (N_4047,N_3757,N_2044);
or U4048 (N_4048,N_3234,N_2346);
nand U4049 (N_4049,N_2101,N_3767);
or U4050 (N_4050,N_3605,N_3483);
or U4051 (N_4051,N_2226,N_3840);
xnor U4052 (N_4052,N_2425,N_2388);
xor U4053 (N_4053,N_2640,N_2957);
nand U4054 (N_4054,N_3724,N_3717);
or U4055 (N_4055,N_3737,N_2683);
nand U4056 (N_4056,N_3881,N_2489);
and U4057 (N_4057,N_2924,N_2423);
xnor U4058 (N_4058,N_3895,N_2845);
and U4059 (N_4059,N_2088,N_3072);
nand U4060 (N_4060,N_3976,N_2457);
nand U4061 (N_4061,N_2169,N_2439);
nor U4062 (N_4062,N_2452,N_3283);
and U4063 (N_4063,N_2664,N_3109);
or U4064 (N_4064,N_3567,N_2450);
and U4065 (N_4065,N_2242,N_2254);
and U4066 (N_4066,N_2157,N_2217);
and U4067 (N_4067,N_3739,N_3776);
and U4068 (N_4068,N_2156,N_3545);
nand U4069 (N_4069,N_2124,N_3718);
or U4070 (N_4070,N_3398,N_2621);
xnor U4071 (N_4071,N_3183,N_3394);
nand U4072 (N_4072,N_2357,N_2819);
or U4073 (N_4073,N_3200,N_3842);
xor U4074 (N_4074,N_3829,N_2099);
and U4075 (N_4075,N_2413,N_2897);
nand U4076 (N_4076,N_3726,N_2697);
nand U4077 (N_4077,N_2497,N_3003);
and U4078 (N_4078,N_3493,N_2522);
nor U4079 (N_4079,N_3067,N_2876);
and U4080 (N_4080,N_2788,N_3702);
nand U4081 (N_4081,N_3729,N_2691);
or U4082 (N_4082,N_2877,N_3278);
and U4083 (N_4083,N_3310,N_2693);
or U4084 (N_4084,N_3867,N_2494);
nand U4085 (N_4085,N_2180,N_2590);
nand U4086 (N_4086,N_2394,N_2348);
xnor U4087 (N_4087,N_2679,N_2549);
nor U4088 (N_4088,N_2557,N_2478);
nor U4089 (N_4089,N_3551,N_3952);
or U4090 (N_4090,N_3350,N_3987);
or U4091 (N_4091,N_2037,N_2023);
xor U4092 (N_4092,N_2849,N_2929);
nand U4093 (N_4093,N_3361,N_3502);
and U4094 (N_4094,N_3178,N_2915);
nor U4095 (N_4095,N_2201,N_3308);
and U4096 (N_4096,N_3962,N_2475);
nand U4097 (N_4097,N_3807,N_2094);
or U4098 (N_4098,N_3295,N_3765);
nor U4099 (N_4099,N_3447,N_2651);
and U4100 (N_4100,N_2505,N_3208);
xnor U4101 (N_4101,N_2466,N_3021);
or U4102 (N_4102,N_3011,N_3956);
xor U4103 (N_4103,N_2002,N_2546);
or U4104 (N_4104,N_3859,N_3552);
and U4105 (N_4105,N_2183,N_2091);
or U4106 (N_4106,N_2230,N_3120);
and U4107 (N_4107,N_2374,N_3532);
or U4108 (N_4108,N_2424,N_3167);
nor U4109 (N_4109,N_3870,N_3675);
nor U4110 (N_4110,N_2336,N_3144);
and U4111 (N_4111,N_3768,N_3988);
or U4112 (N_4112,N_3289,N_2267);
and U4113 (N_4113,N_2892,N_3536);
or U4114 (N_4114,N_2429,N_3917);
nor U4115 (N_4115,N_2868,N_3663);
nor U4116 (N_4116,N_2949,N_2754);
or U4117 (N_4117,N_2012,N_3096);
or U4118 (N_4118,N_2026,N_2438);
and U4119 (N_4119,N_2076,N_3918);
and U4120 (N_4120,N_3916,N_2358);
xnor U4121 (N_4121,N_2378,N_2603);
and U4122 (N_4122,N_2387,N_3479);
and U4123 (N_4123,N_2004,N_3320);
xor U4124 (N_4124,N_2033,N_3754);
or U4125 (N_4125,N_3123,N_2432);
nor U4126 (N_4126,N_3225,N_3570);
xor U4127 (N_4127,N_2453,N_3247);
xor U4128 (N_4128,N_3713,N_2105);
xnor U4129 (N_4129,N_2900,N_2646);
nand U4130 (N_4130,N_3875,N_2532);
or U4131 (N_4131,N_2058,N_2444);
xnor U4132 (N_4132,N_2030,N_2816);
nor U4133 (N_4133,N_3590,N_2882);
or U4134 (N_4134,N_3264,N_2419);
xnor U4135 (N_4135,N_2815,N_3487);
xnor U4136 (N_4136,N_2729,N_3685);
or U4137 (N_4137,N_2096,N_3002);
nor U4138 (N_4138,N_3804,N_2635);
xor U4139 (N_4139,N_2895,N_2339);
xor U4140 (N_4140,N_2027,N_2492);
nor U4141 (N_4141,N_2696,N_3782);
nor U4142 (N_4142,N_3161,N_3470);
xnor U4143 (N_4143,N_3743,N_2663);
xnor U4144 (N_4144,N_3529,N_2331);
xor U4145 (N_4145,N_3110,N_3967);
and U4146 (N_4146,N_3949,N_2270);
nor U4147 (N_4147,N_2263,N_2858);
nand U4148 (N_4148,N_2264,N_2360);
and U4149 (N_4149,N_2885,N_2430);
or U4150 (N_4150,N_3970,N_2786);
xor U4151 (N_4151,N_3336,N_2276);
nor U4152 (N_4152,N_3325,N_3613);
nand U4153 (N_4153,N_3707,N_2446);
nor U4154 (N_4154,N_3747,N_2912);
and U4155 (N_4155,N_2403,N_3077);
nand U4156 (N_4156,N_2657,N_3050);
and U4157 (N_4157,N_2289,N_3338);
and U4158 (N_4158,N_3858,N_2437);
and U4159 (N_4159,N_3353,N_2689);
nor U4160 (N_4160,N_3139,N_2581);
nor U4161 (N_4161,N_2383,N_3423);
or U4162 (N_4162,N_3288,N_3862);
nand U4163 (N_4163,N_3700,N_2483);
or U4164 (N_4164,N_3664,N_3694);
xor U4165 (N_4165,N_3222,N_2593);
or U4166 (N_4166,N_3683,N_3460);
nand U4167 (N_4167,N_2999,N_2108);
nand U4168 (N_4168,N_2735,N_2140);
or U4169 (N_4169,N_2191,N_3083);
nor U4170 (N_4170,N_2409,N_2694);
nor U4171 (N_4171,N_3844,N_2499);
or U4172 (N_4172,N_3039,N_3048);
nand U4173 (N_4173,N_2825,N_3484);
xor U4174 (N_4174,N_3143,N_3367);
xnor U4175 (N_4175,N_3373,N_3272);
nand U4176 (N_4176,N_2846,N_3038);
or U4177 (N_4177,N_2513,N_2698);
xor U4178 (N_4178,N_2523,N_2370);
nand U4179 (N_4179,N_3170,N_3828);
nor U4180 (N_4180,N_2399,N_2606);
nor U4181 (N_4181,N_2928,N_2768);
nor U4182 (N_4182,N_3156,N_3596);
or U4183 (N_4183,N_3131,N_2787);
nand U4184 (N_4184,N_3565,N_3466);
nor U4185 (N_4185,N_3934,N_2995);
or U4186 (N_4186,N_2176,N_3377);
and U4187 (N_4187,N_3327,N_2725);
xor U4188 (N_4188,N_2468,N_3094);
nor U4189 (N_4189,N_2335,N_3731);
nand U4190 (N_4190,N_3207,N_2973);
nand U4191 (N_4191,N_3465,N_3124);
nand U4192 (N_4192,N_3496,N_2185);
or U4193 (N_4193,N_3779,N_2077);
nand U4194 (N_4194,N_2944,N_3195);
and U4195 (N_4195,N_3773,N_2167);
or U4196 (N_4196,N_2962,N_3910);
or U4197 (N_4197,N_3158,N_3518);
and U4198 (N_4198,N_2261,N_2200);
or U4199 (N_4199,N_3929,N_3007);
xnor U4200 (N_4200,N_3191,N_3142);
nor U4201 (N_4201,N_3845,N_3841);
and U4202 (N_4202,N_3175,N_3809);
xor U4203 (N_4203,N_2884,N_2552);
or U4204 (N_4204,N_3643,N_2558);
nor U4205 (N_4205,N_2195,N_3808);
nand U4206 (N_4206,N_3812,N_3482);
and U4207 (N_4207,N_3116,N_3524);
or U4208 (N_4208,N_2607,N_2560);
xor U4209 (N_4209,N_2719,N_3204);
or U4210 (N_4210,N_3271,N_3544);
or U4211 (N_4211,N_2595,N_2332);
or U4212 (N_4212,N_2008,N_2860);
xnor U4213 (N_4213,N_3922,N_3712);
or U4214 (N_4214,N_2642,N_3810);
and U4215 (N_4215,N_2798,N_3185);
xnor U4216 (N_4216,N_3638,N_2009);
nand U4217 (N_4217,N_2040,N_2749);
nor U4218 (N_4218,N_2794,N_3078);
xor U4219 (N_4219,N_2112,N_3266);
or U4220 (N_4220,N_2362,N_2266);
nand U4221 (N_4221,N_2119,N_3965);
nor U4222 (N_4222,N_2155,N_3280);
xnor U4223 (N_4223,N_3081,N_3328);
xnor U4224 (N_4224,N_3117,N_3734);
nor U4225 (N_4225,N_3427,N_3228);
nand U4226 (N_4226,N_3919,N_2278);
nor U4227 (N_4227,N_3589,N_2770);
nor U4228 (N_4228,N_3575,N_2896);
nor U4229 (N_4229,N_3632,N_2334);
nand U4230 (N_4230,N_3212,N_2814);
or U4231 (N_4231,N_3857,N_2216);
and U4232 (N_4232,N_3957,N_2890);
nor U4233 (N_4233,N_3849,N_2926);
nor U4234 (N_4234,N_2193,N_3051);
xor U4235 (N_4235,N_2311,N_3491);
and U4236 (N_4236,N_3236,N_3128);
or U4237 (N_4237,N_2225,N_3762);
or U4238 (N_4238,N_3337,N_3553);
nor U4239 (N_4239,N_3647,N_2934);
or U4240 (N_4240,N_2141,N_3087);
or U4241 (N_4241,N_2032,N_3874);
nand U4242 (N_4242,N_2256,N_3520);
nor U4243 (N_4243,N_3549,N_2467);
nand U4244 (N_4244,N_3885,N_3586);
nor U4245 (N_4245,N_2476,N_2836);
or U4246 (N_4246,N_2946,N_3454);
or U4247 (N_4247,N_2252,N_2114);
and U4248 (N_4248,N_3480,N_3774);
and U4249 (N_4249,N_3221,N_3345);
nand U4250 (N_4250,N_3769,N_2299);
nor U4251 (N_4251,N_3889,N_2960);
nand U4252 (N_4252,N_2609,N_3357);
and U4253 (N_4253,N_2680,N_2007);
nand U4254 (N_4254,N_3371,N_3286);
xnor U4255 (N_4255,N_3751,N_3025);
xor U4256 (N_4256,N_3147,N_3065);
nor U4257 (N_4257,N_3382,N_2474);
xnor U4258 (N_4258,N_3979,N_2104);
nor U4259 (N_4259,N_3187,N_2400);
and U4260 (N_4260,N_3598,N_3940);
nor U4261 (N_4261,N_2420,N_2406);
or U4262 (N_4262,N_3836,N_3854);
nand U4263 (N_4263,N_3610,N_2097);
nand U4264 (N_4264,N_2072,N_2953);
nand U4265 (N_4265,N_2472,N_2737);
xor U4266 (N_4266,N_2843,N_2274);
and U4267 (N_4267,N_3671,N_3323);
nand U4268 (N_4268,N_3219,N_3391);
nor U4269 (N_4269,N_2304,N_3652);
nand U4270 (N_4270,N_3177,N_2213);
xnor U4271 (N_4271,N_2062,N_2171);
or U4272 (N_4272,N_2481,N_3530);
nand U4273 (N_4273,N_3174,N_2792);
xnor U4274 (N_4274,N_2750,N_2748);
xor U4275 (N_4275,N_2716,N_2559);
xnor U4276 (N_4276,N_3068,N_2235);
nand U4277 (N_4277,N_3365,N_3884);
nand U4278 (N_4278,N_3168,N_3151);
nand U4279 (N_4279,N_2553,N_3711);
nand U4280 (N_4280,N_3093,N_3467);
nor U4281 (N_4281,N_2519,N_3559);
nor U4282 (N_4282,N_2521,N_2724);
and U4283 (N_4283,N_3408,N_2580);
nand U4284 (N_4284,N_3604,N_2700);
xor U4285 (N_4285,N_2259,N_2556);
or U4286 (N_4286,N_2395,N_3009);
and U4287 (N_4287,N_2145,N_2630);
nor U4288 (N_4288,N_2340,N_3704);
nand U4289 (N_4289,N_2056,N_3026);
or U4290 (N_4290,N_2298,N_2939);
or U4291 (N_4291,N_3672,N_3145);
xor U4292 (N_4292,N_3425,N_3698);
or U4293 (N_4293,N_2765,N_2533);
xor U4294 (N_4294,N_3714,N_2702);
xor U4295 (N_4295,N_3725,N_3290);
nand U4296 (N_4296,N_3314,N_3625);
or U4297 (N_4297,N_3437,N_3315);
or U4298 (N_4298,N_3888,N_3119);
and U4299 (N_4299,N_2356,N_2070);
or U4300 (N_4300,N_3645,N_3752);
or U4301 (N_4301,N_2703,N_3448);
nor U4302 (N_4302,N_2411,N_2620);
and U4303 (N_4303,N_3481,N_2688);
nor U4304 (N_4304,N_2764,N_3273);
xnor U4305 (N_4305,N_3343,N_3708);
xor U4306 (N_4306,N_2496,N_2582);
or U4307 (N_4307,N_3444,N_2598);
xor U4308 (N_4308,N_3056,N_3364);
nor U4309 (N_4309,N_2535,N_3354);
or U4310 (N_4310,N_3126,N_3497);
nand U4311 (N_4311,N_3413,N_3797);
or U4312 (N_4312,N_2210,N_3378);
and U4313 (N_4313,N_3157,N_3969);
nand U4314 (N_4314,N_3943,N_2078);
and U4315 (N_4315,N_2127,N_2547);
nor U4316 (N_4316,N_3697,N_2526);
xnor U4317 (N_4317,N_3091,N_3393);
and U4318 (N_4318,N_2586,N_3355);
or U4319 (N_4319,N_3803,N_2570);
nor U4320 (N_4320,N_2159,N_3293);
nand U4321 (N_4321,N_2049,N_3637);
nand U4322 (N_4322,N_2726,N_2955);
xnor U4323 (N_4323,N_3710,N_3614);
nor U4324 (N_4324,N_2000,N_2790);
and U4325 (N_4325,N_3538,N_2186);
or U4326 (N_4326,N_2760,N_2612);
nand U4327 (N_4327,N_3503,N_3129);
nor U4328 (N_4328,N_3269,N_2294);
xor U4329 (N_4329,N_2874,N_2385);
xor U4330 (N_4330,N_2913,N_2079);
and U4331 (N_4331,N_2985,N_2020);
and U4332 (N_4332,N_3977,N_2160);
xor U4333 (N_4333,N_3623,N_2555);
xor U4334 (N_4334,N_2269,N_3392);
and U4335 (N_4335,N_2937,N_3612);
nor U4336 (N_4336,N_3557,N_2658);
xnor U4337 (N_4337,N_3102,N_2919);
and U4338 (N_4338,N_2538,N_3347);
and U4339 (N_4339,N_2917,N_2625);
and U4340 (N_4340,N_3326,N_2618);
and U4341 (N_4341,N_2412,N_2279);
xnor U4342 (N_4342,N_2972,N_2158);
xnor U4343 (N_4343,N_2534,N_3396);
or U4344 (N_4344,N_2136,N_2417);
and U4345 (N_4345,N_3303,N_3983);
nand U4346 (N_4346,N_2397,N_2979);
or U4347 (N_4347,N_3738,N_3560);
nand U4348 (N_4348,N_2464,N_2758);
xor U4349 (N_4349,N_2855,N_2268);
and U4350 (N_4350,N_2102,N_3073);
nor U4351 (N_4351,N_3284,N_3505);
and U4352 (N_4352,N_3165,N_2211);
nand U4353 (N_4353,N_3960,N_2498);
nand U4354 (N_4354,N_2375,N_2791);
nand U4355 (N_4355,N_3304,N_3495);
xor U4356 (N_4356,N_2516,N_2194);
xor U4357 (N_4357,N_3903,N_3485);
or U4358 (N_4358,N_3372,N_2143);
and U4359 (N_4359,N_2809,N_2257);
and U4360 (N_4360,N_2650,N_3516);
or U4361 (N_4361,N_2878,N_3978);
or U4362 (N_4362,N_2440,N_2899);
and U4363 (N_4363,N_3334,N_2672);
nor U4364 (N_4364,N_3628,N_2988);
nand U4365 (N_4365,N_2361,N_2774);
and U4366 (N_4366,N_2823,N_3676);
nor U4367 (N_4367,N_3727,N_2525);
or U4368 (N_4368,N_2648,N_3041);
nand U4369 (N_4369,N_3146,N_3591);
nor U4370 (N_4370,N_3861,N_2984);
or U4371 (N_4371,N_3186,N_3968);
nand U4372 (N_4372,N_3180,N_3732);
nand U4373 (N_4373,N_3260,N_2709);
nor U4374 (N_4374,N_2380,N_2321);
or U4375 (N_4375,N_3108,N_2857);
xor U4376 (N_4376,N_3473,N_2142);
nand U4377 (N_4377,N_2057,N_3562);
nor U4378 (N_4378,N_2707,N_3058);
or U4379 (N_4379,N_3179,N_3899);
nand U4380 (N_4380,N_2471,N_2686);
and U4381 (N_4381,N_2347,N_2871);
and U4382 (N_4382,N_3227,N_2569);
or U4383 (N_4383,N_2484,N_2295);
nand U4384 (N_4384,N_2305,N_3576);
nor U4385 (N_4385,N_3439,N_2064);
nand U4386 (N_4386,N_3125,N_2631);
nor U4387 (N_4387,N_2005,N_2879);
nand U4388 (N_4388,N_3730,N_3817);
and U4389 (N_4389,N_2405,N_3457);
nor U4390 (N_4390,N_2222,N_3090);
and U4391 (N_4391,N_2043,N_3886);
nor U4392 (N_4392,N_2956,N_3434);
xor U4393 (N_4393,N_3429,N_2715);
or U4394 (N_4394,N_2998,N_3985);
nand U4395 (N_4395,N_2234,N_3897);
nand U4396 (N_4396,N_2434,N_3931);
or U4397 (N_4397,N_3744,N_2462);
nand U4398 (N_4398,N_3901,N_2923);
nand U4399 (N_4399,N_2113,N_2458);
or U4400 (N_4400,N_2442,N_3385);
and U4401 (N_4401,N_3319,N_3141);
nor U4402 (N_4402,N_3996,N_2435);
or U4403 (N_4403,N_3621,N_3764);
xnor U4404 (N_4404,N_3206,N_3696);
and U4405 (N_4405,N_2859,N_2550);
xor U4406 (N_4406,N_2966,N_3449);
and U4407 (N_4407,N_3923,N_3673);
and U4408 (N_4408,N_3781,N_3397);
or U4409 (N_4409,N_2296,N_2980);
or U4410 (N_4410,N_3510,N_3972);
or U4411 (N_4411,N_3864,N_3046);
nor U4412 (N_4412,N_2316,N_3980);
xnor U4413 (N_4413,N_2742,N_3409);
or U4414 (N_4414,N_2302,N_2647);
nor U4415 (N_4415,N_3907,N_2219);
nor U4416 (N_4416,N_3402,N_2796);
and U4417 (N_4417,N_2908,N_3188);
xnor U4418 (N_4418,N_2118,N_3785);
xor U4419 (N_4419,N_2187,N_2093);
or U4420 (N_4420,N_3276,N_3784);
xnor U4421 (N_4421,N_3646,N_2014);
or U4422 (N_4422,N_3488,N_3196);
and U4423 (N_4423,N_2092,N_2627);
nor U4424 (N_4424,N_2039,N_3525);
nor U4425 (N_4425,N_3593,N_3366);
nand U4426 (N_4426,N_2341,N_2762);
or U4427 (N_4427,N_2585,N_3813);
xnor U4428 (N_4428,N_3153,N_2041);
nand U4429 (N_4429,N_2741,N_2579);
or U4430 (N_4430,N_2753,N_3961);
xnor U4431 (N_4431,N_3703,N_2401);
or U4432 (N_4432,N_2641,N_3459);
nand U4433 (N_4433,N_3013,N_3329);
nand U4434 (N_4434,N_3692,N_3997);
nand U4435 (N_4435,N_2398,N_2454);
xnor U4436 (N_4436,N_3461,N_2643);
xor U4437 (N_4437,N_2530,N_2379);
and U4438 (N_4438,N_3740,N_2354);
xor U4439 (N_4439,N_2368,N_2952);
or U4440 (N_4440,N_3890,N_2515);
nor U4441 (N_4441,N_2418,N_3339);
nor U4442 (N_4442,N_2958,N_3720);
and U4443 (N_4443,N_2003,N_2196);
nand U4444 (N_4444,N_2262,N_3262);
and U4445 (N_4445,N_3937,N_3648);
or U4446 (N_4446,N_2604,N_2671);
and U4447 (N_4447,N_2690,N_2047);
nand U4448 (N_4448,N_3101,N_2001);
nor U4449 (N_4449,N_2837,N_3761);
nor U4450 (N_4450,N_2328,N_3830);
nand U4451 (N_4451,N_3579,N_3259);
or U4452 (N_4452,N_2320,N_2016);
nor U4453 (N_4453,N_3851,N_3311);
nor U4454 (N_4454,N_3455,N_2862);
and U4455 (N_4455,N_3216,N_2965);
and U4456 (N_4456,N_3742,N_2508);
xnor U4457 (N_4457,N_2810,N_3975);
nor U4458 (N_4458,N_2773,N_2327);
nand U4459 (N_4459,N_3537,N_3160);
nand U4460 (N_4460,N_2665,N_3261);
xor U4461 (N_4461,N_2827,N_2051);
xnor U4462 (N_4462,N_3103,N_3352);
nand U4463 (N_4463,N_3556,N_2307);
nand U4464 (N_4464,N_2578,N_3489);
and U4465 (N_4465,N_3063,N_2359);
xnor U4466 (N_4466,N_2066,N_2309);
nor U4467 (N_4467,N_2441,N_2490);
nor U4468 (N_4468,N_3839,N_3686);
nand U4469 (N_4469,N_2733,N_2968);
nand U4470 (N_4470,N_3814,N_2941);
nand U4471 (N_4471,N_3258,N_3332);
nand U4472 (N_4472,N_3309,N_2469);
and U4473 (N_4473,N_3360,N_2861);
and U4474 (N_4474,N_3569,N_2284);
xor U4475 (N_4475,N_2597,N_2539);
nand U4476 (N_4476,N_2682,N_3306);
and U4477 (N_4477,N_2568,N_2218);
nor U4478 (N_4478,N_2248,N_3546);
and U4479 (N_4479,N_2886,N_3535);
xnor U4480 (N_4480,N_3587,N_3148);
nor U4481 (N_4481,N_2329,N_2599);
or U4482 (N_4482,N_2433,N_2486);
nor U4483 (N_4483,N_3383,N_3629);
nand U4484 (N_4484,N_2338,N_3908);
or U4485 (N_4485,N_3816,N_3300);
xor U4486 (N_4486,N_3868,N_3012);
xnor U4487 (N_4487,N_3855,N_3973);
or U4488 (N_4488,N_3341,N_3787);
nand U4489 (N_4489,N_3723,N_2345);
nor U4490 (N_4490,N_3644,N_3420);
xor U4491 (N_4491,N_3974,N_2945);
and U4492 (N_4492,N_3100,N_2121);
or U4493 (N_4493,N_2177,N_3034);
nand U4494 (N_4494,N_2889,N_2129);
or U4495 (N_4495,N_2727,N_2833);
nand U4496 (N_4496,N_3853,N_3057);
nand U4497 (N_4497,N_2847,N_2626);
and U4498 (N_4498,N_3661,N_2826);
nand U4499 (N_4499,N_3432,N_3215);
or U4500 (N_4500,N_3184,N_2427);
xnor U4501 (N_4501,N_3451,N_2322);
nand U4502 (N_4502,N_2706,N_2565);
nor U4503 (N_4503,N_3682,N_2050);
nand U4504 (N_4504,N_3421,N_2745);
and U4505 (N_4505,N_2232,N_3359);
nand U4506 (N_4506,N_3674,N_3181);
nand U4507 (N_4507,N_3049,N_3018);
or U4508 (N_4508,N_2638,N_3154);
nor U4509 (N_4509,N_2314,N_3193);
nand U4510 (N_4510,N_3498,N_2271);
or U4511 (N_4511,N_2624,N_2173);
nor U4512 (N_4512,N_2903,N_2775);
and U4513 (N_4513,N_3202,N_2488);
or U4514 (N_4514,N_2712,N_3879);
or U4515 (N_4515,N_3414,N_2964);
nand U4516 (N_4516,N_3846,N_2111);
or U4517 (N_4517,N_2301,N_2950);
nor U4518 (N_4518,N_3831,N_2408);
and U4519 (N_4519,N_3169,N_3528);
or U4520 (N_4520,N_2520,N_3114);
and U4521 (N_4521,N_3152,N_3641);
and U4522 (N_4522,N_3431,N_3029);
nor U4523 (N_4523,N_2736,N_2482);
and U4524 (N_4524,N_2564,N_2778);
nand U4525 (N_4525,N_2025,N_3217);
and U4526 (N_4526,N_3150,N_2163);
or U4527 (N_4527,N_3758,N_3298);
xor U4528 (N_4528,N_3121,N_2371);
xnor U4529 (N_4529,N_2959,N_2199);
xnor U4530 (N_4530,N_3577,N_3190);
nand U4531 (N_4531,N_3070,N_2615);
xnor U4532 (N_4532,N_2153,N_2828);
or U4533 (N_4533,N_2637,N_3566);
nor U4534 (N_4534,N_3799,N_3171);
nor U4535 (N_4535,N_2824,N_2906);
and U4536 (N_4536,N_2936,N_3571);
or U4537 (N_4537,N_2150,N_2149);
nand U4538 (N_4538,N_2132,N_2838);
nand U4539 (N_4539,N_3035,N_2280);
xnor U4540 (N_4540,N_3416,N_3340);
nand U4541 (N_4541,N_3963,N_2714);
and U4542 (N_4542,N_2713,N_2746);
and U4543 (N_4543,N_2779,N_2139);
and U4544 (N_4544,N_3285,N_2258);
or U4545 (N_4545,N_2873,N_3406);
nand U4546 (N_4546,N_3912,N_3322);
and U4547 (N_4547,N_3380,N_3914);
xnor U4548 (N_4548,N_2841,N_3268);
nand U4549 (N_4549,N_2292,N_2930);
nor U4550 (N_4550,N_3526,N_3265);
nand U4551 (N_4551,N_2933,N_2315);
or U4552 (N_4552,N_3045,N_3871);
nor U4553 (N_4553,N_3232,N_2619);
nor U4554 (N_4554,N_3122,N_3255);
nand U4555 (N_4555,N_2927,N_3500);
nand U4556 (N_4556,N_3004,N_3815);
nand U4557 (N_4557,N_3582,N_3006);
xnor U4558 (N_4558,N_3948,N_2744);
and U4559 (N_4559,N_2431,N_3172);
xnor U4560 (N_4560,N_3238,N_2759);
nor U4561 (N_4561,N_3966,N_3639);
and U4562 (N_4562,N_2137,N_3615);
xnor U4563 (N_4563,N_2059,N_2986);
xor U4564 (N_4564,N_3872,N_2451);
nand U4565 (N_4565,N_2594,N_2035);
and U4566 (N_4566,N_2182,N_3533);
or U4567 (N_4567,N_3820,N_2881);
nand U4568 (N_4568,N_3106,N_2655);
or U4569 (N_4569,N_3920,N_3351);
or U4570 (N_4570,N_3517,N_2783);
nor U4571 (N_4571,N_3954,N_2848);
and U4572 (N_4572,N_3658,N_3294);
nor U4573 (N_4573,N_2584,N_3243);
and U4574 (N_4574,N_2273,N_3602);
and U4575 (N_4575,N_3192,N_3898);
and U4576 (N_4576,N_2850,N_2728);
and U4577 (N_4577,N_2493,N_2633);
and U4578 (N_4578,N_3140,N_3230);
or U4579 (N_4579,N_3990,N_3603);
nor U4580 (N_4580,N_3028,N_3993);
or U4581 (N_4581,N_3401,N_3104);
nor U4582 (N_4582,N_2220,N_3547);
and U4583 (N_4583,N_2789,N_2507);
or U4584 (N_4584,N_3709,N_3446);
or U4585 (N_4585,N_2684,N_3684);
and U4586 (N_4586,N_3302,N_3540);
or U4587 (N_4587,N_2681,N_2148);
nand U4588 (N_4588,N_3660,N_3115);
xnor U4589 (N_4589,N_3032,N_3835);
nand U4590 (N_4590,N_3253,N_2875);
nor U4591 (N_4591,N_2028,N_2291);
or U4592 (N_4592,N_3478,N_2567);
or U4593 (N_4593,N_3281,N_2029);
nor U4594 (N_4594,N_3745,N_2455);
or U4595 (N_4595,N_2531,N_3176);
xnor U4596 (N_4596,N_2052,N_2445);
nor U4597 (N_4597,N_3240,N_2977);
or U4598 (N_4598,N_2456,N_3027);
nand U4599 (N_4599,N_2407,N_2404);
nor U4600 (N_4600,N_2337,N_2543);
nor U4601 (N_4601,N_3941,N_2017);
or U4602 (N_4602,N_2795,N_3932);
xor U4603 (N_4603,N_3079,N_3194);
xnor U4604 (N_4604,N_3054,N_3436);
xnor U4605 (N_4605,N_2544,N_2990);
nand U4606 (N_4606,N_2067,N_3040);
nor U4607 (N_4607,N_3607,N_2781);
nor U4608 (N_4608,N_3802,N_2853);
and U4609 (N_4609,N_3991,N_2250);
and U4610 (N_4610,N_3224,N_3189);
or U4611 (N_4611,N_2246,N_2596);
nor U4612 (N_4612,N_3995,N_2528);
nor U4613 (N_4613,N_3715,N_2154);
nor U4614 (N_4614,N_3695,N_3344);
xnor U4615 (N_4615,N_2610,N_2644);
xnor U4616 (N_4616,N_3159,N_3486);
and U4617 (N_4617,N_2766,N_2021);
nand U4618 (N_4618,N_2524,N_3237);
or U4619 (N_4619,N_2629,N_2685);
and U4620 (N_4620,N_3892,N_3010);
or U4621 (N_4621,N_3893,N_3950);
xor U4622 (N_4622,N_3600,N_3251);
xor U4623 (N_4623,N_2255,N_2969);
and U4624 (N_4624,N_2771,N_3405);
nand U4625 (N_4625,N_3759,N_3928);
nor U4626 (N_4626,N_2061,N_3370);
nor U4627 (N_4627,N_3270,N_2587);
or U4628 (N_4628,N_2504,N_3521);
nor U4629 (N_4629,N_2576,N_2084);
xnor U4630 (N_4630,N_2654,N_2711);
xnor U4631 (N_4631,N_3375,N_2048);
nand U4632 (N_4632,N_2396,N_2529);
xnor U4633 (N_4633,N_2517,N_3736);
xnor U4634 (N_4634,N_3911,N_3331);
xor U4635 (N_4635,N_3805,N_3548);
and U4636 (N_4636,N_3511,N_3583);
and U4637 (N_4637,N_2448,N_2602);
xor U4638 (N_4638,N_2699,N_2573);
and U4639 (N_4639,N_2721,N_3527);
or U4640 (N_4640,N_2805,N_3305);
nand U4641 (N_4641,N_3211,N_3263);
nand U4642 (N_4642,N_3826,N_2804);
nor U4643 (N_4643,N_3792,N_3016);
nand U4644 (N_4644,N_2920,N_3681);
or U4645 (N_4645,N_2287,N_3574);
nor U4646 (N_4646,N_2613,N_2677);
and U4647 (N_4647,N_3887,N_3275);
or U4648 (N_4648,N_3693,N_3749);
and U4649 (N_4649,N_3017,N_3085);
nand U4650 (N_4650,N_3062,N_2073);
xor U4651 (N_4651,N_3424,N_3435);
nand U4652 (N_4652,N_3933,N_2303);
or U4653 (N_4653,N_2835,N_3852);
xor U4654 (N_4654,N_2392,N_3506);
xor U4655 (N_4655,N_2905,N_2352);
xor U4656 (N_4656,N_2366,N_2501);
xor U4657 (N_4657,N_2238,N_3955);
xnor U4658 (N_4658,N_2813,N_2233);
xnor U4659 (N_4659,N_3883,N_3756);
nand U4660 (N_4660,N_2198,N_3760);
xor U4661 (N_4661,N_2202,N_3654);
or U4662 (N_4662,N_3894,N_2367);
and U4663 (N_4663,N_2811,N_3818);
or U4664 (N_4664,N_2174,N_2065);
nand U4665 (N_4665,N_2821,N_2053);
nand U4666 (N_4666,N_3649,N_2013);
nand U4667 (N_4667,N_3620,N_3514);
nor U4668 (N_4668,N_2793,N_2087);
and U4669 (N_4669,N_2554,N_2829);
and U4670 (N_4670,N_2365,N_2856);
nand U4671 (N_4671,N_3627,N_3292);
and U4672 (N_4672,N_3252,N_3542);
or U4673 (N_4673,N_3348,N_2723);
xor U4674 (N_4674,N_2249,N_2982);
or U4675 (N_4675,N_3775,N_2247);
nor U4676 (N_4676,N_2608,N_3395);
nor U4677 (N_4677,N_2993,N_3296);
nor U4678 (N_4678,N_3474,N_2591);
nand U4679 (N_4679,N_2801,N_2909);
nand U4680 (N_4680,N_2080,N_3837);
nor U4681 (N_4681,N_2807,N_3450);
xnor U4682 (N_4682,N_2422,N_2181);
xor U4683 (N_4683,N_2963,N_3452);
and U4684 (N_4684,N_3082,N_3793);
or U4685 (N_4685,N_2800,N_3716);
nor U4686 (N_4686,N_3132,N_2888);
nor U4687 (N_4687,N_2803,N_2931);
xnor U4688 (N_4688,N_3801,N_2616);
or U4689 (N_4689,N_2106,N_2757);
nand U4690 (N_4690,N_3924,N_2083);
or U4691 (N_4691,N_2732,N_2283);
or U4692 (N_4692,N_3651,N_2954);
xor U4693 (N_4693,N_3135,N_3388);
or U4694 (N_4694,N_2710,N_2103);
nand U4695 (N_4695,N_3075,N_3906);
and U4696 (N_4696,N_3786,N_3476);
nor U4697 (N_4697,N_2373,N_2692);
xnor U4698 (N_4698,N_2054,N_3433);
xnor U4699 (N_4699,N_3030,N_3865);
nor U4700 (N_4700,N_3301,N_3036);
and U4701 (N_4701,N_3581,N_3428);
nand U4702 (N_4702,N_3982,N_2503);
nand U4703 (N_4703,N_2751,N_3418);
nand U4704 (N_4704,N_3946,N_3362);
nand U4705 (N_4705,N_2215,N_2231);
nand U4706 (N_4706,N_3964,N_3896);
xnor U4707 (N_4707,N_3453,N_2342);
and U4708 (N_4708,N_3245,N_2743);
xor U4709 (N_4709,N_2018,N_2074);
nand U4710 (N_4710,N_2971,N_3691);
and U4711 (N_4711,N_2904,N_2893);
or U4712 (N_4712,N_2179,N_2364);
nand U4713 (N_4713,N_3880,N_2251);
and U4714 (N_4714,N_3741,N_3513);
nor U4715 (N_4715,N_3791,N_2095);
nand U4716 (N_4716,N_2891,N_2172);
or U4717 (N_4717,N_3984,N_3838);
nor U4718 (N_4718,N_3819,N_3986);
xnor U4719 (N_4719,N_3317,N_2867);
nor U4720 (N_4720,N_2676,N_3592);
or U4721 (N_4721,N_3945,N_2739);
nand U4722 (N_4722,N_2776,N_3936);
nor U4723 (N_4723,N_3939,N_3250);
nor U4724 (N_4724,N_2197,N_2830);
or U4725 (N_4725,N_3074,N_3422);
and U4726 (N_4726,N_3834,N_2740);
xor U4727 (N_4727,N_2865,N_2042);
or U4728 (N_4728,N_2389,N_2872);
nor U4729 (N_4729,N_2011,N_2240);
xor U4730 (N_4730,N_3822,N_3066);
nand U4731 (N_4731,N_3244,N_2541);
and U4732 (N_4732,N_2976,N_2940);
and U4733 (N_4733,N_2802,N_3667);
and U4734 (N_4734,N_2369,N_2323);
or U4735 (N_4735,N_3935,N_3543);
xor U4736 (N_4736,N_2223,N_3105);
nor U4737 (N_4737,N_2901,N_2911);
or U4738 (N_4738,N_2470,N_2632);
nor U4739 (N_4739,N_3800,N_2128);
xor U4740 (N_4740,N_2961,N_3277);
nor U4741 (N_4741,N_3705,N_2506);
and U4742 (N_4742,N_2082,N_2902);
xnor U4743 (N_4743,N_2812,N_3572);
nand U4744 (N_4744,N_2116,N_3248);
xnor U4745 (N_4745,N_3509,N_2734);
or U4746 (N_4746,N_3369,N_3441);
xor U4747 (N_4747,N_2034,N_3541);
nor U4748 (N_4748,N_2673,N_2144);
nor U4749 (N_4749,N_3256,N_2717);
nand U4750 (N_4750,N_2165,N_2575);
or U4751 (N_4751,N_3701,N_3060);
xor U4752 (N_4752,N_3333,N_2126);
nor U4753 (N_4753,N_3490,N_2351);
or U4754 (N_4754,N_3668,N_3882);
nand U4755 (N_4755,N_3573,N_2038);
and U4756 (N_4756,N_3913,N_3233);
and U4757 (N_4757,N_2190,N_3468);
nand U4758 (N_4758,N_3324,N_2854);
and U4759 (N_4759,N_3653,N_2577);
nand U4760 (N_4760,N_3412,N_3064);
and U4761 (N_4761,N_2100,N_3092);
nor U4762 (N_4762,N_2763,N_3863);
nand U4763 (N_4763,N_3735,N_3794);
or U4764 (N_4764,N_2782,N_2060);
nand U4765 (N_4765,N_2844,N_2443);
and U4766 (N_4766,N_3307,N_2207);
or U4767 (N_4767,N_2229,N_2151);
nand U4768 (N_4768,N_3635,N_2834);
nand U4769 (N_4769,N_3274,N_2797);
xnor U4770 (N_4770,N_2312,N_3930);
nand U4771 (N_4771,N_2293,N_2019);
and U4772 (N_4772,N_2666,N_2799);
xor U4773 (N_4773,N_2188,N_2910);
or U4774 (N_4774,N_3609,N_3053);
nand U4775 (N_4775,N_3381,N_2601);
nor U4776 (N_4776,N_3411,N_3772);
nand U4777 (N_4777,N_2069,N_2166);
xor U4778 (N_4778,N_3419,N_2487);
nand U4779 (N_4779,N_2617,N_3387);
nand U4780 (N_4780,N_2527,N_3494);
or U4781 (N_4781,N_3679,N_3076);
nor U4782 (N_4782,N_3297,N_2869);
xor U4783 (N_4783,N_3218,N_2286);
xnor U4784 (N_4784,N_2668,N_2916);
nand U4785 (N_4785,N_2206,N_3798);
nand U4786 (N_4786,N_2611,N_2704);
xor U4787 (N_4787,N_3379,N_2175);
and U4788 (N_4788,N_2614,N_2426);
and U4789 (N_4789,N_3790,N_2634);
and U4790 (N_4790,N_2372,N_3633);
and U4791 (N_4791,N_3636,N_3584);
xor U4792 (N_4792,N_2122,N_3778);
xnor U4793 (N_4793,N_3417,N_3390);
nor U4794 (N_4794,N_2667,N_3138);
nor U4795 (N_4795,N_2416,N_3316);
or U4796 (N_4796,N_2317,N_3241);
nand U4797 (N_4797,N_3951,N_2970);
nor U4798 (N_4798,N_2253,N_2313);
nor U4799 (N_4799,N_2390,N_2123);
and U4800 (N_4800,N_3619,N_2353);
or U4801 (N_4801,N_3597,N_3312);
nor U4802 (N_4802,N_3134,N_2237);
and U4803 (N_4803,N_3052,N_3149);
and U4804 (N_4804,N_3554,N_3728);
nor U4805 (N_4805,N_3464,N_3173);
or U4806 (N_4806,N_2852,N_2989);
xnor U4807 (N_4807,N_2436,N_2914);
and U4808 (N_4808,N_2277,N_2209);
nand U4809 (N_4809,N_2502,N_2147);
xor U4810 (N_4810,N_3777,N_3249);
nand U4811 (N_4811,N_3601,N_3155);
nand U4812 (N_4812,N_2718,N_3374);
xor U4813 (N_4813,N_3848,N_3335);
xnor U4814 (N_4814,N_3833,N_2344);
nand U4815 (N_4815,N_2363,N_3071);
and U4816 (N_4816,N_2391,N_3568);
xor U4817 (N_4817,N_2109,N_2996);
nand U4818 (N_4818,N_3257,N_3267);
nor U4819 (N_4819,N_2135,N_2994);
nand U4820 (N_4820,N_3438,N_3539);
nor U4821 (N_4821,N_2656,N_3022);
nor U4822 (N_4822,N_3825,N_2883);
nor U4823 (N_4823,N_3037,N_3876);
or U4824 (N_4824,N_3622,N_3384);
nand U4825 (N_4825,N_3508,N_3426);
nor U4826 (N_4826,N_3811,N_3788);
nand U4827 (N_4827,N_3127,N_3024);
xnor U4828 (N_4828,N_2592,N_3909);
or U4829 (N_4829,N_3000,N_2325);
and U4830 (N_4830,N_2036,N_2512);
xnor U4831 (N_4831,N_2600,N_2639);
xnor U4832 (N_4832,N_2708,N_3796);
nor U4833 (N_4833,N_2318,N_3363);
and U4834 (N_4834,N_2851,N_3595);
or U4835 (N_4835,N_2473,N_2720);
xor U4836 (N_4836,N_2542,N_2402);
nor U4837 (N_4837,N_2089,N_2319);
nor U4838 (N_4838,N_3721,N_2324);
and U4839 (N_4839,N_2330,N_3650);
xnor U4840 (N_4840,N_2015,N_3618);
nor U4841 (N_4841,N_2333,N_2752);
nand U4842 (N_4842,N_2477,N_3678);
nor U4843 (N_4843,N_2820,N_2832);
and U4844 (N_4844,N_2290,N_2660);
nand U4845 (N_4845,N_3044,N_3136);
or U4846 (N_4846,N_2942,N_2381);
xor U4847 (N_4847,N_3008,N_2178);
xnor U4848 (N_4848,N_2243,N_3927);
xnor U4849 (N_4849,N_2138,N_3971);
nand U4850 (N_4850,N_3349,N_2588);
xnor U4851 (N_4851,N_2306,N_3925);
nand U4852 (N_4852,N_3440,N_3376);
and U4853 (N_4853,N_2653,N_2806);
or U4854 (N_4854,N_2428,N_3611);
xor U4855 (N_4855,N_2645,N_3342);
xnor U4856 (N_4856,N_2421,N_2938);
and U4857 (N_4857,N_3403,N_2943);
nor U4858 (N_4858,N_3130,N_2583);
or U4859 (N_4859,N_2730,N_3860);
and U4860 (N_4860,N_3089,N_2987);
nand U4861 (N_4861,N_3118,N_3588);
nand U4862 (N_4862,N_2622,N_2831);
and U4863 (N_4863,N_2300,N_3162);
xnor U4864 (N_4864,N_2695,N_3291);
xnor U4865 (N_4865,N_2887,N_2551);
nor U4866 (N_4866,N_2326,N_2081);
nand U4867 (N_4867,N_3069,N_3182);
nand U4868 (N_4868,N_2208,N_3005);
or U4869 (N_4869,N_2701,N_2880);
and U4870 (N_4870,N_2777,N_2161);
nand U4871 (N_4871,N_3580,N_3299);
xnor U4872 (N_4872,N_2449,N_3522);
nor U4873 (N_4873,N_3445,N_2203);
xnor U4874 (N_4874,N_3795,N_3055);
and U4875 (N_4875,N_3430,N_2098);
and U4876 (N_4876,N_3492,N_2511);
nor U4877 (N_4877,N_2975,N_2510);
or U4878 (N_4878,N_3023,N_3616);
nand U4879 (N_4879,N_3680,N_3099);
nor U4880 (N_4880,N_3843,N_3750);
or U4881 (N_4881,N_3669,N_3061);
and U4882 (N_4882,N_3015,N_3677);
and U4883 (N_4883,N_3199,N_3958);
and U4884 (N_4884,N_3095,N_3442);
xor U4885 (N_4885,N_2500,N_2343);
nor U4886 (N_4886,N_2628,N_2669);
and U4887 (N_4887,N_3755,N_3642);
xor U4888 (N_4888,N_3501,N_2731);
xnor U4889 (N_4889,N_2245,N_3850);
nor U4890 (N_4890,N_3746,N_3456);
or U4891 (N_4891,N_3287,N_2840);
nor U4892 (N_4892,N_3873,N_3733);
or U4893 (N_4893,N_2414,N_3994);
nor U4894 (N_4894,N_2921,N_2687);
or U4895 (N_4895,N_3763,N_3223);
or U4896 (N_4896,N_2045,N_3205);
xnor U4897 (N_4897,N_2866,N_3687);
and U4898 (N_4898,N_3443,N_2981);
or U4899 (N_4899,N_2146,N_2377);
nand U4900 (N_4900,N_2006,N_3458);
and U4901 (N_4901,N_3719,N_3318);
and U4902 (N_4902,N_2046,N_3475);
nand U4903 (N_4903,N_2224,N_3471);
or U4904 (N_4904,N_2063,N_2085);
or U4905 (N_4905,N_3330,N_3042);
nor U4906 (N_4906,N_3133,N_3992);
xor U4907 (N_4907,N_3998,N_3313);
nor U4908 (N_4908,N_3399,N_2260);
xor U4909 (N_4909,N_3900,N_3279);
xnor U4910 (N_4910,N_3608,N_3624);
and U4911 (N_4911,N_2022,N_3891);
nor U4912 (N_4912,N_3001,N_3019);
xnor U4913 (N_4913,N_3242,N_3904);
nor U4914 (N_4914,N_2491,N_2907);
and U4915 (N_4915,N_2509,N_3959);
nor U4916 (N_4916,N_3463,N_3630);
nand U4917 (N_4917,N_3869,N_2652);
or U4918 (N_4918,N_3938,N_3111);
xor U4919 (N_4919,N_3688,N_2495);
or U4920 (N_4920,N_3321,N_2463);
nor U4921 (N_4921,N_3197,N_3477);
nand U4922 (N_4922,N_3462,N_2376);
or U4923 (N_4923,N_3902,N_2947);
and U4924 (N_4924,N_2722,N_2297);
xnor U4925 (N_4925,N_2518,N_2282);
nand U4926 (N_4926,N_2110,N_2967);
nand U4927 (N_4927,N_3163,N_2170);
nor U4928 (N_4928,N_3389,N_2548);
or U4929 (N_4929,N_3561,N_3112);
xor U4930 (N_4930,N_3088,N_2818);
xor U4931 (N_4931,N_3254,N_2485);
or U4932 (N_4932,N_3631,N_2214);
nor U4933 (N_4933,N_2265,N_2761);
xnor U4934 (N_4934,N_3666,N_3203);
xnor U4935 (N_4935,N_3878,N_2978);
nand U4936 (N_4936,N_2935,N_2839);
xnor U4937 (N_4937,N_3059,N_2281);
nor U4938 (N_4938,N_2212,N_3410);
nand U4939 (N_4939,N_2075,N_3771);
and U4940 (N_4940,N_3877,N_2572);
nor U4941 (N_4941,N_3578,N_2842);
xnor U4942 (N_4942,N_2090,N_2204);
or U4943 (N_4943,N_2992,N_3665);
or U4944 (N_4944,N_2747,N_2162);
xor U4945 (N_4945,N_3515,N_3086);
xnor U4946 (N_4946,N_3519,N_2010);
and U4947 (N_4947,N_2662,N_3656);
and U4948 (N_4948,N_3198,N_2808);
xor U4949 (N_4949,N_2870,N_2974);
nand U4950 (N_4950,N_2545,N_2386);
nor U4951 (N_4951,N_2536,N_2755);
or U4952 (N_4952,N_3246,N_3821);
or U4953 (N_4953,N_3999,N_2355);
nand U4954 (N_4954,N_3098,N_2561);
and U4955 (N_4955,N_3558,N_2349);
nand U4956 (N_4956,N_3856,N_3033);
xnor U4957 (N_4957,N_2864,N_2275);
nor U4958 (N_4958,N_2272,N_3047);
nor U4959 (N_4959,N_3594,N_2055);
nand U4960 (N_4960,N_2574,N_3137);
xnor U4961 (N_4961,N_2674,N_3634);
nor U4962 (N_4962,N_2310,N_2951);
or U4963 (N_4963,N_2024,N_2817);
xnor U4964 (N_4964,N_3472,N_3084);
nor U4965 (N_4965,N_3722,N_2415);
nand U4966 (N_4966,N_2164,N_2991);
xor U4967 (N_4967,N_2117,N_2738);
xnor U4968 (N_4968,N_3655,N_3706);
and U4969 (N_4969,N_3640,N_2894);
nand U4970 (N_4970,N_3226,N_3512);
or U4971 (N_4971,N_3981,N_3690);
nor U4972 (N_4972,N_2393,N_2384);
and U4973 (N_4973,N_3915,N_2784);
nand U4974 (N_4974,N_3626,N_3356);
nor U4975 (N_4975,N_3531,N_2772);
nor U4976 (N_4976,N_2227,N_2670);
and U4977 (N_4977,N_3209,N_3231);
xor U4978 (N_4978,N_3564,N_3662);
xnor U4979 (N_4979,N_3753,N_3832);
nor U4980 (N_4980,N_3020,N_3107);
and U4981 (N_4981,N_3164,N_2068);
or U4982 (N_4982,N_3415,N_2460);
or U4983 (N_4983,N_2184,N_3847);
xor U4984 (N_4984,N_2308,N_3282);
and U4985 (N_4985,N_2285,N_3043);
nor U4986 (N_4986,N_2221,N_2241);
and U4987 (N_4987,N_2780,N_3346);
xor U4988 (N_4988,N_3699,N_2480);
or U4989 (N_4989,N_2925,N_2623);
nand U4990 (N_4990,N_2107,N_3113);
nor U4991 (N_4991,N_2661,N_3235);
nand U4992 (N_4992,N_3469,N_3926);
xor U4993 (N_4993,N_3220,N_3585);
nand U4994 (N_4994,N_2461,N_2239);
nand U4995 (N_4995,N_2756,N_2410);
or U4996 (N_4996,N_3953,N_2192);
or U4997 (N_4997,N_2115,N_2168);
or U4998 (N_4998,N_3905,N_3689);
and U4999 (N_4999,N_2769,N_2228);
xnor U5000 (N_5000,N_2199,N_2283);
nor U5001 (N_5001,N_3614,N_3511);
nor U5002 (N_5002,N_2047,N_3870);
xnor U5003 (N_5003,N_3008,N_2757);
xor U5004 (N_5004,N_3740,N_2615);
xnor U5005 (N_5005,N_2878,N_3869);
and U5006 (N_5006,N_2066,N_2814);
nor U5007 (N_5007,N_3764,N_2857);
xnor U5008 (N_5008,N_2622,N_2774);
nor U5009 (N_5009,N_3617,N_2647);
nor U5010 (N_5010,N_3780,N_2448);
nand U5011 (N_5011,N_3760,N_2333);
nand U5012 (N_5012,N_3793,N_3261);
or U5013 (N_5013,N_3598,N_2203);
or U5014 (N_5014,N_2037,N_2488);
xnor U5015 (N_5015,N_3709,N_3473);
and U5016 (N_5016,N_2721,N_2988);
or U5017 (N_5017,N_2794,N_3471);
and U5018 (N_5018,N_2117,N_2680);
or U5019 (N_5019,N_2410,N_2377);
or U5020 (N_5020,N_3145,N_3353);
and U5021 (N_5021,N_2964,N_3069);
nor U5022 (N_5022,N_2977,N_3074);
and U5023 (N_5023,N_2855,N_2919);
or U5024 (N_5024,N_2582,N_3690);
or U5025 (N_5025,N_2089,N_3038);
or U5026 (N_5026,N_3069,N_3618);
or U5027 (N_5027,N_3260,N_2613);
or U5028 (N_5028,N_2820,N_2180);
or U5029 (N_5029,N_2106,N_2610);
or U5030 (N_5030,N_3237,N_3471);
nand U5031 (N_5031,N_2662,N_2593);
nor U5032 (N_5032,N_3902,N_3023);
and U5033 (N_5033,N_2552,N_2096);
and U5034 (N_5034,N_3234,N_3058);
xnor U5035 (N_5035,N_2814,N_3622);
nand U5036 (N_5036,N_2934,N_2760);
xor U5037 (N_5037,N_3750,N_2594);
nor U5038 (N_5038,N_2541,N_2184);
or U5039 (N_5039,N_2782,N_3956);
nand U5040 (N_5040,N_2185,N_2567);
nor U5041 (N_5041,N_3204,N_2443);
nand U5042 (N_5042,N_3034,N_3064);
xnor U5043 (N_5043,N_2499,N_2064);
nand U5044 (N_5044,N_2968,N_3758);
or U5045 (N_5045,N_2552,N_3437);
and U5046 (N_5046,N_3464,N_2863);
nor U5047 (N_5047,N_2392,N_3584);
and U5048 (N_5048,N_3294,N_2757);
and U5049 (N_5049,N_2582,N_3864);
nor U5050 (N_5050,N_3037,N_2312);
nand U5051 (N_5051,N_3351,N_3159);
xnor U5052 (N_5052,N_3890,N_3535);
xor U5053 (N_5053,N_2918,N_2160);
nor U5054 (N_5054,N_3434,N_2073);
nor U5055 (N_5055,N_3506,N_2703);
and U5056 (N_5056,N_3989,N_3686);
nor U5057 (N_5057,N_3735,N_3978);
nor U5058 (N_5058,N_3078,N_3767);
xor U5059 (N_5059,N_2335,N_3276);
or U5060 (N_5060,N_3969,N_2181);
and U5061 (N_5061,N_2050,N_2687);
nand U5062 (N_5062,N_3121,N_3738);
nand U5063 (N_5063,N_3649,N_2184);
and U5064 (N_5064,N_3825,N_3161);
nand U5065 (N_5065,N_3804,N_3180);
or U5066 (N_5066,N_2295,N_3936);
nand U5067 (N_5067,N_2565,N_3408);
or U5068 (N_5068,N_3025,N_2011);
and U5069 (N_5069,N_2765,N_2565);
nand U5070 (N_5070,N_3781,N_3725);
or U5071 (N_5071,N_3649,N_2036);
nor U5072 (N_5072,N_3607,N_2102);
xor U5073 (N_5073,N_3963,N_3666);
nand U5074 (N_5074,N_2420,N_2197);
nand U5075 (N_5075,N_2667,N_2710);
xor U5076 (N_5076,N_3053,N_2486);
nand U5077 (N_5077,N_3177,N_2532);
or U5078 (N_5078,N_3743,N_2040);
nand U5079 (N_5079,N_3090,N_3209);
xor U5080 (N_5080,N_3740,N_3562);
xnor U5081 (N_5081,N_3472,N_3222);
nand U5082 (N_5082,N_2005,N_3123);
or U5083 (N_5083,N_3797,N_3753);
nor U5084 (N_5084,N_3075,N_2791);
nor U5085 (N_5085,N_2997,N_2389);
nand U5086 (N_5086,N_2691,N_3836);
nand U5087 (N_5087,N_3906,N_3774);
nand U5088 (N_5088,N_3692,N_2463);
nand U5089 (N_5089,N_3502,N_3318);
nand U5090 (N_5090,N_3859,N_2196);
nand U5091 (N_5091,N_2747,N_3332);
nor U5092 (N_5092,N_2534,N_3560);
or U5093 (N_5093,N_2603,N_2463);
or U5094 (N_5094,N_3686,N_2244);
xor U5095 (N_5095,N_3663,N_2360);
and U5096 (N_5096,N_2061,N_2871);
xor U5097 (N_5097,N_3531,N_3045);
nand U5098 (N_5098,N_3617,N_3103);
and U5099 (N_5099,N_2649,N_3409);
nand U5100 (N_5100,N_2964,N_2827);
nand U5101 (N_5101,N_3564,N_2545);
nor U5102 (N_5102,N_3941,N_3577);
and U5103 (N_5103,N_2270,N_3286);
xor U5104 (N_5104,N_3078,N_3884);
and U5105 (N_5105,N_2996,N_3512);
or U5106 (N_5106,N_3983,N_2502);
nand U5107 (N_5107,N_2739,N_2268);
xnor U5108 (N_5108,N_3484,N_2454);
xnor U5109 (N_5109,N_2849,N_2899);
xor U5110 (N_5110,N_3566,N_2418);
nand U5111 (N_5111,N_2556,N_3499);
and U5112 (N_5112,N_3335,N_3351);
nor U5113 (N_5113,N_3889,N_2663);
or U5114 (N_5114,N_3440,N_2506);
nand U5115 (N_5115,N_2499,N_2125);
xor U5116 (N_5116,N_3294,N_3389);
xor U5117 (N_5117,N_3001,N_2245);
xnor U5118 (N_5118,N_3898,N_2048);
xnor U5119 (N_5119,N_2557,N_2144);
nor U5120 (N_5120,N_2831,N_3789);
xnor U5121 (N_5121,N_3231,N_2691);
xor U5122 (N_5122,N_3241,N_3776);
or U5123 (N_5123,N_3107,N_3942);
nor U5124 (N_5124,N_2752,N_2024);
or U5125 (N_5125,N_3560,N_2566);
and U5126 (N_5126,N_2847,N_2748);
nor U5127 (N_5127,N_2426,N_3894);
nand U5128 (N_5128,N_2447,N_2256);
xnor U5129 (N_5129,N_2987,N_3937);
nand U5130 (N_5130,N_2609,N_3141);
xnor U5131 (N_5131,N_2597,N_3727);
nand U5132 (N_5132,N_3253,N_3924);
or U5133 (N_5133,N_3126,N_3654);
nand U5134 (N_5134,N_3540,N_3059);
xor U5135 (N_5135,N_2285,N_2677);
xor U5136 (N_5136,N_3684,N_3846);
nor U5137 (N_5137,N_3929,N_2685);
nand U5138 (N_5138,N_3524,N_2830);
nor U5139 (N_5139,N_2902,N_3477);
xor U5140 (N_5140,N_3032,N_2424);
nand U5141 (N_5141,N_3997,N_2584);
nand U5142 (N_5142,N_3232,N_3038);
nor U5143 (N_5143,N_2408,N_3001);
and U5144 (N_5144,N_3265,N_2485);
xor U5145 (N_5145,N_3832,N_3140);
or U5146 (N_5146,N_3442,N_2635);
nand U5147 (N_5147,N_2134,N_2595);
and U5148 (N_5148,N_3560,N_2654);
nand U5149 (N_5149,N_2241,N_2893);
nand U5150 (N_5150,N_2305,N_3411);
xnor U5151 (N_5151,N_3842,N_3914);
nor U5152 (N_5152,N_3740,N_3552);
nor U5153 (N_5153,N_3011,N_3449);
or U5154 (N_5154,N_3829,N_2335);
xnor U5155 (N_5155,N_2202,N_3880);
or U5156 (N_5156,N_3615,N_2140);
nand U5157 (N_5157,N_2977,N_2774);
xnor U5158 (N_5158,N_3357,N_3540);
nor U5159 (N_5159,N_2500,N_2870);
xor U5160 (N_5160,N_3542,N_3974);
nor U5161 (N_5161,N_3148,N_3097);
or U5162 (N_5162,N_2303,N_2520);
nand U5163 (N_5163,N_3938,N_3086);
nor U5164 (N_5164,N_2980,N_2251);
or U5165 (N_5165,N_2581,N_3807);
or U5166 (N_5166,N_3685,N_2351);
or U5167 (N_5167,N_3241,N_3954);
nand U5168 (N_5168,N_3069,N_3946);
nor U5169 (N_5169,N_2859,N_2311);
xor U5170 (N_5170,N_3973,N_2499);
nor U5171 (N_5171,N_3888,N_3457);
nor U5172 (N_5172,N_2813,N_3691);
nand U5173 (N_5173,N_2869,N_3864);
or U5174 (N_5174,N_3968,N_3560);
or U5175 (N_5175,N_2668,N_2233);
xnor U5176 (N_5176,N_2860,N_3674);
and U5177 (N_5177,N_2557,N_2697);
nor U5178 (N_5178,N_2796,N_3551);
nand U5179 (N_5179,N_3641,N_3734);
nor U5180 (N_5180,N_3068,N_3293);
nor U5181 (N_5181,N_3592,N_2209);
and U5182 (N_5182,N_2511,N_2442);
or U5183 (N_5183,N_2645,N_3232);
and U5184 (N_5184,N_3197,N_2092);
nor U5185 (N_5185,N_3030,N_3171);
nor U5186 (N_5186,N_3811,N_2953);
and U5187 (N_5187,N_3373,N_2724);
nor U5188 (N_5188,N_3545,N_3482);
xor U5189 (N_5189,N_2273,N_2535);
nor U5190 (N_5190,N_3780,N_2439);
nand U5191 (N_5191,N_3436,N_2978);
xor U5192 (N_5192,N_3663,N_3314);
nor U5193 (N_5193,N_2527,N_2803);
or U5194 (N_5194,N_2436,N_3270);
nor U5195 (N_5195,N_3293,N_2824);
nand U5196 (N_5196,N_3647,N_3139);
xnor U5197 (N_5197,N_3928,N_3106);
nor U5198 (N_5198,N_3507,N_2283);
nor U5199 (N_5199,N_2145,N_3319);
nor U5200 (N_5200,N_2578,N_2309);
nand U5201 (N_5201,N_2503,N_2293);
or U5202 (N_5202,N_2382,N_3530);
and U5203 (N_5203,N_2316,N_2389);
and U5204 (N_5204,N_2867,N_2441);
nor U5205 (N_5205,N_2994,N_2208);
nand U5206 (N_5206,N_3156,N_3720);
and U5207 (N_5207,N_3954,N_2329);
xor U5208 (N_5208,N_3439,N_2111);
and U5209 (N_5209,N_3447,N_2383);
and U5210 (N_5210,N_3639,N_3410);
or U5211 (N_5211,N_3399,N_3373);
nor U5212 (N_5212,N_3639,N_3619);
nor U5213 (N_5213,N_3241,N_2822);
or U5214 (N_5214,N_3177,N_2659);
and U5215 (N_5215,N_2480,N_3973);
nor U5216 (N_5216,N_2099,N_3759);
and U5217 (N_5217,N_2057,N_2128);
nor U5218 (N_5218,N_2534,N_3032);
or U5219 (N_5219,N_3812,N_2321);
xnor U5220 (N_5220,N_2029,N_2517);
and U5221 (N_5221,N_2984,N_3852);
xor U5222 (N_5222,N_3842,N_2441);
or U5223 (N_5223,N_3862,N_3255);
or U5224 (N_5224,N_3912,N_3927);
or U5225 (N_5225,N_3114,N_2805);
nor U5226 (N_5226,N_3836,N_2616);
xor U5227 (N_5227,N_3469,N_3474);
nand U5228 (N_5228,N_3636,N_3136);
xor U5229 (N_5229,N_2602,N_3715);
or U5230 (N_5230,N_3278,N_3042);
nor U5231 (N_5231,N_3431,N_3784);
nor U5232 (N_5232,N_3534,N_2211);
nor U5233 (N_5233,N_2771,N_3555);
xor U5234 (N_5234,N_3334,N_3039);
or U5235 (N_5235,N_2750,N_2845);
nor U5236 (N_5236,N_2638,N_2560);
nor U5237 (N_5237,N_3639,N_3367);
and U5238 (N_5238,N_2875,N_3534);
xor U5239 (N_5239,N_2094,N_2234);
nand U5240 (N_5240,N_3749,N_2922);
or U5241 (N_5241,N_2276,N_3361);
or U5242 (N_5242,N_3096,N_2547);
nor U5243 (N_5243,N_2177,N_3327);
nor U5244 (N_5244,N_3418,N_3343);
or U5245 (N_5245,N_3158,N_3467);
and U5246 (N_5246,N_2675,N_3398);
and U5247 (N_5247,N_2311,N_3367);
and U5248 (N_5248,N_3979,N_2692);
nor U5249 (N_5249,N_2791,N_3459);
nor U5250 (N_5250,N_2443,N_2876);
nor U5251 (N_5251,N_2817,N_2777);
and U5252 (N_5252,N_3578,N_2627);
xor U5253 (N_5253,N_2639,N_2585);
nand U5254 (N_5254,N_2623,N_3935);
or U5255 (N_5255,N_2255,N_3590);
nand U5256 (N_5256,N_3752,N_3104);
nand U5257 (N_5257,N_2071,N_3263);
xnor U5258 (N_5258,N_2261,N_3622);
or U5259 (N_5259,N_2796,N_2728);
or U5260 (N_5260,N_2996,N_2965);
and U5261 (N_5261,N_2836,N_2648);
nor U5262 (N_5262,N_3367,N_2079);
nor U5263 (N_5263,N_3742,N_2072);
and U5264 (N_5264,N_3858,N_3112);
or U5265 (N_5265,N_2482,N_3680);
nand U5266 (N_5266,N_2735,N_3488);
nor U5267 (N_5267,N_3273,N_3011);
xor U5268 (N_5268,N_3658,N_2824);
nor U5269 (N_5269,N_3990,N_3829);
nand U5270 (N_5270,N_2402,N_3124);
xor U5271 (N_5271,N_3021,N_2747);
xnor U5272 (N_5272,N_3078,N_2755);
xnor U5273 (N_5273,N_3866,N_3701);
nand U5274 (N_5274,N_2011,N_3935);
nor U5275 (N_5275,N_3336,N_2385);
nand U5276 (N_5276,N_3739,N_2259);
nor U5277 (N_5277,N_3649,N_2045);
and U5278 (N_5278,N_2496,N_3039);
or U5279 (N_5279,N_3594,N_2689);
or U5280 (N_5280,N_3820,N_2466);
nor U5281 (N_5281,N_2517,N_2327);
xor U5282 (N_5282,N_3787,N_3893);
xor U5283 (N_5283,N_3053,N_2599);
nand U5284 (N_5284,N_3594,N_3995);
and U5285 (N_5285,N_3993,N_2444);
and U5286 (N_5286,N_2658,N_2547);
xnor U5287 (N_5287,N_2808,N_3732);
xnor U5288 (N_5288,N_3979,N_2516);
nor U5289 (N_5289,N_2236,N_2024);
nor U5290 (N_5290,N_2405,N_3983);
or U5291 (N_5291,N_2832,N_2333);
xnor U5292 (N_5292,N_2800,N_2967);
and U5293 (N_5293,N_3088,N_3433);
and U5294 (N_5294,N_3489,N_3183);
nand U5295 (N_5295,N_3573,N_2918);
nand U5296 (N_5296,N_3200,N_2806);
and U5297 (N_5297,N_2803,N_2643);
xor U5298 (N_5298,N_3344,N_2473);
and U5299 (N_5299,N_2401,N_2345);
nand U5300 (N_5300,N_3205,N_3857);
nand U5301 (N_5301,N_3440,N_2024);
nand U5302 (N_5302,N_3443,N_2801);
nand U5303 (N_5303,N_2801,N_3225);
nand U5304 (N_5304,N_2732,N_3837);
or U5305 (N_5305,N_3326,N_2064);
and U5306 (N_5306,N_2461,N_3738);
xor U5307 (N_5307,N_2435,N_3376);
nand U5308 (N_5308,N_3592,N_2534);
and U5309 (N_5309,N_2338,N_3242);
nand U5310 (N_5310,N_3124,N_2327);
or U5311 (N_5311,N_2703,N_3272);
nor U5312 (N_5312,N_2189,N_2345);
nor U5313 (N_5313,N_3817,N_3013);
xnor U5314 (N_5314,N_3105,N_3156);
nand U5315 (N_5315,N_3060,N_2807);
and U5316 (N_5316,N_2647,N_3482);
and U5317 (N_5317,N_3048,N_3832);
xor U5318 (N_5318,N_3975,N_3346);
and U5319 (N_5319,N_3461,N_3588);
or U5320 (N_5320,N_3660,N_2454);
xnor U5321 (N_5321,N_2335,N_3187);
nand U5322 (N_5322,N_3956,N_2775);
xnor U5323 (N_5323,N_2944,N_2260);
xor U5324 (N_5324,N_2385,N_2283);
and U5325 (N_5325,N_2291,N_3754);
nand U5326 (N_5326,N_3503,N_3516);
or U5327 (N_5327,N_2585,N_3830);
or U5328 (N_5328,N_3302,N_3830);
or U5329 (N_5329,N_2819,N_2830);
xor U5330 (N_5330,N_2995,N_2518);
xor U5331 (N_5331,N_3455,N_3740);
nand U5332 (N_5332,N_2803,N_3735);
or U5333 (N_5333,N_3981,N_3358);
nand U5334 (N_5334,N_3453,N_3674);
xor U5335 (N_5335,N_3814,N_3805);
nor U5336 (N_5336,N_3709,N_3938);
xnor U5337 (N_5337,N_3407,N_3400);
nor U5338 (N_5338,N_2027,N_3171);
nor U5339 (N_5339,N_3046,N_2399);
or U5340 (N_5340,N_3556,N_2580);
nand U5341 (N_5341,N_3018,N_3255);
nand U5342 (N_5342,N_3338,N_2616);
nor U5343 (N_5343,N_3820,N_2224);
nand U5344 (N_5344,N_2317,N_3494);
nand U5345 (N_5345,N_2359,N_3245);
and U5346 (N_5346,N_3837,N_2936);
and U5347 (N_5347,N_3772,N_2991);
nand U5348 (N_5348,N_2876,N_2818);
or U5349 (N_5349,N_3351,N_3286);
xnor U5350 (N_5350,N_2044,N_3140);
or U5351 (N_5351,N_3260,N_3668);
nand U5352 (N_5352,N_2398,N_3720);
or U5353 (N_5353,N_3164,N_2678);
nand U5354 (N_5354,N_2563,N_3936);
xor U5355 (N_5355,N_2480,N_3202);
xnor U5356 (N_5356,N_3501,N_2014);
nor U5357 (N_5357,N_3918,N_3490);
nand U5358 (N_5358,N_2372,N_3115);
or U5359 (N_5359,N_2188,N_2932);
xor U5360 (N_5360,N_2260,N_3907);
nand U5361 (N_5361,N_2592,N_3320);
and U5362 (N_5362,N_3250,N_2725);
xnor U5363 (N_5363,N_2237,N_2502);
xnor U5364 (N_5364,N_2562,N_3340);
xor U5365 (N_5365,N_3325,N_2845);
and U5366 (N_5366,N_2894,N_2156);
nand U5367 (N_5367,N_2526,N_3051);
xnor U5368 (N_5368,N_2588,N_3800);
nand U5369 (N_5369,N_2138,N_2994);
or U5370 (N_5370,N_2507,N_2694);
or U5371 (N_5371,N_2668,N_3628);
or U5372 (N_5372,N_2054,N_3807);
xnor U5373 (N_5373,N_3534,N_3887);
nor U5374 (N_5374,N_3997,N_2137);
xnor U5375 (N_5375,N_2591,N_2438);
xnor U5376 (N_5376,N_3068,N_3552);
or U5377 (N_5377,N_2975,N_3686);
nor U5378 (N_5378,N_3911,N_3862);
or U5379 (N_5379,N_2123,N_2703);
nand U5380 (N_5380,N_2245,N_2243);
nand U5381 (N_5381,N_2364,N_2523);
nor U5382 (N_5382,N_3510,N_3681);
xor U5383 (N_5383,N_2488,N_2991);
nor U5384 (N_5384,N_3398,N_3313);
nand U5385 (N_5385,N_2762,N_3958);
nor U5386 (N_5386,N_2260,N_2582);
nand U5387 (N_5387,N_3301,N_2204);
nand U5388 (N_5388,N_2147,N_2017);
or U5389 (N_5389,N_3230,N_2350);
xor U5390 (N_5390,N_3095,N_2105);
xor U5391 (N_5391,N_3934,N_2651);
nor U5392 (N_5392,N_2524,N_2888);
and U5393 (N_5393,N_3640,N_3273);
nand U5394 (N_5394,N_2403,N_2115);
and U5395 (N_5395,N_3488,N_2949);
and U5396 (N_5396,N_2844,N_3555);
xor U5397 (N_5397,N_2695,N_3583);
nor U5398 (N_5398,N_3442,N_3459);
nor U5399 (N_5399,N_3426,N_3814);
nor U5400 (N_5400,N_3884,N_3070);
nor U5401 (N_5401,N_3492,N_3531);
nand U5402 (N_5402,N_2806,N_2748);
nand U5403 (N_5403,N_3568,N_3942);
nor U5404 (N_5404,N_3810,N_2724);
nand U5405 (N_5405,N_3746,N_2707);
xnor U5406 (N_5406,N_3470,N_3182);
xor U5407 (N_5407,N_3430,N_3820);
nor U5408 (N_5408,N_3602,N_3435);
nand U5409 (N_5409,N_2805,N_2603);
and U5410 (N_5410,N_2308,N_3468);
xnor U5411 (N_5411,N_2542,N_2208);
or U5412 (N_5412,N_2113,N_3453);
xnor U5413 (N_5413,N_3137,N_3446);
and U5414 (N_5414,N_2432,N_3192);
or U5415 (N_5415,N_2289,N_2061);
and U5416 (N_5416,N_3036,N_3575);
nor U5417 (N_5417,N_2699,N_2214);
nor U5418 (N_5418,N_2175,N_3451);
nand U5419 (N_5419,N_3446,N_2993);
xor U5420 (N_5420,N_2123,N_3260);
or U5421 (N_5421,N_2317,N_3172);
nor U5422 (N_5422,N_2508,N_2361);
xor U5423 (N_5423,N_2546,N_3671);
or U5424 (N_5424,N_2736,N_3990);
xnor U5425 (N_5425,N_3850,N_3764);
nor U5426 (N_5426,N_3144,N_3278);
or U5427 (N_5427,N_2951,N_3428);
or U5428 (N_5428,N_2573,N_2954);
nor U5429 (N_5429,N_2445,N_2141);
and U5430 (N_5430,N_2326,N_2107);
or U5431 (N_5431,N_2454,N_3708);
and U5432 (N_5432,N_2550,N_2924);
xnor U5433 (N_5433,N_3893,N_3549);
nand U5434 (N_5434,N_3634,N_3720);
or U5435 (N_5435,N_2878,N_2338);
or U5436 (N_5436,N_2287,N_3222);
xor U5437 (N_5437,N_2659,N_3770);
or U5438 (N_5438,N_3712,N_2290);
and U5439 (N_5439,N_2921,N_3109);
or U5440 (N_5440,N_2926,N_3256);
nor U5441 (N_5441,N_2709,N_3414);
xor U5442 (N_5442,N_2689,N_2838);
xnor U5443 (N_5443,N_2817,N_2533);
xnor U5444 (N_5444,N_3581,N_3440);
or U5445 (N_5445,N_3432,N_2752);
and U5446 (N_5446,N_2735,N_2137);
and U5447 (N_5447,N_3969,N_2814);
or U5448 (N_5448,N_3395,N_2829);
xnor U5449 (N_5449,N_3004,N_3056);
xor U5450 (N_5450,N_2754,N_3503);
and U5451 (N_5451,N_3987,N_3914);
nor U5452 (N_5452,N_2939,N_3972);
nand U5453 (N_5453,N_3699,N_2519);
or U5454 (N_5454,N_3372,N_3812);
nand U5455 (N_5455,N_3868,N_3623);
xor U5456 (N_5456,N_2520,N_3002);
or U5457 (N_5457,N_3668,N_2690);
xnor U5458 (N_5458,N_3765,N_3130);
xor U5459 (N_5459,N_2395,N_2239);
xnor U5460 (N_5460,N_2673,N_2581);
and U5461 (N_5461,N_2642,N_3897);
nor U5462 (N_5462,N_2607,N_3922);
and U5463 (N_5463,N_2842,N_2944);
nand U5464 (N_5464,N_3489,N_2497);
and U5465 (N_5465,N_3021,N_2081);
xor U5466 (N_5466,N_2701,N_2277);
nand U5467 (N_5467,N_2292,N_3442);
xnor U5468 (N_5468,N_3251,N_3896);
nor U5469 (N_5469,N_3513,N_2301);
nor U5470 (N_5470,N_2760,N_3174);
nand U5471 (N_5471,N_2244,N_2375);
xnor U5472 (N_5472,N_3004,N_2406);
or U5473 (N_5473,N_2324,N_3024);
or U5474 (N_5474,N_2006,N_2069);
nor U5475 (N_5475,N_3473,N_3872);
or U5476 (N_5476,N_3802,N_2474);
nor U5477 (N_5477,N_3642,N_2465);
nor U5478 (N_5478,N_2326,N_3173);
nor U5479 (N_5479,N_3303,N_3972);
and U5480 (N_5480,N_2147,N_3634);
xnor U5481 (N_5481,N_2065,N_3890);
or U5482 (N_5482,N_2756,N_3729);
nor U5483 (N_5483,N_2921,N_3901);
nor U5484 (N_5484,N_2667,N_3855);
and U5485 (N_5485,N_2574,N_2324);
nand U5486 (N_5486,N_3544,N_3414);
xor U5487 (N_5487,N_3012,N_3387);
nand U5488 (N_5488,N_3850,N_2795);
or U5489 (N_5489,N_2167,N_2966);
xor U5490 (N_5490,N_2559,N_3409);
or U5491 (N_5491,N_3727,N_2816);
or U5492 (N_5492,N_3766,N_2547);
xnor U5493 (N_5493,N_2007,N_3698);
xor U5494 (N_5494,N_3174,N_3437);
and U5495 (N_5495,N_2892,N_3380);
or U5496 (N_5496,N_3309,N_2977);
xnor U5497 (N_5497,N_3096,N_3953);
xor U5498 (N_5498,N_2683,N_3212);
or U5499 (N_5499,N_3330,N_3064);
and U5500 (N_5500,N_2647,N_3964);
or U5501 (N_5501,N_2698,N_3440);
nand U5502 (N_5502,N_2810,N_3604);
or U5503 (N_5503,N_2188,N_2178);
nor U5504 (N_5504,N_2492,N_2372);
nor U5505 (N_5505,N_2427,N_2325);
and U5506 (N_5506,N_2622,N_2736);
or U5507 (N_5507,N_2918,N_2087);
and U5508 (N_5508,N_2232,N_3903);
nor U5509 (N_5509,N_3798,N_2003);
nand U5510 (N_5510,N_3454,N_3334);
xor U5511 (N_5511,N_3283,N_3428);
nand U5512 (N_5512,N_3004,N_2510);
or U5513 (N_5513,N_3321,N_2234);
or U5514 (N_5514,N_2991,N_2045);
xnor U5515 (N_5515,N_3464,N_2435);
nand U5516 (N_5516,N_3448,N_2695);
nand U5517 (N_5517,N_3096,N_2334);
nor U5518 (N_5518,N_3250,N_3299);
nand U5519 (N_5519,N_3339,N_3701);
and U5520 (N_5520,N_2815,N_3354);
nor U5521 (N_5521,N_3628,N_3796);
xnor U5522 (N_5522,N_2503,N_3897);
and U5523 (N_5523,N_3901,N_2982);
nand U5524 (N_5524,N_3214,N_2614);
xnor U5525 (N_5525,N_2924,N_2202);
or U5526 (N_5526,N_3016,N_3996);
xor U5527 (N_5527,N_2873,N_2135);
nor U5528 (N_5528,N_2163,N_3029);
nor U5529 (N_5529,N_3031,N_2632);
xor U5530 (N_5530,N_2294,N_2473);
nor U5531 (N_5531,N_2334,N_2698);
nand U5532 (N_5532,N_3279,N_2562);
or U5533 (N_5533,N_3375,N_2964);
nand U5534 (N_5534,N_3489,N_3517);
or U5535 (N_5535,N_2519,N_3723);
nand U5536 (N_5536,N_2526,N_2942);
xor U5537 (N_5537,N_2669,N_3388);
xor U5538 (N_5538,N_2752,N_3449);
nor U5539 (N_5539,N_2508,N_2595);
nor U5540 (N_5540,N_2617,N_3693);
and U5541 (N_5541,N_3091,N_2690);
nand U5542 (N_5542,N_3637,N_2037);
or U5543 (N_5543,N_2111,N_2724);
xor U5544 (N_5544,N_3550,N_2855);
or U5545 (N_5545,N_3260,N_3323);
or U5546 (N_5546,N_3421,N_2467);
and U5547 (N_5547,N_3056,N_2785);
nor U5548 (N_5548,N_2877,N_3489);
nand U5549 (N_5549,N_2327,N_3132);
nor U5550 (N_5550,N_2096,N_3837);
nor U5551 (N_5551,N_3267,N_3780);
and U5552 (N_5552,N_3308,N_2120);
or U5553 (N_5553,N_2418,N_3230);
and U5554 (N_5554,N_3406,N_2894);
and U5555 (N_5555,N_3327,N_3280);
or U5556 (N_5556,N_2677,N_3497);
xor U5557 (N_5557,N_2089,N_3477);
nor U5558 (N_5558,N_2158,N_2872);
or U5559 (N_5559,N_2941,N_3094);
nor U5560 (N_5560,N_2858,N_2927);
nand U5561 (N_5561,N_3917,N_2949);
and U5562 (N_5562,N_3229,N_3210);
and U5563 (N_5563,N_2869,N_3942);
nor U5564 (N_5564,N_2523,N_3092);
nor U5565 (N_5565,N_3659,N_2735);
and U5566 (N_5566,N_3563,N_2958);
and U5567 (N_5567,N_3528,N_3447);
nand U5568 (N_5568,N_3851,N_2738);
nor U5569 (N_5569,N_3880,N_3923);
xnor U5570 (N_5570,N_2974,N_3400);
xnor U5571 (N_5571,N_2931,N_2661);
nor U5572 (N_5572,N_2780,N_2869);
xnor U5573 (N_5573,N_3046,N_2424);
and U5574 (N_5574,N_2089,N_2120);
nor U5575 (N_5575,N_2994,N_3719);
nand U5576 (N_5576,N_3184,N_3608);
nor U5577 (N_5577,N_3671,N_3897);
and U5578 (N_5578,N_3089,N_3975);
and U5579 (N_5579,N_2827,N_2373);
nor U5580 (N_5580,N_2450,N_3484);
and U5581 (N_5581,N_3295,N_3490);
or U5582 (N_5582,N_3785,N_3854);
and U5583 (N_5583,N_3513,N_2068);
nor U5584 (N_5584,N_3333,N_2081);
nand U5585 (N_5585,N_2404,N_3886);
nor U5586 (N_5586,N_2530,N_2762);
or U5587 (N_5587,N_2776,N_2750);
nand U5588 (N_5588,N_2129,N_3683);
xnor U5589 (N_5589,N_3535,N_3418);
nor U5590 (N_5590,N_3445,N_2935);
xnor U5591 (N_5591,N_3835,N_2188);
or U5592 (N_5592,N_2322,N_3770);
nor U5593 (N_5593,N_2043,N_2576);
or U5594 (N_5594,N_3073,N_3865);
nor U5595 (N_5595,N_3898,N_3367);
nand U5596 (N_5596,N_3850,N_2360);
xnor U5597 (N_5597,N_2146,N_3751);
or U5598 (N_5598,N_3686,N_3718);
nand U5599 (N_5599,N_2610,N_3506);
xnor U5600 (N_5600,N_2341,N_2174);
xor U5601 (N_5601,N_2868,N_3816);
nor U5602 (N_5602,N_2911,N_2374);
nand U5603 (N_5603,N_3336,N_3299);
nor U5604 (N_5604,N_2289,N_3005);
or U5605 (N_5605,N_2095,N_2706);
nand U5606 (N_5606,N_3432,N_2054);
nand U5607 (N_5607,N_2858,N_3030);
and U5608 (N_5608,N_2694,N_3018);
nor U5609 (N_5609,N_3145,N_3897);
nor U5610 (N_5610,N_3874,N_2109);
nand U5611 (N_5611,N_2882,N_3208);
xor U5612 (N_5612,N_3306,N_3209);
xnor U5613 (N_5613,N_3325,N_3106);
nor U5614 (N_5614,N_2688,N_3717);
nand U5615 (N_5615,N_2976,N_3888);
nand U5616 (N_5616,N_2894,N_2221);
nor U5617 (N_5617,N_3121,N_3740);
xor U5618 (N_5618,N_3821,N_2292);
xor U5619 (N_5619,N_2007,N_2457);
and U5620 (N_5620,N_2395,N_2347);
or U5621 (N_5621,N_3043,N_3868);
nand U5622 (N_5622,N_2486,N_2091);
or U5623 (N_5623,N_2819,N_2746);
and U5624 (N_5624,N_2012,N_2495);
nand U5625 (N_5625,N_2704,N_2363);
xor U5626 (N_5626,N_2296,N_2193);
nor U5627 (N_5627,N_2957,N_3468);
nor U5628 (N_5628,N_2144,N_2515);
or U5629 (N_5629,N_2290,N_2910);
or U5630 (N_5630,N_2995,N_3024);
and U5631 (N_5631,N_2132,N_2907);
nand U5632 (N_5632,N_3479,N_3060);
nor U5633 (N_5633,N_3086,N_3100);
nand U5634 (N_5634,N_2786,N_2344);
xnor U5635 (N_5635,N_2360,N_2735);
nor U5636 (N_5636,N_2693,N_2041);
xor U5637 (N_5637,N_3507,N_2267);
and U5638 (N_5638,N_2081,N_2664);
nand U5639 (N_5639,N_3489,N_2402);
nand U5640 (N_5640,N_2300,N_3620);
nor U5641 (N_5641,N_2852,N_3122);
nand U5642 (N_5642,N_2588,N_2969);
nand U5643 (N_5643,N_3253,N_2073);
and U5644 (N_5644,N_3961,N_2679);
and U5645 (N_5645,N_2493,N_3451);
xor U5646 (N_5646,N_3576,N_2062);
and U5647 (N_5647,N_2674,N_3984);
or U5648 (N_5648,N_3301,N_2661);
or U5649 (N_5649,N_2815,N_3166);
or U5650 (N_5650,N_3988,N_3855);
xnor U5651 (N_5651,N_2547,N_2791);
nor U5652 (N_5652,N_3150,N_2625);
nor U5653 (N_5653,N_3573,N_3724);
nor U5654 (N_5654,N_2154,N_3753);
nor U5655 (N_5655,N_2184,N_2238);
nand U5656 (N_5656,N_2643,N_3910);
and U5657 (N_5657,N_2211,N_3654);
nor U5658 (N_5658,N_3572,N_3752);
and U5659 (N_5659,N_3776,N_2769);
or U5660 (N_5660,N_2852,N_2478);
nand U5661 (N_5661,N_3066,N_2916);
or U5662 (N_5662,N_3986,N_2178);
nand U5663 (N_5663,N_2784,N_3049);
nor U5664 (N_5664,N_3245,N_3713);
or U5665 (N_5665,N_3122,N_2964);
or U5666 (N_5666,N_2676,N_3017);
nand U5667 (N_5667,N_3468,N_2307);
or U5668 (N_5668,N_3309,N_2684);
or U5669 (N_5669,N_3741,N_2841);
or U5670 (N_5670,N_2188,N_3607);
or U5671 (N_5671,N_2406,N_3887);
nand U5672 (N_5672,N_2615,N_3746);
or U5673 (N_5673,N_3892,N_3352);
nor U5674 (N_5674,N_2159,N_2263);
nor U5675 (N_5675,N_2233,N_2020);
or U5676 (N_5676,N_3106,N_2236);
or U5677 (N_5677,N_2956,N_3642);
xnor U5678 (N_5678,N_2082,N_2157);
xnor U5679 (N_5679,N_2592,N_2638);
nor U5680 (N_5680,N_2886,N_3748);
or U5681 (N_5681,N_2732,N_3218);
xor U5682 (N_5682,N_2633,N_2097);
nor U5683 (N_5683,N_2068,N_2353);
and U5684 (N_5684,N_3182,N_3200);
nand U5685 (N_5685,N_2952,N_2056);
nor U5686 (N_5686,N_2505,N_2660);
nand U5687 (N_5687,N_3422,N_2309);
and U5688 (N_5688,N_3530,N_3351);
nor U5689 (N_5689,N_3025,N_3264);
and U5690 (N_5690,N_2876,N_2039);
or U5691 (N_5691,N_2365,N_2785);
nand U5692 (N_5692,N_3972,N_3809);
xnor U5693 (N_5693,N_2636,N_2397);
nand U5694 (N_5694,N_2478,N_3326);
xor U5695 (N_5695,N_3988,N_3986);
xor U5696 (N_5696,N_3458,N_3360);
nor U5697 (N_5697,N_3620,N_2897);
xnor U5698 (N_5698,N_2240,N_2452);
xor U5699 (N_5699,N_3354,N_2339);
and U5700 (N_5700,N_2478,N_2737);
nand U5701 (N_5701,N_2271,N_3439);
nand U5702 (N_5702,N_2646,N_3488);
and U5703 (N_5703,N_3654,N_3586);
and U5704 (N_5704,N_2409,N_2693);
and U5705 (N_5705,N_3557,N_3576);
nor U5706 (N_5706,N_2946,N_3573);
and U5707 (N_5707,N_3237,N_3987);
nor U5708 (N_5708,N_3686,N_3335);
nor U5709 (N_5709,N_3518,N_2278);
nand U5710 (N_5710,N_3712,N_3130);
and U5711 (N_5711,N_2879,N_2844);
or U5712 (N_5712,N_2611,N_3396);
xor U5713 (N_5713,N_3264,N_2673);
and U5714 (N_5714,N_2467,N_3311);
xor U5715 (N_5715,N_3252,N_3459);
or U5716 (N_5716,N_2592,N_3078);
or U5717 (N_5717,N_2505,N_3464);
and U5718 (N_5718,N_2203,N_3466);
or U5719 (N_5719,N_3190,N_3953);
xor U5720 (N_5720,N_2158,N_3528);
or U5721 (N_5721,N_3779,N_2919);
xor U5722 (N_5722,N_2845,N_2025);
nor U5723 (N_5723,N_2648,N_3760);
xnor U5724 (N_5724,N_2766,N_3910);
nor U5725 (N_5725,N_2854,N_2427);
nand U5726 (N_5726,N_3151,N_2138);
nor U5727 (N_5727,N_3953,N_3502);
nand U5728 (N_5728,N_3797,N_3593);
nor U5729 (N_5729,N_3293,N_2488);
nand U5730 (N_5730,N_2740,N_3995);
nor U5731 (N_5731,N_3630,N_2095);
nor U5732 (N_5732,N_2257,N_2265);
and U5733 (N_5733,N_3581,N_2854);
and U5734 (N_5734,N_3148,N_2840);
nor U5735 (N_5735,N_3566,N_3647);
or U5736 (N_5736,N_2393,N_3535);
nor U5737 (N_5737,N_2533,N_3682);
nor U5738 (N_5738,N_3771,N_3545);
nand U5739 (N_5739,N_3746,N_2259);
xnor U5740 (N_5740,N_3577,N_3224);
xor U5741 (N_5741,N_3629,N_3290);
and U5742 (N_5742,N_3334,N_3846);
xor U5743 (N_5743,N_3772,N_2065);
xor U5744 (N_5744,N_2227,N_3011);
nor U5745 (N_5745,N_2284,N_2001);
nor U5746 (N_5746,N_3592,N_3233);
xor U5747 (N_5747,N_3015,N_3163);
nand U5748 (N_5748,N_3337,N_2582);
nand U5749 (N_5749,N_2677,N_2948);
xnor U5750 (N_5750,N_3303,N_3270);
or U5751 (N_5751,N_3904,N_2908);
nand U5752 (N_5752,N_3321,N_3796);
and U5753 (N_5753,N_2132,N_2484);
and U5754 (N_5754,N_2452,N_3131);
and U5755 (N_5755,N_2734,N_2239);
and U5756 (N_5756,N_3245,N_3797);
or U5757 (N_5757,N_2246,N_2457);
nand U5758 (N_5758,N_3371,N_2955);
or U5759 (N_5759,N_2456,N_2111);
nand U5760 (N_5760,N_3132,N_3603);
xnor U5761 (N_5761,N_2473,N_3716);
xor U5762 (N_5762,N_3034,N_2511);
xor U5763 (N_5763,N_2686,N_2969);
nand U5764 (N_5764,N_3759,N_2920);
and U5765 (N_5765,N_3685,N_3014);
or U5766 (N_5766,N_2960,N_2607);
xnor U5767 (N_5767,N_3076,N_2622);
nor U5768 (N_5768,N_3658,N_2445);
or U5769 (N_5769,N_2317,N_3148);
and U5770 (N_5770,N_3498,N_2674);
nand U5771 (N_5771,N_3538,N_2102);
and U5772 (N_5772,N_3514,N_2894);
or U5773 (N_5773,N_2635,N_3458);
nor U5774 (N_5774,N_3924,N_3008);
nor U5775 (N_5775,N_2022,N_2036);
nand U5776 (N_5776,N_2612,N_2207);
xor U5777 (N_5777,N_3159,N_2051);
nor U5778 (N_5778,N_3689,N_2318);
and U5779 (N_5779,N_3201,N_2365);
xnor U5780 (N_5780,N_2378,N_3108);
or U5781 (N_5781,N_2073,N_3872);
nand U5782 (N_5782,N_2287,N_3625);
xnor U5783 (N_5783,N_2051,N_2918);
nand U5784 (N_5784,N_3291,N_3440);
nor U5785 (N_5785,N_3167,N_3464);
nand U5786 (N_5786,N_3782,N_2833);
xnor U5787 (N_5787,N_3188,N_3901);
or U5788 (N_5788,N_2559,N_3217);
xnor U5789 (N_5789,N_2489,N_2351);
or U5790 (N_5790,N_2186,N_3291);
or U5791 (N_5791,N_2098,N_3339);
and U5792 (N_5792,N_3438,N_3160);
xnor U5793 (N_5793,N_3683,N_2565);
nand U5794 (N_5794,N_2851,N_3075);
xor U5795 (N_5795,N_3781,N_2600);
nand U5796 (N_5796,N_3317,N_3369);
nor U5797 (N_5797,N_2539,N_3783);
nand U5798 (N_5798,N_2737,N_2072);
nor U5799 (N_5799,N_2431,N_2271);
or U5800 (N_5800,N_2053,N_2844);
xor U5801 (N_5801,N_2411,N_3120);
nor U5802 (N_5802,N_2450,N_3251);
nand U5803 (N_5803,N_2397,N_2105);
and U5804 (N_5804,N_3917,N_3148);
or U5805 (N_5805,N_3205,N_3374);
nand U5806 (N_5806,N_3148,N_3140);
xnor U5807 (N_5807,N_2979,N_3389);
or U5808 (N_5808,N_3310,N_2558);
and U5809 (N_5809,N_3512,N_2980);
xnor U5810 (N_5810,N_2102,N_3142);
nand U5811 (N_5811,N_3810,N_2285);
and U5812 (N_5812,N_3723,N_3602);
and U5813 (N_5813,N_2499,N_2332);
xor U5814 (N_5814,N_3183,N_3604);
nor U5815 (N_5815,N_2546,N_3455);
nand U5816 (N_5816,N_2026,N_2740);
xor U5817 (N_5817,N_2330,N_2754);
nand U5818 (N_5818,N_3206,N_3901);
and U5819 (N_5819,N_3172,N_2154);
xor U5820 (N_5820,N_2007,N_3119);
xnor U5821 (N_5821,N_2282,N_2253);
nand U5822 (N_5822,N_2199,N_2698);
or U5823 (N_5823,N_3386,N_2224);
xnor U5824 (N_5824,N_2120,N_2351);
and U5825 (N_5825,N_2042,N_3633);
nor U5826 (N_5826,N_3679,N_2353);
nor U5827 (N_5827,N_2755,N_3617);
nand U5828 (N_5828,N_2816,N_2000);
and U5829 (N_5829,N_2683,N_2179);
xnor U5830 (N_5830,N_3050,N_2462);
nor U5831 (N_5831,N_3027,N_2963);
xnor U5832 (N_5832,N_3633,N_2479);
or U5833 (N_5833,N_3166,N_2856);
nor U5834 (N_5834,N_2765,N_3665);
or U5835 (N_5835,N_3183,N_3156);
nor U5836 (N_5836,N_3030,N_2875);
xor U5837 (N_5837,N_3816,N_2159);
and U5838 (N_5838,N_2610,N_2462);
and U5839 (N_5839,N_3922,N_3896);
nand U5840 (N_5840,N_2716,N_3524);
xor U5841 (N_5841,N_2724,N_2082);
and U5842 (N_5842,N_2924,N_3820);
nand U5843 (N_5843,N_2793,N_3912);
nor U5844 (N_5844,N_3774,N_3734);
xor U5845 (N_5845,N_2737,N_2793);
or U5846 (N_5846,N_3346,N_3668);
xnor U5847 (N_5847,N_2734,N_2430);
or U5848 (N_5848,N_3077,N_2590);
nand U5849 (N_5849,N_3243,N_2851);
and U5850 (N_5850,N_2499,N_3805);
or U5851 (N_5851,N_2492,N_3643);
and U5852 (N_5852,N_3947,N_3476);
nor U5853 (N_5853,N_3932,N_3070);
nand U5854 (N_5854,N_2093,N_2935);
or U5855 (N_5855,N_2304,N_3807);
and U5856 (N_5856,N_3558,N_2255);
nand U5857 (N_5857,N_3739,N_2046);
or U5858 (N_5858,N_2615,N_2522);
or U5859 (N_5859,N_3047,N_3223);
xor U5860 (N_5860,N_2402,N_3532);
and U5861 (N_5861,N_3570,N_3468);
xor U5862 (N_5862,N_3318,N_2502);
or U5863 (N_5863,N_2917,N_2210);
xnor U5864 (N_5864,N_2219,N_2105);
nand U5865 (N_5865,N_2701,N_2030);
xor U5866 (N_5866,N_3966,N_2651);
and U5867 (N_5867,N_3834,N_3111);
or U5868 (N_5868,N_3509,N_3736);
nand U5869 (N_5869,N_2496,N_2937);
nand U5870 (N_5870,N_2465,N_3849);
nand U5871 (N_5871,N_2039,N_2974);
and U5872 (N_5872,N_3982,N_3709);
or U5873 (N_5873,N_3823,N_3305);
and U5874 (N_5874,N_2110,N_3506);
nor U5875 (N_5875,N_2710,N_3757);
xor U5876 (N_5876,N_2987,N_3576);
nand U5877 (N_5877,N_3112,N_3560);
xnor U5878 (N_5878,N_3970,N_2688);
nor U5879 (N_5879,N_3356,N_3434);
nand U5880 (N_5880,N_2439,N_2708);
and U5881 (N_5881,N_3058,N_3459);
nor U5882 (N_5882,N_2668,N_2104);
xnor U5883 (N_5883,N_3287,N_2735);
nand U5884 (N_5884,N_3099,N_3296);
xnor U5885 (N_5885,N_2840,N_3036);
or U5886 (N_5886,N_2619,N_2498);
xnor U5887 (N_5887,N_2975,N_2486);
xnor U5888 (N_5888,N_3632,N_3025);
or U5889 (N_5889,N_3327,N_2994);
nand U5890 (N_5890,N_2252,N_2109);
or U5891 (N_5891,N_2577,N_3141);
and U5892 (N_5892,N_2010,N_3768);
nand U5893 (N_5893,N_2452,N_3974);
nor U5894 (N_5894,N_2938,N_2822);
or U5895 (N_5895,N_3622,N_3615);
nor U5896 (N_5896,N_2904,N_3715);
nand U5897 (N_5897,N_2710,N_3701);
and U5898 (N_5898,N_3843,N_2431);
or U5899 (N_5899,N_2990,N_2679);
nor U5900 (N_5900,N_2746,N_2146);
nand U5901 (N_5901,N_3868,N_3972);
or U5902 (N_5902,N_3312,N_2506);
nor U5903 (N_5903,N_2112,N_3728);
or U5904 (N_5904,N_3489,N_2964);
nor U5905 (N_5905,N_2457,N_3088);
or U5906 (N_5906,N_2433,N_2556);
nand U5907 (N_5907,N_3737,N_3232);
nor U5908 (N_5908,N_2378,N_3643);
nor U5909 (N_5909,N_2348,N_2656);
and U5910 (N_5910,N_3976,N_3509);
nor U5911 (N_5911,N_2571,N_3458);
nor U5912 (N_5912,N_2668,N_3607);
and U5913 (N_5913,N_2907,N_2323);
or U5914 (N_5914,N_3011,N_2590);
nand U5915 (N_5915,N_2554,N_2166);
xor U5916 (N_5916,N_2593,N_2872);
or U5917 (N_5917,N_2908,N_2570);
xor U5918 (N_5918,N_2276,N_3841);
and U5919 (N_5919,N_3964,N_3268);
or U5920 (N_5920,N_2641,N_3770);
xnor U5921 (N_5921,N_2763,N_3407);
nor U5922 (N_5922,N_2184,N_3719);
and U5923 (N_5923,N_3128,N_3547);
xnor U5924 (N_5924,N_3100,N_3601);
nor U5925 (N_5925,N_3148,N_2563);
nand U5926 (N_5926,N_2808,N_2949);
xnor U5927 (N_5927,N_2436,N_2630);
nor U5928 (N_5928,N_3046,N_2026);
xor U5929 (N_5929,N_2157,N_3951);
xnor U5930 (N_5930,N_2018,N_2012);
xnor U5931 (N_5931,N_2516,N_2331);
or U5932 (N_5932,N_3381,N_3218);
and U5933 (N_5933,N_2833,N_2526);
nand U5934 (N_5934,N_2216,N_2227);
nor U5935 (N_5935,N_2875,N_2713);
nor U5936 (N_5936,N_2615,N_2255);
and U5937 (N_5937,N_3487,N_3327);
nor U5938 (N_5938,N_2238,N_3975);
xnor U5939 (N_5939,N_2581,N_2525);
or U5940 (N_5940,N_2696,N_3379);
and U5941 (N_5941,N_2907,N_2540);
and U5942 (N_5942,N_3375,N_2906);
xor U5943 (N_5943,N_3841,N_3896);
or U5944 (N_5944,N_2345,N_2000);
or U5945 (N_5945,N_2446,N_3024);
nand U5946 (N_5946,N_2470,N_2692);
and U5947 (N_5947,N_2553,N_2812);
nand U5948 (N_5948,N_2389,N_3426);
or U5949 (N_5949,N_2550,N_3040);
or U5950 (N_5950,N_2514,N_2820);
xor U5951 (N_5951,N_2969,N_2498);
xor U5952 (N_5952,N_3023,N_2099);
nor U5953 (N_5953,N_3644,N_3097);
xnor U5954 (N_5954,N_2730,N_3117);
nand U5955 (N_5955,N_2054,N_2404);
or U5956 (N_5956,N_3085,N_2742);
nor U5957 (N_5957,N_3125,N_3017);
nor U5958 (N_5958,N_3232,N_3858);
nor U5959 (N_5959,N_2556,N_3334);
nor U5960 (N_5960,N_2489,N_3779);
and U5961 (N_5961,N_3903,N_2774);
nand U5962 (N_5962,N_2902,N_2760);
nand U5963 (N_5963,N_2813,N_2655);
nand U5964 (N_5964,N_2257,N_2762);
nor U5965 (N_5965,N_3020,N_3479);
and U5966 (N_5966,N_3275,N_3656);
xor U5967 (N_5967,N_2561,N_3133);
nand U5968 (N_5968,N_3288,N_2941);
or U5969 (N_5969,N_3279,N_3468);
and U5970 (N_5970,N_2998,N_2375);
nand U5971 (N_5971,N_2363,N_2763);
xnor U5972 (N_5972,N_2737,N_2432);
nor U5973 (N_5973,N_3741,N_3657);
nor U5974 (N_5974,N_3916,N_3945);
xnor U5975 (N_5975,N_2325,N_2602);
xor U5976 (N_5976,N_3792,N_3520);
nor U5977 (N_5977,N_3316,N_2291);
nor U5978 (N_5978,N_2357,N_3505);
xor U5979 (N_5979,N_3784,N_2230);
and U5980 (N_5980,N_3521,N_2954);
nand U5981 (N_5981,N_2513,N_2665);
nand U5982 (N_5982,N_2568,N_2459);
or U5983 (N_5983,N_2040,N_3723);
and U5984 (N_5984,N_3509,N_3960);
or U5985 (N_5985,N_2778,N_2079);
or U5986 (N_5986,N_3385,N_3011);
nand U5987 (N_5987,N_2936,N_2040);
xor U5988 (N_5988,N_3286,N_2170);
nand U5989 (N_5989,N_3174,N_3937);
nor U5990 (N_5990,N_2087,N_2695);
nor U5991 (N_5991,N_3899,N_2563);
xnor U5992 (N_5992,N_2111,N_3105);
nor U5993 (N_5993,N_2634,N_2337);
xor U5994 (N_5994,N_2186,N_2488);
xor U5995 (N_5995,N_3372,N_3760);
nand U5996 (N_5996,N_3229,N_3938);
or U5997 (N_5997,N_3198,N_3133);
or U5998 (N_5998,N_2012,N_3990);
nand U5999 (N_5999,N_3666,N_2725);
xnor U6000 (N_6000,N_5337,N_5628);
xor U6001 (N_6001,N_4413,N_5631);
xnor U6002 (N_6002,N_5253,N_5466);
nand U6003 (N_6003,N_4454,N_5285);
nand U6004 (N_6004,N_5187,N_4075);
xnor U6005 (N_6005,N_4110,N_5735);
nand U6006 (N_6006,N_4305,N_5299);
nor U6007 (N_6007,N_4577,N_4743);
and U6008 (N_6008,N_5484,N_4631);
or U6009 (N_6009,N_5852,N_5641);
and U6010 (N_6010,N_5159,N_5661);
xnor U6011 (N_6011,N_5806,N_5205);
and U6012 (N_6012,N_5600,N_5164);
or U6013 (N_6013,N_5987,N_5734);
nor U6014 (N_6014,N_5040,N_5390);
or U6015 (N_6015,N_5448,N_4938);
or U6016 (N_6016,N_4544,N_5167);
or U6017 (N_6017,N_5956,N_5842);
xor U6018 (N_6018,N_4490,N_4291);
and U6019 (N_6019,N_4258,N_5589);
nor U6020 (N_6020,N_4031,N_4330);
nor U6021 (N_6021,N_5787,N_4590);
xor U6022 (N_6022,N_4396,N_4777);
nand U6023 (N_6023,N_4340,N_5036);
nand U6024 (N_6024,N_4520,N_5217);
nor U6025 (N_6025,N_4083,N_4939);
nor U6026 (N_6026,N_4072,N_4355);
xnor U6027 (N_6027,N_4346,N_5720);
or U6028 (N_6028,N_4232,N_5096);
nor U6029 (N_6029,N_4806,N_4391);
nand U6030 (N_6030,N_5612,N_5312);
xnor U6031 (N_6031,N_4662,N_5882);
nor U6032 (N_6032,N_5634,N_4036);
and U6033 (N_6033,N_5707,N_5537);
or U6034 (N_6034,N_4090,N_5408);
nand U6035 (N_6035,N_5302,N_4148);
nor U6036 (N_6036,N_4261,N_5026);
and U6037 (N_6037,N_4143,N_4804);
and U6038 (N_6038,N_5608,N_4485);
nor U6039 (N_6039,N_4989,N_5913);
nand U6040 (N_6040,N_5199,N_4023);
or U6041 (N_6041,N_5982,N_4648);
nand U6042 (N_6042,N_5535,N_4367);
and U6043 (N_6043,N_4913,N_5386);
or U6044 (N_6044,N_5581,N_5170);
nor U6045 (N_6045,N_4762,N_4280);
xnor U6046 (N_6046,N_5635,N_5498);
nand U6047 (N_6047,N_4242,N_5795);
and U6048 (N_6048,N_5186,N_4224);
nand U6049 (N_6049,N_5437,N_5737);
or U6050 (N_6050,N_5878,N_4877);
nand U6051 (N_6051,N_4755,N_4271);
nand U6052 (N_6052,N_4741,N_5945);
nor U6053 (N_6053,N_4898,N_5381);
xor U6054 (N_6054,N_5942,N_5998);
and U6055 (N_6055,N_4178,N_5176);
nor U6056 (N_6056,N_5823,N_4293);
nor U6057 (N_6057,N_5695,N_5680);
or U6058 (N_6058,N_5478,N_5816);
xor U6059 (N_6059,N_4265,N_4596);
nand U6060 (N_6060,N_4501,N_4526);
or U6061 (N_6061,N_5221,N_5065);
and U6062 (N_6062,N_4095,N_4449);
and U6063 (N_6063,N_4558,N_5659);
and U6064 (N_6064,N_5469,N_4444);
nor U6065 (N_6065,N_4248,N_4792);
nor U6066 (N_6066,N_5952,N_4870);
nand U6067 (N_6067,N_5201,N_4331);
xnor U6068 (N_6068,N_5836,N_5841);
nor U6069 (N_6069,N_5772,N_5446);
nor U6070 (N_6070,N_5260,N_4519);
nand U6071 (N_6071,N_5939,N_4781);
and U6072 (N_6072,N_5003,N_5980);
and U6073 (N_6073,N_4298,N_5012);
nor U6074 (N_6074,N_5997,N_5403);
and U6075 (N_6075,N_5563,N_4254);
xnor U6076 (N_6076,N_5413,N_4619);
nor U6077 (N_6077,N_5528,N_5968);
nor U6078 (N_6078,N_5145,N_4687);
and U6079 (N_6079,N_5568,N_4187);
xor U6080 (N_6080,N_4494,N_4883);
nand U6081 (N_6081,N_4848,N_5226);
or U6082 (N_6082,N_4982,N_5066);
or U6083 (N_6083,N_4015,N_5276);
or U6084 (N_6084,N_4216,N_5499);
or U6085 (N_6085,N_5678,N_5101);
xor U6086 (N_6086,N_5778,N_5726);
and U6087 (N_6087,N_5219,N_5874);
or U6088 (N_6088,N_5231,N_5307);
xor U6089 (N_6089,N_5214,N_5188);
and U6090 (N_6090,N_5870,N_4556);
xor U6091 (N_6091,N_4711,N_4948);
xnor U6092 (N_6092,N_5995,N_4991);
nor U6093 (N_6093,N_4112,N_4719);
xnor U6094 (N_6094,N_5564,N_4124);
and U6095 (N_6095,N_5704,N_4056);
xor U6096 (N_6096,N_5783,N_5367);
and U6097 (N_6097,N_5906,N_4260);
xor U6098 (N_6098,N_4397,N_4003);
or U6099 (N_6099,N_5027,N_5570);
nor U6100 (N_6100,N_5712,N_4040);
nand U6101 (N_6101,N_4239,N_5890);
xor U6102 (N_6102,N_5593,N_4165);
nor U6103 (N_6103,N_4591,N_5742);
xor U6104 (N_6104,N_5494,N_4632);
nor U6105 (N_6105,N_5429,N_5780);
nor U6106 (N_6106,N_4096,N_4757);
xnor U6107 (N_6107,N_5001,N_4303);
and U6108 (N_6108,N_5122,N_4094);
nand U6109 (N_6109,N_4332,N_4973);
nand U6110 (N_6110,N_4790,N_5179);
nand U6111 (N_6111,N_4195,N_4155);
nor U6112 (N_6112,N_4339,N_5895);
or U6113 (N_6113,N_4814,N_4552);
xnor U6114 (N_6114,N_5846,N_4512);
nand U6115 (N_6115,N_5769,N_5690);
nor U6116 (N_6116,N_4884,N_5308);
nand U6117 (N_6117,N_4000,N_4177);
nor U6118 (N_6118,N_5309,N_4442);
nor U6119 (N_6119,N_5082,N_4925);
nand U6120 (N_6120,N_5002,N_5043);
nor U6121 (N_6121,N_5433,N_4764);
xor U6122 (N_6122,N_5149,N_4680);
or U6123 (N_6123,N_5228,N_5625);
nand U6124 (N_6124,N_5809,N_5211);
and U6125 (N_6125,N_5957,N_4841);
and U6126 (N_6126,N_5965,N_4933);
and U6127 (N_6127,N_5472,N_5586);
nor U6128 (N_6128,N_5165,N_5288);
nand U6129 (N_6129,N_4770,N_4162);
nor U6130 (N_6130,N_4447,N_4601);
nand U6131 (N_6131,N_5834,N_5732);
xor U6132 (N_6132,N_4381,N_5120);
and U6133 (N_6133,N_4364,N_5792);
or U6134 (N_6134,N_5985,N_4759);
or U6135 (N_6135,N_5407,N_5021);
and U6136 (N_6136,N_4076,N_4021);
and U6137 (N_6137,N_4459,N_5166);
xnor U6138 (N_6138,N_4725,N_5766);
nand U6139 (N_6139,N_5454,N_5422);
nand U6140 (N_6140,N_5453,N_4477);
xor U6141 (N_6141,N_4557,N_5526);
nand U6142 (N_6142,N_5130,N_4935);
or U6143 (N_6143,N_5767,N_5688);
xor U6144 (N_6144,N_5303,N_4789);
nor U6145 (N_6145,N_4312,N_5281);
and U6146 (N_6146,N_4820,N_5329);
xor U6147 (N_6147,N_4218,N_5632);
xnor U6148 (N_6148,N_5046,N_5610);
nor U6149 (N_6149,N_4536,N_5860);
xnor U6150 (N_6150,N_5833,N_4409);
and U6151 (N_6151,N_5497,N_5404);
xor U6152 (N_6152,N_5960,N_5639);
or U6153 (N_6153,N_4832,N_4361);
and U6154 (N_6154,N_5547,N_4173);
or U6155 (N_6155,N_5335,N_4726);
and U6156 (N_6156,N_5022,N_5738);
nand U6157 (N_6157,N_4852,N_5590);
nor U6158 (N_6158,N_4943,N_5934);
and U6159 (N_6159,N_4105,N_4425);
nor U6160 (N_6160,N_5949,N_4069);
nor U6161 (N_6161,N_4139,N_5669);
xor U6162 (N_6162,N_5891,N_5668);
and U6163 (N_6163,N_5902,N_4588);
or U6164 (N_6164,N_4844,N_4290);
nand U6165 (N_6165,N_4585,N_4829);
or U6166 (N_6166,N_4629,N_5810);
and U6167 (N_6167,N_4567,N_5579);
nand U6168 (N_6168,N_5677,N_4412);
nand U6169 (N_6169,N_4869,N_5693);
nor U6170 (N_6170,N_5592,N_4862);
xnor U6171 (N_6171,N_4666,N_5121);
or U6172 (N_6172,N_4059,N_4300);
and U6173 (N_6173,N_5443,N_4845);
nand U6174 (N_6174,N_5277,N_5162);
or U6175 (N_6175,N_5585,N_4915);
or U6176 (N_6176,N_5378,N_5627);
nand U6177 (N_6177,N_4754,N_4240);
nor U6178 (N_6178,N_5648,N_4380);
and U6179 (N_6179,N_4058,N_4984);
xnor U6180 (N_6180,N_5931,N_5831);
and U6181 (N_6181,N_5969,N_5030);
and U6182 (N_6182,N_5054,N_4209);
and U6183 (N_6183,N_4448,N_5575);
xnor U6184 (N_6184,N_4524,N_4694);
nand U6185 (N_6185,N_5553,N_4227);
and U6186 (N_6186,N_4568,N_4768);
xor U6187 (N_6187,N_5966,N_4854);
nor U6188 (N_6188,N_4182,N_5333);
nand U6189 (N_6189,N_5624,N_4100);
and U6190 (N_6190,N_4663,N_4326);
or U6191 (N_6191,N_5081,N_5658);
nor U6192 (N_6192,N_4795,N_5896);
xnor U6193 (N_6193,N_5743,N_4198);
nor U6194 (N_6194,N_5527,N_4233);
xnor U6195 (N_6195,N_4476,N_4065);
and U6196 (N_6196,N_5311,N_5605);
nand U6197 (N_6197,N_4295,N_4267);
nand U6198 (N_6198,N_4263,N_5353);
nand U6199 (N_6199,N_4462,N_4583);
or U6200 (N_6200,N_5153,N_5572);
xor U6201 (N_6201,N_5866,N_5576);
nor U6202 (N_6202,N_5758,N_4002);
nand U6203 (N_6203,N_5880,N_5935);
and U6204 (N_6204,N_5999,N_4342);
nor U6205 (N_6205,N_4019,N_5394);
xnor U6206 (N_6206,N_5824,N_4866);
nand U6207 (N_6207,N_4780,N_5349);
or U6208 (N_6208,N_5932,N_4990);
nor U6209 (N_6209,N_5273,N_4273);
and U6210 (N_6210,N_4902,N_4861);
xor U6211 (N_6211,N_5215,N_5033);
nor U6212 (N_6212,N_4199,N_5936);
nand U6213 (N_6213,N_5405,N_5974);
xor U6214 (N_6214,N_4064,N_4615);
nor U6215 (N_6215,N_4788,N_4562);
nand U6216 (N_6216,N_4471,N_5198);
nand U6217 (N_6217,N_4049,N_4977);
and U6218 (N_6218,N_4801,N_5267);
xnor U6219 (N_6219,N_5068,N_5609);
xor U6220 (N_6220,N_5334,N_5976);
and U6221 (N_6221,N_5280,N_4377);
or U6222 (N_6222,N_4424,N_5583);
and U6223 (N_6223,N_4289,N_4665);
and U6224 (N_6224,N_4167,N_5750);
nor U6225 (N_6225,N_5723,N_5079);
or U6226 (N_6226,N_4513,N_5284);
xnor U6227 (N_6227,N_4621,N_5197);
or U6228 (N_6228,N_4658,N_5072);
or U6229 (N_6229,N_5924,N_5943);
and U6230 (N_6230,N_4613,N_5561);
or U6231 (N_6231,N_4466,N_5200);
or U6232 (N_6232,N_4288,N_4134);
and U6233 (N_6233,N_5252,N_5045);
nor U6234 (N_6234,N_5416,N_5460);
xnor U6235 (N_6235,N_5613,N_4537);
or U6236 (N_6236,N_5191,N_4472);
xor U6237 (N_6237,N_5293,N_4231);
or U6238 (N_6238,N_4484,N_4246);
nor U6239 (N_6239,N_5623,N_5569);
nor U6240 (N_6240,N_5811,N_4128);
nor U6241 (N_6241,N_5319,N_5463);
nor U6242 (N_6242,N_4661,N_4098);
nor U6243 (N_6243,N_4111,N_5438);
nor U6244 (N_6244,N_4219,N_4256);
and U6245 (N_6245,N_5470,N_5055);
and U6246 (N_6246,N_4153,N_4529);
and U6247 (N_6247,N_5173,N_5837);
nand U6248 (N_6248,N_5944,N_4971);
nand U6249 (N_6249,N_4318,N_4509);
nand U6250 (N_6250,N_4132,N_4835);
nand U6251 (N_6251,N_5289,N_5981);
xnor U6252 (N_6252,N_5315,N_4214);
and U6253 (N_6253,N_4878,N_5971);
nand U6254 (N_6254,N_4565,N_4699);
nor U6255 (N_6255,N_4874,N_4099);
or U6256 (N_6256,N_4463,N_5243);
and U6257 (N_6257,N_5141,N_4994);
and U6258 (N_6258,N_5958,N_5522);
or U6259 (N_6259,N_4030,N_5377);
or U6260 (N_6260,N_5611,N_5951);
nor U6261 (N_6261,N_5004,N_4718);
and U6262 (N_6262,N_5414,N_4088);
and U6263 (N_6263,N_4491,N_4388);
or U6264 (N_6264,N_4993,N_5886);
nor U6265 (N_6265,N_4347,N_4196);
nand U6266 (N_6266,N_5941,N_5139);
nor U6267 (N_6267,N_4838,N_5914);
xnor U6268 (N_6268,N_4394,N_5113);
xnor U6269 (N_6269,N_5975,N_4249);
or U6270 (N_6270,N_4603,N_4037);
nor U6271 (N_6271,N_4976,N_4504);
nand U6272 (N_6272,N_4321,N_5946);
xor U6273 (N_6273,N_5389,N_4539);
and U6274 (N_6274,N_5967,N_5269);
and U6275 (N_6275,N_5530,N_5227);
nor U6276 (N_6276,N_5133,N_5274);
nor U6277 (N_6277,N_5229,N_5395);
or U6278 (N_6278,N_4079,N_4287);
xnor U6279 (N_6279,N_4437,N_5323);
xnor U6280 (N_6280,N_4840,N_5222);
and U6281 (N_6281,N_4825,N_5480);
nor U6282 (N_6282,N_4296,N_5571);
nor U6283 (N_6283,N_5005,N_4488);
xor U6284 (N_6284,N_4348,N_5889);
xor U6285 (N_6285,N_5250,N_4275);
xor U6286 (N_6286,N_5451,N_4607);
nand U6287 (N_6287,N_5447,N_4510);
nand U6288 (N_6288,N_5468,N_4882);
nor U6289 (N_6289,N_5616,N_4220);
and U6290 (N_6290,N_4681,N_4356);
nand U6291 (N_6291,N_4434,N_4368);
or U6292 (N_6292,N_5092,N_5800);
nand U6293 (N_6293,N_5794,N_5597);
xnor U6294 (N_6294,N_5711,N_5341);
and U6295 (N_6295,N_5925,N_4432);
and U6296 (N_6296,N_4149,N_5247);
or U6297 (N_6297,N_4691,N_4783);
nor U6298 (N_6298,N_5304,N_5788);
nor U6299 (N_6299,N_4033,N_5691);
and U6300 (N_6300,N_4404,N_5441);
xnor U6301 (N_6301,N_5491,N_4604);
nor U6302 (N_6302,N_4039,N_4888);
or U6303 (N_6303,N_4235,N_4980);
or U6304 (N_6304,N_4113,N_4589);
and U6305 (N_6305,N_5393,N_5015);
xor U6306 (N_6306,N_5235,N_4673);
xnor U6307 (N_6307,N_5556,N_4257);
nand U6308 (N_6308,N_5916,N_5595);
xnor U6309 (N_6309,N_5348,N_5671);
and U6310 (N_6310,N_4086,N_4074);
nand U6311 (N_6311,N_4084,N_5127);
nor U6312 (N_6312,N_5410,N_5764);
or U6313 (N_6313,N_4638,N_5128);
nor U6314 (N_6314,N_4778,N_4237);
nand U6315 (N_6315,N_5444,N_5102);
nand U6316 (N_6316,N_5427,N_5209);
or U6317 (N_6317,N_5655,N_4057);
and U6318 (N_6318,N_5701,N_5099);
nand U6319 (N_6319,N_4334,N_4353);
or U6320 (N_6320,N_4495,N_5970);
nor U6321 (N_6321,N_4954,N_4011);
or U6322 (N_6322,N_4244,N_5821);
or U6323 (N_6323,N_5850,N_4439);
or U6324 (N_6324,N_4677,N_4891);
nor U6325 (N_6325,N_5119,N_5014);
or U6326 (N_6326,N_4749,N_5336);
nor U6327 (N_6327,N_4934,N_4910);
nand U6328 (N_6328,N_5620,N_5032);
xor U6329 (N_6329,N_5955,N_4478);
xor U6330 (N_6330,N_4761,N_5483);
xnor U6331 (N_6331,N_5859,N_4507);
or U6332 (N_6332,N_5884,N_5700);
nor U6333 (N_6333,N_5351,N_5291);
nor U6334 (N_6334,N_4630,N_5430);
or U6335 (N_6335,N_4929,N_4742);
nor U6336 (N_6336,N_4587,N_5069);
or U6337 (N_6337,N_4390,N_5324);
and U6338 (N_6338,N_5512,N_4206);
or U6339 (N_6339,N_4483,N_5086);
nand U6340 (N_6340,N_5445,N_5724);
xor U6341 (N_6341,N_5630,N_5013);
nor U6342 (N_6342,N_4774,N_4194);
xnor U6343 (N_6343,N_5802,N_5440);
and U6344 (N_6344,N_4532,N_5155);
and U6345 (N_6345,N_4593,N_5727);
and U6346 (N_6346,N_5134,N_4685);
and U6347 (N_6347,N_5617,N_5555);
nor U6348 (N_6348,N_5224,N_5398);
xnor U6349 (N_6349,N_5557,N_4890);
or U6350 (N_6350,N_4160,N_5047);
nand U6351 (N_6351,N_4461,N_4894);
nor U6352 (N_6352,N_4414,N_5718);
nor U6353 (N_6353,N_4701,N_4422);
nor U6354 (N_6354,N_4516,N_4606);
or U6355 (N_6355,N_5116,N_4141);
and U6356 (N_6356,N_5278,N_4947);
nor U6357 (N_6357,N_5305,N_4895);
and U6358 (N_6358,N_4705,N_4129);
nand U6359 (N_6359,N_4995,N_4335);
nor U6360 (N_6360,N_4714,N_4530);
nand U6361 (N_6361,N_4972,N_4497);
nor U6362 (N_6362,N_5851,N_4833);
or U6363 (N_6363,N_5744,N_4395);
nand U6364 (N_6364,N_5708,N_4174);
and U6365 (N_6365,N_5790,N_5301);
and U6366 (N_6366,N_5763,N_4012);
and U6367 (N_6367,N_5423,N_5584);
nand U6368 (N_6368,N_4286,N_5652);
and U6369 (N_6369,N_4161,N_4570);
nor U6370 (N_6370,N_5596,N_5492);
nor U6371 (N_6371,N_4837,N_4842);
xor U6372 (N_6372,N_4796,N_5129);
or U6373 (N_6373,N_4406,N_5515);
nor U6374 (N_6374,N_5745,N_5843);
or U6375 (N_6375,N_4121,N_4091);
xor U6376 (N_6376,N_4763,N_4078);
or U6377 (N_6377,N_5136,N_5401);
xor U6378 (N_6378,N_5911,N_5255);
nand U6379 (N_6379,N_4575,N_5431);
nor U6380 (N_6380,N_5773,N_5748);
nand U6381 (N_6381,N_4253,N_4944);
xnor U6382 (N_6382,N_5747,N_4435);
nand U6383 (N_6383,N_5504,N_5832);
nand U6384 (N_6384,N_4281,N_5684);
and U6385 (N_6385,N_4952,N_4370);
nor U6386 (N_6386,N_4758,N_4965);
and U6387 (N_6387,N_4085,N_4600);
or U6388 (N_6388,N_5070,N_5805);
or U6389 (N_6389,N_4533,N_5959);
or U6390 (N_6390,N_4736,N_5485);
and U6391 (N_6391,N_5867,N_5900);
nand U6392 (N_6392,N_5674,N_5223);
xnor U6393 (N_6393,N_5318,N_4745);
nand U6394 (N_6394,N_5044,N_4077);
xor U6395 (N_6395,N_4465,N_5779);
or U6396 (N_6396,N_4545,N_5118);
xor U6397 (N_6397,N_5031,N_4297);
nor U6398 (N_6398,N_5412,N_4067);
nor U6399 (N_6399,N_5785,N_4492);
and U6400 (N_6400,N_4211,N_4150);
nor U6401 (N_6401,N_5741,N_4051);
xor U6402 (N_6402,N_4986,N_4304);
or U6403 (N_6403,N_5272,N_5213);
nand U6404 (N_6404,N_5245,N_4359);
and U6405 (N_6405,N_4423,N_5169);
nor U6406 (N_6406,N_5927,N_4264);
xor U6407 (N_6407,N_4928,N_4203);
xnor U6408 (N_6408,N_5713,N_4418);
nand U6409 (N_6409,N_5760,N_4400);
nor U6410 (N_6410,N_4357,N_5095);
xor U6411 (N_6411,N_5543,N_4816);
nand U6412 (N_6412,N_4614,N_4847);
xor U6413 (N_6413,N_4176,N_5518);
or U6414 (N_6414,N_5513,N_4865);
xnor U6415 (N_6415,N_5037,N_5567);
nor U6416 (N_6416,N_5479,N_5885);
nand U6417 (N_6417,N_5195,N_4133);
nand U6418 (N_6418,N_5464,N_4311);
and U6419 (N_6419,N_4698,N_5409);
and U6420 (N_6420,N_4744,N_4171);
and U6421 (N_6421,N_5722,N_5275);
nand U6422 (N_6422,N_5108,N_5230);
xor U6423 (N_6423,N_4554,N_4292);
nor U6424 (N_6424,N_4333,N_4351);
xnor U6425 (N_6425,N_5042,N_5481);
nor U6426 (N_6426,N_5534,N_4323);
nand U6427 (N_6427,N_4120,N_5524);
or U6428 (N_6428,N_5715,N_4987);
and U6429 (N_6429,N_4066,N_4896);
nor U6430 (N_6430,N_5877,N_4366);
and U6431 (N_6431,N_4158,N_4169);
or U6432 (N_6432,N_4043,N_5771);
or U6433 (N_6433,N_4103,N_4889);
nand U6434 (N_6434,N_5117,N_5150);
and U6435 (N_6435,N_5604,N_5125);
or U6436 (N_6436,N_5915,N_4779);
nand U6437 (N_6437,N_4908,N_4616);
and U6438 (N_6438,N_5112,N_4953);
nand U6439 (N_6439,N_4416,N_4563);
nor U6440 (N_6440,N_4608,N_5057);
nor U6441 (N_6441,N_5808,N_5190);
xor U6442 (N_6442,N_4876,N_5158);
and U6443 (N_6443,N_4301,N_5918);
xnor U6444 (N_6444,N_5283,N_5905);
or U6445 (N_6445,N_5626,N_4401);
and U6446 (N_6446,N_5849,N_4654);
xnor U6447 (N_6447,N_5131,N_5689);
xnor U6448 (N_6448,N_5539,N_5177);
and U6449 (N_6449,N_5819,N_5007);
and U6450 (N_6450,N_4486,N_5178);
xnor U6451 (N_6451,N_5574,N_4598);
xor U6452 (N_6452,N_5257,N_5362);
and U6453 (N_6453,N_4785,N_4345);
nand U6454 (N_6454,N_5107,N_4481);
nor U6455 (N_6455,N_4893,N_4317);
xor U6456 (N_6456,N_4753,N_4159);
xnor U6457 (N_6457,N_5872,N_5551);
or U6458 (N_6458,N_4923,N_4542);
and U6459 (N_6459,N_4398,N_5651);
xnor U6460 (N_6460,N_4147,N_5418);
nor U6461 (N_6461,N_4146,N_5084);
xor U6462 (N_6462,N_5582,N_4875);
nand U6463 (N_6463,N_4032,N_5799);
nor U6464 (N_6464,N_4467,N_5937);
xor U6465 (N_6465,N_5922,N_5168);
xnor U6466 (N_6466,N_4702,N_5034);
and U6467 (N_6467,N_4070,N_4389);
or U6468 (N_6468,N_4371,N_5238);
and U6469 (N_6469,N_4383,N_5725);
nand U6470 (N_6470,N_4784,N_5203);
and U6471 (N_6471,N_5558,N_4081);
xor U6472 (N_6472,N_4046,N_4712);
or U6473 (N_6473,N_5262,N_5369);
or U6474 (N_6474,N_5853,N_4863);
nor U6475 (N_6475,N_5672,N_4341);
nor U6476 (N_6476,N_5008,N_4999);
nor U6477 (N_6477,N_5899,N_4071);
and U6478 (N_6478,N_5598,N_4215);
and U6479 (N_6479,N_4722,N_5338);
nor U6480 (N_6480,N_4584,N_5873);
nor U6481 (N_6481,N_5379,N_4140);
nand U6482 (N_6482,N_4252,N_4322);
or U6483 (N_6483,N_4005,N_4352);
xor U6484 (N_6484,N_5840,N_5415);
xor U6485 (N_6485,N_5983,N_5023);
nor U6486 (N_6486,N_5554,N_4041);
nand U6487 (N_6487,N_5370,N_5820);
xor U6488 (N_6488,N_4184,N_4234);
nor U6489 (N_6489,N_5477,N_4101);
or U6490 (N_6490,N_5220,N_5105);
nand U6491 (N_6491,N_4279,N_4599);
or U6492 (N_6492,N_5088,N_5384);
nor U6493 (N_6493,N_4365,N_5344);
and U6494 (N_6494,N_5160,N_4793);
nor U6495 (N_6495,N_4669,N_5656);
nor U6496 (N_6496,N_5920,N_4560);
and U6497 (N_6497,N_5452,N_5455);
and U6498 (N_6498,N_5077,N_4411);
and U6499 (N_6499,N_5666,N_4752);
nand U6500 (N_6500,N_5664,N_4746);
or U6501 (N_6501,N_5080,N_4044);
nand U6502 (N_6502,N_4922,N_4968);
nor U6503 (N_6503,N_4962,N_5685);
or U6504 (N_6504,N_4873,N_5270);
and U6505 (N_6505,N_4975,N_5019);
xnor U6506 (N_6506,N_5368,N_4107);
nand U6507 (N_6507,N_4731,N_5986);
and U6508 (N_6508,N_4482,N_5897);
or U6509 (N_6509,N_4429,N_5109);
nand U6510 (N_6510,N_5565,N_4750);
xnor U6511 (N_6511,N_4941,N_5114);
nor U6512 (N_6512,N_5347,N_4142);
xnor U6513 (N_6513,N_5244,N_5350);
or U6514 (N_6514,N_4737,N_4931);
nand U6515 (N_6515,N_4453,N_5545);
or U6516 (N_6516,N_5954,N_5011);
nor U6517 (N_6517,N_4548,N_4255);
nor U6518 (N_6518,N_5420,N_4399);
nor U6519 (N_6519,N_5016,N_5298);
xnor U6520 (N_6520,N_4498,N_4826);
nor U6521 (N_6521,N_4468,N_5754);
nor U6522 (N_6522,N_4385,N_4799);
or U6523 (N_6523,N_5864,N_5049);
and U6524 (N_6524,N_4500,N_4885);
xor U6525 (N_6525,N_4727,N_4868);
and U6526 (N_6526,N_5580,N_5402);
and U6527 (N_6527,N_4946,N_5665);
or U6528 (N_6528,N_4791,N_5181);
and U6529 (N_6529,N_5061,N_4671);
xor U6530 (N_6530,N_5450,N_5041);
xor U6531 (N_6531,N_4960,N_5364);
nor U6532 (N_6532,N_5888,N_4183);
or U6533 (N_6533,N_4329,N_4642);
and U6534 (N_6534,N_4152,N_4028);
xor U6535 (N_6535,N_5206,N_5560);
nand U6536 (N_6536,N_4054,N_4170);
nor U6537 (N_6537,N_5812,N_5856);
and U6538 (N_6538,N_5822,N_5775);
and U6539 (N_6539,N_5559,N_4914);
or U6540 (N_6540,N_4052,N_5089);
nor U6541 (N_6541,N_4867,N_5894);
xor U6542 (N_6542,N_5660,N_4903);
xnor U6543 (N_6543,N_4909,N_5514);
or U6544 (N_6544,N_5928,N_4949);
nor U6545 (N_6545,N_4082,N_5717);
nor U6546 (N_6546,N_5039,N_4858);
or U6547 (N_6547,N_5074,N_5903);
nor U6548 (N_6548,N_4407,N_5050);
xnor U6549 (N_6549,N_4821,N_5901);
or U6550 (N_6550,N_4967,N_5266);
xor U6551 (N_6551,N_4733,N_5517);
nand U6552 (N_6552,N_4859,N_4628);
xor U6553 (N_6553,N_4228,N_5144);
nor U6554 (N_6554,N_5752,N_4786);
and U6555 (N_6555,N_4541,N_5509);
and U6556 (N_6556,N_5439,N_5239);
or U6557 (N_6557,N_5146,N_5059);
nand U6558 (N_6558,N_4667,N_4625);
and U6559 (N_6559,N_4551,N_5879);
nand U6560 (N_6560,N_4800,N_4480);
xnor U6561 (N_6561,N_5520,N_5359);
xor U6562 (N_6562,N_4327,N_5829);
xnor U6563 (N_6563,N_4245,N_4940);
or U6564 (N_6564,N_4458,N_4164);
and U6565 (N_6565,N_5372,N_5355);
xor U6566 (N_6566,N_5465,N_4721);
nand U6567 (N_6567,N_5496,N_4307);
or U6568 (N_6568,N_5171,N_4916);
xnor U6569 (N_6569,N_4724,N_5048);
nor U6570 (N_6570,N_4269,N_4125);
xnor U6571 (N_6571,N_5679,N_5320);
or U6572 (N_6572,N_4586,N_5774);
nand U6573 (N_6573,N_5898,N_4595);
nand U6574 (N_6574,N_5544,N_5621);
or U6575 (N_6575,N_4470,N_5352);
nand U6576 (N_6576,N_5332,N_5321);
and U6577 (N_6577,N_4415,N_4156);
xnor U6578 (N_6578,N_4650,N_5185);
xnor U6579 (N_6579,N_5432,N_5071);
or U6580 (N_6580,N_4168,N_5813);
or U6581 (N_6581,N_5791,N_5692);
or U6582 (N_6582,N_4363,N_5075);
nand U6583 (N_6583,N_5435,N_5588);
nor U6584 (N_6584,N_5417,N_5297);
xor U6585 (N_6585,N_5038,N_4266);
nand U6586 (N_6586,N_5529,N_5825);
xor U6587 (N_6587,N_5115,N_5279);
or U6588 (N_6588,N_5110,N_4145);
nor U6589 (N_6589,N_4338,N_4649);
and U6590 (N_6590,N_5411,N_5755);
nand U6591 (N_6591,N_5210,N_5506);
nor U6592 (N_6592,N_5532,N_4523);
and U6593 (N_6593,N_4229,N_4426);
nand U6594 (N_6594,N_4605,N_4201);
nand U6595 (N_6595,N_4284,N_4887);
xnor U6596 (N_6596,N_4626,N_5855);
xnor U6597 (N_6597,N_5657,N_5424);
nor U6598 (N_6598,N_4243,N_5067);
or U6599 (N_6599,N_5374,N_4299);
xor U6600 (N_6600,N_5531,N_4376);
and U6601 (N_6601,N_4897,N_4921);
nand U6602 (N_6602,N_5241,N_5719);
xnor U6603 (N_6603,N_4350,N_4904);
and U6604 (N_6604,N_5457,N_5993);
and U6605 (N_6605,N_4707,N_5702);
and U6606 (N_6606,N_5521,N_5881);
nor U6607 (N_6607,N_5653,N_4729);
and U6608 (N_6608,N_4042,N_4251);
xor U6609 (N_6609,N_4728,N_5018);
xor U6610 (N_6610,N_4427,N_4782);
and U6611 (N_6611,N_4020,N_5933);
xor U6612 (N_6612,N_4362,N_4672);
nor U6613 (N_6613,N_4978,N_5844);
nand U6614 (N_6614,N_4643,N_4817);
xnor U6615 (N_6615,N_4696,N_5919);
and U6616 (N_6616,N_4807,N_4703);
nor U6617 (N_6617,N_4812,N_4818);
nand U6618 (N_6618,N_4535,N_4963);
nand U6619 (N_6619,N_5646,N_5237);
or U6620 (N_6620,N_4566,N_5449);
nor U6621 (N_6621,N_4851,N_5124);
or U6622 (N_6622,N_4217,N_5212);
nand U6623 (N_6623,N_4428,N_5459);
xor U6624 (N_6624,N_4457,N_5803);
or U6625 (N_6625,N_4580,N_4907);
nor U6626 (N_6626,N_4060,N_5342);
nor U6627 (N_6627,N_5286,N_5428);
nor U6628 (N_6628,N_5271,N_4372);
and U6629 (N_6629,N_5363,N_5151);
or U6630 (N_6630,N_4634,N_4709);
and U6631 (N_6631,N_4639,N_4766);
nand U6632 (N_6632,N_4617,N_4652);
and U6633 (N_6633,N_4319,N_5263);
nand U6634 (N_6634,N_5140,N_4794);
or U6635 (N_6635,N_5204,N_4751);
or U6636 (N_6636,N_4942,N_5977);
xor U6637 (N_6637,N_4200,N_4937);
or U6638 (N_6638,N_4983,N_4670);
or U6639 (N_6639,N_4018,N_5388);
or U6640 (N_6640,N_4739,N_5006);
nand U6641 (N_6641,N_5759,N_4204);
xor U6642 (N_6642,N_4274,N_4911);
or U6643 (N_6643,N_5686,N_4208);
xnor U6644 (N_6644,N_4905,N_5817);
nand U6645 (N_6645,N_4225,N_5830);
xnor U6646 (N_6646,N_5929,N_4118);
or U6647 (N_6647,N_4917,N_4123);
xor U6648 (N_6648,N_4278,N_5083);
xnor U6649 (N_6649,N_5599,N_4316);
or U6650 (N_6650,N_4210,N_4460);
and U6651 (N_6651,N_4930,N_5541);
or U6652 (N_6652,N_5490,N_5287);
and U6653 (N_6653,N_4964,N_4561);
nor U6654 (N_6654,N_4309,N_4469);
xor U6655 (N_6655,N_5662,N_4676);
and U6656 (N_6656,N_4102,N_4572);
nand U6657 (N_6657,N_4543,N_4010);
and U6658 (N_6658,N_4131,N_4700);
and U6659 (N_6659,N_4027,N_5192);
or U6660 (N_6660,N_4180,N_4511);
xnor U6661 (N_6661,N_4247,N_4387);
or U6662 (N_6662,N_4880,N_4578);
or U6663 (N_6663,N_5087,N_5607);
nor U6664 (N_6664,N_5940,N_4958);
nand U6665 (N_6665,N_4104,N_4564);
nand U6666 (N_6666,N_5594,N_4646);
nand U6667 (N_6667,N_4354,N_5839);
xor U6668 (N_6668,N_4310,N_5962);
xor U6669 (N_6669,N_5781,N_5984);
nand U6670 (N_6670,N_4597,N_5699);
nor U6671 (N_6671,N_5912,N_4864);
nor U6672 (N_6672,N_5996,N_4689);
xor U6673 (N_6673,N_4063,N_4576);
xor U6674 (N_6674,N_4527,N_5591);
or U6675 (N_6675,N_4277,N_4130);
or U6676 (N_6676,N_4645,N_5549);
nor U6677 (N_6677,N_4349,N_5325);
xor U6678 (N_6678,N_5078,N_4730);
or U6679 (N_6679,N_5765,N_5373);
nand U6680 (N_6680,N_4828,N_5815);
and U6681 (N_6681,N_5328,N_4270);
nor U6682 (N_6682,N_4222,N_5675);
nand U6683 (N_6683,N_4014,N_4506);
nand U6684 (N_6684,N_5989,N_5062);
or U6685 (N_6685,N_4855,N_4272);
nand U6686 (N_6686,N_4047,N_4117);
xor U6687 (N_6687,N_4479,N_4573);
or U6688 (N_6688,N_5383,N_5854);
or U6689 (N_6689,N_5904,N_4185);
nand U6690 (N_6690,N_4686,N_4172);
or U6691 (N_6691,N_5098,N_5797);
xnor U6692 (N_6692,N_5573,N_4212);
xor U6693 (N_6693,N_5796,N_5295);
or U6694 (N_6694,N_4981,N_4979);
nor U6695 (N_6695,N_5473,N_4996);
nand U6696 (N_6696,N_4384,N_4306);
nor U6697 (N_6697,N_4386,N_5157);
nand U6698 (N_6698,N_4450,N_4382);
or U6699 (N_6699,N_4061,N_5603);
nor U6700 (N_6700,N_4122,N_4119);
and U6701 (N_6701,N_4811,N_4956);
nand U6702 (N_6702,N_4106,N_4710);
or U6703 (N_6703,N_4114,N_5858);
and U6704 (N_6704,N_5687,N_5218);
xor U6705 (N_6705,N_5093,N_4966);
nor U6706 (N_6706,N_5489,N_4029);
nand U6707 (N_6707,N_5024,N_5868);
or U6708 (N_6708,N_4116,N_5994);
nand U6709 (N_6709,N_5893,N_5908);
nand U6710 (N_6710,N_4959,N_5063);
nor U6711 (N_6711,N_4734,N_4517);
nor U6712 (N_6712,N_5519,N_5501);
and U6713 (N_6713,N_4927,N_4241);
nor U6714 (N_6714,N_4769,N_5256);
nor U6715 (N_6715,N_5391,N_5029);
and U6716 (N_6716,N_5892,N_5838);
or U6717 (N_6717,N_4945,N_4827);
or U6718 (N_6718,N_5663,N_4618);
or U6719 (N_6719,N_5052,N_4682);
xor U6720 (N_6720,N_5510,N_5871);
or U6721 (N_6721,N_4693,N_4776);
nor U6722 (N_6722,N_4431,N_4857);
and U6723 (N_6723,N_4489,N_5097);
or U6724 (N_6724,N_4610,N_4899);
nand U6725 (N_6725,N_5845,N_5807);
nand U6726 (N_6726,N_4684,N_5804);
and U6727 (N_6727,N_4824,N_4226);
and U6728 (N_6728,N_4004,N_4001);
or U6729 (N_6729,N_5090,N_5777);
and U6730 (N_6730,N_4651,N_4697);
nor U6731 (N_6731,N_4555,N_5644);
and U6732 (N_6732,N_4708,N_4135);
nand U6733 (N_6733,N_5857,N_5236);
or U6734 (N_6734,N_5776,N_5523);
xnor U6735 (N_6735,N_5618,N_4007);
nor U6736 (N_6736,N_4087,N_4268);
and U6737 (N_6737,N_4419,N_5736);
or U6738 (N_6738,N_5380,N_4538);
nand U6739 (N_6739,N_5317,N_4451);
nor U6740 (N_6740,N_5292,N_5733);
or U6741 (N_6741,N_4024,N_5647);
xnor U6742 (N_6742,N_4836,N_4823);
nand U6743 (N_6743,N_5930,N_5399);
or U6744 (N_6744,N_5835,N_5265);
or U6745 (N_6745,N_5000,N_5184);
and U6746 (N_6746,N_4343,N_5330);
nand U6747 (N_6747,N_4464,N_5009);
xnor U6748 (N_6748,N_5721,N_4505);
nand U6749 (N_6749,N_4314,N_4276);
or U6750 (N_6750,N_5240,N_4985);
nor U6751 (N_6751,N_4221,N_4189);
nand U6752 (N_6752,N_5442,N_4624);
xor U6753 (N_6753,N_4961,N_4970);
nand U6754 (N_6754,N_4912,N_4640);
or U6755 (N_6755,N_4773,N_5972);
and U6756 (N_6756,N_5340,N_5106);
or U6757 (N_6757,N_5073,N_4006);
or U6758 (N_6758,N_5261,N_5296);
or U6759 (N_6759,N_5180,N_5358);
or U6760 (N_6760,N_4025,N_5577);
nor U6761 (N_6761,N_5566,N_5847);
nor U6762 (N_6762,N_4262,N_5175);
and U6763 (N_6763,N_4421,N_4787);
and U6764 (N_6764,N_4860,N_4474);
and U6765 (N_6765,N_4765,N_4974);
nand U6766 (N_6766,N_4822,N_5503);
nor U6767 (N_6767,N_5462,N_5474);
nand U6768 (N_6768,N_4518,N_4315);
xor U6769 (N_6769,N_4259,N_5147);
and U6770 (N_6770,N_4360,N_5208);
or U6771 (N_6771,N_4320,N_5248);
and U6772 (N_6772,N_5300,N_4664);
nand U6773 (N_6773,N_5682,N_4402);
xnor U6774 (N_6774,N_5917,N_5716);
xor U6775 (N_6775,N_5493,N_5233);
nor U6776 (N_6776,N_5731,N_4108);
or U6777 (N_6777,N_4571,N_4408);
nand U6778 (N_6778,N_5028,N_5863);
nor U6779 (N_6779,N_5216,N_5990);
and U6780 (N_6780,N_5676,N_5533);
nor U6781 (N_6781,N_4109,N_4988);
and U6782 (N_6782,N_5642,N_5782);
and U6783 (N_6783,N_5978,N_4055);
nand U6784 (N_6784,N_5331,N_5705);
and U6785 (N_6785,N_4053,N_5282);
and U6786 (N_6786,N_4230,N_5546);
nor U6787 (N_6787,N_4016,N_4853);
or U6788 (N_6788,N_5182,N_5346);
nor U6789 (N_6789,N_5798,N_5696);
xnor U6790 (N_6790,N_5728,N_5487);
nor U6791 (N_6791,N_5132,N_5339);
nand U6792 (N_6792,N_5910,N_4157);
and U6793 (N_6793,N_4798,N_5875);
nor U6794 (N_6794,N_5154,N_4926);
xnor U6795 (N_6795,N_5681,N_4515);
and U6796 (N_6796,N_5207,N_5793);
nand U6797 (N_6797,N_4436,N_4738);
nor U6798 (N_6798,N_4205,N_4127);
or U6799 (N_6799,N_5654,N_5753);
and U6800 (N_6800,N_5550,N_4647);
or U6801 (N_6801,N_5251,N_5876);
or U6802 (N_6802,N_4692,N_4546);
or U6803 (N_6803,N_4808,N_5562);
nand U6804 (N_6804,N_5476,N_4900);
or U6805 (N_6805,N_5697,N_5104);
xor U6806 (N_6806,N_4772,N_4369);
and U6807 (N_6807,N_4657,N_4594);
and U6808 (N_6808,N_5058,N_4175);
and U6809 (N_6809,N_4850,N_5400);
and U6810 (N_6810,N_5540,N_5387);
or U6811 (N_6811,N_4547,N_5313);
or U6812 (N_6812,N_4740,N_5500);
and U6813 (N_6813,N_4487,N_5163);
and U6814 (N_6814,N_5749,N_4093);
nand U6815 (N_6815,N_4846,N_5761);
or U6816 (N_6816,N_5382,N_5137);
and U6817 (N_6817,N_5667,N_5643);
xor U6818 (N_6818,N_4704,N_4830);
nand U6819 (N_6819,N_5746,N_5035);
and U6820 (N_6820,N_4611,N_5085);
or U6821 (N_6821,N_4748,N_5973);
nor U6822 (N_6822,N_5174,N_4635);
xor U6823 (N_6823,N_5979,N_4879);
and U6824 (N_6824,N_5505,N_5148);
xnor U6825 (N_6825,N_4068,N_5601);
xor U6826 (N_6826,N_5051,N_4213);
xor U6827 (N_6827,N_5706,N_4433);
or U6828 (N_6828,N_5486,N_5017);
nand U6829 (N_6829,N_4553,N_5947);
nand U6830 (N_6830,N_5360,N_5094);
or U6831 (N_6831,N_4950,N_5784);
nor U6832 (N_6832,N_5602,N_5683);
nand U6833 (N_6833,N_5991,N_4592);
xor U6834 (N_6834,N_4690,N_5757);
nor U6835 (N_6835,N_5848,N_4932);
nand U6836 (N_6836,N_5818,N_4834);
nand U6837 (N_6837,N_4508,N_4810);
xnor U6838 (N_6838,N_4344,N_5536);
or U6839 (N_6839,N_5964,N_5138);
nand U6840 (N_6840,N_5123,N_4013);
or U6841 (N_6841,N_5458,N_4531);
or U6842 (N_6842,N_4192,N_4771);
nor U6843 (N_6843,N_4581,N_5615);
and U6844 (N_6844,N_4767,N_5234);
xor U6845 (N_6845,N_5143,N_5343);
and U6846 (N_6846,N_4534,N_5196);
and U6847 (N_6847,N_4716,N_5064);
nand U6848 (N_6848,N_4550,N_5827);
xnor U6849 (N_6849,N_4373,N_4336);
nand U6850 (N_6850,N_4097,N_4715);
and U6851 (N_6851,N_5988,N_4473);
or U6852 (N_6852,N_5619,N_5645);
or U6853 (N_6853,N_4446,N_4906);
nor U6854 (N_6854,N_4438,N_4154);
nand U6855 (N_6855,N_4136,N_4528);
xor U6856 (N_6856,N_5950,N_5698);
nor U6857 (N_6857,N_5242,N_5548);
xor U6858 (N_6858,N_4163,N_4901);
xor U6859 (N_6859,N_4223,N_5756);
and U6860 (N_6860,N_4137,N_5436);
or U6861 (N_6861,N_5637,N_4856);
or U6862 (N_6862,N_4918,N_4641);
and U6863 (N_6863,N_4417,N_5103);
and U6864 (N_6864,N_5640,N_5406);
xor U6865 (N_6865,N_5552,N_5326);
and U6866 (N_6866,N_5507,N_5953);
xor U6867 (N_6867,N_5152,N_4569);
or U6868 (N_6868,N_4813,N_4839);
and U6869 (N_6869,N_4138,N_4202);
nand U6870 (N_6870,N_5614,N_4441);
xor U6871 (N_6871,N_4892,N_4375);
and U6872 (N_6872,N_4499,N_4636);
and U6873 (N_6873,N_5730,N_4633);
and U6874 (N_6874,N_4957,N_5948);
and U6875 (N_6875,N_5471,N_4073);
or U6876 (N_6876,N_4358,N_4393);
or U6877 (N_6877,N_5709,N_4881);
nor U6878 (N_6878,N_5861,N_4992);
or U6879 (N_6879,N_5327,N_4521);
and U6880 (N_6880,N_4668,N_4655);
nand U6881 (N_6881,N_5264,N_5397);
or U6882 (N_6882,N_5425,N_4440);
nor U6883 (N_6883,N_4475,N_5862);
xor U6884 (N_6884,N_5963,N_5310);
xnor U6885 (N_6885,N_4048,N_4186);
and U6886 (N_6886,N_5010,N_5053);
and U6887 (N_6887,N_5670,N_4179);
and U6888 (N_6888,N_4035,N_5869);
xnor U6889 (N_6889,N_5907,N_5258);
and U6890 (N_6890,N_4308,N_4193);
nand U6891 (N_6891,N_5762,N_4525);
and U6892 (N_6892,N_5202,N_4430);
xnor U6893 (N_6893,N_4735,N_5714);
or U6894 (N_6894,N_5142,N_5508);
nand U6895 (N_6895,N_5371,N_4197);
or U6896 (N_6896,N_5385,N_5786);
or U6897 (N_6897,N_4713,N_4420);
nor U6898 (N_6898,N_5739,N_4062);
nor U6899 (N_6899,N_4849,N_4579);
nand U6900 (N_6900,N_4313,N_4017);
xor U6901 (N_6901,N_5100,N_4609);
or U6902 (N_6902,N_4924,N_4582);
or U6903 (N_6903,N_4378,N_4540);
nor U6904 (N_6904,N_5650,N_4181);
or U6905 (N_6905,N_4092,N_5926);
nor U6906 (N_6906,N_5992,N_4496);
nor U6907 (N_6907,N_5375,N_4126);
and U6908 (N_6908,N_4679,N_4805);
xnor U6909 (N_6909,N_4623,N_4574);
xnor U6910 (N_6910,N_4683,N_4802);
nor U6911 (N_6911,N_4045,N_4282);
or U6912 (N_6912,N_4653,N_5694);
or U6913 (N_6913,N_4678,N_5633);
and U6914 (N_6914,N_5909,N_5306);
and U6915 (N_6915,N_5887,N_4238);
or U6916 (N_6916,N_4283,N_4674);
nor U6917 (N_6917,N_4549,N_4207);
and U6918 (N_6918,N_4951,N_4144);
xor U6919 (N_6919,N_4919,N_5883);
or U6920 (N_6920,N_4720,N_4747);
or U6921 (N_6921,N_4656,N_5801);
and U6922 (N_6922,N_5710,N_5649);
and U6923 (N_6923,N_4236,N_4166);
and U6924 (N_6924,N_5770,N_4026);
or U6925 (N_6925,N_5740,N_5345);
nor U6926 (N_6926,N_5516,N_4756);
nor U6927 (N_6927,N_5768,N_4452);
xnor U6928 (N_6928,N_4089,N_5020);
nand U6929 (N_6929,N_5314,N_4843);
and U6930 (N_6930,N_4871,N_4456);
and U6931 (N_6931,N_4445,N_5456);
or U6932 (N_6932,N_4324,N_5365);
nor U6933 (N_6933,N_4775,N_4115);
nand U6934 (N_6934,N_4325,N_5376);
xnor U6935 (N_6935,N_4285,N_5475);
xor U6936 (N_6936,N_5419,N_5921);
xnor U6937 (N_6937,N_4190,N_4659);
nand U6938 (N_6938,N_4760,N_5294);
nand U6939 (N_6939,N_4080,N_4514);
nand U6940 (N_6940,N_4695,N_5434);
or U6941 (N_6941,N_5511,N_4337);
or U6942 (N_6942,N_4809,N_5268);
and U6943 (N_6943,N_4559,N_4803);
nor U6944 (N_6944,N_5814,N_4050);
xnor U6945 (N_6945,N_5232,N_4688);
and U6946 (N_6946,N_4998,N_5183);
nand U6947 (N_6947,N_5126,N_5467);
or U6948 (N_6948,N_5193,N_4502);
nor U6949 (N_6949,N_5189,N_5361);
or U6950 (N_6950,N_4815,N_5488);
or U6951 (N_6951,N_5606,N_5578);
and U6952 (N_6952,N_5322,N_5076);
and U6953 (N_6953,N_5542,N_4151);
and U6954 (N_6954,N_5502,N_4443);
and U6955 (N_6955,N_5622,N_4732);
xor U6956 (N_6956,N_4602,N_5636);
or U6957 (N_6957,N_5111,N_5156);
xnor U6958 (N_6958,N_4675,N_4955);
xnor U6959 (N_6959,N_4493,N_5396);
and U6960 (N_6960,N_5290,N_5056);
nor U6961 (N_6961,N_5703,N_4622);
and U6962 (N_6962,N_5461,N_5426);
nor U6963 (N_6963,N_5421,N_5751);
and U6964 (N_6964,N_5225,N_4405);
or U6965 (N_6965,N_4886,N_4831);
or U6966 (N_6966,N_4009,N_5356);
nor U6967 (N_6967,N_5673,N_4969);
and U6968 (N_6968,N_4410,N_5525);
and U6969 (N_6969,N_5828,N_5025);
or U6970 (N_6970,N_5316,N_4819);
xor U6971 (N_6971,N_4522,N_5249);
nand U6972 (N_6972,N_5354,N_5246);
and U6973 (N_6973,N_4022,N_4188);
and U6974 (N_6974,N_5392,N_5629);
nor U6975 (N_6975,N_5495,N_4872);
nand U6976 (N_6976,N_4797,N_4191);
nor U6977 (N_6977,N_4392,N_4374);
nor U6978 (N_6978,N_4717,N_4936);
and U6979 (N_6979,N_4660,N_5826);
and U6980 (N_6980,N_4644,N_5587);
xnor U6981 (N_6981,N_4920,N_5366);
or U6982 (N_6982,N_5923,N_5172);
and U6983 (N_6983,N_5194,N_4302);
xor U6984 (N_6984,N_4328,N_4455);
or U6985 (N_6985,N_5638,N_5060);
xnor U6986 (N_6986,N_4620,N_5259);
or U6987 (N_6987,N_4294,N_4379);
nor U6988 (N_6988,N_4997,N_5254);
and U6989 (N_6989,N_5357,N_5729);
or U6990 (N_6990,N_5789,N_5538);
nor U6991 (N_6991,N_4250,N_4034);
nor U6992 (N_6992,N_4637,N_5865);
nor U6993 (N_6993,N_5161,N_4627);
nand U6994 (N_6994,N_5938,N_4503);
xor U6995 (N_6995,N_5135,N_4723);
and U6996 (N_6996,N_4038,N_5482);
and U6997 (N_6997,N_4612,N_4706);
or U6998 (N_6998,N_4008,N_5091);
xor U6999 (N_6999,N_4403,N_5961);
xor U7000 (N_7000,N_4414,N_4070);
nor U7001 (N_7001,N_5661,N_4735);
or U7002 (N_7002,N_5279,N_5687);
or U7003 (N_7003,N_4716,N_4216);
and U7004 (N_7004,N_4233,N_5859);
nand U7005 (N_7005,N_5107,N_5879);
and U7006 (N_7006,N_4358,N_4629);
xor U7007 (N_7007,N_5714,N_5804);
nand U7008 (N_7008,N_5751,N_4415);
nand U7009 (N_7009,N_5250,N_4676);
xor U7010 (N_7010,N_4757,N_4655);
and U7011 (N_7011,N_4297,N_5443);
nor U7012 (N_7012,N_5941,N_5609);
xnor U7013 (N_7013,N_4638,N_4204);
xnor U7014 (N_7014,N_5886,N_5591);
nor U7015 (N_7015,N_4573,N_4791);
nor U7016 (N_7016,N_5639,N_4587);
nor U7017 (N_7017,N_4748,N_4836);
and U7018 (N_7018,N_4936,N_5636);
xnor U7019 (N_7019,N_5593,N_4296);
nor U7020 (N_7020,N_4889,N_5330);
and U7021 (N_7021,N_4001,N_4176);
nor U7022 (N_7022,N_4049,N_4289);
xnor U7023 (N_7023,N_4055,N_4610);
or U7024 (N_7024,N_5028,N_5106);
nor U7025 (N_7025,N_5939,N_5054);
or U7026 (N_7026,N_5721,N_5975);
and U7027 (N_7027,N_5909,N_4600);
nand U7028 (N_7028,N_4826,N_5618);
xnor U7029 (N_7029,N_4209,N_5493);
and U7030 (N_7030,N_5647,N_4256);
and U7031 (N_7031,N_4215,N_5545);
nand U7032 (N_7032,N_4498,N_5107);
nand U7033 (N_7033,N_5847,N_4028);
and U7034 (N_7034,N_4379,N_5573);
nor U7035 (N_7035,N_4706,N_5902);
or U7036 (N_7036,N_5342,N_5014);
and U7037 (N_7037,N_5900,N_5556);
nand U7038 (N_7038,N_5131,N_5003);
nand U7039 (N_7039,N_4195,N_4286);
nand U7040 (N_7040,N_4531,N_4645);
xor U7041 (N_7041,N_4995,N_4182);
xor U7042 (N_7042,N_5829,N_5303);
and U7043 (N_7043,N_5439,N_4499);
xor U7044 (N_7044,N_5600,N_4299);
xor U7045 (N_7045,N_5819,N_5483);
or U7046 (N_7046,N_5940,N_5759);
xor U7047 (N_7047,N_5599,N_5808);
or U7048 (N_7048,N_5265,N_5991);
or U7049 (N_7049,N_4770,N_4140);
or U7050 (N_7050,N_5593,N_5899);
nor U7051 (N_7051,N_4403,N_5527);
nor U7052 (N_7052,N_4994,N_4775);
or U7053 (N_7053,N_4985,N_5501);
nor U7054 (N_7054,N_4583,N_5876);
nand U7055 (N_7055,N_4853,N_4788);
nand U7056 (N_7056,N_4392,N_4586);
xnor U7057 (N_7057,N_4362,N_4398);
nand U7058 (N_7058,N_5453,N_4376);
nor U7059 (N_7059,N_5275,N_4809);
or U7060 (N_7060,N_5392,N_4717);
xnor U7061 (N_7061,N_5211,N_5193);
and U7062 (N_7062,N_4964,N_4545);
and U7063 (N_7063,N_5395,N_4580);
xnor U7064 (N_7064,N_4556,N_4174);
nor U7065 (N_7065,N_5091,N_5575);
xor U7066 (N_7066,N_4908,N_4528);
xor U7067 (N_7067,N_5443,N_5369);
xnor U7068 (N_7068,N_5146,N_5623);
nor U7069 (N_7069,N_4510,N_5091);
nand U7070 (N_7070,N_4123,N_5405);
and U7071 (N_7071,N_4262,N_4059);
and U7072 (N_7072,N_5035,N_5755);
and U7073 (N_7073,N_5583,N_4763);
xor U7074 (N_7074,N_5285,N_5358);
and U7075 (N_7075,N_5955,N_4790);
xnor U7076 (N_7076,N_5531,N_4228);
xnor U7077 (N_7077,N_5386,N_5250);
nor U7078 (N_7078,N_5285,N_4858);
xnor U7079 (N_7079,N_5820,N_4754);
nand U7080 (N_7080,N_4586,N_5328);
xnor U7081 (N_7081,N_4729,N_5032);
nor U7082 (N_7082,N_5732,N_4353);
or U7083 (N_7083,N_5656,N_5020);
nor U7084 (N_7084,N_5394,N_4225);
and U7085 (N_7085,N_4746,N_5872);
xnor U7086 (N_7086,N_4726,N_5612);
xor U7087 (N_7087,N_4043,N_4002);
nor U7088 (N_7088,N_4938,N_5116);
or U7089 (N_7089,N_5663,N_5245);
and U7090 (N_7090,N_5568,N_5482);
nor U7091 (N_7091,N_4996,N_5218);
xor U7092 (N_7092,N_4376,N_5268);
nand U7093 (N_7093,N_5040,N_4742);
xor U7094 (N_7094,N_4800,N_4172);
nor U7095 (N_7095,N_5353,N_5398);
nor U7096 (N_7096,N_5015,N_4541);
or U7097 (N_7097,N_4766,N_4108);
nor U7098 (N_7098,N_5437,N_4412);
xor U7099 (N_7099,N_5902,N_4240);
xor U7100 (N_7100,N_5132,N_4495);
or U7101 (N_7101,N_4158,N_5300);
and U7102 (N_7102,N_5311,N_4571);
and U7103 (N_7103,N_5447,N_4472);
nor U7104 (N_7104,N_5428,N_5184);
and U7105 (N_7105,N_4675,N_4222);
nand U7106 (N_7106,N_5141,N_4699);
xor U7107 (N_7107,N_4432,N_4437);
xnor U7108 (N_7108,N_5290,N_5498);
and U7109 (N_7109,N_4107,N_4197);
and U7110 (N_7110,N_5542,N_5397);
nor U7111 (N_7111,N_5430,N_5099);
and U7112 (N_7112,N_5458,N_5847);
nor U7113 (N_7113,N_4145,N_5522);
xnor U7114 (N_7114,N_4576,N_5339);
and U7115 (N_7115,N_5484,N_4147);
or U7116 (N_7116,N_5050,N_4228);
and U7117 (N_7117,N_5422,N_4802);
or U7118 (N_7118,N_5777,N_5237);
or U7119 (N_7119,N_5884,N_5265);
nand U7120 (N_7120,N_5654,N_4689);
or U7121 (N_7121,N_5711,N_4713);
nor U7122 (N_7122,N_5683,N_5817);
and U7123 (N_7123,N_4291,N_4690);
nand U7124 (N_7124,N_4548,N_4698);
nand U7125 (N_7125,N_4501,N_4180);
xnor U7126 (N_7126,N_5634,N_5832);
nor U7127 (N_7127,N_4913,N_5452);
nor U7128 (N_7128,N_5490,N_4256);
xor U7129 (N_7129,N_5779,N_5361);
nand U7130 (N_7130,N_5235,N_4254);
and U7131 (N_7131,N_4002,N_4211);
xor U7132 (N_7132,N_4664,N_4073);
nor U7133 (N_7133,N_4792,N_4781);
nor U7134 (N_7134,N_4632,N_5870);
or U7135 (N_7135,N_5187,N_4077);
xnor U7136 (N_7136,N_4881,N_5595);
xnor U7137 (N_7137,N_4744,N_5016);
or U7138 (N_7138,N_4512,N_5942);
nor U7139 (N_7139,N_5879,N_5474);
and U7140 (N_7140,N_4599,N_5635);
xnor U7141 (N_7141,N_4713,N_4272);
and U7142 (N_7142,N_4217,N_4307);
or U7143 (N_7143,N_4780,N_4541);
or U7144 (N_7144,N_4319,N_4129);
nor U7145 (N_7145,N_5776,N_5321);
xor U7146 (N_7146,N_4842,N_4587);
nor U7147 (N_7147,N_5251,N_5200);
nor U7148 (N_7148,N_4550,N_4564);
and U7149 (N_7149,N_5077,N_4874);
nand U7150 (N_7150,N_4246,N_4783);
or U7151 (N_7151,N_5809,N_4175);
xnor U7152 (N_7152,N_5374,N_4736);
xor U7153 (N_7153,N_4759,N_4762);
or U7154 (N_7154,N_5191,N_4666);
xor U7155 (N_7155,N_4702,N_4437);
nand U7156 (N_7156,N_5983,N_5453);
or U7157 (N_7157,N_4739,N_5573);
nor U7158 (N_7158,N_5187,N_5597);
nor U7159 (N_7159,N_4160,N_5626);
nand U7160 (N_7160,N_4165,N_4761);
xnor U7161 (N_7161,N_4617,N_5887);
or U7162 (N_7162,N_5639,N_4341);
or U7163 (N_7163,N_4456,N_5582);
nand U7164 (N_7164,N_5581,N_4339);
nor U7165 (N_7165,N_5458,N_5386);
or U7166 (N_7166,N_4898,N_5669);
and U7167 (N_7167,N_5486,N_4618);
or U7168 (N_7168,N_5551,N_4139);
and U7169 (N_7169,N_5873,N_4105);
nand U7170 (N_7170,N_4453,N_5208);
nor U7171 (N_7171,N_5399,N_4545);
nand U7172 (N_7172,N_4571,N_4573);
and U7173 (N_7173,N_4819,N_4613);
nor U7174 (N_7174,N_4223,N_4458);
nand U7175 (N_7175,N_4723,N_4139);
xnor U7176 (N_7176,N_5832,N_4313);
or U7177 (N_7177,N_4625,N_4369);
or U7178 (N_7178,N_4712,N_5310);
and U7179 (N_7179,N_5757,N_5542);
xor U7180 (N_7180,N_4815,N_5465);
or U7181 (N_7181,N_4267,N_5417);
or U7182 (N_7182,N_4975,N_5250);
nor U7183 (N_7183,N_5897,N_5323);
xor U7184 (N_7184,N_5026,N_4644);
nor U7185 (N_7185,N_4454,N_4666);
nand U7186 (N_7186,N_4888,N_5533);
or U7187 (N_7187,N_4793,N_5261);
nor U7188 (N_7188,N_5027,N_4279);
nand U7189 (N_7189,N_4240,N_4644);
xnor U7190 (N_7190,N_5681,N_5028);
and U7191 (N_7191,N_4485,N_4869);
nand U7192 (N_7192,N_5197,N_4342);
nor U7193 (N_7193,N_5095,N_4801);
nand U7194 (N_7194,N_4995,N_4313);
nand U7195 (N_7195,N_5392,N_5468);
nor U7196 (N_7196,N_4175,N_4618);
and U7197 (N_7197,N_5098,N_5885);
nor U7198 (N_7198,N_5220,N_5125);
and U7199 (N_7199,N_5475,N_5756);
and U7200 (N_7200,N_4471,N_4811);
and U7201 (N_7201,N_4594,N_4441);
nor U7202 (N_7202,N_4004,N_5311);
nor U7203 (N_7203,N_4778,N_5489);
nand U7204 (N_7204,N_4122,N_5298);
nor U7205 (N_7205,N_5713,N_4249);
xnor U7206 (N_7206,N_5747,N_4391);
nor U7207 (N_7207,N_5187,N_5267);
or U7208 (N_7208,N_5979,N_4211);
or U7209 (N_7209,N_5666,N_5218);
or U7210 (N_7210,N_5122,N_5154);
nor U7211 (N_7211,N_5158,N_4684);
or U7212 (N_7212,N_4372,N_4704);
nand U7213 (N_7213,N_5142,N_4513);
nand U7214 (N_7214,N_4332,N_5147);
xnor U7215 (N_7215,N_4601,N_5329);
or U7216 (N_7216,N_4122,N_4579);
xnor U7217 (N_7217,N_4151,N_4291);
or U7218 (N_7218,N_4962,N_5883);
nor U7219 (N_7219,N_4672,N_5009);
nand U7220 (N_7220,N_5148,N_5086);
and U7221 (N_7221,N_5035,N_5918);
or U7222 (N_7222,N_4869,N_5176);
xor U7223 (N_7223,N_5058,N_4354);
and U7224 (N_7224,N_4197,N_5927);
and U7225 (N_7225,N_4877,N_4517);
or U7226 (N_7226,N_4663,N_5527);
nand U7227 (N_7227,N_4330,N_4494);
nor U7228 (N_7228,N_5650,N_4235);
and U7229 (N_7229,N_5005,N_5894);
and U7230 (N_7230,N_4047,N_4103);
and U7231 (N_7231,N_5178,N_4164);
xnor U7232 (N_7232,N_4450,N_5144);
or U7233 (N_7233,N_5881,N_4683);
or U7234 (N_7234,N_5266,N_4405);
or U7235 (N_7235,N_5585,N_4743);
nand U7236 (N_7236,N_5156,N_4226);
nand U7237 (N_7237,N_4454,N_4023);
nor U7238 (N_7238,N_5622,N_5755);
or U7239 (N_7239,N_5703,N_5995);
and U7240 (N_7240,N_4847,N_4256);
nand U7241 (N_7241,N_5500,N_4182);
or U7242 (N_7242,N_4468,N_5440);
nor U7243 (N_7243,N_5724,N_5470);
or U7244 (N_7244,N_4251,N_5122);
nor U7245 (N_7245,N_4827,N_4519);
nor U7246 (N_7246,N_5877,N_5429);
nor U7247 (N_7247,N_4225,N_4748);
and U7248 (N_7248,N_5646,N_5459);
or U7249 (N_7249,N_5539,N_4257);
or U7250 (N_7250,N_5071,N_5093);
and U7251 (N_7251,N_5370,N_4680);
nand U7252 (N_7252,N_5028,N_5718);
nor U7253 (N_7253,N_5262,N_4531);
or U7254 (N_7254,N_4838,N_4699);
nor U7255 (N_7255,N_4700,N_5004);
nand U7256 (N_7256,N_5434,N_4198);
nand U7257 (N_7257,N_4263,N_5895);
nand U7258 (N_7258,N_5832,N_4355);
xnor U7259 (N_7259,N_5921,N_4484);
xor U7260 (N_7260,N_5667,N_5899);
nand U7261 (N_7261,N_4991,N_4600);
xor U7262 (N_7262,N_5437,N_5144);
nand U7263 (N_7263,N_5467,N_5902);
nor U7264 (N_7264,N_4676,N_4282);
xnor U7265 (N_7265,N_4608,N_4309);
nand U7266 (N_7266,N_5523,N_5918);
xnor U7267 (N_7267,N_5362,N_5758);
or U7268 (N_7268,N_5296,N_4931);
nor U7269 (N_7269,N_4169,N_5937);
nor U7270 (N_7270,N_5570,N_5702);
or U7271 (N_7271,N_4854,N_5625);
or U7272 (N_7272,N_5075,N_4891);
or U7273 (N_7273,N_4185,N_5058);
or U7274 (N_7274,N_5529,N_5020);
nand U7275 (N_7275,N_4931,N_4029);
xor U7276 (N_7276,N_4654,N_4841);
nor U7277 (N_7277,N_4486,N_5965);
nand U7278 (N_7278,N_5864,N_4454);
nor U7279 (N_7279,N_5735,N_5333);
and U7280 (N_7280,N_5491,N_5673);
and U7281 (N_7281,N_5941,N_4318);
xnor U7282 (N_7282,N_4503,N_4217);
nor U7283 (N_7283,N_4434,N_4782);
nor U7284 (N_7284,N_4135,N_5495);
xnor U7285 (N_7285,N_4613,N_5874);
and U7286 (N_7286,N_5917,N_5114);
or U7287 (N_7287,N_5076,N_4512);
xor U7288 (N_7288,N_4133,N_4112);
xnor U7289 (N_7289,N_5188,N_5061);
xnor U7290 (N_7290,N_4673,N_4708);
and U7291 (N_7291,N_4841,N_5111);
and U7292 (N_7292,N_4223,N_5033);
xor U7293 (N_7293,N_4633,N_4166);
xnor U7294 (N_7294,N_5980,N_5430);
or U7295 (N_7295,N_4412,N_4171);
and U7296 (N_7296,N_5721,N_4080);
and U7297 (N_7297,N_5320,N_5427);
nand U7298 (N_7298,N_5916,N_5883);
or U7299 (N_7299,N_5586,N_5321);
xor U7300 (N_7300,N_4549,N_5073);
nand U7301 (N_7301,N_5033,N_5763);
nor U7302 (N_7302,N_5851,N_5222);
and U7303 (N_7303,N_5428,N_4645);
xor U7304 (N_7304,N_4313,N_4789);
xnor U7305 (N_7305,N_5606,N_5229);
or U7306 (N_7306,N_4639,N_5427);
and U7307 (N_7307,N_4273,N_5726);
and U7308 (N_7308,N_4493,N_5732);
nor U7309 (N_7309,N_4293,N_5795);
or U7310 (N_7310,N_5160,N_4904);
or U7311 (N_7311,N_5826,N_5778);
nor U7312 (N_7312,N_4187,N_4036);
nand U7313 (N_7313,N_5385,N_4277);
or U7314 (N_7314,N_5742,N_5015);
and U7315 (N_7315,N_5519,N_5628);
or U7316 (N_7316,N_4127,N_5678);
nor U7317 (N_7317,N_4816,N_4436);
nor U7318 (N_7318,N_5194,N_4167);
nand U7319 (N_7319,N_4360,N_5352);
nand U7320 (N_7320,N_5293,N_4673);
xnor U7321 (N_7321,N_5147,N_5849);
nand U7322 (N_7322,N_5340,N_5915);
or U7323 (N_7323,N_5683,N_5803);
nand U7324 (N_7324,N_4602,N_4642);
xnor U7325 (N_7325,N_5709,N_4271);
nand U7326 (N_7326,N_5624,N_5194);
nor U7327 (N_7327,N_4778,N_5332);
xnor U7328 (N_7328,N_4503,N_4307);
xor U7329 (N_7329,N_4054,N_5536);
and U7330 (N_7330,N_4892,N_5451);
and U7331 (N_7331,N_5447,N_5942);
or U7332 (N_7332,N_5600,N_4072);
xnor U7333 (N_7333,N_4328,N_4220);
nor U7334 (N_7334,N_5570,N_4815);
or U7335 (N_7335,N_5374,N_5001);
xnor U7336 (N_7336,N_4102,N_4426);
and U7337 (N_7337,N_5894,N_4645);
or U7338 (N_7338,N_5909,N_5871);
or U7339 (N_7339,N_5922,N_4686);
nand U7340 (N_7340,N_5303,N_5414);
nand U7341 (N_7341,N_5882,N_5709);
or U7342 (N_7342,N_5259,N_4731);
nor U7343 (N_7343,N_4786,N_5288);
xor U7344 (N_7344,N_4237,N_4275);
and U7345 (N_7345,N_4263,N_5794);
nor U7346 (N_7346,N_5806,N_4950);
and U7347 (N_7347,N_5355,N_4281);
and U7348 (N_7348,N_4638,N_4347);
and U7349 (N_7349,N_5516,N_5651);
nor U7350 (N_7350,N_4824,N_5631);
xor U7351 (N_7351,N_4538,N_5894);
nor U7352 (N_7352,N_5253,N_4426);
xor U7353 (N_7353,N_4197,N_5870);
and U7354 (N_7354,N_5512,N_4035);
xnor U7355 (N_7355,N_4222,N_4256);
and U7356 (N_7356,N_4379,N_5203);
xnor U7357 (N_7357,N_5535,N_4446);
nor U7358 (N_7358,N_4123,N_5744);
nand U7359 (N_7359,N_4061,N_4823);
and U7360 (N_7360,N_4196,N_5288);
or U7361 (N_7361,N_4869,N_5045);
and U7362 (N_7362,N_4517,N_4483);
and U7363 (N_7363,N_4753,N_4569);
and U7364 (N_7364,N_4121,N_4954);
or U7365 (N_7365,N_4547,N_5884);
nor U7366 (N_7366,N_4790,N_4911);
nand U7367 (N_7367,N_4353,N_4970);
nor U7368 (N_7368,N_4448,N_4995);
and U7369 (N_7369,N_5473,N_5937);
xnor U7370 (N_7370,N_5479,N_5553);
nand U7371 (N_7371,N_5943,N_4208);
xnor U7372 (N_7372,N_5538,N_5360);
and U7373 (N_7373,N_5983,N_4395);
nand U7374 (N_7374,N_4605,N_5447);
nand U7375 (N_7375,N_4685,N_4642);
nor U7376 (N_7376,N_4305,N_5361);
xnor U7377 (N_7377,N_5790,N_5652);
nor U7378 (N_7378,N_4393,N_5829);
nand U7379 (N_7379,N_4794,N_5437);
and U7380 (N_7380,N_4711,N_5510);
nand U7381 (N_7381,N_5251,N_5572);
and U7382 (N_7382,N_5167,N_4121);
xnor U7383 (N_7383,N_4356,N_5913);
and U7384 (N_7384,N_5423,N_4234);
xor U7385 (N_7385,N_4815,N_4722);
nor U7386 (N_7386,N_4944,N_4432);
and U7387 (N_7387,N_5639,N_4698);
nand U7388 (N_7388,N_5565,N_5575);
and U7389 (N_7389,N_4218,N_5558);
nand U7390 (N_7390,N_5047,N_5954);
nor U7391 (N_7391,N_4438,N_5188);
nand U7392 (N_7392,N_5679,N_5251);
or U7393 (N_7393,N_4752,N_4026);
and U7394 (N_7394,N_5564,N_5881);
nor U7395 (N_7395,N_5065,N_5591);
nand U7396 (N_7396,N_5829,N_5967);
and U7397 (N_7397,N_5786,N_5365);
xor U7398 (N_7398,N_5224,N_5197);
nor U7399 (N_7399,N_4104,N_4001);
xor U7400 (N_7400,N_5117,N_4275);
or U7401 (N_7401,N_5921,N_4188);
and U7402 (N_7402,N_4885,N_5880);
or U7403 (N_7403,N_5058,N_5075);
xor U7404 (N_7404,N_5880,N_5019);
and U7405 (N_7405,N_4367,N_5453);
nor U7406 (N_7406,N_5039,N_4067);
xor U7407 (N_7407,N_5701,N_4923);
nand U7408 (N_7408,N_5675,N_4019);
and U7409 (N_7409,N_4785,N_4387);
nand U7410 (N_7410,N_4313,N_5933);
nor U7411 (N_7411,N_4897,N_5243);
or U7412 (N_7412,N_5421,N_4808);
nand U7413 (N_7413,N_5055,N_5353);
and U7414 (N_7414,N_5624,N_5799);
nor U7415 (N_7415,N_5274,N_5764);
nor U7416 (N_7416,N_4886,N_4641);
and U7417 (N_7417,N_5389,N_5400);
nand U7418 (N_7418,N_4323,N_5567);
nand U7419 (N_7419,N_4868,N_5057);
xor U7420 (N_7420,N_5136,N_4760);
and U7421 (N_7421,N_5664,N_4367);
xor U7422 (N_7422,N_5951,N_4461);
xor U7423 (N_7423,N_5299,N_5213);
nand U7424 (N_7424,N_5124,N_4338);
and U7425 (N_7425,N_4915,N_4377);
and U7426 (N_7426,N_4248,N_5046);
nand U7427 (N_7427,N_4677,N_4719);
and U7428 (N_7428,N_4942,N_4734);
or U7429 (N_7429,N_4780,N_5540);
and U7430 (N_7430,N_5245,N_4109);
xor U7431 (N_7431,N_4315,N_4663);
nand U7432 (N_7432,N_5433,N_4935);
or U7433 (N_7433,N_5222,N_5766);
or U7434 (N_7434,N_4930,N_5421);
and U7435 (N_7435,N_4965,N_4835);
and U7436 (N_7436,N_4185,N_5733);
nor U7437 (N_7437,N_4379,N_5995);
xnor U7438 (N_7438,N_5085,N_4064);
nand U7439 (N_7439,N_4256,N_4172);
nor U7440 (N_7440,N_5235,N_5767);
and U7441 (N_7441,N_5139,N_4622);
xnor U7442 (N_7442,N_4884,N_5948);
and U7443 (N_7443,N_4922,N_4398);
and U7444 (N_7444,N_4866,N_5107);
xor U7445 (N_7445,N_4251,N_4082);
nand U7446 (N_7446,N_5640,N_4137);
nand U7447 (N_7447,N_4118,N_4661);
or U7448 (N_7448,N_4854,N_5431);
nand U7449 (N_7449,N_4727,N_4606);
or U7450 (N_7450,N_5236,N_5792);
or U7451 (N_7451,N_4395,N_5177);
or U7452 (N_7452,N_5217,N_4942);
xor U7453 (N_7453,N_5708,N_5797);
nor U7454 (N_7454,N_5187,N_5318);
and U7455 (N_7455,N_5369,N_5486);
xor U7456 (N_7456,N_5633,N_4004);
xor U7457 (N_7457,N_5839,N_4523);
nand U7458 (N_7458,N_5334,N_5955);
nor U7459 (N_7459,N_4468,N_5528);
and U7460 (N_7460,N_5495,N_5721);
nor U7461 (N_7461,N_4001,N_4665);
nor U7462 (N_7462,N_5777,N_5023);
xnor U7463 (N_7463,N_4803,N_4398);
xnor U7464 (N_7464,N_5817,N_4208);
or U7465 (N_7465,N_5606,N_4682);
and U7466 (N_7466,N_4598,N_4289);
nand U7467 (N_7467,N_4271,N_5407);
xnor U7468 (N_7468,N_5387,N_4626);
nand U7469 (N_7469,N_5542,N_4527);
nand U7470 (N_7470,N_4040,N_5222);
or U7471 (N_7471,N_4133,N_5454);
nor U7472 (N_7472,N_4946,N_4468);
nand U7473 (N_7473,N_4748,N_5645);
nor U7474 (N_7474,N_5205,N_4770);
xor U7475 (N_7475,N_5875,N_5365);
nand U7476 (N_7476,N_4917,N_4192);
or U7477 (N_7477,N_5198,N_4494);
and U7478 (N_7478,N_4986,N_4894);
and U7479 (N_7479,N_5626,N_4400);
xor U7480 (N_7480,N_5899,N_4261);
or U7481 (N_7481,N_5438,N_5856);
and U7482 (N_7482,N_4394,N_5657);
xor U7483 (N_7483,N_4490,N_4357);
nor U7484 (N_7484,N_4216,N_4338);
xnor U7485 (N_7485,N_5802,N_5162);
xor U7486 (N_7486,N_5598,N_5285);
xnor U7487 (N_7487,N_4546,N_4950);
or U7488 (N_7488,N_4152,N_5496);
nor U7489 (N_7489,N_4904,N_5046);
xor U7490 (N_7490,N_5272,N_5650);
xnor U7491 (N_7491,N_5116,N_4130);
and U7492 (N_7492,N_4969,N_4337);
and U7493 (N_7493,N_5878,N_4926);
nand U7494 (N_7494,N_5165,N_5164);
and U7495 (N_7495,N_5017,N_5609);
nand U7496 (N_7496,N_4056,N_4000);
nand U7497 (N_7497,N_5936,N_5157);
nand U7498 (N_7498,N_5162,N_5456);
and U7499 (N_7499,N_5121,N_5228);
and U7500 (N_7500,N_4915,N_4052);
or U7501 (N_7501,N_4123,N_4281);
and U7502 (N_7502,N_5282,N_5617);
xor U7503 (N_7503,N_5425,N_4269);
or U7504 (N_7504,N_5672,N_5496);
xor U7505 (N_7505,N_4999,N_4270);
xnor U7506 (N_7506,N_5997,N_4343);
or U7507 (N_7507,N_5236,N_4132);
or U7508 (N_7508,N_5263,N_4029);
and U7509 (N_7509,N_4664,N_4498);
xnor U7510 (N_7510,N_5689,N_5936);
or U7511 (N_7511,N_5208,N_5102);
nor U7512 (N_7512,N_5875,N_5281);
or U7513 (N_7513,N_4561,N_4338);
nand U7514 (N_7514,N_5999,N_4813);
nand U7515 (N_7515,N_5009,N_5925);
nor U7516 (N_7516,N_4880,N_5718);
or U7517 (N_7517,N_5923,N_5775);
nor U7518 (N_7518,N_5705,N_4679);
or U7519 (N_7519,N_4504,N_4298);
nor U7520 (N_7520,N_4821,N_4219);
or U7521 (N_7521,N_4521,N_5191);
nor U7522 (N_7522,N_4511,N_4376);
or U7523 (N_7523,N_5376,N_4785);
xor U7524 (N_7524,N_4709,N_5582);
or U7525 (N_7525,N_5229,N_5460);
and U7526 (N_7526,N_5629,N_4769);
nor U7527 (N_7527,N_4079,N_5865);
xor U7528 (N_7528,N_5614,N_4713);
nor U7529 (N_7529,N_4141,N_4632);
xor U7530 (N_7530,N_4343,N_5752);
or U7531 (N_7531,N_5314,N_5685);
xnor U7532 (N_7532,N_4861,N_5601);
and U7533 (N_7533,N_5068,N_5809);
nor U7534 (N_7534,N_5181,N_5975);
or U7535 (N_7535,N_4337,N_5917);
nand U7536 (N_7536,N_4568,N_4952);
xor U7537 (N_7537,N_5599,N_4041);
and U7538 (N_7538,N_5695,N_4946);
nor U7539 (N_7539,N_5409,N_5248);
nand U7540 (N_7540,N_5109,N_4437);
and U7541 (N_7541,N_4658,N_4942);
and U7542 (N_7542,N_4060,N_4699);
nand U7543 (N_7543,N_5234,N_5345);
nand U7544 (N_7544,N_5474,N_4154);
and U7545 (N_7545,N_5607,N_5451);
and U7546 (N_7546,N_4355,N_4707);
xor U7547 (N_7547,N_5264,N_4532);
nand U7548 (N_7548,N_5234,N_4246);
and U7549 (N_7549,N_5066,N_4747);
and U7550 (N_7550,N_4755,N_4674);
nand U7551 (N_7551,N_4956,N_5657);
xnor U7552 (N_7552,N_5786,N_5661);
nor U7553 (N_7553,N_5416,N_5762);
nand U7554 (N_7554,N_4719,N_4517);
or U7555 (N_7555,N_5394,N_4822);
xnor U7556 (N_7556,N_4709,N_4763);
and U7557 (N_7557,N_5284,N_4915);
xor U7558 (N_7558,N_4829,N_4179);
xor U7559 (N_7559,N_5548,N_5867);
xnor U7560 (N_7560,N_4650,N_4014);
xnor U7561 (N_7561,N_5923,N_5731);
or U7562 (N_7562,N_4504,N_4187);
nor U7563 (N_7563,N_4486,N_5709);
nor U7564 (N_7564,N_5075,N_4742);
or U7565 (N_7565,N_5298,N_5053);
xor U7566 (N_7566,N_5312,N_4486);
or U7567 (N_7567,N_4669,N_5864);
and U7568 (N_7568,N_5122,N_4686);
xnor U7569 (N_7569,N_5745,N_4847);
and U7570 (N_7570,N_4400,N_5603);
nand U7571 (N_7571,N_5288,N_5687);
and U7572 (N_7572,N_5878,N_4410);
or U7573 (N_7573,N_4921,N_5999);
and U7574 (N_7574,N_5865,N_5477);
nand U7575 (N_7575,N_4928,N_4709);
and U7576 (N_7576,N_5598,N_4752);
and U7577 (N_7577,N_4051,N_5421);
nand U7578 (N_7578,N_4795,N_5138);
and U7579 (N_7579,N_5458,N_4762);
and U7580 (N_7580,N_5841,N_5146);
nand U7581 (N_7581,N_4053,N_4196);
and U7582 (N_7582,N_4390,N_5069);
xnor U7583 (N_7583,N_5843,N_5597);
nor U7584 (N_7584,N_4600,N_5675);
nor U7585 (N_7585,N_5088,N_5019);
and U7586 (N_7586,N_5176,N_5465);
and U7587 (N_7587,N_4572,N_4405);
and U7588 (N_7588,N_5511,N_5010);
or U7589 (N_7589,N_5089,N_4048);
nand U7590 (N_7590,N_4119,N_4989);
and U7591 (N_7591,N_4290,N_4436);
or U7592 (N_7592,N_4794,N_5986);
xnor U7593 (N_7593,N_5046,N_5152);
nor U7594 (N_7594,N_4301,N_4395);
and U7595 (N_7595,N_4150,N_5681);
and U7596 (N_7596,N_4134,N_4059);
xor U7597 (N_7597,N_5656,N_4640);
or U7598 (N_7598,N_4410,N_5578);
nor U7599 (N_7599,N_4560,N_4758);
or U7600 (N_7600,N_4419,N_4258);
nand U7601 (N_7601,N_4411,N_5366);
nand U7602 (N_7602,N_5538,N_4203);
and U7603 (N_7603,N_5145,N_4377);
nand U7604 (N_7604,N_5779,N_5945);
and U7605 (N_7605,N_5972,N_5638);
and U7606 (N_7606,N_4587,N_4126);
xnor U7607 (N_7607,N_4219,N_4371);
and U7608 (N_7608,N_5100,N_5942);
xor U7609 (N_7609,N_5910,N_4958);
nor U7610 (N_7610,N_5639,N_5964);
nand U7611 (N_7611,N_5713,N_5962);
and U7612 (N_7612,N_4654,N_5777);
or U7613 (N_7613,N_5766,N_4379);
nand U7614 (N_7614,N_4353,N_5528);
nand U7615 (N_7615,N_5602,N_4933);
or U7616 (N_7616,N_5399,N_4288);
xor U7617 (N_7617,N_4636,N_5780);
or U7618 (N_7618,N_5725,N_4808);
nor U7619 (N_7619,N_5582,N_4338);
and U7620 (N_7620,N_5000,N_4177);
or U7621 (N_7621,N_4139,N_5963);
xnor U7622 (N_7622,N_5675,N_4971);
nor U7623 (N_7623,N_5560,N_5793);
nand U7624 (N_7624,N_4318,N_5890);
nor U7625 (N_7625,N_4219,N_4591);
and U7626 (N_7626,N_4822,N_4637);
nor U7627 (N_7627,N_4476,N_5953);
nor U7628 (N_7628,N_4425,N_5951);
and U7629 (N_7629,N_4767,N_4842);
xnor U7630 (N_7630,N_4657,N_5090);
and U7631 (N_7631,N_5647,N_5786);
and U7632 (N_7632,N_4753,N_4245);
and U7633 (N_7633,N_5377,N_5672);
nand U7634 (N_7634,N_4394,N_4873);
xor U7635 (N_7635,N_4717,N_5955);
nand U7636 (N_7636,N_4578,N_5084);
xor U7637 (N_7637,N_4329,N_4726);
nand U7638 (N_7638,N_5415,N_5998);
and U7639 (N_7639,N_5669,N_5307);
nor U7640 (N_7640,N_4260,N_5585);
nor U7641 (N_7641,N_5640,N_4706);
xnor U7642 (N_7642,N_4886,N_5919);
nor U7643 (N_7643,N_4728,N_4418);
nand U7644 (N_7644,N_4223,N_4326);
or U7645 (N_7645,N_5214,N_4658);
and U7646 (N_7646,N_5914,N_4115);
or U7647 (N_7647,N_4032,N_5986);
nor U7648 (N_7648,N_4105,N_5266);
xor U7649 (N_7649,N_5237,N_4010);
and U7650 (N_7650,N_5407,N_4643);
nor U7651 (N_7651,N_4219,N_5013);
or U7652 (N_7652,N_4393,N_5585);
xnor U7653 (N_7653,N_5152,N_4964);
xnor U7654 (N_7654,N_5633,N_5921);
nand U7655 (N_7655,N_4936,N_5368);
and U7656 (N_7656,N_5157,N_5071);
and U7657 (N_7657,N_4913,N_4497);
or U7658 (N_7658,N_5977,N_5248);
or U7659 (N_7659,N_5636,N_5385);
nand U7660 (N_7660,N_4253,N_5708);
xnor U7661 (N_7661,N_4125,N_4434);
nand U7662 (N_7662,N_4244,N_4820);
or U7663 (N_7663,N_5222,N_4401);
or U7664 (N_7664,N_4747,N_4454);
nor U7665 (N_7665,N_5464,N_4928);
and U7666 (N_7666,N_5352,N_4149);
xor U7667 (N_7667,N_4836,N_4463);
nor U7668 (N_7668,N_5343,N_5353);
nor U7669 (N_7669,N_4933,N_5405);
nor U7670 (N_7670,N_5173,N_5236);
and U7671 (N_7671,N_4498,N_4913);
and U7672 (N_7672,N_4251,N_5929);
nor U7673 (N_7673,N_4288,N_4552);
nor U7674 (N_7674,N_4181,N_5591);
nor U7675 (N_7675,N_5144,N_4864);
nor U7676 (N_7676,N_4420,N_5543);
and U7677 (N_7677,N_5494,N_5998);
nor U7678 (N_7678,N_5678,N_4451);
or U7679 (N_7679,N_4868,N_5486);
and U7680 (N_7680,N_4640,N_4184);
or U7681 (N_7681,N_5912,N_5052);
nand U7682 (N_7682,N_5293,N_5949);
or U7683 (N_7683,N_4624,N_5918);
and U7684 (N_7684,N_5552,N_4234);
or U7685 (N_7685,N_4027,N_5522);
nor U7686 (N_7686,N_4575,N_4459);
nand U7687 (N_7687,N_5030,N_4702);
nor U7688 (N_7688,N_5556,N_4304);
nand U7689 (N_7689,N_4901,N_5214);
nor U7690 (N_7690,N_4567,N_4312);
nor U7691 (N_7691,N_5477,N_5875);
or U7692 (N_7692,N_4535,N_5422);
xnor U7693 (N_7693,N_4552,N_5126);
nand U7694 (N_7694,N_4418,N_4595);
nor U7695 (N_7695,N_5530,N_4975);
and U7696 (N_7696,N_5010,N_5669);
and U7697 (N_7697,N_5509,N_5673);
or U7698 (N_7698,N_5380,N_4043);
nand U7699 (N_7699,N_5697,N_4293);
xnor U7700 (N_7700,N_5976,N_5855);
nand U7701 (N_7701,N_5680,N_4287);
xor U7702 (N_7702,N_4607,N_5859);
xor U7703 (N_7703,N_5647,N_5500);
or U7704 (N_7704,N_5594,N_5444);
nand U7705 (N_7705,N_5274,N_4946);
or U7706 (N_7706,N_5633,N_4450);
and U7707 (N_7707,N_5041,N_5397);
or U7708 (N_7708,N_4730,N_4813);
and U7709 (N_7709,N_4535,N_4280);
nor U7710 (N_7710,N_4990,N_4533);
or U7711 (N_7711,N_4703,N_4503);
nand U7712 (N_7712,N_5680,N_5435);
or U7713 (N_7713,N_4219,N_5455);
or U7714 (N_7714,N_5286,N_4390);
nand U7715 (N_7715,N_4813,N_5326);
nand U7716 (N_7716,N_4783,N_4101);
nor U7717 (N_7717,N_4028,N_5334);
or U7718 (N_7718,N_5713,N_4687);
nor U7719 (N_7719,N_4842,N_5648);
or U7720 (N_7720,N_4189,N_4318);
nand U7721 (N_7721,N_5792,N_4538);
nand U7722 (N_7722,N_5393,N_4344);
nand U7723 (N_7723,N_5194,N_4535);
and U7724 (N_7724,N_4909,N_4696);
or U7725 (N_7725,N_4536,N_4418);
nand U7726 (N_7726,N_4337,N_4749);
and U7727 (N_7727,N_4715,N_5863);
nand U7728 (N_7728,N_4164,N_5494);
and U7729 (N_7729,N_4430,N_4543);
nor U7730 (N_7730,N_5344,N_4530);
nand U7731 (N_7731,N_5790,N_5533);
and U7732 (N_7732,N_5423,N_5947);
nand U7733 (N_7733,N_4190,N_4361);
and U7734 (N_7734,N_5644,N_5023);
nor U7735 (N_7735,N_4440,N_4050);
xnor U7736 (N_7736,N_5241,N_5413);
xor U7737 (N_7737,N_4946,N_4709);
and U7738 (N_7738,N_5607,N_4615);
xnor U7739 (N_7739,N_4792,N_4996);
nor U7740 (N_7740,N_5814,N_4587);
nand U7741 (N_7741,N_5570,N_4589);
nand U7742 (N_7742,N_4663,N_4902);
nor U7743 (N_7743,N_5464,N_4044);
nor U7744 (N_7744,N_4095,N_4300);
and U7745 (N_7745,N_5975,N_4323);
nand U7746 (N_7746,N_4460,N_4758);
nand U7747 (N_7747,N_4175,N_4892);
nand U7748 (N_7748,N_4057,N_5965);
or U7749 (N_7749,N_4447,N_5518);
and U7750 (N_7750,N_5509,N_5833);
or U7751 (N_7751,N_4051,N_4129);
or U7752 (N_7752,N_4605,N_4398);
and U7753 (N_7753,N_5750,N_5446);
nor U7754 (N_7754,N_4429,N_4194);
nor U7755 (N_7755,N_5290,N_5324);
nand U7756 (N_7756,N_5534,N_4279);
nand U7757 (N_7757,N_5056,N_5893);
or U7758 (N_7758,N_5262,N_4652);
or U7759 (N_7759,N_5463,N_5197);
nand U7760 (N_7760,N_5102,N_4998);
and U7761 (N_7761,N_5450,N_4289);
nand U7762 (N_7762,N_4621,N_5791);
nor U7763 (N_7763,N_4369,N_5452);
nand U7764 (N_7764,N_4122,N_4439);
nand U7765 (N_7765,N_4075,N_5904);
and U7766 (N_7766,N_4863,N_4516);
and U7767 (N_7767,N_4438,N_4164);
and U7768 (N_7768,N_4978,N_5073);
or U7769 (N_7769,N_4343,N_4305);
or U7770 (N_7770,N_5660,N_4504);
or U7771 (N_7771,N_5006,N_4245);
nor U7772 (N_7772,N_5635,N_5079);
nand U7773 (N_7773,N_4003,N_4258);
or U7774 (N_7774,N_4683,N_4451);
xor U7775 (N_7775,N_5446,N_4279);
or U7776 (N_7776,N_5046,N_4783);
or U7777 (N_7777,N_4617,N_4629);
nor U7778 (N_7778,N_5349,N_5744);
nand U7779 (N_7779,N_5761,N_5260);
nand U7780 (N_7780,N_4754,N_4746);
xor U7781 (N_7781,N_4324,N_5181);
nor U7782 (N_7782,N_4329,N_5638);
or U7783 (N_7783,N_4251,N_5008);
xnor U7784 (N_7784,N_4055,N_5107);
or U7785 (N_7785,N_4887,N_5929);
nand U7786 (N_7786,N_5538,N_4531);
nor U7787 (N_7787,N_5482,N_4751);
or U7788 (N_7788,N_4583,N_4846);
nor U7789 (N_7789,N_4599,N_4361);
nor U7790 (N_7790,N_4581,N_5016);
nand U7791 (N_7791,N_5580,N_5846);
nand U7792 (N_7792,N_4219,N_5230);
or U7793 (N_7793,N_5510,N_5539);
nand U7794 (N_7794,N_4566,N_5416);
xor U7795 (N_7795,N_4878,N_5677);
xor U7796 (N_7796,N_4458,N_4462);
and U7797 (N_7797,N_5323,N_5569);
nand U7798 (N_7798,N_4376,N_4800);
or U7799 (N_7799,N_4242,N_5183);
xnor U7800 (N_7800,N_4226,N_5850);
and U7801 (N_7801,N_5135,N_5281);
and U7802 (N_7802,N_5625,N_4297);
nand U7803 (N_7803,N_5835,N_4151);
and U7804 (N_7804,N_4274,N_5260);
nor U7805 (N_7805,N_4736,N_5357);
and U7806 (N_7806,N_4718,N_5687);
nor U7807 (N_7807,N_4411,N_4927);
nor U7808 (N_7808,N_4454,N_5146);
or U7809 (N_7809,N_5484,N_5862);
and U7810 (N_7810,N_5520,N_5671);
nand U7811 (N_7811,N_5611,N_5147);
nor U7812 (N_7812,N_5924,N_5472);
or U7813 (N_7813,N_4794,N_4975);
and U7814 (N_7814,N_4661,N_4986);
xor U7815 (N_7815,N_5309,N_4727);
or U7816 (N_7816,N_5463,N_4877);
or U7817 (N_7817,N_4243,N_4817);
xnor U7818 (N_7818,N_5554,N_5083);
and U7819 (N_7819,N_5611,N_4918);
and U7820 (N_7820,N_5045,N_5626);
nand U7821 (N_7821,N_4957,N_5628);
or U7822 (N_7822,N_5370,N_4912);
xnor U7823 (N_7823,N_4193,N_4030);
and U7824 (N_7824,N_4426,N_4180);
or U7825 (N_7825,N_4211,N_4775);
or U7826 (N_7826,N_5714,N_5813);
nand U7827 (N_7827,N_4988,N_5776);
and U7828 (N_7828,N_5586,N_4743);
nor U7829 (N_7829,N_4092,N_5795);
nor U7830 (N_7830,N_5000,N_5919);
or U7831 (N_7831,N_4401,N_5577);
nor U7832 (N_7832,N_4024,N_4292);
nand U7833 (N_7833,N_5728,N_5134);
or U7834 (N_7834,N_5417,N_4549);
nor U7835 (N_7835,N_5339,N_4625);
and U7836 (N_7836,N_4045,N_5285);
nand U7837 (N_7837,N_5828,N_5253);
xnor U7838 (N_7838,N_4797,N_4307);
xnor U7839 (N_7839,N_5243,N_4653);
nor U7840 (N_7840,N_4339,N_4202);
xor U7841 (N_7841,N_4818,N_4236);
xnor U7842 (N_7842,N_4591,N_4872);
and U7843 (N_7843,N_5643,N_5449);
and U7844 (N_7844,N_5096,N_4467);
or U7845 (N_7845,N_4687,N_4832);
nor U7846 (N_7846,N_4499,N_4706);
nor U7847 (N_7847,N_5316,N_5760);
and U7848 (N_7848,N_4048,N_5022);
xor U7849 (N_7849,N_5789,N_5377);
or U7850 (N_7850,N_5347,N_5556);
xnor U7851 (N_7851,N_4536,N_4782);
nand U7852 (N_7852,N_5986,N_5108);
nor U7853 (N_7853,N_4999,N_4988);
and U7854 (N_7854,N_5771,N_4565);
nand U7855 (N_7855,N_4602,N_4036);
nand U7856 (N_7856,N_5546,N_4737);
xor U7857 (N_7857,N_5853,N_5427);
nor U7858 (N_7858,N_5081,N_4072);
xor U7859 (N_7859,N_4038,N_4428);
nor U7860 (N_7860,N_5149,N_4873);
nand U7861 (N_7861,N_4865,N_5082);
or U7862 (N_7862,N_4882,N_5259);
xor U7863 (N_7863,N_5478,N_4742);
or U7864 (N_7864,N_5929,N_4497);
xor U7865 (N_7865,N_4970,N_4275);
nor U7866 (N_7866,N_5950,N_5075);
or U7867 (N_7867,N_4742,N_5849);
or U7868 (N_7868,N_5999,N_5798);
nor U7869 (N_7869,N_5478,N_5376);
xor U7870 (N_7870,N_5706,N_4174);
xor U7871 (N_7871,N_4852,N_4402);
and U7872 (N_7872,N_5999,N_5486);
and U7873 (N_7873,N_4889,N_5672);
and U7874 (N_7874,N_5958,N_5093);
xnor U7875 (N_7875,N_4120,N_5274);
nor U7876 (N_7876,N_5501,N_4129);
and U7877 (N_7877,N_4175,N_4913);
nor U7878 (N_7878,N_4337,N_5706);
nor U7879 (N_7879,N_5530,N_4370);
or U7880 (N_7880,N_4850,N_4857);
or U7881 (N_7881,N_4208,N_4099);
xor U7882 (N_7882,N_4864,N_5926);
xnor U7883 (N_7883,N_4999,N_5729);
xor U7884 (N_7884,N_4437,N_4181);
or U7885 (N_7885,N_5326,N_4143);
and U7886 (N_7886,N_5413,N_4200);
and U7887 (N_7887,N_5422,N_5248);
nor U7888 (N_7888,N_5358,N_4357);
nor U7889 (N_7889,N_5590,N_5659);
nand U7890 (N_7890,N_5156,N_5514);
nor U7891 (N_7891,N_5980,N_4615);
and U7892 (N_7892,N_4198,N_5333);
or U7893 (N_7893,N_4371,N_5416);
nand U7894 (N_7894,N_4038,N_5842);
and U7895 (N_7895,N_5934,N_4758);
xnor U7896 (N_7896,N_4686,N_4354);
nand U7897 (N_7897,N_5178,N_4970);
or U7898 (N_7898,N_4963,N_4799);
and U7899 (N_7899,N_5619,N_4450);
and U7900 (N_7900,N_4248,N_4042);
or U7901 (N_7901,N_5017,N_5507);
xnor U7902 (N_7902,N_4292,N_5128);
and U7903 (N_7903,N_5848,N_5062);
nand U7904 (N_7904,N_4355,N_4043);
nand U7905 (N_7905,N_5296,N_5615);
or U7906 (N_7906,N_4974,N_5184);
or U7907 (N_7907,N_4694,N_5990);
or U7908 (N_7908,N_4932,N_5242);
nor U7909 (N_7909,N_4404,N_5907);
nor U7910 (N_7910,N_4067,N_5656);
nand U7911 (N_7911,N_4593,N_4733);
xnor U7912 (N_7912,N_4692,N_4052);
and U7913 (N_7913,N_4300,N_4617);
and U7914 (N_7914,N_5573,N_5078);
nand U7915 (N_7915,N_4573,N_4480);
or U7916 (N_7916,N_4686,N_5514);
and U7917 (N_7917,N_4896,N_4445);
nand U7918 (N_7918,N_4810,N_5420);
nor U7919 (N_7919,N_4799,N_5292);
and U7920 (N_7920,N_4109,N_5252);
xor U7921 (N_7921,N_4860,N_5496);
nand U7922 (N_7922,N_4118,N_4616);
nor U7923 (N_7923,N_4330,N_4794);
xor U7924 (N_7924,N_4514,N_5897);
nor U7925 (N_7925,N_4104,N_4291);
and U7926 (N_7926,N_4928,N_5180);
nor U7927 (N_7927,N_4391,N_5988);
xnor U7928 (N_7928,N_5737,N_5179);
or U7929 (N_7929,N_4028,N_4123);
or U7930 (N_7930,N_5672,N_4558);
nand U7931 (N_7931,N_4825,N_4574);
nand U7932 (N_7932,N_4303,N_5362);
xor U7933 (N_7933,N_4416,N_4286);
nor U7934 (N_7934,N_4527,N_5550);
or U7935 (N_7935,N_4334,N_4882);
nand U7936 (N_7936,N_5715,N_5246);
and U7937 (N_7937,N_5585,N_4931);
or U7938 (N_7938,N_4608,N_4724);
xnor U7939 (N_7939,N_4086,N_5080);
or U7940 (N_7940,N_4502,N_5451);
nor U7941 (N_7941,N_5682,N_5852);
or U7942 (N_7942,N_4890,N_4097);
and U7943 (N_7943,N_4862,N_4754);
nand U7944 (N_7944,N_5685,N_4700);
nor U7945 (N_7945,N_5358,N_4253);
xnor U7946 (N_7946,N_5481,N_5737);
nand U7947 (N_7947,N_5075,N_5343);
xnor U7948 (N_7948,N_5202,N_5062);
nand U7949 (N_7949,N_5888,N_4906);
xnor U7950 (N_7950,N_4183,N_5925);
and U7951 (N_7951,N_4478,N_5159);
and U7952 (N_7952,N_4037,N_5434);
or U7953 (N_7953,N_5234,N_4184);
nor U7954 (N_7954,N_4639,N_4334);
or U7955 (N_7955,N_5853,N_4561);
nor U7956 (N_7956,N_5685,N_4325);
and U7957 (N_7957,N_4594,N_4952);
or U7958 (N_7958,N_5818,N_4908);
or U7959 (N_7959,N_5141,N_5939);
xnor U7960 (N_7960,N_5988,N_5286);
nand U7961 (N_7961,N_4759,N_4901);
or U7962 (N_7962,N_4754,N_5536);
and U7963 (N_7963,N_4579,N_5519);
and U7964 (N_7964,N_5861,N_5205);
nand U7965 (N_7965,N_5830,N_5268);
and U7966 (N_7966,N_4443,N_5584);
nand U7967 (N_7967,N_5556,N_4140);
and U7968 (N_7968,N_5635,N_4901);
and U7969 (N_7969,N_4942,N_4427);
and U7970 (N_7970,N_5678,N_4462);
xor U7971 (N_7971,N_5858,N_4018);
nand U7972 (N_7972,N_4002,N_4403);
or U7973 (N_7973,N_4790,N_5079);
or U7974 (N_7974,N_4697,N_4815);
nor U7975 (N_7975,N_5322,N_4454);
and U7976 (N_7976,N_5424,N_5200);
and U7977 (N_7977,N_5545,N_4464);
nor U7978 (N_7978,N_5907,N_5659);
nor U7979 (N_7979,N_5641,N_5002);
xor U7980 (N_7980,N_5644,N_5407);
and U7981 (N_7981,N_4672,N_5773);
or U7982 (N_7982,N_5091,N_4933);
nand U7983 (N_7983,N_4436,N_4806);
nand U7984 (N_7984,N_5547,N_4440);
xnor U7985 (N_7985,N_4983,N_5222);
nand U7986 (N_7986,N_5290,N_5604);
or U7987 (N_7987,N_5120,N_5492);
xnor U7988 (N_7988,N_5945,N_4160);
nor U7989 (N_7989,N_4742,N_4257);
or U7990 (N_7990,N_4299,N_5631);
nor U7991 (N_7991,N_4246,N_5751);
nor U7992 (N_7992,N_5645,N_5766);
nand U7993 (N_7993,N_5204,N_4612);
or U7994 (N_7994,N_4225,N_5657);
nor U7995 (N_7995,N_5868,N_5350);
nor U7996 (N_7996,N_5457,N_5598);
nor U7997 (N_7997,N_4885,N_4367);
nor U7998 (N_7998,N_4309,N_4270);
nor U7999 (N_7999,N_5157,N_4318);
xor U8000 (N_8000,N_7003,N_7442);
or U8001 (N_8001,N_6774,N_7853);
or U8002 (N_8002,N_6164,N_6423);
xor U8003 (N_8003,N_6606,N_7649);
xnor U8004 (N_8004,N_7790,N_6247);
xnor U8005 (N_8005,N_6386,N_7400);
nand U8006 (N_8006,N_6492,N_7960);
or U8007 (N_8007,N_7584,N_6540);
xnor U8008 (N_8008,N_7633,N_6822);
and U8009 (N_8009,N_7217,N_7388);
and U8010 (N_8010,N_7177,N_6958);
or U8011 (N_8011,N_6017,N_6257);
nor U8012 (N_8012,N_7076,N_7865);
xor U8013 (N_8013,N_7377,N_6404);
xnor U8014 (N_8014,N_6767,N_7618);
xnor U8015 (N_8015,N_6996,N_6148);
xor U8016 (N_8016,N_7834,N_7372);
xor U8017 (N_8017,N_7472,N_6376);
nand U8018 (N_8018,N_6915,N_6782);
or U8019 (N_8019,N_6760,N_7815);
and U8020 (N_8020,N_6664,N_6648);
and U8021 (N_8021,N_7830,N_6738);
or U8022 (N_8022,N_7084,N_7260);
or U8023 (N_8023,N_6904,N_6413);
xor U8024 (N_8024,N_6117,N_7765);
and U8025 (N_8025,N_7926,N_6443);
nor U8026 (N_8026,N_6687,N_7886);
nor U8027 (N_8027,N_7548,N_6455);
xor U8028 (N_8028,N_7513,N_7857);
nand U8029 (N_8029,N_6133,N_6512);
and U8030 (N_8030,N_6937,N_6167);
or U8031 (N_8031,N_6088,N_7862);
xnor U8032 (N_8032,N_7007,N_6977);
xnor U8033 (N_8033,N_7892,N_7957);
and U8034 (N_8034,N_6861,N_6938);
xor U8035 (N_8035,N_7622,N_6106);
nor U8036 (N_8036,N_6182,N_7060);
or U8037 (N_8037,N_7360,N_7514);
nand U8038 (N_8038,N_6896,N_6297);
or U8039 (N_8039,N_7778,N_6195);
xnor U8040 (N_8040,N_6199,N_6175);
xor U8041 (N_8041,N_7574,N_7030);
nand U8042 (N_8042,N_7614,N_7565);
xor U8043 (N_8043,N_7329,N_7215);
or U8044 (N_8044,N_7621,N_7443);
nor U8045 (N_8045,N_7594,N_6322);
nor U8046 (N_8046,N_6038,N_7365);
nand U8047 (N_8047,N_6976,N_7236);
nor U8048 (N_8048,N_7698,N_6342);
and U8049 (N_8049,N_7558,N_6232);
or U8050 (N_8050,N_6672,N_7560);
or U8051 (N_8051,N_6373,N_7688);
xnor U8052 (N_8052,N_6995,N_6962);
nand U8053 (N_8053,N_6029,N_7160);
and U8054 (N_8054,N_6170,N_6629);
nor U8055 (N_8055,N_6523,N_7982);
xor U8056 (N_8056,N_6318,N_7283);
or U8057 (N_8057,N_6266,N_6625);
nor U8058 (N_8058,N_7635,N_7937);
xor U8059 (N_8059,N_7351,N_6168);
nor U8060 (N_8060,N_6281,N_6790);
nor U8061 (N_8061,N_6985,N_6589);
or U8062 (N_8062,N_6713,N_7879);
xnor U8063 (N_8063,N_6476,N_7952);
nand U8064 (N_8064,N_7122,N_6360);
nand U8065 (N_8065,N_7252,N_7569);
nand U8066 (N_8066,N_6399,N_6803);
and U8067 (N_8067,N_6426,N_7014);
or U8068 (N_8068,N_6953,N_7034);
nor U8069 (N_8069,N_7304,N_6220);
nand U8070 (N_8070,N_7518,N_7657);
nand U8071 (N_8071,N_7470,N_7191);
or U8072 (N_8072,N_6372,N_6341);
nand U8073 (N_8073,N_6216,N_6747);
or U8074 (N_8074,N_7495,N_7451);
and U8075 (N_8075,N_7093,N_7496);
nand U8076 (N_8076,N_7972,N_7728);
and U8077 (N_8077,N_7586,N_7025);
nand U8078 (N_8078,N_6115,N_7298);
nand U8079 (N_8079,N_7146,N_6223);
or U8080 (N_8080,N_6273,N_6241);
or U8081 (N_8081,N_7918,N_7804);
nand U8082 (N_8082,N_7666,N_7132);
or U8083 (N_8083,N_6789,N_6152);
nand U8084 (N_8084,N_6003,N_7978);
and U8085 (N_8085,N_6946,N_7747);
nand U8086 (N_8086,N_7411,N_6569);
xor U8087 (N_8087,N_7224,N_6974);
nor U8088 (N_8088,N_7986,N_6181);
xor U8089 (N_8089,N_7788,N_7955);
xnor U8090 (N_8090,N_6304,N_7038);
and U8091 (N_8091,N_6661,N_7259);
or U8092 (N_8092,N_6296,N_6428);
or U8093 (N_8093,N_6650,N_7282);
nand U8094 (N_8094,N_7017,N_6440);
and U8095 (N_8095,N_7683,N_7433);
nor U8096 (N_8096,N_7350,N_6781);
xor U8097 (N_8097,N_6514,N_7416);
xnor U8098 (N_8098,N_6303,N_6327);
or U8099 (N_8099,N_6785,N_7418);
nand U8100 (N_8100,N_7032,N_6603);
and U8101 (N_8101,N_6993,N_7202);
and U8102 (N_8102,N_6353,N_7602);
and U8103 (N_8103,N_7846,N_6343);
and U8104 (N_8104,N_7041,N_6775);
or U8105 (N_8105,N_7860,N_7627);
and U8106 (N_8106,N_7968,N_6513);
nand U8107 (N_8107,N_6936,N_7048);
and U8108 (N_8108,N_6599,N_6555);
xor U8109 (N_8109,N_6809,N_7992);
or U8110 (N_8110,N_6808,N_7225);
nand U8111 (N_8111,N_6464,N_6568);
nand U8112 (N_8112,N_6483,N_6082);
xnor U8113 (N_8113,N_7634,N_7258);
and U8114 (N_8114,N_6224,N_7254);
and U8115 (N_8115,N_6971,N_7744);
nand U8116 (N_8116,N_6816,N_7151);
and U8117 (N_8117,N_6312,N_6352);
nor U8118 (N_8118,N_7150,N_6330);
nand U8119 (N_8119,N_6099,N_7587);
or U8120 (N_8120,N_6856,N_7425);
nand U8121 (N_8121,N_7381,N_6132);
and U8122 (N_8122,N_7042,N_7953);
nor U8123 (N_8123,N_6313,N_6729);
and U8124 (N_8124,N_6592,N_7000);
nor U8125 (N_8125,N_7813,N_6897);
xor U8126 (N_8126,N_6023,N_7534);
and U8127 (N_8127,N_7616,N_7553);
or U8128 (N_8128,N_6157,N_7674);
and U8129 (N_8129,N_7148,N_6588);
xnor U8130 (N_8130,N_6584,N_7168);
and U8131 (N_8131,N_7913,N_6585);
or U8132 (N_8132,N_6316,N_7905);
or U8133 (N_8133,N_6145,N_6143);
xor U8134 (N_8134,N_6005,N_6609);
or U8135 (N_8135,N_6300,N_6931);
nor U8136 (N_8136,N_6965,N_6979);
and U8137 (N_8137,N_6255,N_7228);
nor U8138 (N_8138,N_6138,N_7783);
and U8139 (N_8139,N_6587,N_6722);
xor U8140 (N_8140,N_7803,N_6857);
nor U8141 (N_8141,N_7682,N_7091);
xor U8142 (N_8142,N_6048,N_6825);
xor U8143 (N_8143,N_6642,N_7625);
and U8144 (N_8144,N_6819,N_7904);
and U8145 (N_8145,N_7467,N_6626);
and U8146 (N_8146,N_7178,N_7863);
xor U8147 (N_8147,N_7916,N_7872);
xnor U8148 (N_8148,N_6154,N_6004);
or U8149 (N_8149,N_7592,N_6100);
nor U8150 (N_8150,N_6914,N_7535);
xor U8151 (N_8151,N_7566,N_7099);
nand U8152 (N_8152,N_7339,N_7741);
or U8153 (N_8153,N_7531,N_7510);
and U8154 (N_8154,N_6689,N_6185);
or U8155 (N_8155,N_6743,N_6955);
xor U8156 (N_8156,N_6957,N_6545);
and U8157 (N_8157,N_6449,N_7907);
xnor U8158 (N_8158,N_6416,N_7998);
nand U8159 (N_8159,N_7573,N_6524);
nand U8160 (N_8160,N_7869,N_6668);
nor U8161 (N_8161,N_6470,N_7071);
or U8162 (N_8162,N_6657,N_6007);
nor U8163 (N_8163,N_7476,N_6260);
nor U8164 (N_8164,N_6293,N_7727);
nor U8165 (N_8165,N_6594,N_6261);
and U8166 (N_8166,N_6102,N_7811);
xnor U8167 (N_8167,N_6471,N_6705);
or U8168 (N_8168,N_6410,N_6282);
nand U8169 (N_8169,N_6405,N_7367);
or U8170 (N_8170,N_6579,N_7434);
xor U8171 (N_8171,N_6395,N_7735);
nand U8172 (N_8172,N_6206,N_6299);
nand U8173 (N_8173,N_6964,N_6961);
nand U8174 (N_8174,N_6806,N_6541);
nand U8175 (N_8175,N_7988,N_6735);
xor U8176 (N_8176,N_6285,N_7662);
nand U8177 (N_8177,N_7948,N_7082);
and U8178 (N_8178,N_7250,N_7393);
nand U8179 (N_8179,N_6120,N_7423);
nor U8180 (N_8180,N_6187,N_7792);
and U8181 (N_8181,N_6800,N_6051);
nor U8182 (N_8182,N_6277,N_7827);
or U8183 (N_8183,N_6928,N_6639);
nand U8184 (N_8184,N_7340,N_6338);
or U8185 (N_8185,N_7800,N_7361);
or U8186 (N_8186,N_6892,N_6901);
and U8187 (N_8187,N_7873,N_6876);
nor U8188 (N_8188,N_7711,N_6383);
xnor U8189 (N_8189,N_7094,N_6786);
and U8190 (N_8190,N_7113,N_7563);
and U8191 (N_8191,N_6880,N_7519);
nor U8192 (N_8192,N_7248,N_7856);
nor U8193 (N_8193,N_7319,N_6848);
xor U8194 (N_8194,N_7723,N_6254);
nand U8195 (N_8195,N_6717,N_6250);
and U8196 (N_8196,N_7737,N_6994);
xnor U8197 (N_8197,N_7922,N_6403);
or U8198 (N_8198,N_7874,N_6918);
xnor U8199 (N_8199,N_6814,N_6991);
or U8200 (N_8200,N_7058,N_7362);
nor U8201 (N_8201,N_6943,N_6539);
or U8202 (N_8202,N_7687,N_6560);
or U8203 (N_8203,N_7703,N_7753);
xor U8204 (N_8204,N_6675,N_6022);
nand U8205 (N_8205,N_6952,N_7516);
nor U8206 (N_8206,N_7110,N_6577);
nand U8207 (N_8207,N_6565,N_7305);
or U8208 (N_8208,N_7368,N_6724);
nor U8209 (N_8209,N_6114,N_6663);
and U8210 (N_8210,N_7520,N_6150);
nand U8211 (N_8211,N_7095,N_7855);
xor U8212 (N_8212,N_6497,N_6721);
xor U8213 (N_8213,N_6110,N_7709);
nor U8214 (N_8214,N_7129,N_6796);
xor U8215 (N_8215,N_7257,N_7983);
or U8216 (N_8216,N_7161,N_6496);
nor U8217 (N_8217,N_6354,N_6611);
nand U8218 (N_8218,N_7100,N_6841);
and U8219 (N_8219,N_7130,N_7775);
nor U8220 (N_8220,N_7581,N_6001);
or U8221 (N_8221,N_6718,N_7359);
nand U8222 (N_8222,N_6368,N_7175);
and U8223 (N_8223,N_6791,N_7133);
nand U8224 (N_8224,N_6845,N_6380);
nand U8225 (N_8225,N_7655,N_7890);
or U8226 (N_8226,N_7118,N_6381);
and U8227 (N_8227,N_7432,N_7567);
xor U8228 (N_8228,N_6667,N_6046);
and U8229 (N_8229,N_7936,N_6863);
and U8230 (N_8230,N_7457,N_6212);
nand U8231 (N_8231,N_7426,N_7836);
nor U8232 (N_8232,N_7525,N_7200);
xor U8233 (N_8233,N_7664,N_7600);
nor U8234 (N_8234,N_6094,N_6369);
and U8235 (N_8235,N_7826,N_7522);
nor U8236 (N_8236,N_7773,N_6419);
nor U8237 (N_8237,N_6367,N_6484);
and U8238 (N_8238,N_6923,N_6548);
nor U8239 (N_8239,N_7185,N_6475);
nand U8240 (N_8240,N_6479,N_7090);
nand U8241 (N_8241,N_6235,N_6549);
and U8242 (N_8242,N_6087,N_6425);
and U8243 (N_8243,N_7256,N_6927);
nor U8244 (N_8244,N_6502,N_6888);
xnor U8245 (N_8245,N_7067,N_7139);
or U8246 (N_8246,N_6163,N_6018);
nor U8247 (N_8247,N_6093,N_7291);
xor U8248 (N_8248,N_6237,N_7170);
and U8249 (N_8249,N_6495,N_6509);
or U8250 (N_8250,N_6446,N_7288);
nor U8251 (N_8251,N_7754,N_7849);
or U8252 (N_8252,N_7341,N_6109);
nor U8253 (N_8253,N_7552,N_6238);
and U8254 (N_8254,N_7537,N_6086);
xnor U8255 (N_8255,N_7669,N_7375);
or U8256 (N_8256,N_6628,N_7561);
xor U8257 (N_8257,N_7240,N_7821);
xnor U8258 (N_8258,N_6151,N_6983);
or U8259 (N_8259,N_7736,N_7493);
xor U8260 (N_8260,N_7578,N_6008);
nand U8261 (N_8261,N_7541,N_6695);
and U8262 (N_8262,N_6391,N_7412);
xnor U8263 (N_8263,N_7019,N_6614);
or U8264 (N_8264,N_7290,N_6634);
or U8265 (N_8265,N_7123,N_6412);
or U8266 (N_8266,N_6337,N_7712);
nand U8267 (N_8267,N_7508,N_6144);
nand U8268 (N_8268,N_7689,N_6477);
or U8269 (N_8269,N_7546,N_7352);
nor U8270 (N_8270,N_7239,N_6456);
xor U8271 (N_8271,N_7731,N_6838);
or U8272 (N_8272,N_6457,N_7805);
nand U8273 (N_8273,N_6417,N_6101);
and U8274 (N_8274,N_7387,N_7061);
xnor U8275 (N_8275,N_7384,N_6392);
nand U8276 (N_8276,N_6503,N_6286);
nand U8277 (N_8277,N_6956,N_6068);
xnor U8278 (N_8278,N_7956,N_6287);
or U8279 (N_8279,N_6319,N_7987);
nand U8280 (N_8280,N_6486,N_7121);
nor U8281 (N_8281,N_6111,N_7029);
and U8282 (N_8282,N_7422,N_6314);
or U8283 (N_8283,N_7023,N_6720);
nor U8284 (N_8284,N_7392,N_6044);
nand U8285 (N_8285,N_7929,N_7624);
or U8286 (N_8286,N_7613,N_6184);
xnor U8287 (N_8287,N_6362,N_7571);
or U8288 (N_8288,N_7464,N_7994);
or U8289 (N_8289,N_6619,N_7278);
nor U8290 (N_8290,N_7866,N_6610);
xor U8291 (N_8291,N_7538,N_7167);
xor U8292 (N_8292,N_6894,N_7509);
nor U8293 (N_8293,N_7149,N_6307);
nor U8294 (N_8294,N_6968,N_7701);
and U8295 (N_8295,N_6649,N_6990);
or U8296 (N_8296,N_7162,N_7889);
or U8297 (N_8297,N_6409,N_7763);
or U8298 (N_8298,N_7072,N_7066);
xor U8299 (N_8299,N_7801,N_6079);
or U8300 (N_8300,N_7532,N_7734);
or U8301 (N_8301,N_7414,N_6561);
or U8302 (N_8302,N_6732,N_7626);
and U8303 (N_8303,N_6701,N_7771);
nand U8304 (N_8304,N_6128,N_6518);
nor U8305 (N_8305,N_7906,N_7745);
nor U8306 (N_8306,N_6351,N_6234);
and U8307 (N_8307,N_6877,N_7715);
xor U8308 (N_8308,N_7272,N_7658);
nor U8309 (N_8309,N_7249,N_7310);
xor U8310 (N_8310,N_6700,N_6719);
or U8311 (N_8311,N_7762,N_7793);
xor U8312 (N_8312,N_6836,N_7279);
xor U8313 (N_8313,N_7659,N_7394);
nand U8314 (N_8314,N_7446,N_6014);
and U8315 (N_8315,N_7297,N_7124);
or U8316 (N_8316,N_7458,N_7164);
nor U8317 (N_8317,N_6766,N_7366);
nand U8318 (N_8318,N_6842,N_7995);
and U8319 (N_8319,N_6728,N_7979);
or U8320 (N_8320,N_6658,N_7852);
and U8321 (N_8321,N_6393,N_7229);
and U8322 (N_8322,N_6834,N_7511);
xor U8323 (N_8323,N_7065,N_7833);
nor U8324 (N_8324,N_6792,N_7219);
xnor U8325 (N_8325,N_6349,N_6229);
or U8326 (N_8326,N_7544,N_7222);
nor U8327 (N_8327,N_6306,N_7266);
or U8328 (N_8328,N_6978,N_6815);
nand U8329 (N_8329,N_7647,N_6414);
nand U8330 (N_8330,N_6358,N_6580);
or U8331 (N_8331,N_7932,N_6438);
and U8332 (N_8332,N_7410,N_6704);
or U8333 (N_8333,N_7925,N_7596);
xnor U8334 (N_8334,N_6744,N_7812);
nor U8335 (N_8335,N_7115,N_7742);
nand U8336 (N_8336,N_7299,N_7027);
nand U8337 (N_8337,N_7501,N_7880);
and U8338 (N_8338,N_6777,N_7105);
and U8339 (N_8339,N_6214,N_7631);
and U8340 (N_8340,N_7606,N_6301);
or U8341 (N_8341,N_6010,N_7996);
xor U8342 (N_8342,N_7981,N_7453);
or U8343 (N_8343,N_6450,N_6058);
or U8344 (N_8344,N_6715,N_7894);
nor U8345 (N_8345,N_6315,N_6666);
nor U8346 (N_8346,N_6105,N_7088);
nand U8347 (N_8347,N_6481,N_6630);
nor U8348 (N_8348,N_6334,N_7172);
xnor U8349 (N_8349,N_7335,N_7895);
xor U8350 (N_8350,N_7136,N_6552);
nand U8351 (N_8351,N_7656,N_7902);
or U8352 (N_8352,N_6291,N_7026);
nor U8353 (N_8353,N_7636,N_6252);
and U8354 (N_8354,N_6573,N_7840);
nor U8355 (N_8355,N_7246,N_7308);
and U8356 (N_8356,N_6787,N_7818);
nor U8357 (N_8357,N_7764,N_6849);
and U8358 (N_8358,N_6253,N_6180);
nand U8359 (N_8359,N_6275,N_6544);
nand U8360 (N_8360,N_6467,N_6890);
or U8361 (N_8361,N_7238,N_7802);
nor U8362 (N_8362,N_7106,N_7370);
nand U8363 (N_8363,N_6294,N_7369);
nand U8364 (N_8364,N_6770,N_6829);
or U8365 (N_8365,N_6156,N_7749);
and U8366 (N_8366,N_7171,N_7678);
and U8367 (N_8367,N_7331,N_7280);
nor U8368 (N_8368,N_6067,N_6908);
nand U8369 (N_8369,N_7439,N_6601);
nor U8370 (N_8370,N_7967,N_6116);
nor U8371 (N_8371,N_6763,N_7975);
nor U8372 (N_8372,N_7379,N_7796);
xor U8373 (N_8373,N_6759,N_7112);
and U8374 (N_8374,N_6274,N_6272);
nand U8375 (N_8375,N_7214,N_6853);
or U8376 (N_8376,N_7490,N_7482);
xor U8377 (N_8377,N_7402,N_6171);
and U8378 (N_8378,N_7730,N_7134);
and U8379 (N_8379,N_7022,N_6696);
nand U8380 (N_8380,N_7407,N_6948);
xnor U8381 (N_8381,N_6903,N_7009);
xor U8382 (N_8382,N_6525,N_7469);
and U8383 (N_8383,N_6563,N_7449);
nor U8384 (N_8384,N_6246,N_6574);
or U8385 (N_8385,N_7062,N_6060);
and U8386 (N_8386,N_7896,N_7864);
or U8387 (N_8387,N_7323,N_7403);
and U8388 (N_8388,N_6726,N_6289);
nor U8389 (N_8389,N_6651,N_6325);
and U8390 (N_8390,N_7440,N_7502);
nand U8391 (N_8391,N_7670,N_7216);
and U8392 (N_8392,N_6571,N_6828);
nand U8393 (N_8393,N_6269,N_7914);
and U8394 (N_8394,N_7884,N_6427);
nor U8395 (N_8395,N_6487,N_7054);
nand U8396 (N_8396,N_6783,N_7585);
and U8397 (N_8397,N_7477,N_7582);
nor U8398 (N_8398,N_7770,N_6802);
xnor U8399 (N_8399,N_6041,N_6714);
nor U8400 (N_8400,N_7642,N_6681);
and U8401 (N_8401,N_7119,N_7390);
or U8402 (N_8402,N_6632,N_7244);
and U8403 (N_8403,N_7938,N_6531);
or U8404 (N_8404,N_7004,N_6776);
or U8405 (N_8405,N_6702,N_7506);
nor U8406 (N_8406,N_6207,N_6424);
or U8407 (N_8407,N_6934,N_6075);
xnor U8408 (N_8408,N_6764,N_7499);
nand U8409 (N_8409,N_6329,N_7980);
xnor U8410 (N_8410,N_7623,N_6134);
or U8411 (N_8411,N_6799,N_7317);
nand U8412 (N_8412,N_6895,N_6685);
or U8413 (N_8413,N_7523,N_7611);
or U8414 (N_8414,N_6462,N_7590);
or U8415 (N_8415,N_7144,N_7958);
or U8416 (N_8416,N_7485,N_7312);
and U8417 (N_8417,N_7145,N_7740);
nand U8418 (N_8418,N_7281,N_7521);
and U8419 (N_8419,N_6429,N_6846);
nor U8420 (N_8420,N_6244,N_7718);
and U8421 (N_8421,N_6731,N_6081);
nor U8422 (N_8422,N_6543,N_6448);
nor U8423 (N_8423,N_7111,N_7868);
or U8424 (N_8424,N_6501,N_7756);
xnor U8425 (N_8425,N_7823,N_7315);
nand U8426 (N_8426,N_6118,N_6401);
xnor U8427 (N_8427,N_7463,N_6750);
or U8428 (N_8428,N_6056,N_7210);
xor U8429 (N_8429,N_7448,N_6375);
and U8430 (N_8430,N_7679,N_6966);
and U8431 (N_8431,N_6711,N_6420);
or U8432 (N_8432,N_6366,N_6872);
nand U8433 (N_8433,N_7924,N_7719);
or U8434 (N_8434,N_6878,N_7181);
xnor U8435 (N_8435,N_6998,N_7651);
xor U8436 (N_8436,N_6737,N_6478);
nor U8437 (N_8437,N_7713,N_6902);
nand U8438 (N_8438,N_7640,N_7069);
xor U8439 (N_8439,N_6465,N_6408);
or U8440 (N_8440,N_7031,N_6442);
nor U8441 (N_8441,N_6177,N_6365);
nor U8442 (N_8442,N_6122,N_7057);
and U8443 (N_8443,N_6941,N_7555);
and U8444 (N_8444,N_6925,N_6745);
xor U8445 (N_8445,N_7841,N_6640);
nor U8446 (N_8446,N_7013,N_7292);
xnor U8447 (N_8447,N_7505,N_6546);
xnor U8448 (N_8448,N_6139,N_6454);
and U8449 (N_8449,N_7269,N_6582);
nor U8450 (N_8450,N_7504,N_6499);
xor U8451 (N_8451,N_6169,N_7660);
or U8452 (N_8452,N_6875,N_6485);
xor U8453 (N_8453,N_7438,N_7699);
nor U8454 (N_8454,N_7908,N_7005);
or U8455 (N_8455,N_6665,N_6891);
and U8456 (N_8456,N_6027,N_6521);
nor U8457 (N_8457,N_7743,N_6248);
nand U8458 (N_8458,N_7053,N_6359);
nor U8459 (N_8459,N_6371,N_7706);
nor U8460 (N_8460,N_7708,N_7166);
xor U8461 (N_8461,N_7417,N_6510);
nand U8462 (N_8462,N_7819,N_7714);
xor U8463 (N_8463,N_7646,N_7475);
nor U8464 (N_8464,N_6959,N_6765);
xnor U8465 (N_8465,N_7524,N_7990);
or U8466 (N_8466,N_6336,N_6221);
nand U8467 (N_8467,N_7073,N_7309);
nor U8468 (N_8468,N_7615,N_7915);
nor U8469 (N_8469,N_6581,N_7489);
and U8470 (N_8470,N_7445,N_6859);
or U8471 (N_8471,N_6703,N_7720);
xor U8472 (N_8472,N_6335,N_7338);
or U8473 (N_8473,N_7944,N_7081);
nand U8474 (N_8474,N_6140,N_6204);
or U8475 (N_8475,N_6707,N_6647);
xor U8476 (N_8476,N_7055,N_6203);
xor U8477 (N_8477,N_7243,N_6862);
nand U8478 (N_8478,N_7398,N_7012);
and U8479 (N_8479,N_7404,N_6604);
xnor U8480 (N_8480,N_6070,N_6388);
and U8481 (N_8481,N_7461,N_6166);
xor U8482 (N_8482,N_7389,N_6797);
nor U8483 (N_8483,N_6328,N_7933);
nand U8484 (N_8484,N_6988,N_7630);
nor U8485 (N_8485,N_6437,N_7809);
or U8486 (N_8486,N_6095,N_6921);
nor U8487 (N_8487,N_6951,N_6141);
xor U8488 (N_8488,N_6520,N_6762);
and U8489 (N_8489,N_6473,N_6679);
xnor U8490 (N_8490,N_7854,N_7748);
and U8491 (N_8491,N_6490,N_6680);
nand U8492 (N_8492,N_7492,N_7786);
or U8493 (N_8493,N_6062,N_7010);
xnor U8494 (N_8494,N_7421,N_6500);
nor U8495 (N_8495,N_7676,N_7087);
nand U8496 (N_8496,N_7861,N_6769);
nor U8497 (N_8497,N_6772,N_6239);
nor U8498 (N_8498,N_6635,N_6542);
nor U8499 (N_8499,N_7702,N_6034);
and U8500 (N_8500,N_7568,N_7301);
nand U8501 (N_8501,N_7126,N_7080);
nand U8502 (N_8502,N_6305,N_6910);
nor U8503 (N_8503,N_7966,N_7479);
nor U8504 (N_8504,N_6554,N_7086);
xnor U8505 (N_8505,N_7314,N_7816);
nand U8506 (N_8506,N_6407,N_7002);
and U8507 (N_8507,N_7935,N_7233);
and U8508 (N_8508,N_7580,N_7320);
nand U8509 (N_8509,N_6071,N_7313);
and U8510 (N_8510,N_6489,N_7900);
nor U8511 (N_8511,N_7188,N_7406);
and U8512 (N_8512,N_7638,N_7491);
and U8513 (N_8513,N_6378,N_7083);
or U8514 (N_8514,N_6159,N_7887);
nor U8515 (N_8515,N_6472,N_7074);
or U8516 (N_8516,N_7722,N_6522);
nand U8517 (N_8517,N_7194,N_6989);
and U8518 (N_8518,N_6411,N_7549);
and U8519 (N_8519,N_6740,N_6033);
and U8520 (N_8520,N_6655,N_6137);
and U8521 (N_8521,N_6659,N_7295);
nor U8522 (N_8522,N_7044,N_6259);
and U8523 (N_8523,N_6669,N_7104);
nand U8524 (N_8524,N_6126,N_6215);
nor U8525 (N_8525,N_6432,N_7456);
and U8526 (N_8526,N_7693,N_6992);
nor U8527 (N_8527,N_7355,N_7668);
nand U8528 (N_8528,N_7364,N_7294);
nor U8529 (N_8529,N_6227,N_6466);
and U8530 (N_8530,N_7893,N_7620);
nand U8531 (N_8531,N_6085,N_6645);
xnor U8532 (N_8532,N_6256,N_6055);
nand U8533 (N_8533,N_7311,N_6865);
nor U8534 (N_8534,N_7059,N_7503);
and U8535 (N_8535,N_7147,N_7385);
nand U8536 (N_8536,N_7671,N_7721);
or U8537 (N_8537,N_7353,N_6972);
xor U8538 (N_8538,N_6179,N_7075);
xor U8539 (N_8539,N_7046,N_6688);
and U8540 (N_8540,N_7478,N_6019);
nand U8541 (N_8541,N_7079,N_6135);
nand U8542 (N_8542,N_6127,N_6698);
or U8543 (N_8543,N_6905,N_7198);
or U8544 (N_8544,N_6572,N_6801);
or U8545 (N_8545,N_7942,N_7428);
nand U8546 (N_8546,N_6192,N_7971);
nor U8547 (N_8547,N_6973,N_6643);
xnor U8548 (N_8548,N_6123,N_7481);
and U8549 (N_8549,N_6047,N_7700);
or U8550 (N_8550,N_7930,N_6321);
or U8551 (N_8551,N_7020,N_7401);
nand U8552 (N_8552,N_7951,N_6226);
and U8553 (N_8553,N_7536,N_6954);
xor U8554 (N_8554,N_6771,N_6831);
nor U8555 (N_8555,N_7036,N_7817);
nand U8556 (N_8556,N_6037,N_6015);
and U8557 (N_8557,N_7444,N_6379);
or U8558 (N_8558,N_7777,N_6463);
or U8559 (N_8559,N_6885,N_7337);
xnor U8560 (N_8560,N_7825,N_7692);
xor U8561 (N_8561,N_6197,N_7820);
and U8562 (N_8562,N_7455,N_6866);
xnor U8563 (N_8563,N_7324,N_7551);
nor U8564 (N_8564,N_6827,N_7661);
xor U8565 (N_8565,N_7539,N_7102);
or U8566 (N_8566,N_6190,N_6821);
or U8567 (N_8567,N_6433,N_6909);
xnor U8568 (N_8568,N_6331,N_6710);
nor U8569 (N_8569,N_6874,N_7776);
nor U8570 (N_8570,N_6860,N_6339);
or U8571 (N_8571,N_7497,N_6493);
and U8572 (N_8572,N_7397,N_7431);
xnor U8573 (N_8573,N_6887,N_7358);
xor U8574 (N_8574,N_6355,N_7675);
nand U8575 (N_8575,N_7964,N_7760);
xor U8576 (N_8576,N_6778,N_6131);
nand U8577 (N_8577,N_6302,N_6868);
nand U8578 (N_8578,N_6621,N_7380);
nand U8579 (N_8579,N_6533,N_7570);
or U8580 (N_8580,N_6439,N_6756);
nand U8581 (N_8581,N_6491,N_7289);
nor U8582 (N_8582,N_6146,N_7427);
or U8583 (N_8583,N_6986,N_6673);
xor U8584 (N_8584,N_7650,N_6323);
and U8585 (N_8585,N_6980,N_6893);
xnor U8586 (N_8586,N_6508,N_7273);
xnor U8587 (N_8587,N_6686,N_6900);
or U8588 (N_8588,N_7395,N_6623);
xor U8589 (N_8589,N_7654,N_7962);
nor U8590 (N_8590,N_7556,N_7336);
xor U8591 (N_8591,N_7345,N_6566);
nand U8592 (N_8592,N_7286,N_7970);
nand U8593 (N_8593,N_6225,N_6149);
or U8594 (N_8594,N_7176,N_7867);
nand U8595 (N_8595,N_6434,N_6929);
or U8596 (N_8596,N_7131,N_7755);
xnor U8597 (N_8597,N_7333,N_6852);
xor U8598 (N_8598,N_7858,N_7483);
and U8599 (N_8599,N_6279,N_7576);
nor U8600 (N_8600,N_6920,N_7037);
nor U8601 (N_8601,N_7985,N_7460);
nor U8602 (N_8602,N_7917,N_7976);
nand U8603 (N_8603,N_6600,N_6057);
nand U8604 (N_8604,N_7845,N_6240);
nor U8605 (N_8605,N_6377,N_6363);
and U8606 (N_8606,N_7881,N_7050);
or U8607 (N_8607,N_7774,N_7265);
and U8608 (N_8608,N_6347,N_6124);
and U8609 (N_8609,N_7437,N_6692);
or U8610 (N_8610,N_7726,N_6000);
or U8611 (N_8611,N_6361,N_6595);
or U8612 (N_8612,N_6881,N_6677);
nand U8613 (N_8613,N_6045,N_7382);
or U8614 (N_8614,N_6108,N_7791);
xnor U8615 (N_8615,N_7089,N_7117);
or U8616 (N_8616,N_7097,N_7686);
xor U8617 (N_8617,N_7751,N_7237);
nand U8618 (N_8618,N_6265,N_6233);
and U8619 (N_8619,N_6208,N_6222);
and U8620 (N_8620,N_7910,N_6209);
and U8621 (N_8621,N_7373,N_7045);
or U8622 (N_8622,N_6054,N_6012);
nor U8623 (N_8623,N_6249,N_6231);
nor U8624 (N_8624,N_7203,N_7182);
nand U8625 (N_8625,N_7159,N_7589);
xnor U8626 (N_8626,N_7617,N_6091);
xnor U8627 (N_8627,N_7533,N_7705);
and U8628 (N_8628,N_6656,N_7468);
nand U8629 (N_8629,N_7604,N_7120);
or U8630 (N_8630,N_7696,N_7593);
xnor U8631 (N_8631,N_6939,N_7261);
xnor U8632 (N_8632,N_6708,N_6557);
xor U8633 (N_8633,N_7772,N_7785);
nand U8634 (N_8634,N_7205,N_7142);
nor U8635 (N_8635,N_6804,N_6295);
xor U8636 (N_8636,N_7832,N_6912);
xor U8637 (N_8637,N_7949,N_6823);
nor U8638 (N_8638,N_7838,N_7782);
or U8639 (N_8639,N_6662,N_7847);
nor U8640 (N_8640,N_7190,N_7494);
xnor U8641 (N_8641,N_7040,N_6924);
nand U8642 (N_8642,N_6078,N_6883);
or U8643 (N_8643,N_7270,N_7950);
and U8644 (N_8644,N_6228,N_7346);
nor U8645 (N_8645,N_7835,N_6755);
and U8646 (N_8646,N_7920,N_7767);
nand U8647 (N_8647,N_6011,N_6529);
or U8648 (N_8648,N_7143,N_7579);
xor U8649 (N_8649,N_7135,N_7885);
or U8650 (N_8650,N_7844,N_6830);
xor U8651 (N_8651,N_7595,N_6061);
and U8652 (N_8652,N_7223,N_7218);
and U8653 (N_8653,N_7694,N_6967);
and U8654 (N_8654,N_7206,N_7989);
xor U8655 (N_8655,N_6576,N_7474);
or U8656 (N_8656,N_6693,N_6390);
nor U8657 (N_8657,N_6092,N_6788);
or U8658 (N_8658,N_6009,N_7954);
or U8659 (N_8659,N_6553,N_7184);
xnor U8660 (N_8660,N_7898,N_6674);
xnor U8661 (N_8661,N_7963,N_6591);
and U8662 (N_8662,N_7138,N_7107);
nand U8663 (N_8663,N_7934,N_6867);
nor U8664 (N_8664,N_6683,N_7947);
and U8665 (N_8665,N_7334,N_6210);
or U8666 (N_8666,N_6607,N_7564);
nor U8667 (N_8667,N_6242,N_6873);
or U8668 (N_8668,N_6652,N_6271);
xnor U8669 (N_8669,N_6090,N_6276);
xor U8670 (N_8670,N_6201,N_7199);
and U8671 (N_8671,N_7408,N_6387);
nor U8672 (N_8672,N_7943,N_7921);
nor U8673 (N_8673,N_6536,N_7550);
xnor U8674 (N_8674,N_6851,N_6620);
nor U8675 (N_8675,N_6024,N_7140);
xor U8676 (N_8676,N_6480,N_6911);
nand U8677 (N_8677,N_7409,N_7209);
and U8678 (N_8678,N_6613,N_7326);
or U8679 (N_8679,N_7665,N_6940);
or U8680 (N_8680,N_7192,N_6944);
xnor U8681 (N_8681,N_7739,N_6050);
xor U8682 (N_8682,N_7941,N_6748);
nor U8683 (N_8683,N_6590,N_7851);
xnor U8684 (N_8684,N_6188,N_6236);
and U8685 (N_8685,N_7859,N_7419);
and U8686 (N_8686,N_6538,N_7752);
or U8687 (N_8687,N_7557,N_7806);
nand U8688 (N_8688,N_7681,N_6564);
nand U8689 (N_8689,N_7285,N_6535);
nand U8690 (N_8690,N_6646,N_6072);
xor U8691 (N_8691,N_6400,N_6430);
nor U8692 (N_8692,N_6739,N_6602);
or U8693 (N_8693,N_6879,N_7997);
or U8694 (N_8694,N_7116,N_6690);
and U8695 (N_8695,N_6129,N_6734);
nor U8696 (N_8696,N_6723,N_6172);
nor U8697 (N_8697,N_7405,N_7644);
and U8698 (N_8698,N_6886,N_6415);
and U8699 (N_8699,N_6583,N_6418);
nand U8700 (N_8700,N_6077,N_7984);
xnor U8701 (N_8701,N_7064,N_7349);
or U8702 (N_8702,N_7766,N_6691);
nand U8703 (N_8703,N_6488,N_6036);
or U8704 (N_8704,N_7264,N_6112);
or U8705 (N_8705,N_6746,N_6984);
and U8706 (N_8706,N_7931,N_6326);
xor U8707 (N_8707,N_6198,N_6963);
xor U8708 (N_8708,N_7253,N_6230);
and U8709 (N_8709,N_7163,N_7277);
xnor U8710 (N_8710,N_7543,N_7945);
xnor U8711 (N_8711,N_6615,N_7577);
nor U8712 (N_8712,N_7498,N_7242);
or U8713 (N_8713,N_6064,N_7035);
nor U8714 (N_8714,N_6835,N_7837);
nand U8715 (N_8715,N_6709,N_6043);
and U8716 (N_8716,N_7610,N_6780);
nand U8717 (N_8717,N_6660,N_6751);
and U8718 (N_8718,N_6173,N_7347);
nand U8719 (N_8719,N_7321,N_7746);
xnor U8720 (N_8720,N_6671,N_7154);
or U8721 (N_8721,N_6451,N_6807);
or U8722 (N_8722,N_7197,N_7378);
nand U8723 (N_8723,N_6882,N_6727);
nand U8724 (N_8724,N_6435,N_6042);
nand U8725 (N_8725,N_7653,N_7758);
xor U8726 (N_8726,N_7441,N_6817);
xnor U8727 (N_8727,N_7928,N_6076);
or U8728 (N_8728,N_6810,N_7648);
xnor U8729 (N_8729,N_7612,N_6053);
nand U8730 (N_8730,N_7241,N_6311);
and U8731 (N_8731,N_6459,N_6389);
nand U8732 (N_8732,N_7262,N_6854);
nor U8733 (N_8733,N_6113,N_7787);
and U8734 (N_8734,N_6575,N_6969);
nor U8735 (N_8735,N_7180,N_6987);
nand U8736 (N_8736,N_7667,N_7940);
and U8737 (N_8737,N_6562,N_6999);
or U8738 (N_8738,N_7527,N_7109);
and U8739 (N_8739,N_6982,N_6461);
nand U8740 (N_8740,N_7114,N_7267);
and U8741 (N_8741,N_6263,N_6178);
and U8742 (N_8742,N_7637,N_7605);
nor U8743 (N_8743,N_6730,N_7784);
and U8744 (N_8744,N_7911,N_7342);
nor U8745 (N_8745,N_6422,N_7685);
nor U8746 (N_8746,N_6453,N_7609);
and U8747 (N_8747,N_7750,N_7293);
nor U8748 (N_8748,N_6397,N_6837);
and U8749 (N_8749,N_7780,N_7652);
nand U8750 (N_8750,N_7973,N_7643);
xnor U8751 (N_8751,N_7230,N_6742);
or U8752 (N_8752,N_6506,N_7016);
or U8753 (N_8753,N_6858,N_7540);
and U8754 (N_8754,N_6813,N_7070);
nor U8755 (N_8755,N_7824,N_6712);
xnor U8756 (N_8756,N_7063,N_7348);
xor U8757 (N_8757,N_7959,N_6505);
nand U8758 (N_8758,N_6532,N_7186);
nand U8759 (N_8759,N_7213,N_7101);
nor U8760 (N_8760,N_7255,N_6697);
nor U8761 (N_8761,N_7695,N_7245);
nor U8762 (N_8762,N_6080,N_7562);
or U8763 (N_8763,N_7645,N_7251);
or U8764 (N_8764,N_7383,N_7220);
xnor U8765 (N_8765,N_6637,N_7354);
xor U8766 (N_8766,N_6083,N_6384);
and U8767 (N_8767,N_6016,N_6217);
and U8768 (N_8768,N_6283,N_7454);
or U8769 (N_8769,N_6753,N_6292);
and U8770 (N_8770,N_6155,N_6761);
and U8771 (N_8771,N_7946,N_7814);
and U8772 (N_8772,N_6243,N_7871);
and U8773 (N_8773,N_6494,N_6933);
and U8774 (N_8774,N_7068,N_7663);
nand U8775 (N_8775,N_6020,N_6926);
and U8776 (N_8776,N_7158,N_6218);
xor U8777 (N_8777,N_7526,N_7529);
nand U8778 (N_8778,N_6975,N_7704);
or U8779 (N_8779,N_6638,N_6482);
or U8780 (N_8780,N_7465,N_7156);
xor U8781 (N_8781,N_7234,N_6200);
nand U8782 (N_8782,N_6622,N_7386);
and U8783 (N_8783,N_7052,N_7165);
or U8784 (N_8784,N_7629,N_6605);
or U8785 (N_8785,N_6812,N_7691);
and U8786 (N_8786,N_6608,N_6847);
or U8787 (N_8787,N_6864,N_7883);
nand U8788 (N_8788,N_7274,N_6333);
or U8789 (N_8789,N_6385,N_6165);
nand U8790 (N_8790,N_7322,N_7512);
and U8791 (N_8791,N_7919,N_6245);
or U8792 (N_8792,N_6441,N_7303);
or U8793 (N_8793,N_7043,N_7376);
and U8794 (N_8794,N_7227,N_6211);
xnor U8795 (N_8795,N_7991,N_7420);
nor U8796 (N_8796,N_6103,N_7296);
or U8797 (N_8797,N_6586,N_7808);
xor U8798 (N_8798,N_7697,N_7850);
and U8799 (N_8799,N_7729,N_6356);
nor U8800 (N_8800,N_7204,N_7795);
nand U8801 (N_8801,N_6516,N_6332);
or U8802 (N_8802,N_7601,N_7588);
or U8803 (N_8803,N_6189,N_7415);
or U8804 (N_8804,N_7033,N_6550);
nor U8805 (N_8805,N_7607,N_7429);
or U8806 (N_8806,N_6578,N_6089);
and U8807 (N_8807,N_7545,N_6396);
and U8808 (N_8808,N_6833,N_6932);
or U8809 (N_8809,N_6121,N_6290);
xnor U8810 (N_8810,N_7891,N_7343);
xor U8811 (N_8811,N_6618,N_6906);
or U8812 (N_8812,N_6186,N_6612);
and U8813 (N_8813,N_6288,N_6507);
nand U8814 (N_8814,N_7307,N_6194);
xnor U8815 (N_8815,N_7810,N_7424);
or U8816 (N_8816,N_7572,N_6469);
nand U8817 (N_8817,N_7287,N_6205);
and U8818 (N_8818,N_7848,N_6251);
nand U8819 (N_8819,N_6431,N_6364);
nor U8820 (N_8820,N_6757,N_7575);
nand U8821 (N_8821,N_6025,N_7757);
nor U8822 (N_8822,N_7436,N_7542);
xnor U8823 (N_8823,N_6031,N_7797);
xnor U8824 (N_8824,N_7300,N_7530);
xor U8825 (N_8825,N_7974,N_6162);
or U8826 (N_8826,N_7356,N_7779);
nand U8827 (N_8827,N_6032,N_6559);
or U8828 (N_8828,N_6593,N_6006);
xor U8829 (N_8829,N_7330,N_7008);
nand U8830 (N_8830,N_7232,N_6002);
xor U8831 (N_8831,N_6818,N_6570);
nor U8832 (N_8832,N_7923,N_6310);
and U8833 (N_8833,N_6694,N_7127);
xnor U8834 (N_8834,N_6268,N_6768);
xnor U8835 (N_8835,N_7108,N_7977);
or U8836 (N_8836,N_6096,N_6345);
and U8837 (N_8837,N_6551,N_6947);
or U8838 (N_8838,N_6468,N_7212);
and U8839 (N_8839,N_6636,N_7677);
or U8840 (N_8840,N_6158,N_6063);
or U8841 (N_8841,N_6065,N_6160);
xor U8842 (N_8842,N_7435,N_7462);
xnor U8843 (N_8843,N_6452,N_7173);
or U8844 (N_8844,N_7517,N_6474);
or U8845 (N_8845,N_6370,N_6997);
or U8846 (N_8846,N_7583,N_7235);
nand U8847 (N_8847,N_6317,N_6898);
nand U8848 (N_8848,N_7842,N_7707);
nand U8849 (N_8849,N_6213,N_6125);
nor U8850 (N_8850,N_7909,N_7769);
and U8851 (N_8851,N_7641,N_6644);
nor U8852 (N_8852,N_6706,N_6039);
nor U8853 (N_8853,N_7899,N_6074);
nor U8854 (N_8854,N_6950,N_7077);
nor U8855 (N_8855,N_6119,N_6832);
or U8856 (N_8856,N_6558,N_6824);
or U8857 (N_8857,N_7268,N_6193);
and U8858 (N_8858,N_6107,N_7969);
nor U8859 (N_8859,N_7325,N_7927);
nor U8860 (N_8860,N_6357,N_7328);
and U8861 (N_8861,N_6444,N_6309);
and U8862 (N_8862,N_7829,N_7363);
nand U8863 (N_8863,N_6035,N_7738);
and U8864 (N_8864,N_6596,N_6374);
and U8865 (N_8865,N_6202,N_7912);
nand U8866 (N_8866,N_6556,N_6308);
nand U8867 (N_8867,N_6130,N_6930);
nor U8868 (N_8868,N_7684,N_7473);
or U8869 (N_8869,N_7761,N_7597);
xor U8870 (N_8870,N_6794,N_6981);
and U8871 (N_8871,N_7137,N_6298);
nand U8872 (N_8872,N_7085,N_6320);
and U8873 (N_8873,N_6284,N_6684);
nand U8874 (N_8874,N_6754,N_7271);
nor U8875 (N_8875,N_7450,N_7877);
nand U8876 (N_8876,N_6398,N_7201);
nor U8877 (N_8877,N_6084,N_6907);
nand U8878 (N_8878,N_6052,N_7807);
nor U8879 (N_8879,N_7680,N_7452);
and U8880 (N_8880,N_7961,N_7716);
xnor U8881 (N_8881,N_7306,N_7901);
nor U8882 (N_8882,N_7789,N_7327);
xor U8883 (N_8883,N_7554,N_7193);
nor U8884 (N_8884,N_7732,N_7302);
nand U8885 (N_8885,N_6889,N_6219);
nor U8886 (N_8886,N_7207,N_7870);
nor U8887 (N_8887,N_7781,N_7488);
and U8888 (N_8888,N_7371,N_7056);
or U8889 (N_8889,N_6676,N_7263);
nor U8890 (N_8890,N_6869,N_6030);
or U8891 (N_8891,N_6394,N_6960);
nor U8892 (N_8892,N_7598,N_6725);
or U8893 (N_8893,N_6653,N_7047);
nor U8894 (N_8894,N_7189,N_7798);
nand U8895 (N_8895,N_6641,N_6741);
nor U8896 (N_8896,N_7413,N_7487);
and U8897 (N_8897,N_6270,N_6406);
xnor U8898 (N_8898,N_7015,N_7759);
or U8899 (N_8899,N_7098,N_6850);
nor U8900 (N_8900,N_7374,N_7221);
and U8901 (N_8901,N_7559,N_6733);
nor U8902 (N_8902,N_6436,N_7226);
nor U8903 (N_8903,N_6136,N_6527);
nor U8904 (N_8904,N_7672,N_7725);
nand U8905 (N_8905,N_7430,N_7051);
xnor U8906 (N_8906,N_6916,N_6026);
nand U8907 (N_8907,N_6519,N_6526);
and U8908 (N_8908,N_7515,N_6073);
xor U8909 (N_8909,N_6382,N_6616);
or U8910 (N_8910,N_6278,N_7011);
xnor U8911 (N_8911,N_7591,N_6191);
nand U8912 (N_8912,N_7316,N_6264);
and U8913 (N_8913,N_6820,N_6498);
nor U8914 (N_8914,N_7396,N_7078);
or U8915 (N_8915,N_7018,N_6749);
nand U8916 (N_8916,N_6183,N_7724);
xnor U8917 (N_8917,N_6534,N_6805);
or U8918 (N_8918,N_7174,N_7939);
xor U8919 (N_8919,N_7878,N_6511);
and U8920 (N_8920,N_6340,N_6142);
xnor U8921 (N_8921,N_7179,N_6793);
nor U8922 (N_8922,N_7187,N_6627);
and U8923 (N_8923,N_7195,N_6040);
nor U8924 (N_8924,N_7001,N_6196);
nor U8925 (N_8925,N_7275,N_7507);
nand U8926 (N_8926,N_7128,N_6174);
or U8927 (N_8927,N_6515,N_7710);
nand U8928 (N_8928,N_6258,N_7284);
xor U8929 (N_8929,N_7965,N_7673);
nor U8930 (N_8930,N_6917,N_7183);
and U8931 (N_8931,N_7153,N_7399);
nand U8932 (N_8932,N_7828,N_6682);
and U8933 (N_8933,N_6344,N_6945);
nor U8934 (N_8934,N_7888,N_6460);
or U8935 (N_8935,N_6458,N_6066);
xor U8936 (N_8936,N_7717,N_7480);
or U8937 (N_8937,N_6826,N_6153);
xnor U8938 (N_8938,N_7882,N_7391);
xor U8939 (N_8939,N_7875,N_6617);
nand U8940 (N_8940,N_6567,N_7831);
nor U8941 (N_8941,N_6517,N_6919);
nor U8942 (N_8942,N_7628,N_6348);
and U8943 (N_8943,N_7619,N_6779);
and U8944 (N_8944,N_7799,N_6654);
xor U8945 (N_8945,N_6884,N_6811);
and U8946 (N_8946,N_7211,N_7603);
and U8947 (N_8947,N_7028,N_7447);
xnor U8948 (N_8948,N_6402,N_6537);
nor U8949 (N_8949,N_7276,N_6970);
nor U8950 (N_8950,N_6773,N_7794);
and U8951 (N_8951,N_6844,N_6280);
nand U8952 (N_8952,N_7486,N_7231);
xnor U8953 (N_8953,N_6147,N_6758);
nand U8954 (N_8954,N_7897,N_7049);
and U8955 (N_8955,N_7332,N_7141);
nor U8956 (N_8956,N_7466,N_6547);
and U8957 (N_8957,N_6421,N_7096);
or U8958 (N_8958,N_7357,N_7208);
nand U8959 (N_8959,N_7547,N_7733);
or U8960 (N_8960,N_6839,N_6870);
xor U8961 (N_8961,N_6267,N_6716);
xor U8962 (N_8962,N_6528,N_6678);
xor U8963 (N_8963,N_7839,N_7039);
and U8964 (N_8964,N_6597,N_6631);
xnor U8965 (N_8965,N_7639,N_7103);
nor U8966 (N_8966,N_7768,N_7528);
and U8967 (N_8967,N_7318,N_6752);
or U8968 (N_8968,N_7993,N_6840);
nor U8969 (N_8969,N_6736,N_6942);
nor U8970 (N_8970,N_6069,N_7632);
and U8971 (N_8971,N_7599,N_7092);
xnor U8972 (N_8972,N_7344,N_7843);
nor U8973 (N_8973,N_7024,N_6935);
nand U8974 (N_8974,N_6013,N_6855);
xnor U8975 (N_8975,N_7006,N_7608);
nand U8976 (N_8976,N_6871,N_6699);
nand U8977 (N_8977,N_6899,N_6624);
nor U8978 (N_8978,N_6922,N_7903);
or U8979 (N_8979,N_6346,N_7196);
nand U8980 (N_8980,N_7876,N_6598);
and U8981 (N_8981,N_6670,N_6104);
nand U8982 (N_8982,N_6445,N_6028);
nor U8983 (N_8983,N_6504,N_6021);
nor U8984 (N_8984,N_6530,N_7157);
and U8985 (N_8985,N_6098,N_6049);
nor U8986 (N_8986,N_7500,N_6350);
nor U8987 (N_8987,N_6324,N_6798);
nor U8988 (N_8988,N_7021,N_6843);
or U8989 (N_8989,N_7822,N_6059);
nand U8990 (N_8990,N_7459,N_7247);
and U8991 (N_8991,N_6913,N_7999);
and U8992 (N_8992,N_7152,N_6633);
nand U8993 (N_8993,N_7169,N_6161);
or U8994 (N_8994,N_7471,N_6784);
nand U8995 (N_8995,N_6176,N_6949);
or U8996 (N_8996,N_6447,N_6262);
nor U8997 (N_8997,N_6795,N_6097);
or U8998 (N_8998,N_7690,N_7484);
nand U8999 (N_8999,N_7125,N_7155);
xor U9000 (N_9000,N_7259,N_6950);
xor U9001 (N_9001,N_6214,N_7694);
xnor U9002 (N_9002,N_7324,N_7616);
or U9003 (N_9003,N_7906,N_7712);
nand U9004 (N_9004,N_7765,N_6671);
xor U9005 (N_9005,N_6994,N_7862);
or U9006 (N_9006,N_7544,N_7765);
and U9007 (N_9007,N_6798,N_6420);
xor U9008 (N_9008,N_7827,N_7511);
or U9009 (N_9009,N_7971,N_7581);
or U9010 (N_9010,N_6933,N_6939);
nand U9011 (N_9011,N_7888,N_6606);
or U9012 (N_9012,N_6764,N_7645);
or U9013 (N_9013,N_6869,N_6293);
nand U9014 (N_9014,N_7901,N_6238);
or U9015 (N_9015,N_7970,N_6244);
or U9016 (N_9016,N_7704,N_6034);
and U9017 (N_9017,N_7941,N_7292);
nor U9018 (N_9018,N_7871,N_6254);
and U9019 (N_9019,N_7000,N_7811);
xnor U9020 (N_9020,N_7682,N_6608);
or U9021 (N_9021,N_7361,N_7005);
nor U9022 (N_9022,N_7271,N_6463);
nor U9023 (N_9023,N_7281,N_6142);
nand U9024 (N_9024,N_7837,N_6669);
xor U9025 (N_9025,N_7228,N_6460);
nand U9026 (N_9026,N_6639,N_7988);
and U9027 (N_9027,N_6378,N_6257);
or U9028 (N_9028,N_7065,N_7647);
or U9029 (N_9029,N_6375,N_6204);
nand U9030 (N_9030,N_6242,N_6813);
nor U9031 (N_9031,N_6989,N_6721);
and U9032 (N_9032,N_7291,N_7975);
xor U9033 (N_9033,N_7582,N_6621);
nand U9034 (N_9034,N_6579,N_6753);
or U9035 (N_9035,N_7154,N_7278);
xnor U9036 (N_9036,N_6169,N_6681);
nor U9037 (N_9037,N_6198,N_7122);
nor U9038 (N_9038,N_7510,N_7761);
and U9039 (N_9039,N_6022,N_6398);
xor U9040 (N_9040,N_6757,N_6701);
nand U9041 (N_9041,N_7500,N_7934);
nor U9042 (N_9042,N_6705,N_7703);
and U9043 (N_9043,N_7648,N_6826);
nor U9044 (N_9044,N_6754,N_7372);
xor U9045 (N_9045,N_7471,N_7934);
and U9046 (N_9046,N_7913,N_7829);
nand U9047 (N_9047,N_6713,N_6123);
nand U9048 (N_9048,N_7812,N_6992);
nor U9049 (N_9049,N_7661,N_7084);
or U9050 (N_9050,N_7609,N_7380);
xnor U9051 (N_9051,N_6704,N_7574);
xor U9052 (N_9052,N_6485,N_6145);
or U9053 (N_9053,N_7373,N_6713);
and U9054 (N_9054,N_7231,N_7736);
and U9055 (N_9055,N_6439,N_7910);
nand U9056 (N_9056,N_7478,N_7311);
or U9057 (N_9057,N_6465,N_6837);
xor U9058 (N_9058,N_7745,N_7300);
nor U9059 (N_9059,N_7824,N_6126);
and U9060 (N_9060,N_6245,N_7569);
and U9061 (N_9061,N_7557,N_6561);
and U9062 (N_9062,N_7837,N_7344);
and U9063 (N_9063,N_7893,N_7199);
nand U9064 (N_9064,N_7943,N_6825);
and U9065 (N_9065,N_7423,N_7275);
nor U9066 (N_9066,N_7529,N_6298);
or U9067 (N_9067,N_7476,N_6195);
nor U9068 (N_9068,N_6518,N_6927);
nor U9069 (N_9069,N_7218,N_7177);
xor U9070 (N_9070,N_6203,N_7934);
or U9071 (N_9071,N_6705,N_6609);
or U9072 (N_9072,N_7040,N_6372);
or U9073 (N_9073,N_7570,N_7812);
and U9074 (N_9074,N_6145,N_6612);
or U9075 (N_9075,N_6244,N_7927);
nor U9076 (N_9076,N_6225,N_6680);
xor U9077 (N_9077,N_7745,N_7081);
or U9078 (N_9078,N_6708,N_7249);
or U9079 (N_9079,N_6803,N_7839);
xnor U9080 (N_9080,N_6905,N_6156);
or U9081 (N_9081,N_6518,N_7569);
and U9082 (N_9082,N_6774,N_6434);
nand U9083 (N_9083,N_7866,N_6616);
or U9084 (N_9084,N_6315,N_7605);
or U9085 (N_9085,N_7749,N_7790);
and U9086 (N_9086,N_7714,N_6263);
nor U9087 (N_9087,N_7469,N_6354);
xnor U9088 (N_9088,N_6939,N_6965);
nor U9089 (N_9089,N_7699,N_7005);
or U9090 (N_9090,N_7807,N_6166);
and U9091 (N_9091,N_7811,N_6930);
and U9092 (N_9092,N_7947,N_6949);
and U9093 (N_9093,N_7326,N_7062);
and U9094 (N_9094,N_7663,N_6361);
and U9095 (N_9095,N_7509,N_6094);
xor U9096 (N_9096,N_7452,N_7503);
xor U9097 (N_9097,N_7221,N_7098);
nand U9098 (N_9098,N_7899,N_6968);
and U9099 (N_9099,N_7338,N_7655);
and U9100 (N_9100,N_6069,N_6358);
nor U9101 (N_9101,N_7835,N_6398);
and U9102 (N_9102,N_6655,N_6009);
and U9103 (N_9103,N_7837,N_6902);
or U9104 (N_9104,N_7067,N_7706);
nor U9105 (N_9105,N_6734,N_7038);
xor U9106 (N_9106,N_6687,N_6086);
xnor U9107 (N_9107,N_6667,N_6861);
or U9108 (N_9108,N_6792,N_7501);
and U9109 (N_9109,N_6208,N_6847);
nor U9110 (N_9110,N_7409,N_7348);
or U9111 (N_9111,N_6983,N_6477);
or U9112 (N_9112,N_6344,N_7809);
nor U9113 (N_9113,N_7549,N_7639);
xnor U9114 (N_9114,N_7656,N_6317);
xnor U9115 (N_9115,N_7323,N_7955);
xor U9116 (N_9116,N_6294,N_6906);
nor U9117 (N_9117,N_6477,N_7447);
and U9118 (N_9118,N_6076,N_6280);
xnor U9119 (N_9119,N_6238,N_7434);
nand U9120 (N_9120,N_6990,N_6060);
nand U9121 (N_9121,N_7769,N_6780);
and U9122 (N_9122,N_7324,N_7411);
nor U9123 (N_9123,N_7955,N_6696);
xnor U9124 (N_9124,N_6073,N_6006);
xnor U9125 (N_9125,N_6386,N_6888);
nor U9126 (N_9126,N_6681,N_6304);
and U9127 (N_9127,N_6431,N_7821);
and U9128 (N_9128,N_7378,N_7977);
xor U9129 (N_9129,N_6030,N_6603);
or U9130 (N_9130,N_6822,N_6494);
and U9131 (N_9131,N_7906,N_6832);
nand U9132 (N_9132,N_7191,N_7490);
or U9133 (N_9133,N_6955,N_7298);
nor U9134 (N_9134,N_7483,N_6105);
and U9135 (N_9135,N_6369,N_6669);
and U9136 (N_9136,N_6890,N_6922);
and U9137 (N_9137,N_6102,N_6020);
nand U9138 (N_9138,N_6417,N_6585);
or U9139 (N_9139,N_7007,N_7355);
nand U9140 (N_9140,N_6626,N_6146);
nand U9141 (N_9141,N_7042,N_7350);
nand U9142 (N_9142,N_6531,N_6411);
nand U9143 (N_9143,N_6912,N_6932);
or U9144 (N_9144,N_6866,N_6570);
and U9145 (N_9145,N_6697,N_6935);
xor U9146 (N_9146,N_6774,N_7603);
xor U9147 (N_9147,N_7262,N_6702);
xnor U9148 (N_9148,N_7482,N_6330);
nand U9149 (N_9149,N_7394,N_7490);
and U9150 (N_9150,N_6815,N_6648);
xor U9151 (N_9151,N_7848,N_7797);
nand U9152 (N_9152,N_7674,N_6160);
xor U9153 (N_9153,N_7799,N_6643);
nor U9154 (N_9154,N_7558,N_6087);
nand U9155 (N_9155,N_7855,N_6171);
nor U9156 (N_9156,N_6129,N_6882);
nand U9157 (N_9157,N_7760,N_7218);
or U9158 (N_9158,N_6896,N_6878);
xnor U9159 (N_9159,N_7075,N_6842);
xnor U9160 (N_9160,N_6096,N_7863);
nor U9161 (N_9161,N_7988,N_7964);
nor U9162 (N_9162,N_6804,N_6303);
xor U9163 (N_9163,N_6357,N_7192);
nand U9164 (N_9164,N_7033,N_6686);
or U9165 (N_9165,N_7879,N_7245);
nand U9166 (N_9166,N_7424,N_6499);
and U9167 (N_9167,N_7657,N_6337);
and U9168 (N_9168,N_7366,N_7192);
or U9169 (N_9169,N_6448,N_6342);
nor U9170 (N_9170,N_7379,N_7160);
nand U9171 (N_9171,N_7784,N_7430);
and U9172 (N_9172,N_7600,N_6360);
xnor U9173 (N_9173,N_6113,N_6318);
and U9174 (N_9174,N_6546,N_7628);
or U9175 (N_9175,N_6928,N_7719);
xor U9176 (N_9176,N_6234,N_6027);
or U9177 (N_9177,N_7210,N_7949);
nand U9178 (N_9178,N_6052,N_7966);
nor U9179 (N_9179,N_6170,N_7754);
or U9180 (N_9180,N_7171,N_7712);
or U9181 (N_9181,N_7453,N_6030);
nor U9182 (N_9182,N_7178,N_7119);
nor U9183 (N_9183,N_6155,N_7541);
nor U9184 (N_9184,N_6529,N_6632);
xnor U9185 (N_9185,N_7390,N_6487);
xor U9186 (N_9186,N_6350,N_7310);
xor U9187 (N_9187,N_6925,N_7014);
nand U9188 (N_9188,N_7120,N_6814);
xor U9189 (N_9189,N_7584,N_6362);
nand U9190 (N_9190,N_6763,N_7998);
nor U9191 (N_9191,N_6583,N_6138);
nor U9192 (N_9192,N_7600,N_6885);
xor U9193 (N_9193,N_6478,N_6063);
xnor U9194 (N_9194,N_7292,N_6265);
nand U9195 (N_9195,N_7570,N_7197);
and U9196 (N_9196,N_6157,N_6654);
and U9197 (N_9197,N_6836,N_6150);
xnor U9198 (N_9198,N_6824,N_6292);
nor U9199 (N_9199,N_7578,N_7639);
or U9200 (N_9200,N_7048,N_6367);
and U9201 (N_9201,N_7642,N_7819);
and U9202 (N_9202,N_6910,N_7780);
nand U9203 (N_9203,N_7949,N_6101);
nand U9204 (N_9204,N_6437,N_7021);
xnor U9205 (N_9205,N_6160,N_6823);
nor U9206 (N_9206,N_6327,N_7335);
nor U9207 (N_9207,N_7750,N_7566);
or U9208 (N_9208,N_7340,N_6626);
or U9209 (N_9209,N_7672,N_7611);
nor U9210 (N_9210,N_7104,N_7247);
nor U9211 (N_9211,N_6960,N_7159);
or U9212 (N_9212,N_7860,N_7388);
nand U9213 (N_9213,N_7806,N_7596);
or U9214 (N_9214,N_7281,N_7944);
or U9215 (N_9215,N_6277,N_6621);
xnor U9216 (N_9216,N_6716,N_6631);
nor U9217 (N_9217,N_7167,N_6348);
or U9218 (N_9218,N_7838,N_6566);
nor U9219 (N_9219,N_6716,N_6574);
and U9220 (N_9220,N_7693,N_7864);
nand U9221 (N_9221,N_6465,N_6739);
nand U9222 (N_9222,N_6506,N_6364);
nor U9223 (N_9223,N_6009,N_7158);
nand U9224 (N_9224,N_6841,N_7458);
nor U9225 (N_9225,N_6457,N_6009);
xnor U9226 (N_9226,N_6430,N_7140);
nor U9227 (N_9227,N_7165,N_7962);
or U9228 (N_9228,N_7665,N_7988);
and U9229 (N_9229,N_7173,N_7190);
and U9230 (N_9230,N_6941,N_7071);
nand U9231 (N_9231,N_7821,N_7003);
xnor U9232 (N_9232,N_6606,N_6593);
xor U9233 (N_9233,N_7141,N_7854);
and U9234 (N_9234,N_6471,N_7958);
xnor U9235 (N_9235,N_6232,N_6600);
xnor U9236 (N_9236,N_7688,N_7058);
nor U9237 (N_9237,N_6378,N_7115);
nor U9238 (N_9238,N_6489,N_6977);
and U9239 (N_9239,N_6425,N_6206);
nand U9240 (N_9240,N_7654,N_6372);
or U9241 (N_9241,N_6001,N_6391);
xnor U9242 (N_9242,N_6918,N_7000);
nand U9243 (N_9243,N_6555,N_6049);
nand U9244 (N_9244,N_7678,N_7817);
nor U9245 (N_9245,N_6444,N_6715);
nor U9246 (N_9246,N_7566,N_7124);
or U9247 (N_9247,N_7013,N_6741);
xor U9248 (N_9248,N_6098,N_6308);
nor U9249 (N_9249,N_6011,N_6493);
and U9250 (N_9250,N_6916,N_7840);
nor U9251 (N_9251,N_6798,N_6962);
and U9252 (N_9252,N_7874,N_6653);
nor U9253 (N_9253,N_7235,N_7883);
and U9254 (N_9254,N_7924,N_7531);
xor U9255 (N_9255,N_7878,N_7096);
nor U9256 (N_9256,N_7814,N_7248);
or U9257 (N_9257,N_7582,N_7485);
and U9258 (N_9258,N_7631,N_6599);
and U9259 (N_9259,N_6928,N_6700);
nor U9260 (N_9260,N_6717,N_6368);
and U9261 (N_9261,N_6794,N_6942);
or U9262 (N_9262,N_7553,N_6331);
or U9263 (N_9263,N_6862,N_7765);
xor U9264 (N_9264,N_7074,N_7343);
nand U9265 (N_9265,N_6341,N_6778);
nor U9266 (N_9266,N_7165,N_6575);
nand U9267 (N_9267,N_7694,N_6389);
nor U9268 (N_9268,N_7530,N_7077);
and U9269 (N_9269,N_6651,N_6812);
nor U9270 (N_9270,N_7366,N_6227);
or U9271 (N_9271,N_6792,N_7563);
nor U9272 (N_9272,N_7382,N_7772);
xor U9273 (N_9273,N_6168,N_7623);
nor U9274 (N_9274,N_7215,N_6796);
and U9275 (N_9275,N_7352,N_7582);
or U9276 (N_9276,N_6054,N_6297);
or U9277 (N_9277,N_6071,N_7358);
nor U9278 (N_9278,N_7017,N_6730);
xnor U9279 (N_9279,N_6561,N_7336);
or U9280 (N_9280,N_7943,N_6687);
and U9281 (N_9281,N_6319,N_7076);
or U9282 (N_9282,N_7965,N_6086);
and U9283 (N_9283,N_6382,N_6887);
nand U9284 (N_9284,N_7264,N_7484);
or U9285 (N_9285,N_6376,N_6193);
or U9286 (N_9286,N_7689,N_7882);
xnor U9287 (N_9287,N_7176,N_6048);
and U9288 (N_9288,N_7583,N_7523);
xor U9289 (N_9289,N_7877,N_6534);
and U9290 (N_9290,N_6208,N_7503);
or U9291 (N_9291,N_6707,N_7790);
xor U9292 (N_9292,N_6992,N_6299);
or U9293 (N_9293,N_7924,N_7778);
or U9294 (N_9294,N_7012,N_6128);
nand U9295 (N_9295,N_6822,N_7306);
xnor U9296 (N_9296,N_7708,N_7702);
nand U9297 (N_9297,N_7651,N_7617);
nor U9298 (N_9298,N_6646,N_7899);
nor U9299 (N_9299,N_6892,N_6801);
and U9300 (N_9300,N_6020,N_6973);
or U9301 (N_9301,N_7731,N_6609);
and U9302 (N_9302,N_7867,N_6163);
or U9303 (N_9303,N_7702,N_6004);
xnor U9304 (N_9304,N_6076,N_7572);
and U9305 (N_9305,N_7269,N_7578);
nand U9306 (N_9306,N_7157,N_6658);
xnor U9307 (N_9307,N_6165,N_7885);
nor U9308 (N_9308,N_6874,N_6341);
nand U9309 (N_9309,N_7530,N_7359);
or U9310 (N_9310,N_7833,N_6111);
xnor U9311 (N_9311,N_7847,N_7320);
nor U9312 (N_9312,N_7896,N_6766);
nor U9313 (N_9313,N_7349,N_6197);
or U9314 (N_9314,N_7131,N_6275);
nor U9315 (N_9315,N_7992,N_7212);
nand U9316 (N_9316,N_7059,N_7390);
and U9317 (N_9317,N_6778,N_6477);
xor U9318 (N_9318,N_7136,N_7545);
nor U9319 (N_9319,N_7650,N_7534);
and U9320 (N_9320,N_7552,N_6370);
xor U9321 (N_9321,N_6824,N_7819);
nand U9322 (N_9322,N_6218,N_7285);
nor U9323 (N_9323,N_7946,N_7886);
nand U9324 (N_9324,N_7569,N_6411);
and U9325 (N_9325,N_7161,N_7432);
or U9326 (N_9326,N_7688,N_6378);
xor U9327 (N_9327,N_6901,N_6095);
and U9328 (N_9328,N_6261,N_7435);
xnor U9329 (N_9329,N_7309,N_6174);
and U9330 (N_9330,N_7545,N_7179);
or U9331 (N_9331,N_6168,N_6627);
and U9332 (N_9332,N_7630,N_7685);
and U9333 (N_9333,N_7504,N_6902);
nand U9334 (N_9334,N_7126,N_7770);
or U9335 (N_9335,N_6622,N_7868);
nor U9336 (N_9336,N_6675,N_6188);
or U9337 (N_9337,N_7305,N_6978);
nor U9338 (N_9338,N_7799,N_6212);
and U9339 (N_9339,N_6196,N_6559);
or U9340 (N_9340,N_6147,N_7665);
and U9341 (N_9341,N_7378,N_6286);
nor U9342 (N_9342,N_7590,N_7051);
nor U9343 (N_9343,N_6616,N_6069);
nor U9344 (N_9344,N_7322,N_6838);
nand U9345 (N_9345,N_6381,N_6134);
and U9346 (N_9346,N_7038,N_7742);
xnor U9347 (N_9347,N_6500,N_6292);
or U9348 (N_9348,N_6487,N_6639);
nor U9349 (N_9349,N_6623,N_7203);
nand U9350 (N_9350,N_6500,N_7030);
nor U9351 (N_9351,N_7943,N_7556);
xnor U9352 (N_9352,N_7580,N_7210);
or U9353 (N_9353,N_6820,N_6349);
nor U9354 (N_9354,N_7347,N_7909);
and U9355 (N_9355,N_6652,N_6443);
xor U9356 (N_9356,N_6419,N_7624);
xnor U9357 (N_9357,N_7273,N_6836);
xor U9358 (N_9358,N_7144,N_6884);
nor U9359 (N_9359,N_6877,N_6215);
and U9360 (N_9360,N_6590,N_6673);
and U9361 (N_9361,N_6290,N_7877);
xnor U9362 (N_9362,N_6086,N_7956);
and U9363 (N_9363,N_6584,N_7190);
nand U9364 (N_9364,N_7350,N_7490);
and U9365 (N_9365,N_7442,N_7659);
and U9366 (N_9366,N_7566,N_7453);
nor U9367 (N_9367,N_7593,N_7829);
nor U9368 (N_9368,N_7079,N_6466);
xor U9369 (N_9369,N_6562,N_6915);
xnor U9370 (N_9370,N_7095,N_7406);
or U9371 (N_9371,N_7469,N_7142);
or U9372 (N_9372,N_7575,N_6560);
or U9373 (N_9373,N_6512,N_7477);
or U9374 (N_9374,N_6650,N_6117);
and U9375 (N_9375,N_7556,N_7326);
and U9376 (N_9376,N_7486,N_7717);
nand U9377 (N_9377,N_6995,N_7471);
nor U9378 (N_9378,N_7812,N_6020);
nand U9379 (N_9379,N_6582,N_6004);
xor U9380 (N_9380,N_6616,N_7739);
xnor U9381 (N_9381,N_6138,N_6710);
xnor U9382 (N_9382,N_7899,N_6598);
and U9383 (N_9383,N_7123,N_6334);
or U9384 (N_9384,N_6305,N_6932);
xor U9385 (N_9385,N_7730,N_7578);
nand U9386 (N_9386,N_7718,N_6389);
xor U9387 (N_9387,N_7230,N_7163);
or U9388 (N_9388,N_7189,N_6622);
and U9389 (N_9389,N_6044,N_6515);
xor U9390 (N_9390,N_7293,N_6648);
xnor U9391 (N_9391,N_6491,N_7197);
and U9392 (N_9392,N_7311,N_7179);
and U9393 (N_9393,N_7782,N_6368);
nand U9394 (N_9394,N_6172,N_6214);
xnor U9395 (N_9395,N_7339,N_7496);
xnor U9396 (N_9396,N_6603,N_7264);
nor U9397 (N_9397,N_7806,N_6083);
or U9398 (N_9398,N_7275,N_6636);
or U9399 (N_9399,N_6714,N_7866);
nor U9400 (N_9400,N_6794,N_6870);
and U9401 (N_9401,N_7685,N_7397);
xnor U9402 (N_9402,N_6935,N_6791);
and U9403 (N_9403,N_6587,N_6026);
or U9404 (N_9404,N_7073,N_7411);
nor U9405 (N_9405,N_6911,N_6625);
or U9406 (N_9406,N_6351,N_7776);
or U9407 (N_9407,N_6723,N_6210);
xor U9408 (N_9408,N_6160,N_7907);
xnor U9409 (N_9409,N_6640,N_6629);
xnor U9410 (N_9410,N_7340,N_7215);
or U9411 (N_9411,N_7340,N_6172);
nand U9412 (N_9412,N_7978,N_7508);
nor U9413 (N_9413,N_7895,N_7210);
or U9414 (N_9414,N_6016,N_7983);
nand U9415 (N_9415,N_6792,N_7105);
xor U9416 (N_9416,N_7094,N_6938);
nand U9417 (N_9417,N_7108,N_7033);
nor U9418 (N_9418,N_7502,N_7915);
xnor U9419 (N_9419,N_6968,N_7957);
or U9420 (N_9420,N_7849,N_6365);
xnor U9421 (N_9421,N_7572,N_7258);
nor U9422 (N_9422,N_7325,N_7233);
nor U9423 (N_9423,N_7580,N_7857);
or U9424 (N_9424,N_7590,N_7380);
nand U9425 (N_9425,N_6298,N_7121);
and U9426 (N_9426,N_6859,N_6665);
xnor U9427 (N_9427,N_7481,N_6219);
nand U9428 (N_9428,N_6299,N_6502);
or U9429 (N_9429,N_7174,N_7283);
nand U9430 (N_9430,N_7360,N_7574);
or U9431 (N_9431,N_7706,N_7252);
or U9432 (N_9432,N_6931,N_7425);
nor U9433 (N_9433,N_7894,N_7608);
nor U9434 (N_9434,N_6029,N_6709);
nand U9435 (N_9435,N_7537,N_6526);
nand U9436 (N_9436,N_7596,N_6454);
nand U9437 (N_9437,N_7302,N_6069);
xnor U9438 (N_9438,N_7934,N_6931);
or U9439 (N_9439,N_6958,N_7995);
nor U9440 (N_9440,N_6933,N_7299);
nand U9441 (N_9441,N_7708,N_7369);
nor U9442 (N_9442,N_7752,N_7659);
xor U9443 (N_9443,N_7995,N_6611);
nand U9444 (N_9444,N_6056,N_6522);
xnor U9445 (N_9445,N_7824,N_6893);
nor U9446 (N_9446,N_6572,N_6540);
nor U9447 (N_9447,N_6829,N_7137);
xnor U9448 (N_9448,N_6654,N_6705);
or U9449 (N_9449,N_7141,N_6108);
nand U9450 (N_9450,N_6138,N_7300);
nor U9451 (N_9451,N_6646,N_7839);
nand U9452 (N_9452,N_6261,N_7395);
nand U9453 (N_9453,N_6251,N_7878);
nor U9454 (N_9454,N_7054,N_6148);
nand U9455 (N_9455,N_6398,N_6460);
and U9456 (N_9456,N_6665,N_7237);
nor U9457 (N_9457,N_7697,N_6641);
xor U9458 (N_9458,N_6675,N_7122);
xnor U9459 (N_9459,N_7538,N_7707);
xnor U9460 (N_9460,N_7536,N_6515);
nand U9461 (N_9461,N_7004,N_7877);
xor U9462 (N_9462,N_7026,N_6019);
xor U9463 (N_9463,N_7074,N_7193);
or U9464 (N_9464,N_6220,N_7111);
xor U9465 (N_9465,N_7585,N_6529);
nor U9466 (N_9466,N_7434,N_6316);
and U9467 (N_9467,N_7749,N_7349);
xnor U9468 (N_9468,N_7994,N_7827);
nand U9469 (N_9469,N_6765,N_7329);
xor U9470 (N_9470,N_6360,N_6096);
xor U9471 (N_9471,N_6650,N_6203);
or U9472 (N_9472,N_7229,N_6955);
nand U9473 (N_9473,N_6397,N_6166);
and U9474 (N_9474,N_6987,N_7975);
nand U9475 (N_9475,N_6643,N_6275);
xor U9476 (N_9476,N_7757,N_7218);
and U9477 (N_9477,N_6381,N_7473);
or U9478 (N_9478,N_7886,N_7018);
nor U9479 (N_9479,N_6890,N_7575);
xnor U9480 (N_9480,N_6738,N_7447);
nand U9481 (N_9481,N_7080,N_6252);
xnor U9482 (N_9482,N_6620,N_7674);
and U9483 (N_9483,N_7933,N_7247);
or U9484 (N_9484,N_6153,N_6924);
and U9485 (N_9485,N_7468,N_7489);
or U9486 (N_9486,N_6946,N_7377);
nor U9487 (N_9487,N_7645,N_7779);
and U9488 (N_9488,N_6609,N_6434);
or U9489 (N_9489,N_6312,N_6973);
xnor U9490 (N_9490,N_6705,N_6989);
xor U9491 (N_9491,N_7784,N_6782);
xor U9492 (N_9492,N_6978,N_7841);
and U9493 (N_9493,N_7582,N_7166);
xnor U9494 (N_9494,N_6171,N_7027);
and U9495 (N_9495,N_7470,N_6938);
nor U9496 (N_9496,N_7888,N_7818);
or U9497 (N_9497,N_7649,N_6869);
nor U9498 (N_9498,N_6855,N_6223);
xor U9499 (N_9499,N_6397,N_7757);
nor U9500 (N_9500,N_6626,N_7618);
or U9501 (N_9501,N_6575,N_6671);
nor U9502 (N_9502,N_6375,N_7635);
xor U9503 (N_9503,N_7227,N_7975);
nor U9504 (N_9504,N_7375,N_6358);
nor U9505 (N_9505,N_6961,N_6915);
xor U9506 (N_9506,N_6935,N_6035);
xnor U9507 (N_9507,N_6615,N_6383);
nand U9508 (N_9508,N_7593,N_6811);
nand U9509 (N_9509,N_7277,N_7505);
xnor U9510 (N_9510,N_7356,N_6330);
or U9511 (N_9511,N_7271,N_6414);
and U9512 (N_9512,N_7262,N_6497);
or U9513 (N_9513,N_6223,N_6986);
or U9514 (N_9514,N_6836,N_6311);
or U9515 (N_9515,N_7818,N_6402);
xor U9516 (N_9516,N_7707,N_6174);
nand U9517 (N_9517,N_7791,N_6424);
and U9518 (N_9518,N_6518,N_7377);
nand U9519 (N_9519,N_7928,N_7736);
nand U9520 (N_9520,N_7406,N_7999);
and U9521 (N_9521,N_7802,N_7776);
nor U9522 (N_9522,N_7789,N_7670);
or U9523 (N_9523,N_7683,N_7220);
nand U9524 (N_9524,N_6898,N_7304);
xnor U9525 (N_9525,N_7934,N_6736);
nor U9526 (N_9526,N_6393,N_7796);
and U9527 (N_9527,N_6040,N_6419);
nor U9528 (N_9528,N_7760,N_7883);
and U9529 (N_9529,N_6514,N_7030);
and U9530 (N_9530,N_7239,N_7496);
xor U9531 (N_9531,N_6941,N_7638);
and U9532 (N_9532,N_7490,N_6251);
xnor U9533 (N_9533,N_7069,N_7115);
xor U9534 (N_9534,N_7092,N_7304);
and U9535 (N_9535,N_7405,N_7056);
and U9536 (N_9536,N_7043,N_7622);
nor U9537 (N_9537,N_7214,N_7811);
xor U9538 (N_9538,N_7164,N_7456);
nor U9539 (N_9539,N_6405,N_7064);
and U9540 (N_9540,N_7106,N_7286);
xor U9541 (N_9541,N_7364,N_7832);
and U9542 (N_9542,N_6764,N_6398);
and U9543 (N_9543,N_7000,N_7448);
and U9544 (N_9544,N_7129,N_6289);
xor U9545 (N_9545,N_7384,N_7884);
xor U9546 (N_9546,N_6947,N_7614);
xor U9547 (N_9547,N_6953,N_7859);
nor U9548 (N_9548,N_6268,N_7494);
xnor U9549 (N_9549,N_7582,N_6152);
and U9550 (N_9550,N_7663,N_6000);
or U9551 (N_9551,N_6085,N_6394);
nor U9552 (N_9552,N_6082,N_7399);
xnor U9553 (N_9553,N_7160,N_7521);
or U9554 (N_9554,N_7310,N_7065);
nand U9555 (N_9555,N_7437,N_7721);
nor U9556 (N_9556,N_6034,N_6310);
xor U9557 (N_9557,N_7599,N_7914);
nor U9558 (N_9558,N_7839,N_6840);
xor U9559 (N_9559,N_6307,N_6530);
or U9560 (N_9560,N_6064,N_6156);
and U9561 (N_9561,N_6944,N_7973);
and U9562 (N_9562,N_7149,N_7014);
nor U9563 (N_9563,N_7703,N_7317);
xor U9564 (N_9564,N_7798,N_7459);
or U9565 (N_9565,N_7678,N_7281);
xnor U9566 (N_9566,N_7967,N_7445);
and U9567 (N_9567,N_7593,N_6822);
and U9568 (N_9568,N_6018,N_7700);
xnor U9569 (N_9569,N_7255,N_6023);
and U9570 (N_9570,N_6947,N_7682);
xnor U9571 (N_9571,N_7670,N_7942);
and U9572 (N_9572,N_7887,N_7987);
nand U9573 (N_9573,N_7966,N_7324);
or U9574 (N_9574,N_7908,N_6397);
and U9575 (N_9575,N_7540,N_6162);
xor U9576 (N_9576,N_6585,N_6230);
or U9577 (N_9577,N_7737,N_6303);
and U9578 (N_9578,N_7490,N_6482);
or U9579 (N_9579,N_7680,N_6271);
nor U9580 (N_9580,N_7833,N_6321);
xnor U9581 (N_9581,N_7634,N_7941);
and U9582 (N_9582,N_7905,N_6832);
xor U9583 (N_9583,N_7800,N_7887);
and U9584 (N_9584,N_6102,N_7999);
nand U9585 (N_9585,N_6853,N_6386);
and U9586 (N_9586,N_6944,N_6000);
nor U9587 (N_9587,N_6316,N_6518);
nor U9588 (N_9588,N_7577,N_6809);
nor U9589 (N_9589,N_6068,N_7905);
nor U9590 (N_9590,N_6491,N_7588);
and U9591 (N_9591,N_6295,N_6255);
nor U9592 (N_9592,N_7585,N_7713);
and U9593 (N_9593,N_7352,N_7066);
nor U9594 (N_9594,N_6937,N_7964);
nand U9595 (N_9595,N_7092,N_6348);
or U9596 (N_9596,N_7470,N_6432);
and U9597 (N_9597,N_7211,N_7403);
nand U9598 (N_9598,N_7726,N_7730);
nor U9599 (N_9599,N_6125,N_7684);
nand U9600 (N_9600,N_6013,N_6860);
nand U9601 (N_9601,N_6786,N_6639);
xor U9602 (N_9602,N_6681,N_6648);
nand U9603 (N_9603,N_7604,N_6845);
and U9604 (N_9604,N_7149,N_6560);
and U9605 (N_9605,N_7139,N_7348);
or U9606 (N_9606,N_6282,N_6580);
nand U9607 (N_9607,N_7686,N_7743);
xnor U9608 (N_9608,N_6900,N_7183);
and U9609 (N_9609,N_6623,N_6033);
nand U9610 (N_9610,N_7746,N_7173);
xor U9611 (N_9611,N_6658,N_7834);
xnor U9612 (N_9612,N_6928,N_6362);
and U9613 (N_9613,N_6223,N_7550);
nand U9614 (N_9614,N_7923,N_7025);
xor U9615 (N_9615,N_6478,N_7583);
xor U9616 (N_9616,N_7797,N_7616);
or U9617 (N_9617,N_7301,N_6840);
nand U9618 (N_9618,N_7697,N_6629);
xnor U9619 (N_9619,N_6804,N_6442);
nor U9620 (N_9620,N_6161,N_7184);
nor U9621 (N_9621,N_6211,N_7917);
or U9622 (N_9622,N_6949,N_6516);
and U9623 (N_9623,N_7427,N_6970);
nor U9624 (N_9624,N_6913,N_6125);
nor U9625 (N_9625,N_7140,N_7116);
nor U9626 (N_9626,N_7988,N_6689);
nor U9627 (N_9627,N_7878,N_6454);
xnor U9628 (N_9628,N_7188,N_7977);
nor U9629 (N_9629,N_6204,N_7490);
nor U9630 (N_9630,N_6871,N_6623);
and U9631 (N_9631,N_7058,N_7867);
or U9632 (N_9632,N_7832,N_7387);
nor U9633 (N_9633,N_6007,N_6083);
nor U9634 (N_9634,N_6624,N_7833);
nand U9635 (N_9635,N_6825,N_7959);
or U9636 (N_9636,N_7240,N_7022);
xor U9637 (N_9637,N_7341,N_7673);
and U9638 (N_9638,N_6935,N_6851);
or U9639 (N_9639,N_6646,N_7177);
xor U9640 (N_9640,N_6344,N_6085);
nand U9641 (N_9641,N_6579,N_6832);
xnor U9642 (N_9642,N_7341,N_7898);
xor U9643 (N_9643,N_7271,N_7074);
nand U9644 (N_9644,N_7931,N_6014);
and U9645 (N_9645,N_7847,N_6840);
or U9646 (N_9646,N_7632,N_7183);
or U9647 (N_9647,N_6695,N_7417);
nand U9648 (N_9648,N_7446,N_6450);
xor U9649 (N_9649,N_6526,N_7108);
xor U9650 (N_9650,N_7211,N_7206);
xnor U9651 (N_9651,N_7830,N_7549);
or U9652 (N_9652,N_6717,N_6226);
and U9653 (N_9653,N_7674,N_6264);
nor U9654 (N_9654,N_6203,N_7703);
and U9655 (N_9655,N_6636,N_6815);
or U9656 (N_9656,N_6804,N_7146);
xnor U9657 (N_9657,N_7532,N_7705);
nor U9658 (N_9658,N_7869,N_6400);
or U9659 (N_9659,N_7610,N_6192);
nor U9660 (N_9660,N_7976,N_7834);
or U9661 (N_9661,N_6041,N_6275);
and U9662 (N_9662,N_6657,N_6536);
nand U9663 (N_9663,N_6447,N_6855);
nand U9664 (N_9664,N_6979,N_6539);
or U9665 (N_9665,N_6237,N_7569);
or U9666 (N_9666,N_7714,N_6676);
xnor U9667 (N_9667,N_7663,N_6986);
and U9668 (N_9668,N_7313,N_6911);
or U9669 (N_9669,N_6121,N_6014);
nand U9670 (N_9670,N_7114,N_7586);
nand U9671 (N_9671,N_6184,N_6236);
nor U9672 (N_9672,N_7772,N_6339);
or U9673 (N_9673,N_6219,N_7399);
or U9674 (N_9674,N_7261,N_6294);
nand U9675 (N_9675,N_6936,N_7828);
or U9676 (N_9676,N_6667,N_7201);
nand U9677 (N_9677,N_6997,N_7396);
or U9678 (N_9678,N_6650,N_6511);
xor U9679 (N_9679,N_6255,N_7546);
nand U9680 (N_9680,N_7614,N_7314);
nor U9681 (N_9681,N_6118,N_6698);
nand U9682 (N_9682,N_6947,N_7913);
xor U9683 (N_9683,N_7346,N_6672);
nor U9684 (N_9684,N_6509,N_6742);
nor U9685 (N_9685,N_7610,N_6934);
xor U9686 (N_9686,N_7937,N_7389);
and U9687 (N_9687,N_6615,N_7317);
xor U9688 (N_9688,N_6310,N_7374);
or U9689 (N_9689,N_7632,N_7362);
xor U9690 (N_9690,N_6347,N_7005);
nor U9691 (N_9691,N_6291,N_6528);
nor U9692 (N_9692,N_7107,N_7342);
or U9693 (N_9693,N_6200,N_7254);
or U9694 (N_9694,N_6323,N_6470);
nor U9695 (N_9695,N_7009,N_6587);
nor U9696 (N_9696,N_7071,N_6815);
nor U9697 (N_9697,N_7846,N_7728);
or U9698 (N_9698,N_6824,N_6541);
or U9699 (N_9699,N_7075,N_6163);
and U9700 (N_9700,N_6452,N_6227);
nor U9701 (N_9701,N_7348,N_6058);
nand U9702 (N_9702,N_7069,N_7328);
nor U9703 (N_9703,N_7469,N_7185);
xor U9704 (N_9704,N_6189,N_6782);
or U9705 (N_9705,N_7424,N_6890);
xnor U9706 (N_9706,N_6041,N_7708);
or U9707 (N_9707,N_6791,N_6514);
nand U9708 (N_9708,N_6352,N_6197);
and U9709 (N_9709,N_7482,N_6358);
nor U9710 (N_9710,N_7980,N_7829);
nand U9711 (N_9711,N_7262,N_7977);
nand U9712 (N_9712,N_6497,N_6255);
nand U9713 (N_9713,N_6282,N_7265);
xor U9714 (N_9714,N_6476,N_6927);
or U9715 (N_9715,N_7986,N_6903);
or U9716 (N_9716,N_7429,N_7219);
xor U9717 (N_9717,N_6689,N_6519);
nor U9718 (N_9718,N_7446,N_7507);
nor U9719 (N_9719,N_7423,N_6572);
and U9720 (N_9720,N_7869,N_7414);
and U9721 (N_9721,N_6575,N_7541);
nand U9722 (N_9722,N_6718,N_6200);
xor U9723 (N_9723,N_7225,N_6948);
nor U9724 (N_9724,N_7959,N_6344);
and U9725 (N_9725,N_6079,N_7122);
nor U9726 (N_9726,N_7557,N_7627);
nand U9727 (N_9727,N_7348,N_6779);
and U9728 (N_9728,N_6832,N_7807);
xnor U9729 (N_9729,N_7282,N_6475);
or U9730 (N_9730,N_7976,N_6511);
xnor U9731 (N_9731,N_6756,N_6924);
nor U9732 (N_9732,N_7482,N_7008);
and U9733 (N_9733,N_6700,N_6116);
and U9734 (N_9734,N_7030,N_6052);
xnor U9735 (N_9735,N_6597,N_6087);
nand U9736 (N_9736,N_7274,N_7188);
xnor U9737 (N_9737,N_6387,N_7889);
or U9738 (N_9738,N_7490,N_7241);
and U9739 (N_9739,N_7259,N_7204);
or U9740 (N_9740,N_6862,N_7884);
and U9741 (N_9741,N_6608,N_7991);
nor U9742 (N_9742,N_7932,N_6249);
nor U9743 (N_9743,N_6966,N_6442);
nand U9744 (N_9744,N_7463,N_7988);
or U9745 (N_9745,N_6549,N_6047);
nand U9746 (N_9746,N_7511,N_6749);
nor U9747 (N_9747,N_6978,N_7732);
nor U9748 (N_9748,N_6961,N_7084);
nor U9749 (N_9749,N_6126,N_6491);
nand U9750 (N_9750,N_6230,N_7346);
nor U9751 (N_9751,N_7742,N_7305);
nor U9752 (N_9752,N_7867,N_7370);
or U9753 (N_9753,N_7642,N_7856);
xnor U9754 (N_9754,N_7988,N_7241);
or U9755 (N_9755,N_7910,N_7437);
nand U9756 (N_9756,N_7001,N_6491);
xor U9757 (N_9757,N_7980,N_6129);
nor U9758 (N_9758,N_7031,N_7116);
and U9759 (N_9759,N_6760,N_7807);
nor U9760 (N_9760,N_6022,N_7221);
xor U9761 (N_9761,N_7766,N_7701);
nor U9762 (N_9762,N_6968,N_7768);
nor U9763 (N_9763,N_6685,N_6458);
and U9764 (N_9764,N_7628,N_6307);
and U9765 (N_9765,N_6466,N_6117);
nand U9766 (N_9766,N_7998,N_7049);
nor U9767 (N_9767,N_7219,N_7267);
or U9768 (N_9768,N_6377,N_7941);
xor U9769 (N_9769,N_7422,N_7352);
and U9770 (N_9770,N_7839,N_6303);
and U9771 (N_9771,N_6526,N_7420);
xor U9772 (N_9772,N_6916,N_6178);
nand U9773 (N_9773,N_6033,N_6158);
nor U9774 (N_9774,N_6818,N_7278);
xor U9775 (N_9775,N_7497,N_6194);
and U9776 (N_9776,N_7061,N_6060);
and U9777 (N_9777,N_6366,N_6014);
nor U9778 (N_9778,N_7698,N_7659);
and U9779 (N_9779,N_6407,N_7410);
or U9780 (N_9780,N_6449,N_6720);
and U9781 (N_9781,N_7691,N_6703);
nand U9782 (N_9782,N_6359,N_6978);
and U9783 (N_9783,N_7670,N_7732);
and U9784 (N_9784,N_6148,N_7761);
nor U9785 (N_9785,N_7475,N_6536);
or U9786 (N_9786,N_7345,N_7060);
or U9787 (N_9787,N_6854,N_6990);
and U9788 (N_9788,N_7238,N_7109);
and U9789 (N_9789,N_7955,N_7146);
and U9790 (N_9790,N_6984,N_7807);
nand U9791 (N_9791,N_6404,N_7804);
nor U9792 (N_9792,N_7527,N_6804);
and U9793 (N_9793,N_7052,N_6540);
or U9794 (N_9794,N_7678,N_7298);
and U9795 (N_9795,N_7189,N_7533);
or U9796 (N_9796,N_6801,N_6162);
nor U9797 (N_9797,N_7679,N_6468);
nor U9798 (N_9798,N_7261,N_6758);
or U9799 (N_9799,N_6322,N_6687);
and U9800 (N_9800,N_6466,N_6880);
or U9801 (N_9801,N_6091,N_7813);
and U9802 (N_9802,N_7823,N_6504);
and U9803 (N_9803,N_7704,N_6266);
or U9804 (N_9804,N_6620,N_6613);
or U9805 (N_9805,N_7167,N_6033);
or U9806 (N_9806,N_7836,N_7210);
or U9807 (N_9807,N_6312,N_6000);
xnor U9808 (N_9808,N_6435,N_6897);
and U9809 (N_9809,N_6160,N_7681);
or U9810 (N_9810,N_6757,N_6792);
or U9811 (N_9811,N_6427,N_7274);
xor U9812 (N_9812,N_6980,N_6372);
nand U9813 (N_9813,N_6770,N_6398);
nand U9814 (N_9814,N_6489,N_6179);
nor U9815 (N_9815,N_6903,N_6250);
and U9816 (N_9816,N_6666,N_7062);
or U9817 (N_9817,N_7730,N_7937);
or U9818 (N_9818,N_7834,N_7989);
nor U9819 (N_9819,N_7778,N_6541);
nand U9820 (N_9820,N_6577,N_6735);
nor U9821 (N_9821,N_7027,N_6235);
xor U9822 (N_9822,N_7557,N_7772);
or U9823 (N_9823,N_6515,N_6976);
or U9824 (N_9824,N_7550,N_7357);
xnor U9825 (N_9825,N_7221,N_6588);
and U9826 (N_9826,N_7165,N_7116);
nand U9827 (N_9827,N_6117,N_7350);
and U9828 (N_9828,N_6817,N_7850);
and U9829 (N_9829,N_7569,N_7255);
xnor U9830 (N_9830,N_6323,N_7663);
or U9831 (N_9831,N_7371,N_6085);
nor U9832 (N_9832,N_7259,N_7636);
and U9833 (N_9833,N_7363,N_6887);
or U9834 (N_9834,N_7366,N_7312);
or U9835 (N_9835,N_6572,N_7795);
and U9836 (N_9836,N_7365,N_6505);
or U9837 (N_9837,N_6075,N_7549);
nand U9838 (N_9838,N_6548,N_6301);
nor U9839 (N_9839,N_7573,N_7505);
nor U9840 (N_9840,N_7414,N_7297);
nor U9841 (N_9841,N_6645,N_6151);
xnor U9842 (N_9842,N_6592,N_6725);
and U9843 (N_9843,N_6304,N_6486);
xnor U9844 (N_9844,N_7253,N_7543);
or U9845 (N_9845,N_7291,N_6734);
nand U9846 (N_9846,N_7676,N_7266);
nand U9847 (N_9847,N_7451,N_6936);
or U9848 (N_9848,N_7492,N_7628);
and U9849 (N_9849,N_6780,N_6421);
nand U9850 (N_9850,N_6834,N_7877);
and U9851 (N_9851,N_7069,N_7723);
xor U9852 (N_9852,N_6139,N_7232);
and U9853 (N_9853,N_6138,N_6640);
nor U9854 (N_9854,N_7120,N_7790);
nor U9855 (N_9855,N_6082,N_7628);
nand U9856 (N_9856,N_7739,N_7783);
and U9857 (N_9857,N_7137,N_7101);
xor U9858 (N_9858,N_6148,N_6865);
and U9859 (N_9859,N_7825,N_7980);
xor U9860 (N_9860,N_7144,N_7635);
and U9861 (N_9861,N_7659,N_6549);
xor U9862 (N_9862,N_6712,N_6114);
nand U9863 (N_9863,N_6411,N_7633);
and U9864 (N_9864,N_6423,N_7939);
nand U9865 (N_9865,N_6433,N_7681);
or U9866 (N_9866,N_6609,N_6703);
or U9867 (N_9867,N_6940,N_6433);
or U9868 (N_9868,N_6734,N_6814);
xnor U9869 (N_9869,N_6705,N_7532);
nand U9870 (N_9870,N_7971,N_7830);
nor U9871 (N_9871,N_6259,N_7246);
nor U9872 (N_9872,N_6580,N_7969);
nor U9873 (N_9873,N_6385,N_6237);
and U9874 (N_9874,N_6419,N_6746);
or U9875 (N_9875,N_7673,N_7845);
xor U9876 (N_9876,N_6248,N_7586);
or U9877 (N_9877,N_7729,N_6115);
and U9878 (N_9878,N_7605,N_6285);
nor U9879 (N_9879,N_6337,N_6232);
nand U9880 (N_9880,N_6086,N_7047);
xor U9881 (N_9881,N_7932,N_7853);
nand U9882 (N_9882,N_6876,N_7228);
nor U9883 (N_9883,N_7457,N_7273);
or U9884 (N_9884,N_6138,N_6126);
xor U9885 (N_9885,N_6931,N_7286);
or U9886 (N_9886,N_7789,N_7541);
nor U9887 (N_9887,N_6950,N_7473);
and U9888 (N_9888,N_6652,N_7723);
nor U9889 (N_9889,N_6978,N_6308);
nor U9890 (N_9890,N_7119,N_7920);
nand U9891 (N_9891,N_6545,N_6676);
or U9892 (N_9892,N_7092,N_6462);
and U9893 (N_9893,N_6372,N_6654);
or U9894 (N_9894,N_6075,N_6890);
nor U9895 (N_9895,N_6007,N_7713);
and U9896 (N_9896,N_7334,N_6013);
and U9897 (N_9897,N_6365,N_6104);
and U9898 (N_9898,N_7103,N_7632);
xnor U9899 (N_9899,N_6310,N_6773);
or U9900 (N_9900,N_6345,N_7127);
nand U9901 (N_9901,N_6061,N_6953);
or U9902 (N_9902,N_7717,N_7625);
or U9903 (N_9903,N_7645,N_7011);
xor U9904 (N_9904,N_6276,N_6164);
xor U9905 (N_9905,N_6474,N_7800);
nor U9906 (N_9906,N_6212,N_6754);
and U9907 (N_9907,N_7090,N_7038);
or U9908 (N_9908,N_7564,N_6279);
xor U9909 (N_9909,N_6454,N_6584);
xor U9910 (N_9910,N_7548,N_6596);
or U9911 (N_9911,N_7447,N_6714);
or U9912 (N_9912,N_6620,N_6789);
and U9913 (N_9913,N_6720,N_6874);
or U9914 (N_9914,N_7932,N_6675);
and U9915 (N_9915,N_7004,N_6654);
nor U9916 (N_9916,N_6394,N_7316);
xor U9917 (N_9917,N_6514,N_7322);
or U9918 (N_9918,N_6246,N_7782);
xnor U9919 (N_9919,N_7399,N_7283);
nor U9920 (N_9920,N_6932,N_7919);
and U9921 (N_9921,N_6242,N_6117);
or U9922 (N_9922,N_6782,N_6460);
nand U9923 (N_9923,N_7758,N_7915);
or U9924 (N_9924,N_6268,N_7058);
nor U9925 (N_9925,N_7719,N_6090);
xor U9926 (N_9926,N_6703,N_7651);
nand U9927 (N_9927,N_7571,N_6084);
xnor U9928 (N_9928,N_6396,N_6927);
or U9929 (N_9929,N_7268,N_7636);
nor U9930 (N_9930,N_6215,N_6578);
or U9931 (N_9931,N_6850,N_6239);
or U9932 (N_9932,N_6027,N_7915);
nor U9933 (N_9933,N_6953,N_7279);
nand U9934 (N_9934,N_6268,N_7750);
xor U9935 (N_9935,N_6948,N_7410);
nand U9936 (N_9936,N_7620,N_7261);
nand U9937 (N_9937,N_7003,N_7030);
nor U9938 (N_9938,N_7747,N_6793);
nand U9939 (N_9939,N_7971,N_7181);
nor U9940 (N_9940,N_6840,N_7289);
xnor U9941 (N_9941,N_6969,N_6023);
or U9942 (N_9942,N_7040,N_7951);
nor U9943 (N_9943,N_7146,N_7472);
nor U9944 (N_9944,N_7017,N_7762);
and U9945 (N_9945,N_7129,N_7031);
nand U9946 (N_9946,N_7066,N_7243);
nand U9947 (N_9947,N_6296,N_6644);
nor U9948 (N_9948,N_6314,N_7386);
nor U9949 (N_9949,N_6648,N_7136);
nor U9950 (N_9950,N_6341,N_7197);
nand U9951 (N_9951,N_6996,N_7913);
xor U9952 (N_9952,N_6007,N_7642);
or U9953 (N_9953,N_7568,N_7929);
xor U9954 (N_9954,N_6021,N_6568);
xor U9955 (N_9955,N_7097,N_6592);
nor U9956 (N_9956,N_7420,N_7613);
nand U9957 (N_9957,N_7801,N_6508);
and U9958 (N_9958,N_7464,N_6908);
nor U9959 (N_9959,N_7958,N_6399);
xor U9960 (N_9960,N_6724,N_7019);
or U9961 (N_9961,N_7407,N_7371);
or U9962 (N_9962,N_6547,N_6054);
and U9963 (N_9963,N_7850,N_6509);
xnor U9964 (N_9964,N_7732,N_7396);
and U9965 (N_9965,N_6658,N_6698);
xnor U9966 (N_9966,N_6546,N_6797);
nor U9967 (N_9967,N_6252,N_7828);
xnor U9968 (N_9968,N_7551,N_7829);
or U9969 (N_9969,N_6001,N_7756);
nor U9970 (N_9970,N_7504,N_7408);
or U9971 (N_9971,N_6231,N_7612);
or U9972 (N_9972,N_6838,N_7661);
nor U9973 (N_9973,N_7423,N_7728);
and U9974 (N_9974,N_7979,N_7474);
nor U9975 (N_9975,N_6804,N_6130);
and U9976 (N_9976,N_6050,N_6977);
nand U9977 (N_9977,N_6104,N_6935);
nand U9978 (N_9978,N_6495,N_7609);
nor U9979 (N_9979,N_7029,N_7683);
xnor U9980 (N_9980,N_6407,N_7565);
nor U9981 (N_9981,N_6736,N_6105);
and U9982 (N_9982,N_6480,N_6879);
nand U9983 (N_9983,N_6868,N_6889);
and U9984 (N_9984,N_7909,N_6054);
xor U9985 (N_9985,N_7649,N_7491);
nand U9986 (N_9986,N_7466,N_7468);
xor U9987 (N_9987,N_6023,N_6447);
or U9988 (N_9988,N_7060,N_6596);
nor U9989 (N_9989,N_6814,N_6975);
xnor U9990 (N_9990,N_6688,N_7062);
nor U9991 (N_9991,N_7356,N_7993);
nor U9992 (N_9992,N_6184,N_6457);
or U9993 (N_9993,N_6617,N_7443);
and U9994 (N_9994,N_7336,N_6893);
nand U9995 (N_9995,N_7896,N_7879);
and U9996 (N_9996,N_6840,N_7264);
xnor U9997 (N_9997,N_6221,N_6655);
xnor U9998 (N_9998,N_7122,N_6608);
and U9999 (N_9999,N_7092,N_6963);
and UO_0 (O_0,N_8585,N_9615);
xnor UO_1 (O_1,N_9285,N_9466);
or UO_2 (O_2,N_9268,N_9757);
and UO_3 (O_3,N_8476,N_9951);
or UO_4 (O_4,N_8578,N_8520);
and UO_5 (O_5,N_8496,N_9525);
or UO_6 (O_6,N_9270,N_8523);
or UO_7 (O_7,N_9831,N_8437);
nand UO_8 (O_8,N_9988,N_9290);
and UO_9 (O_9,N_8226,N_8161);
and UO_10 (O_10,N_8868,N_8611);
or UO_11 (O_11,N_9494,N_9950);
nor UO_12 (O_12,N_9942,N_9987);
and UO_13 (O_13,N_9781,N_8512);
nand UO_14 (O_14,N_9884,N_9720);
and UO_15 (O_15,N_8278,N_9899);
nor UO_16 (O_16,N_9046,N_9262);
xnor UO_17 (O_17,N_8786,N_8613);
nand UO_18 (O_18,N_9275,N_9581);
nand UO_19 (O_19,N_8045,N_9598);
xnor UO_20 (O_20,N_9177,N_9080);
and UO_21 (O_21,N_9448,N_8475);
xor UO_22 (O_22,N_9964,N_9040);
and UO_23 (O_23,N_9733,N_8406);
nand UO_24 (O_24,N_9149,N_9137);
or UO_25 (O_25,N_9447,N_8127);
or UO_26 (O_26,N_8194,N_9308);
xor UO_27 (O_27,N_9032,N_8415);
and UO_28 (O_28,N_9976,N_8261);
and UO_29 (O_29,N_8183,N_9963);
or UO_30 (O_30,N_8800,N_8925);
nor UO_31 (O_31,N_8423,N_8486);
or UO_32 (O_32,N_8900,N_8802);
xor UO_33 (O_33,N_8279,N_9854);
xor UO_34 (O_34,N_9572,N_9990);
or UO_35 (O_35,N_9858,N_9147);
nor UO_36 (O_36,N_9370,N_8391);
xnor UO_37 (O_37,N_8402,N_9979);
or UO_38 (O_38,N_8084,N_9485);
nand UO_39 (O_39,N_9429,N_9413);
or UO_40 (O_40,N_9744,N_9315);
nand UO_41 (O_41,N_8690,N_8990);
and UO_42 (O_42,N_8721,N_9240);
nand UO_43 (O_43,N_9197,N_8381);
nand UO_44 (O_44,N_8352,N_8844);
nand UO_45 (O_45,N_9484,N_9419);
and UO_46 (O_46,N_8995,N_8787);
xnor UO_47 (O_47,N_8228,N_8292);
xnor UO_48 (O_48,N_8389,N_9341);
xnor UO_49 (O_49,N_8846,N_9031);
or UO_50 (O_50,N_9168,N_8863);
xnor UO_51 (O_51,N_8707,N_8098);
nor UO_52 (O_52,N_8984,N_8674);
xor UO_53 (O_53,N_9667,N_9521);
nand UO_54 (O_54,N_8448,N_8068);
and UO_55 (O_55,N_9300,N_8086);
and UO_56 (O_56,N_8621,N_8688);
nor UO_57 (O_57,N_8174,N_9456);
or UO_58 (O_58,N_8092,N_9420);
xnor UO_59 (O_59,N_8275,N_9391);
or UO_60 (O_60,N_9029,N_9962);
nor UO_61 (O_61,N_9365,N_8967);
or UO_62 (O_62,N_9647,N_8972);
and UO_63 (O_63,N_9425,N_8214);
xor UO_64 (O_64,N_9575,N_8701);
xor UO_65 (O_65,N_8359,N_8249);
nor UO_66 (O_66,N_8252,N_9444);
and UO_67 (O_67,N_9739,N_8923);
nor UO_68 (O_68,N_8162,N_8399);
and UO_69 (O_69,N_8042,N_8717);
nand UO_70 (O_70,N_9660,N_9296);
nor UO_71 (O_71,N_8499,N_9714);
or UO_72 (O_72,N_8041,N_8856);
and UO_73 (O_73,N_9779,N_9941);
or UO_74 (O_74,N_9056,N_9504);
and UO_75 (O_75,N_9669,N_9401);
and UO_76 (O_76,N_8273,N_8792);
nand UO_77 (O_77,N_9167,N_8341);
and UO_78 (O_78,N_9001,N_8811);
nand UO_79 (O_79,N_8977,N_8747);
or UO_80 (O_80,N_9568,N_8938);
or UO_81 (O_81,N_8016,N_8114);
and UO_82 (O_82,N_9061,N_8018);
nor UO_83 (O_83,N_9476,N_8675);
or UO_84 (O_84,N_9576,N_8858);
xnor UO_85 (O_85,N_8372,N_9299);
nand UO_86 (O_86,N_8227,N_8011);
nor UO_87 (O_87,N_8907,N_8232);
xnor UO_88 (O_88,N_8693,N_9938);
nand UO_89 (O_89,N_9688,N_9074);
and UO_90 (O_90,N_8122,N_9919);
nor UO_91 (O_91,N_9491,N_9678);
or UO_92 (O_92,N_8049,N_9666);
xnor UO_93 (O_93,N_8366,N_8296);
nor UO_94 (O_94,N_8681,N_8460);
xnor UO_95 (O_95,N_9217,N_9064);
and UO_96 (O_96,N_8013,N_8036);
and UO_97 (O_97,N_8123,N_8766);
xor UO_98 (O_98,N_8739,N_9821);
xnor UO_99 (O_99,N_9828,N_8742);
or UO_100 (O_100,N_8009,N_8640);
xor UO_101 (O_101,N_8764,N_9418);
nand UO_102 (O_102,N_8582,N_9057);
or UO_103 (O_103,N_9215,N_9993);
xor UO_104 (O_104,N_8875,N_9120);
xor UO_105 (O_105,N_9743,N_9742);
nor UO_106 (O_106,N_9297,N_8153);
and UO_107 (O_107,N_8477,N_9354);
xor UO_108 (O_108,N_8973,N_9277);
xor UO_109 (O_109,N_9642,N_9664);
nor UO_110 (O_110,N_8978,N_9923);
and UO_111 (O_111,N_9550,N_8994);
and UO_112 (O_112,N_9211,N_9780);
and UO_113 (O_113,N_9819,N_8403);
nand UO_114 (O_114,N_8132,N_9195);
and UO_115 (O_115,N_9128,N_9477);
or UO_116 (O_116,N_9981,N_9972);
or UO_117 (O_117,N_9661,N_9908);
nor UO_118 (O_118,N_8697,N_8609);
and UO_119 (O_119,N_8720,N_9247);
xnor UO_120 (O_120,N_9105,N_8119);
nor UO_121 (O_121,N_9018,N_8788);
xor UO_122 (O_122,N_9059,N_9327);
nand UO_123 (O_123,N_9827,N_9852);
and UO_124 (O_124,N_9912,N_8926);
xnor UO_125 (O_125,N_9102,N_8861);
or UO_126 (O_126,N_8615,N_9515);
and UO_127 (O_127,N_8441,N_8628);
nor UO_128 (O_128,N_9547,N_9324);
and UO_129 (O_129,N_8625,N_8173);
and UO_130 (O_130,N_9857,N_8506);
xnor UO_131 (O_131,N_8083,N_8418);
xnor UO_132 (O_132,N_9383,N_8446);
nor UO_133 (O_133,N_8427,N_8121);
or UO_134 (O_134,N_8837,N_9362);
nand UO_135 (O_135,N_9233,N_8223);
nand UO_136 (O_136,N_8367,N_9999);
or UO_137 (O_137,N_8558,N_8789);
or UO_138 (O_138,N_8111,N_9797);
or UO_139 (O_139,N_9850,N_9088);
xnor UO_140 (O_140,N_9093,N_8642);
nor UO_141 (O_141,N_8164,N_8224);
nand UO_142 (O_142,N_8708,N_9148);
nand UO_143 (O_143,N_8833,N_9288);
and UO_144 (O_144,N_9124,N_8037);
xor UO_145 (O_145,N_9493,N_9529);
nor UO_146 (O_146,N_8234,N_9778);
and UO_147 (O_147,N_8646,N_8565);
or UO_148 (O_148,N_9690,N_9470);
nor UO_149 (O_149,N_9867,N_8159);
or UO_150 (O_150,N_9671,N_8516);
and UO_151 (O_151,N_9198,N_9263);
xnor UO_152 (O_152,N_8485,N_8848);
xnor UO_153 (O_153,N_9414,N_8716);
nand UO_154 (O_154,N_8061,N_9075);
and UO_155 (O_155,N_8665,N_8313);
xnor UO_156 (O_156,N_9335,N_8482);
nand UO_157 (O_157,N_8746,N_8768);
nand UO_158 (O_158,N_8257,N_9980);
nor UO_159 (O_159,N_8942,N_8650);
nor UO_160 (O_160,N_8364,N_9604);
xnor UO_161 (O_161,N_8745,N_9675);
xnor UO_162 (O_162,N_8535,N_8094);
nand UO_163 (O_163,N_9531,N_8656);
nand UO_164 (O_164,N_8350,N_8060);
or UO_165 (O_165,N_8566,N_9767);
and UO_166 (O_166,N_8019,N_9726);
nor UO_167 (O_167,N_8553,N_9936);
xor UO_168 (O_168,N_9388,N_8479);
xor UO_169 (O_169,N_9738,N_9874);
nor UO_170 (O_170,N_9906,N_8731);
or UO_171 (O_171,N_8758,N_8100);
nor UO_172 (O_172,N_9127,N_9013);
or UO_173 (O_173,N_9573,N_8362);
or UO_174 (O_174,N_9756,N_8825);
or UO_175 (O_175,N_8304,N_9792);
and UO_176 (O_176,N_8443,N_8300);
or UO_177 (O_177,N_8102,N_8676);
or UO_178 (O_178,N_8073,N_9620);
and UO_179 (O_179,N_9537,N_8927);
xor UO_180 (O_180,N_9848,N_9161);
and UO_181 (O_181,N_9344,N_9927);
nor UO_182 (O_182,N_8895,N_9452);
xnor UO_183 (O_183,N_9788,N_9928);
and UO_184 (O_184,N_9823,N_9995);
and UO_185 (O_185,N_8408,N_9037);
xor UO_186 (O_186,N_9350,N_8230);
and UO_187 (O_187,N_9238,N_9814);
xnor UO_188 (O_188,N_8673,N_9321);
nor UO_189 (O_189,N_9378,N_9184);
nor UO_190 (O_190,N_9183,N_9934);
or UO_191 (O_191,N_8590,N_9665);
nor UO_192 (O_192,N_9041,N_9699);
and UO_193 (O_193,N_8751,N_9313);
nor UO_194 (O_194,N_9891,N_8547);
or UO_195 (O_195,N_8954,N_9440);
nand UO_196 (O_196,N_9503,N_8556);
nor UO_197 (O_197,N_8879,N_9248);
or UO_198 (O_198,N_8712,N_8635);
nor UO_199 (O_199,N_9935,N_8149);
nand UO_200 (O_200,N_8729,N_8039);
nor UO_201 (O_201,N_9106,N_8644);
xor UO_202 (O_202,N_9385,N_9036);
or UO_203 (O_203,N_8333,N_9500);
nand UO_204 (O_204,N_8892,N_8245);
or UO_205 (O_205,N_9379,N_9600);
xor UO_206 (O_206,N_9333,N_8597);
nor UO_207 (O_207,N_9276,N_8189);
or UO_208 (O_208,N_8065,N_8794);
nor UO_209 (O_209,N_9790,N_8284);
nand UO_210 (O_210,N_8532,N_9367);
or UO_211 (O_211,N_8078,N_9880);
nand UO_212 (O_212,N_8821,N_9191);
and UO_213 (O_213,N_9117,N_9955);
and UO_214 (O_214,N_9317,N_9212);
or UO_215 (O_215,N_9736,N_8269);
or UO_216 (O_216,N_9590,N_9110);
or UO_217 (O_217,N_8006,N_9092);
nor UO_218 (O_218,N_9395,N_9178);
nor UO_219 (O_219,N_9889,N_8904);
nor UO_220 (O_220,N_8015,N_9325);
or UO_221 (O_221,N_8259,N_9314);
nand UO_222 (O_222,N_9236,N_9989);
nand UO_223 (O_223,N_8407,N_8434);
or UO_224 (O_224,N_9358,N_9833);
nand UO_225 (O_225,N_9023,N_9490);
xor UO_226 (O_226,N_9599,N_8891);
or UO_227 (O_227,N_8250,N_8521);
xor UO_228 (O_228,N_8812,N_8495);
nand UO_229 (O_229,N_8360,N_9707);
xor UO_230 (O_230,N_9614,N_8085);
and UO_231 (O_231,N_8680,N_9246);
xor UO_232 (O_232,N_8209,N_8193);
or UO_233 (O_233,N_8303,N_9312);
or UO_234 (O_234,N_8345,N_8283);
and UO_235 (O_235,N_8614,N_8822);
xor UO_236 (O_236,N_9230,N_9111);
and UO_237 (O_237,N_9291,N_8116);
nor UO_238 (O_238,N_8291,N_9533);
nor UO_239 (O_239,N_9301,N_8583);
nor UO_240 (O_240,N_8494,N_8139);
and UO_241 (O_241,N_8988,N_8101);
or UO_242 (O_242,N_9510,N_9638);
nand UO_243 (O_243,N_9925,N_8450);
nor UO_244 (O_244,N_8991,N_9557);
or UO_245 (O_245,N_9280,N_9498);
nand UO_246 (O_246,N_8975,N_8658);
and UO_247 (O_247,N_8603,N_9479);
and UO_248 (O_248,N_8809,N_8401);
nand UO_249 (O_249,N_9210,N_8574);
and UO_250 (O_250,N_8498,N_8618);
xnor UO_251 (O_251,N_8405,N_8157);
nand UO_252 (O_252,N_8593,N_8736);
xnor UO_253 (O_253,N_9715,N_9000);
xor UO_254 (O_254,N_8946,N_9135);
and UO_255 (O_255,N_8952,N_9794);
or UO_256 (O_256,N_9643,N_9644);
nor UO_257 (O_257,N_8976,N_9446);
nand UO_258 (O_258,N_8782,N_8480);
nand UO_259 (O_259,N_8150,N_8133);
xnor UO_260 (O_260,N_9645,N_9777);
xnor UO_261 (O_261,N_8236,N_9910);
xnor UO_262 (O_262,N_8726,N_9151);
or UO_263 (O_263,N_9108,N_9156);
nor UO_264 (O_264,N_9593,N_8957);
xnor UO_265 (O_265,N_9104,N_9534);
nand UO_266 (O_266,N_8217,N_8240);
nand UO_267 (O_267,N_8616,N_8444);
xor UO_268 (O_268,N_9261,N_8435);
or UO_269 (O_269,N_9454,N_8206);
nand UO_270 (O_270,N_9727,N_8519);
xor UO_271 (O_271,N_8033,N_9189);
or UO_272 (O_272,N_9766,N_9409);
or UO_273 (O_273,N_8177,N_8369);
and UO_274 (O_274,N_8666,N_8274);
nor UO_275 (O_275,N_8796,N_9250);
xnor UO_276 (O_276,N_9783,N_8867);
xor UO_277 (O_277,N_8180,N_8572);
nand UO_278 (O_278,N_8817,N_8562);
or UO_279 (O_279,N_8106,N_9750);
nor UO_280 (O_280,N_8000,N_8436);
or UO_281 (O_281,N_9795,N_9589);
nor UO_282 (O_282,N_9163,N_8327);
or UO_283 (O_283,N_9882,N_8508);
and UO_284 (O_284,N_8383,N_8513);
xor UO_285 (O_285,N_9602,N_8043);
nor UO_286 (O_286,N_8823,N_9706);
xnor UO_287 (O_287,N_9134,N_9641);
nor UO_288 (O_288,N_9451,N_9115);
or UO_289 (O_289,N_9509,N_8473);
xor UO_290 (O_290,N_9435,N_8683);
nand UO_291 (O_291,N_9588,N_8511);
and UO_292 (O_292,N_8373,N_9488);
nand UO_293 (O_293,N_9190,N_9810);
xnor UO_294 (O_294,N_8761,N_8564);
xnor UO_295 (O_295,N_9752,N_9754);
or UO_296 (O_296,N_8131,N_9540);
and UO_297 (O_297,N_8493,N_8312);
nand UO_298 (O_298,N_8467,N_9931);
nand UO_299 (O_299,N_9613,N_9621);
or UO_300 (O_300,N_9890,N_8941);
or UO_301 (O_301,N_9798,N_9293);
xnor UO_302 (O_302,N_9406,N_9961);
or UO_303 (O_303,N_9791,N_9186);
or UO_304 (O_304,N_8514,N_9911);
nand UO_305 (O_305,N_9717,N_9711);
nand UO_306 (O_306,N_8400,N_8134);
or UO_307 (O_307,N_9020,N_9450);
nor UO_308 (O_308,N_9097,N_8280);
nand UO_309 (O_309,N_8771,N_8687);
nand UO_310 (O_310,N_8035,N_9695);
and UO_311 (O_311,N_9465,N_8502);
xor UO_312 (O_312,N_9782,N_8798);
xnor UO_313 (O_313,N_9352,N_9216);
and UO_314 (O_314,N_9303,N_9787);
nor UO_315 (O_315,N_8357,N_8830);
nand UO_316 (O_316,N_9058,N_8982);
xor UO_317 (O_317,N_9486,N_9507);
or UO_318 (O_318,N_9357,N_8913);
xnor UO_319 (O_319,N_8810,N_9524);
or UO_320 (O_320,N_8202,N_8864);
xnor UO_321 (O_321,N_9812,N_8963);
or UO_322 (O_322,N_9400,N_9815);
nand UO_323 (O_323,N_8243,N_8774);
nor UO_324 (O_324,N_9753,N_8622);
or UO_325 (O_325,N_9996,N_9553);
nand UO_326 (O_326,N_8989,N_9121);
and UO_327 (O_327,N_8026,N_9703);
nor UO_328 (O_328,N_9868,N_9998);
or UO_329 (O_329,N_9326,N_9837);
nand UO_330 (O_330,N_9652,N_8933);
or UO_331 (O_331,N_8376,N_8860);
nor UO_332 (O_332,N_9086,N_8544);
nor UO_333 (O_333,N_9089,N_8432);
nand UO_334 (O_334,N_9113,N_8058);
nand UO_335 (O_335,N_9940,N_9763);
nor UO_336 (O_336,N_9271,N_9402);
or UO_337 (O_337,N_9255,N_9603);
or UO_338 (O_338,N_9079,N_9829);
and UO_339 (O_339,N_8417,N_8797);
and UO_340 (O_340,N_8152,N_8987);
nand UO_341 (O_341,N_8937,N_8072);
and UO_342 (O_342,N_9225,N_9471);
xor UO_343 (O_343,N_9719,N_8097);
xor UO_344 (O_344,N_8816,N_8487);
or UO_345 (O_345,N_8439,N_9294);
nand UO_346 (O_346,N_8874,N_8619);
nand UO_347 (O_347,N_9309,N_9208);
nand UO_348 (O_348,N_9244,N_9898);
or UO_349 (O_349,N_9519,N_8667);
xnor UO_350 (O_350,N_8067,N_9260);
nor UO_351 (O_351,N_8694,N_8002);
nand UO_352 (O_352,N_9251,N_9307);
or UO_353 (O_353,N_9234,N_8231);
xor UO_354 (O_354,N_9207,N_8958);
or UO_355 (O_355,N_9606,N_9655);
or UO_356 (O_356,N_9332,N_9144);
xor UO_357 (O_357,N_8679,N_9343);
and UO_358 (O_358,N_9626,N_9453);
xor UO_359 (O_359,N_9653,N_9336);
xnor UO_360 (O_360,N_8143,N_8470);
nor UO_361 (O_361,N_9501,N_8299);
or UO_362 (O_362,N_9619,N_8524);
nor UO_363 (O_363,N_8393,N_9202);
nor UO_364 (O_364,N_9571,N_8509);
or UO_365 (O_365,N_8354,N_8272);
xnor UO_366 (O_366,N_8428,N_9570);
nor UO_367 (O_367,N_8461,N_8997);
and UO_368 (O_368,N_9340,N_9813);
nand UO_369 (O_369,N_8375,N_9824);
or UO_370 (O_370,N_9939,N_8293);
and UO_371 (O_371,N_8160,N_8242);
nand UO_372 (O_372,N_9239,N_9683);
or UO_373 (O_373,N_9226,N_8754);
and UO_374 (O_374,N_9592,N_9982);
and UO_375 (O_375,N_9012,N_8331);
and UO_376 (O_376,N_8491,N_8251);
xor UO_377 (O_377,N_8749,N_8763);
nand UO_378 (O_378,N_9381,N_9607);
xnor UO_379 (O_379,N_8355,N_8709);
or UO_380 (O_380,N_9836,N_9895);
and UO_381 (O_381,N_9915,N_8192);
xor UO_382 (O_382,N_9055,N_8826);
nand UO_383 (O_383,N_9072,N_9970);
xor UO_384 (O_384,N_8268,N_9746);
nor UO_385 (O_385,N_9253,N_8843);
and UO_386 (O_386,N_9584,N_8090);
and UO_387 (O_387,N_9017,N_8539);
nand UO_388 (O_388,N_8911,N_8901);
nand UO_389 (O_389,N_8741,N_8145);
xnor UO_390 (O_390,N_8263,N_8993);
or UO_391 (O_391,N_9583,N_8713);
or UO_392 (O_392,N_8710,N_9944);
xnor UO_393 (O_393,N_8069,N_9424);
or UO_394 (O_394,N_9489,N_9724);
nor UO_395 (O_395,N_8244,N_8725);
nor UO_396 (O_396,N_8239,N_8641);
and UO_397 (O_397,N_8056,N_9081);
and UO_398 (O_398,N_8971,N_8914);
or UO_399 (O_399,N_8155,N_8657);
xor UO_400 (O_400,N_9769,N_9974);
or UO_401 (O_401,N_8865,N_9881);
and UO_402 (O_402,N_9803,N_8271);
or UO_403 (O_403,N_8610,N_9434);
and UO_404 (O_404,N_9920,N_8651);
nand UO_405 (O_405,N_8605,N_8334);
xnor UO_406 (O_406,N_9863,N_8385);
or UO_407 (O_407,N_9482,N_8536);
nor UO_408 (O_408,N_9096,N_9917);
nand UO_409 (O_409,N_8653,N_9070);
and UO_410 (O_410,N_8020,N_8528);
and UO_411 (O_411,N_9449,N_8141);
and UO_412 (O_412,N_8305,N_8216);
and UO_413 (O_413,N_9991,N_8107);
nor UO_414 (O_414,N_9580,N_9983);
xor UO_415 (O_415,N_8801,N_8440);
or UO_416 (O_416,N_9696,N_8577);
xnor UO_417 (O_417,N_8940,N_8778);
and UO_418 (O_418,N_8607,N_8596);
xor UO_419 (O_419,N_8307,N_9464);
or UO_420 (O_420,N_8265,N_8395);
and UO_421 (O_421,N_9003,N_9199);
nand UO_422 (O_422,N_9805,N_9807);
or UO_423 (O_423,N_9279,N_9608);
and UO_424 (O_424,N_8897,N_8003);
nand UO_425 (O_425,N_9337,N_9133);
nand UO_426 (O_426,N_8104,N_9052);
nand UO_427 (O_427,N_9822,N_8219);
xnor UO_428 (O_428,N_8735,N_8526);
or UO_429 (O_429,N_9461,N_8589);
and UO_430 (O_430,N_9249,N_8371);
nor UO_431 (O_431,N_9901,N_8627);
and UO_432 (O_432,N_8624,N_8581);
and UO_433 (O_433,N_8126,N_8483);
nor UO_434 (O_434,N_8256,N_9684);
nand UO_435 (O_435,N_8808,N_8178);
and UO_436 (O_436,N_9019,N_8733);
nor UO_437 (O_437,N_8167,N_9834);
or UO_438 (O_438,N_9138,N_8096);
xnor UO_439 (O_439,N_9832,N_9334);
xnor UO_440 (O_440,N_8636,N_9404);
nand UO_441 (O_441,N_8820,N_8884);
or UO_442 (O_442,N_8815,N_9508);
and UO_443 (O_443,N_8105,N_9705);
or UO_444 (O_444,N_8842,N_8422);
nor UO_445 (O_445,N_9038,N_9043);
nand UO_446 (O_446,N_9967,N_9897);
or UO_447 (O_447,N_8322,N_9241);
and UO_448 (O_448,N_9560,N_8113);
nor UO_449 (O_449,N_8617,N_8429);
xnor UO_450 (O_450,N_9468,N_8337);
or UO_451 (O_451,N_8248,N_8956);
or UO_452 (O_452,N_9549,N_9229);
and UO_453 (O_453,N_9126,N_8057);
nand UO_454 (O_454,N_8459,N_9100);
nand UO_455 (O_455,N_8790,N_8325);
or UO_456 (O_456,N_9558,N_8387);
and UO_457 (O_457,N_9725,N_8738);
nand UO_458 (O_458,N_9094,N_8108);
and UO_459 (O_459,N_8414,N_9264);
or UO_460 (O_460,N_8430,N_8534);
and UO_461 (O_461,N_9339,N_8919);
xnor UO_462 (O_462,N_8361,N_8246);
nor UO_463 (O_463,N_9016,N_8005);
nand UO_464 (O_464,N_9087,N_9994);
xnor UO_465 (O_465,N_8862,N_9789);
xor UO_466 (O_466,N_8876,N_8336);
nor UO_467 (O_467,N_9078,N_9235);
xor UO_468 (O_468,N_9188,N_8438);
or UO_469 (O_469,N_8445,N_8397);
and UO_470 (O_470,N_9033,N_8545);
and UO_471 (O_471,N_9160,N_8306);
nand UO_472 (O_472,N_9513,N_8503);
and UO_473 (O_473,N_9316,N_9165);
nor UO_474 (O_474,N_9693,N_8510);
and UO_475 (O_475,N_9022,N_9747);
nand UO_476 (O_476,N_9065,N_8970);
xor UO_477 (O_477,N_9745,N_9492);
and UO_478 (O_478,N_9103,N_9181);
or UO_479 (O_479,N_8260,N_8088);
nor UO_480 (O_480,N_9948,N_8222);
and UO_481 (O_481,N_8229,N_9728);
nor UO_482 (O_482,N_8922,N_8871);
xor UO_483 (O_483,N_9864,N_9310);
and UO_484 (O_484,N_8504,N_8158);
nand UO_485 (O_485,N_9770,N_8677);
nand UO_486 (O_486,N_8103,N_8267);
or UO_487 (O_487,N_8453,N_8968);
xnor UO_488 (O_488,N_8047,N_9953);
xor UO_489 (O_489,N_8686,N_9281);
nor UO_490 (O_490,N_8238,N_9755);
nor UO_491 (O_491,N_9194,N_8813);
xnor UO_492 (O_492,N_8320,N_9662);
or UO_493 (O_493,N_8527,N_9806);
nor UO_494 (O_494,N_9722,N_8398);
or UO_495 (O_495,N_8023,N_9616);
nand UO_496 (O_496,N_9286,N_8118);
nor UO_497 (O_497,N_8744,N_8087);
or UO_498 (O_498,N_8918,N_9349);
or UO_499 (O_499,N_8255,N_9390);
nor UO_500 (O_500,N_9629,N_8165);
xor UO_501 (O_501,N_8166,N_9839);
and UO_502 (O_502,N_9364,N_9360);
nand UO_503 (O_503,N_9257,N_9594);
nor UO_504 (O_504,N_9730,N_9201);
xnor UO_505 (O_505,N_9992,N_9909);
nand UO_506 (O_506,N_9030,N_8311);
and UO_507 (O_507,N_8814,N_9259);
nor UO_508 (O_508,N_9578,N_9841);
and UO_509 (O_509,N_9382,N_8404);
nand UO_510 (O_510,N_9222,N_8870);
xor UO_511 (O_511,N_8780,N_8253);
or UO_512 (O_512,N_9947,N_9816);
and UO_513 (O_513,N_9015,N_9353);
nand UO_514 (O_514,N_8386,N_9213);
and UO_515 (O_515,N_8384,N_8314);
and UO_516 (O_516,N_9430,N_9497);
and UO_517 (O_517,N_9691,N_9680);
xnor UO_518 (O_518,N_9760,N_9118);
or UO_519 (O_519,N_8038,N_8140);
and UO_520 (O_520,N_8835,N_8567);
or UO_521 (O_521,N_8481,N_8329);
or UO_522 (O_522,N_9496,N_8643);
nand UO_523 (O_523,N_8807,N_8136);
and UO_524 (O_524,N_9145,N_8601);
or UO_525 (O_525,N_8568,N_8916);
xnor UO_526 (O_526,N_9522,N_9157);
nand UO_527 (O_527,N_9623,N_9067);
nor UO_528 (O_528,N_8120,N_9597);
or UO_529 (O_529,N_8866,N_9021);
or UO_530 (O_530,N_9562,N_9505);
xnor UO_531 (O_531,N_9957,N_9826);
and UO_532 (O_532,N_9676,N_9702);
or UO_533 (O_533,N_8629,N_9221);
xor UO_534 (O_534,N_8454,N_9393);
xnor UO_535 (O_535,N_8203,N_8571);
nor UO_536 (O_536,N_8700,N_9502);
and UO_537 (O_537,N_9527,N_9267);
xnor UO_538 (O_538,N_8378,N_8929);
or UO_539 (O_539,N_9793,N_9320);
xnor UO_540 (O_540,N_8723,N_8237);
and UO_541 (O_541,N_8082,N_8775);
nand UO_542 (O_542,N_8760,N_8541);
or UO_543 (O_543,N_8670,N_8877);
or UO_544 (O_544,N_8080,N_9735);
or UO_545 (O_545,N_8351,N_9460);
nor UO_546 (O_546,N_8902,N_9376);
nor UO_547 (O_547,N_9561,N_8910);
nor UO_548 (O_548,N_9131,N_9929);
and UO_549 (O_549,N_8207,N_9532);
and UO_550 (O_550,N_9682,N_8301);
or UO_551 (O_551,N_8996,N_8550);
xnor UO_552 (O_552,N_8779,N_9687);
nor UO_553 (O_553,N_8623,N_9749);
nand UO_554 (O_554,N_9169,N_9965);
nand UO_555 (O_555,N_8962,N_9209);
or UO_556 (O_556,N_9526,N_9457);
nor UO_557 (O_557,N_8659,N_8594);
xor UO_558 (O_558,N_9069,N_9564);
xnor UO_559 (O_559,N_8769,N_9411);
xor UO_560 (O_560,N_8752,N_8648);
nor UO_561 (O_561,N_8580,N_9624);
nor UO_562 (O_562,N_9342,N_9175);
nor UO_563 (O_563,N_8287,N_9060);
nor UO_564 (O_564,N_9499,N_9002);
xor UO_565 (O_565,N_8053,N_9924);
and UO_566 (O_566,N_8295,N_8182);
nand UO_567 (O_567,N_9506,N_9997);
nor UO_568 (O_568,N_9851,N_8187);
xnor UO_569 (O_569,N_9164,N_8999);
nor UO_570 (O_570,N_9090,N_9764);
nor UO_571 (O_571,N_9116,N_8950);
and UO_572 (O_572,N_8592,N_9784);
nor UO_573 (O_573,N_8324,N_8330);
xnor UO_574 (O_574,N_8684,N_9761);
nor UO_575 (O_575,N_8409,N_9008);
or UO_576 (O_576,N_8947,N_8899);
nor UO_577 (O_577,N_9511,N_8290);
and UO_578 (O_578,N_8772,N_9563);
nor UO_579 (O_579,N_8691,N_8948);
nor UO_580 (O_580,N_9853,N_8767);
nor UO_581 (O_581,N_9254,N_9439);
xor UO_582 (O_582,N_8718,N_9284);
and UO_583 (O_583,N_8599,N_8606);
or UO_584 (O_584,N_8887,N_9265);
or UO_585 (O_585,N_9516,N_8965);
nor UO_586 (O_586,N_9896,N_8953);
nand UO_587 (O_587,N_8930,N_8492);
xnor UO_588 (O_588,N_8850,N_8678);
or UO_589 (O_589,N_8620,N_9886);
and UO_590 (O_590,N_9475,N_8579);
xor UO_591 (O_591,N_8420,N_9759);
xnor UO_592 (O_592,N_9258,N_8356);
nor UO_593 (O_593,N_9283,N_9952);
nor UO_594 (O_594,N_8457,N_9141);
xor UO_595 (O_595,N_9586,N_9182);
nor UO_596 (O_596,N_9883,N_9774);
or UO_597 (O_597,N_8734,N_9154);
nor UO_598 (O_598,N_8685,N_9099);
nor UO_599 (O_599,N_8264,N_8819);
and UO_600 (O_600,N_8791,N_9066);
or UO_601 (O_601,N_8980,N_9173);
nor UO_602 (O_602,N_9034,N_9407);
xor UO_603 (O_603,N_9956,N_8022);
or UO_604 (O_604,N_8829,N_9377);
and UO_605 (O_605,N_8600,N_8765);
nand UO_606 (O_606,N_9966,N_9921);
nor UO_607 (O_607,N_9721,N_9347);
or UO_608 (O_608,N_9845,N_9930);
xor UO_609 (O_609,N_8706,N_8878);
and UO_610 (O_610,N_9838,N_8931);
xnor UO_611 (O_611,N_9187,N_9051);
xnor UO_612 (O_612,N_9811,N_9129);
and UO_613 (O_613,N_9673,N_9818);
xnor UO_614 (O_614,N_8469,N_8185);
or UO_615 (O_615,N_9443,N_8591);
nand UO_616 (O_616,N_9926,N_9132);
nand UO_617 (O_617,N_8186,N_9885);
nand UO_618 (O_618,N_8818,N_9637);
or UO_619 (O_619,N_9905,N_9954);
nand UO_620 (O_620,N_9085,N_9656);
and UO_621 (O_621,N_8638,N_8692);
or UO_622 (O_622,N_8724,N_8235);
nor UO_623 (O_623,N_9101,N_9123);
xor UO_624 (O_624,N_8117,N_8655);
nor UO_625 (O_625,N_9958,N_8266);
nor UO_626 (O_626,N_9846,N_9577);
nor UO_627 (O_627,N_9681,N_8634);
or UO_628 (O_628,N_9716,N_9050);
nor UO_629 (O_629,N_9859,N_9668);
or UO_630 (O_630,N_8546,N_9762);
nand UO_631 (O_631,N_8955,N_8961);
nand UO_632 (O_632,N_9567,N_8233);
nand UO_633 (O_633,N_9847,N_8298);
xor UO_634 (O_634,N_8630,N_8944);
and UO_635 (O_635,N_8201,N_8560);
and UO_636 (O_636,N_8569,N_9609);
nand UO_637 (O_637,N_9801,N_9894);
xnor UO_638 (O_638,N_8063,N_9480);
xnor UO_639 (O_639,N_8943,N_9649);
nor UO_640 (O_640,N_8896,N_8317);
xnor UO_641 (O_641,N_9977,N_8985);
nand UO_642 (O_642,N_9916,N_8573);
xor UO_643 (O_643,N_8785,N_8054);
nor UO_644 (O_644,N_8857,N_9748);
or UO_645 (O_645,N_9605,N_9968);
nor UO_646 (O_646,N_8964,N_9266);
nand UO_647 (O_647,N_8890,N_9338);
nand UO_648 (O_648,N_9657,N_9758);
xor UO_649 (O_649,N_8012,N_9319);
xnor UO_650 (O_650,N_9635,N_8880);
nand UO_651 (O_651,N_9224,N_9799);
and UO_652 (O_652,N_8608,N_9692);
or UO_653 (O_653,N_9005,N_9463);
xnor UO_654 (O_654,N_9596,N_9196);
nor UO_655 (O_655,N_9566,N_8294);
nor UO_656 (O_656,N_9694,N_9306);
and UO_657 (O_657,N_9723,N_9913);
nand UO_658 (O_658,N_9933,N_9677);
xnor UO_659 (O_659,N_9304,N_8598);
and UO_660 (O_660,N_9904,N_8849);
and UO_661 (O_661,N_8631,N_9902);
nand UO_662 (O_662,N_9731,N_8932);
nor UO_663 (O_663,N_9751,N_8169);
and UO_664 (O_664,N_9384,N_8497);
nor UO_665 (O_665,N_8413,N_8342);
and UO_666 (O_666,N_9083,N_8066);
or UO_667 (O_667,N_8753,N_9467);
or UO_668 (O_668,N_9617,N_9119);
and UO_669 (O_669,N_9960,N_9672);
nand UO_670 (O_670,N_8431,N_9729);
and UO_671 (O_671,N_8200,N_9713);
nand UO_672 (O_672,N_9329,N_8840);
or UO_673 (O_673,N_8557,N_9025);
or UO_674 (O_674,N_9701,N_8883);
and UO_675 (O_675,N_8554,N_9945);
nand UO_676 (O_676,N_8211,N_8044);
nand UO_677 (O_677,N_9487,N_9146);
xnor UO_678 (O_678,N_9269,N_8008);
nor UO_679 (O_679,N_8172,N_8525);
nor UO_680 (O_680,N_8394,N_9223);
or UO_681 (O_681,N_8452,N_9473);
and UO_682 (O_682,N_9422,N_9245);
nor UO_683 (O_683,N_9098,N_8949);
xor UO_684 (O_684,N_8392,N_8834);
or UO_685 (O_685,N_8335,N_8176);
nor UO_686 (O_686,N_9875,N_9800);
xnor UO_687 (O_687,N_9455,N_8010);
or UO_688 (O_688,N_8258,N_8945);
nor UO_689 (O_689,N_8549,N_8208);
nand UO_690 (O_690,N_9469,N_9535);
nand UO_691 (O_691,N_8115,N_8456);
xnor UO_692 (O_692,N_9252,N_9205);
and UO_693 (O_693,N_8832,N_8129);
nand UO_694 (O_694,N_8110,N_8587);
and UO_695 (O_695,N_8076,N_8468);
and UO_696 (O_696,N_9459,N_9585);
nor UO_697 (O_697,N_9625,N_8478);
nand UO_698 (O_698,N_8522,N_8869);
nor UO_699 (O_699,N_8455,N_9785);
xor UO_700 (O_700,N_9943,N_9530);
xnor UO_701 (O_701,N_8847,N_9375);
and UO_702 (O_702,N_8951,N_8377);
nand UO_703 (O_703,N_8872,N_8204);
and UO_704 (O_704,N_8032,N_9185);
or UO_705 (O_705,N_8348,N_9172);
or UO_706 (O_706,N_9786,N_8770);
nand UO_707 (O_707,N_8489,N_8030);
xor UO_708 (O_708,N_9423,N_8966);
xnor UO_709 (O_709,N_8633,N_8500);
or UO_710 (O_710,N_9387,N_9416);
nor UO_711 (O_711,N_8934,N_8649);
xnor UO_712 (O_712,N_8270,N_9077);
and UO_713 (O_713,N_9441,N_8992);
xnor UO_714 (O_714,N_8125,N_8889);
xnor UO_715 (O_715,N_9273,N_8353);
xnor UO_716 (O_716,N_8714,N_9227);
or UO_717 (O_717,N_9830,N_8652);
nand UO_718 (O_718,N_8986,N_9219);
and UO_719 (O_719,N_9179,N_9523);
and UO_720 (O_720,N_8882,N_8803);
and UO_721 (O_721,N_9436,N_8836);
nor UO_722 (O_722,N_8028,N_9569);
xnor UO_723 (O_723,N_9361,N_8289);
xor UO_724 (O_724,N_8029,N_9840);
xnor UO_725 (O_725,N_8737,N_8390);
nor UO_726 (O_726,N_8905,N_8703);
nand UO_727 (O_727,N_8442,N_8969);
nand UO_728 (O_728,N_9289,N_9011);
nor UO_729 (O_729,N_8175,N_8668);
nand UO_730 (O_730,N_8388,N_8859);
or UO_731 (O_731,N_8205,N_8762);
and UO_732 (O_732,N_8663,N_9351);
nor UO_733 (O_733,N_9392,N_8750);
or UO_734 (O_734,N_8365,N_8612);
and UO_735 (O_735,N_9345,N_9355);
nor UO_736 (O_736,N_8077,N_8001);
nand UO_737 (O_737,N_9975,N_9796);
and UO_738 (O_738,N_8698,N_8024);
nand UO_739 (O_739,N_8755,N_9363);
nand UO_740 (O_740,N_9125,N_9866);
xnor UO_741 (O_741,N_8112,N_9171);
nand UO_742 (O_742,N_9618,N_8109);
xnor UO_743 (O_743,N_8757,N_9768);
nand UO_744 (O_744,N_8124,N_8059);
xnor UO_745 (O_745,N_9698,N_9428);
and UO_746 (O_746,N_9091,N_9552);
or UO_747 (O_747,N_8885,N_9663);
or UO_748 (O_748,N_9180,N_9408);
xor UO_749 (O_749,N_9394,N_9554);
and UO_750 (O_750,N_8433,N_9228);
and UO_751 (O_751,N_8898,N_8979);
or UO_752 (O_752,N_8715,N_8484);
nand UO_753 (O_753,N_8682,N_9368);
nand UO_754 (O_754,N_9495,N_9969);
and UO_755 (O_755,N_8091,N_8315);
or UO_756 (O_756,N_9685,N_9632);
and UO_757 (O_757,N_9399,N_9574);
and UO_758 (O_758,N_8179,N_8743);
xor UO_759 (O_759,N_9071,N_8505);
xor UO_760 (O_760,N_8894,N_8705);
nor UO_761 (O_761,N_8824,N_9591);
or UO_762 (O_762,N_8046,N_9143);
and UO_763 (O_763,N_9518,N_8382);
and UO_764 (O_764,N_8732,N_9674);
xnor UO_765 (O_765,N_8282,N_8841);
nand UO_766 (O_766,N_9914,N_8021);
nor UO_767 (O_767,N_8297,N_8286);
and UO_768 (O_768,N_9302,N_8696);
nor UO_769 (O_769,N_9879,N_8128);
xnor UO_770 (O_770,N_9073,N_9323);
xor UO_771 (O_771,N_9155,N_8912);
nand UO_772 (O_772,N_8586,N_8576);
nor UO_773 (O_773,N_8308,N_8570);
xor UO_774 (O_774,N_8854,N_8888);
or UO_775 (O_775,N_9538,N_8338);
xnor UO_776 (O_776,N_9842,N_9024);
nand UO_777 (O_777,N_8637,N_9712);
xor UO_778 (O_778,N_8146,N_8199);
and UO_779 (O_779,N_9174,N_9776);
nand UO_780 (O_780,N_9686,N_8472);
xor UO_781 (O_781,N_9348,N_9918);
or UO_782 (O_782,N_9802,N_8277);
and UO_783 (O_783,N_8773,N_8626);
or UO_784 (O_784,N_8561,N_8276);
nand UO_785 (O_785,N_9765,N_8669);
and UO_786 (O_786,N_9042,N_8380);
and UO_787 (O_787,N_9631,N_8349);
xor UO_788 (O_788,N_8421,N_8288);
xor UO_789 (O_789,N_9622,N_8368);
nor UO_790 (O_790,N_8181,N_8632);
and UO_791 (O_791,N_8419,N_9478);
nor UO_792 (O_792,N_8533,N_8447);
and UO_793 (O_793,N_9417,N_9373);
nand UO_794 (O_794,N_9380,N_9718);
nand UO_795 (O_795,N_8645,N_8704);
nand UO_796 (O_796,N_8154,N_8254);
xnor UO_797 (O_797,N_9432,N_9130);
nand UO_798 (O_798,N_8310,N_8551);
nor UO_799 (O_799,N_8424,N_8191);
and UO_800 (O_800,N_8981,N_9648);
or UO_801 (O_801,N_9405,N_8806);
nor UO_802 (O_802,N_9231,N_8783);
nand UO_803 (O_803,N_8346,N_8071);
xnor UO_804 (O_804,N_9062,N_8501);
and UO_805 (O_805,N_8689,N_8924);
nor UO_806 (O_806,N_9481,N_9545);
nor UO_807 (O_807,N_8488,N_9371);
and UO_808 (O_808,N_9542,N_9176);
or UO_809 (O_809,N_8917,N_9082);
nand UO_810 (O_810,N_8095,N_8396);
or UO_811 (O_811,N_8070,N_9318);
nand UO_812 (O_812,N_9192,N_9109);
and UO_813 (O_813,N_8828,N_9860);
and UO_814 (O_814,N_8881,N_8074);
and UO_815 (O_815,N_9601,N_8171);
nand UO_816 (O_816,N_8748,N_9809);
xor UO_817 (O_817,N_9937,N_9544);
nor UO_818 (O_818,N_9835,N_8699);
nand UO_819 (O_819,N_8855,N_9458);
nor UO_820 (O_820,N_9272,N_8014);
or UO_821 (O_821,N_9517,N_9978);
or UO_822 (O_822,N_9541,N_9292);
nor UO_823 (O_823,N_8089,N_8695);
nand UO_824 (O_824,N_8662,N_8727);
xnor UO_825 (O_825,N_9410,N_9870);
and UO_826 (O_826,N_8144,N_8142);
nand UO_827 (O_827,N_8332,N_8886);
nand UO_828 (O_828,N_8838,N_8664);
nor UO_829 (O_829,N_9565,N_9295);
nand UO_830 (O_830,N_9627,N_9817);
xnor UO_831 (O_831,N_9328,N_8425);
nand UO_832 (O_832,N_9804,N_9112);
xnor UO_833 (O_833,N_9872,N_9865);
or UO_834 (O_834,N_9878,N_9855);
xor UO_835 (O_835,N_8563,N_8363);
or UO_836 (O_836,N_9876,N_8326);
xor UO_837 (O_837,N_9546,N_9442);
and UO_838 (O_838,N_9053,N_9514);
or UO_839 (O_839,N_9305,N_8702);
nor UO_840 (O_840,N_8075,N_9734);
nand UO_841 (O_841,N_9214,N_9398);
nor UO_842 (O_842,N_9932,N_8048);
nand UO_843 (O_843,N_8017,N_8064);
nor UO_844 (O_844,N_8983,N_9232);
xor UO_845 (O_845,N_9959,N_9282);
nor UO_846 (O_846,N_8960,N_8052);
nor UO_847 (O_847,N_9374,N_9049);
nor UO_848 (O_848,N_8466,N_8604);
nor UO_849 (O_849,N_9483,N_8756);
nor UO_850 (O_850,N_8412,N_8552);
nor UO_851 (O_851,N_9322,N_9415);
xnor UO_852 (O_852,N_8220,N_8795);
and UO_853 (O_853,N_8465,N_8839);
nand UO_854 (O_854,N_9704,N_9612);
or UO_855 (O_855,N_8831,N_8218);
and UO_856 (O_856,N_9871,N_9651);
nand UO_857 (O_857,N_9737,N_9014);
or UO_858 (O_858,N_9862,N_9559);
or UO_859 (O_859,N_9035,N_8759);
and UO_860 (O_860,N_9331,N_9142);
nor UO_861 (O_861,N_8081,N_9640);
xor UO_862 (O_862,N_8374,N_9710);
nand UO_863 (O_863,N_8518,N_9139);
nand UO_864 (O_864,N_9548,N_9856);
or UO_865 (O_865,N_9206,N_8147);
nor UO_866 (O_866,N_8654,N_8318);
and UO_867 (O_867,N_9741,N_8170);
nor UO_868 (O_868,N_8247,N_9063);
nand UO_869 (O_869,N_8959,N_9039);
nand UO_870 (O_870,N_9274,N_9010);
nor UO_871 (O_871,N_9536,N_9204);
or UO_872 (O_872,N_9922,N_8212);
xnor UO_873 (O_873,N_8050,N_9330);
and UO_874 (O_874,N_8163,N_9437);
and UO_875 (O_875,N_8285,N_8805);
nor UO_876 (O_876,N_9412,N_9843);
nor UO_877 (O_877,N_8148,N_9159);
nand UO_878 (O_878,N_9359,N_8575);
xor UO_879 (O_879,N_8893,N_8462);
nand UO_880 (O_880,N_9004,N_9218);
nor UO_881 (O_881,N_8464,N_9709);
nand UO_882 (O_882,N_8711,N_9166);
or UO_883 (O_883,N_8559,N_8471);
nand UO_884 (O_884,N_9372,N_8004);
and UO_885 (O_885,N_8316,N_8340);
nand UO_886 (O_886,N_8661,N_9006);
and UO_887 (O_887,N_9122,N_9543);
and UO_888 (O_888,N_9985,N_9170);
nand UO_889 (O_889,N_8168,N_8034);
xor UO_890 (O_890,N_8776,N_9150);
and UO_891 (O_891,N_9877,N_8793);
xnor UO_892 (O_892,N_9474,N_8555);
nand UO_893 (O_893,N_9048,N_9421);
xnor UO_894 (O_894,N_8719,N_9009);
nand UO_895 (O_895,N_9027,N_8542);
and UO_896 (O_896,N_8908,N_8920);
and UO_897 (O_897,N_9949,N_9825);
nand UO_898 (O_898,N_9670,N_8660);
and UO_899 (O_899,N_9659,N_8671);
nor UO_900 (O_900,N_9431,N_9873);
and UO_901 (O_901,N_8529,N_9628);
nor UO_902 (O_902,N_8426,N_9869);
xor UO_903 (O_903,N_9888,N_9849);
nand UO_904 (O_904,N_8309,N_9973);
and UO_905 (O_905,N_9861,N_8730);
or UO_906 (O_906,N_9287,N_8099);
xnor UO_907 (O_907,N_9068,N_9026);
and UO_908 (O_908,N_9587,N_8135);
xor UO_909 (O_909,N_8928,N_8138);
nor UO_910 (O_910,N_9771,N_8936);
nand UO_911 (O_911,N_8647,N_9582);
xnor UO_912 (O_912,N_9611,N_9512);
nand UO_913 (O_913,N_9426,N_8463);
xor UO_914 (O_914,N_9389,N_8221);
nand UO_915 (O_915,N_9427,N_8537);
xor UO_916 (O_916,N_8921,N_8906);
and UO_917 (O_917,N_9551,N_9356);
nor UO_918 (O_918,N_8196,N_9153);
and UO_919 (O_919,N_9900,N_9095);
nor UO_920 (O_920,N_8531,N_9700);
nand UO_921 (O_921,N_8851,N_9971);
xor UO_922 (O_922,N_8130,N_8370);
and UO_923 (O_923,N_9775,N_9472);
and UO_924 (O_924,N_8588,N_9054);
nor UO_925 (O_925,N_9907,N_8198);
and UO_926 (O_926,N_9243,N_9903);
nand UO_927 (O_927,N_9237,N_9366);
xor UO_928 (O_928,N_9689,N_8903);
nor UO_929 (O_929,N_9654,N_8602);
and UO_930 (O_930,N_9242,N_8915);
and UO_931 (O_931,N_9433,N_9403);
xnor UO_932 (O_932,N_9152,N_8672);
or UO_933 (O_933,N_9679,N_8804);
xnor UO_934 (O_934,N_8781,N_8939);
xor UO_935 (O_935,N_9438,N_8358);
or UO_936 (O_936,N_9708,N_8051);
nand UO_937 (O_937,N_8639,N_8007);
nor UO_938 (O_938,N_9397,N_9140);
nor UO_939 (O_939,N_8784,N_8530);
or UO_940 (O_940,N_9773,N_9893);
xnor UO_941 (O_941,N_9045,N_8262);
nor UO_942 (O_942,N_9579,N_9946);
xnor UO_943 (O_943,N_8025,N_8827);
nand UO_944 (O_944,N_9650,N_8449);
or UO_945 (O_945,N_8740,N_8595);
or UO_946 (O_946,N_9044,N_9256);
or UO_947 (O_947,N_9346,N_8458);
nor UO_948 (O_948,N_8197,N_8241);
or UO_949 (O_949,N_9740,N_8213);
nand UO_950 (O_950,N_8451,N_8909);
or UO_951 (O_951,N_8344,N_9658);
and UO_952 (O_952,N_9386,N_9084);
nor UO_953 (O_953,N_8507,N_8974);
or UO_954 (O_954,N_8410,N_9610);
or UO_955 (O_955,N_8799,N_8190);
or UO_956 (O_956,N_8515,N_8543);
xnor UO_957 (O_957,N_8474,N_8517);
and UO_958 (O_958,N_9298,N_8853);
xor UO_959 (O_959,N_8281,N_8873);
xor UO_960 (O_960,N_9634,N_9556);
xor UO_961 (O_961,N_8540,N_9887);
nand UO_962 (O_962,N_8031,N_8411);
nor UO_963 (O_963,N_9028,N_8379);
or UO_964 (O_964,N_8215,N_8490);
nor UO_965 (O_965,N_8040,N_8137);
and UO_966 (O_966,N_9203,N_9311);
or UO_967 (O_967,N_8323,N_9076);
nor UO_968 (O_968,N_8998,N_8210);
and UO_969 (O_969,N_9772,N_8728);
xor UO_970 (O_970,N_9136,N_8151);
and UO_971 (O_971,N_8845,N_9007);
nand UO_972 (O_972,N_9107,N_8184);
or UO_973 (O_973,N_9396,N_9892);
or UO_974 (O_974,N_9278,N_8777);
and UO_975 (O_975,N_8319,N_8852);
xnor UO_976 (O_976,N_8079,N_9193);
nor UO_977 (O_977,N_9445,N_9633);
nor UO_978 (O_978,N_8722,N_8347);
and UO_979 (O_979,N_9636,N_8548);
nand UO_980 (O_980,N_9047,N_8328);
nor UO_981 (O_981,N_9732,N_9630);
nor UO_982 (O_982,N_8339,N_8321);
xnor UO_983 (O_983,N_8188,N_8935);
and UO_984 (O_984,N_9162,N_9697);
nor UO_985 (O_985,N_8027,N_9200);
xnor UO_986 (O_986,N_8093,N_9844);
xor UO_987 (O_987,N_9462,N_9528);
or UO_988 (O_988,N_9158,N_9646);
nand UO_989 (O_989,N_9539,N_8195);
nor UO_990 (O_990,N_8416,N_8343);
and UO_991 (O_991,N_9984,N_9555);
and UO_992 (O_992,N_8156,N_9639);
or UO_993 (O_993,N_9369,N_9820);
or UO_994 (O_994,N_9986,N_9520);
and UO_995 (O_995,N_9114,N_9808);
nor UO_996 (O_996,N_9220,N_8225);
or UO_997 (O_997,N_8055,N_9595);
or UO_998 (O_998,N_8584,N_8538);
nor UO_999 (O_999,N_8062,N_8302);
xnor UO_1000 (O_1000,N_8100,N_8497);
and UO_1001 (O_1001,N_8214,N_9923);
xnor UO_1002 (O_1002,N_8004,N_8218);
xnor UO_1003 (O_1003,N_9478,N_8694);
and UO_1004 (O_1004,N_8923,N_8383);
xnor UO_1005 (O_1005,N_8772,N_9699);
and UO_1006 (O_1006,N_8030,N_9900);
or UO_1007 (O_1007,N_8958,N_8259);
nand UO_1008 (O_1008,N_9524,N_8058);
and UO_1009 (O_1009,N_8186,N_9209);
or UO_1010 (O_1010,N_9048,N_8980);
nor UO_1011 (O_1011,N_9978,N_9033);
nand UO_1012 (O_1012,N_8010,N_8074);
nand UO_1013 (O_1013,N_9542,N_9053);
and UO_1014 (O_1014,N_9085,N_8938);
and UO_1015 (O_1015,N_8844,N_9256);
nand UO_1016 (O_1016,N_8229,N_9842);
and UO_1017 (O_1017,N_9354,N_9727);
nand UO_1018 (O_1018,N_8197,N_9216);
and UO_1019 (O_1019,N_8440,N_9020);
or UO_1020 (O_1020,N_9393,N_8464);
nor UO_1021 (O_1021,N_9563,N_8996);
and UO_1022 (O_1022,N_9447,N_8304);
nand UO_1023 (O_1023,N_8569,N_8345);
or UO_1024 (O_1024,N_8038,N_8247);
xor UO_1025 (O_1025,N_8863,N_8285);
xor UO_1026 (O_1026,N_9117,N_9752);
or UO_1027 (O_1027,N_9929,N_9689);
xor UO_1028 (O_1028,N_9781,N_9082);
xor UO_1029 (O_1029,N_9419,N_8192);
or UO_1030 (O_1030,N_8799,N_8061);
nor UO_1031 (O_1031,N_8405,N_9391);
nand UO_1032 (O_1032,N_9146,N_9962);
and UO_1033 (O_1033,N_9624,N_9783);
xnor UO_1034 (O_1034,N_8030,N_8802);
nor UO_1035 (O_1035,N_8147,N_8579);
xnor UO_1036 (O_1036,N_9964,N_8537);
or UO_1037 (O_1037,N_9548,N_8364);
and UO_1038 (O_1038,N_8791,N_8686);
nand UO_1039 (O_1039,N_9581,N_8845);
nand UO_1040 (O_1040,N_8321,N_8847);
and UO_1041 (O_1041,N_9759,N_9646);
nor UO_1042 (O_1042,N_9902,N_9798);
xor UO_1043 (O_1043,N_9623,N_8731);
nand UO_1044 (O_1044,N_8367,N_9486);
and UO_1045 (O_1045,N_9313,N_9281);
xor UO_1046 (O_1046,N_9497,N_8725);
and UO_1047 (O_1047,N_8705,N_8754);
and UO_1048 (O_1048,N_8509,N_8311);
and UO_1049 (O_1049,N_9571,N_8067);
nor UO_1050 (O_1050,N_8416,N_9817);
nor UO_1051 (O_1051,N_9782,N_8876);
and UO_1052 (O_1052,N_8398,N_9983);
xnor UO_1053 (O_1053,N_8982,N_9404);
nand UO_1054 (O_1054,N_9345,N_8810);
xor UO_1055 (O_1055,N_9337,N_9102);
nand UO_1056 (O_1056,N_8746,N_8797);
or UO_1057 (O_1057,N_8159,N_8321);
nor UO_1058 (O_1058,N_9644,N_8248);
nand UO_1059 (O_1059,N_9201,N_9919);
or UO_1060 (O_1060,N_9082,N_9763);
nand UO_1061 (O_1061,N_9653,N_9704);
or UO_1062 (O_1062,N_9738,N_9278);
nor UO_1063 (O_1063,N_9641,N_9813);
xnor UO_1064 (O_1064,N_8236,N_8634);
nor UO_1065 (O_1065,N_8342,N_9050);
nor UO_1066 (O_1066,N_9887,N_8008);
or UO_1067 (O_1067,N_8491,N_8763);
xor UO_1068 (O_1068,N_9621,N_8867);
nor UO_1069 (O_1069,N_8072,N_8910);
nor UO_1070 (O_1070,N_9883,N_9431);
nand UO_1071 (O_1071,N_9141,N_8347);
and UO_1072 (O_1072,N_9433,N_9219);
or UO_1073 (O_1073,N_9745,N_9135);
xnor UO_1074 (O_1074,N_9608,N_8405);
nand UO_1075 (O_1075,N_9772,N_9351);
nor UO_1076 (O_1076,N_8426,N_8779);
nor UO_1077 (O_1077,N_9298,N_8153);
nor UO_1078 (O_1078,N_9685,N_8404);
and UO_1079 (O_1079,N_9393,N_8739);
xor UO_1080 (O_1080,N_8288,N_8946);
or UO_1081 (O_1081,N_8283,N_8224);
xnor UO_1082 (O_1082,N_8390,N_8001);
or UO_1083 (O_1083,N_8262,N_8274);
or UO_1084 (O_1084,N_9595,N_9580);
or UO_1085 (O_1085,N_8454,N_8752);
or UO_1086 (O_1086,N_9965,N_9575);
or UO_1087 (O_1087,N_8803,N_9995);
and UO_1088 (O_1088,N_9956,N_8384);
and UO_1089 (O_1089,N_9702,N_9820);
nand UO_1090 (O_1090,N_8872,N_9838);
nand UO_1091 (O_1091,N_9176,N_8759);
and UO_1092 (O_1092,N_9307,N_9655);
and UO_1093 (O_1093,N_8622,N_8374);
or UO_1094 (O_1094,N_8559,N_9618);
nand UO_1095 (O_1095,N_9546,N_8282);
nor UO_1096 (O_1096,N_9900,N_9595);
and UO_1097 (O_1097,N_8460,N_8857);
or UO_1098 (O_1098,N_8741,N_9539);
nor UO_1099 (O_1099,N_8032,N_9454);
nand UO_1100 (O_1100,N_9971,N_8444);
and UO_1101 (O_1101,N_9879,N_9551);
nand UO_1102 (O_1102,N_9168,N_9408);
and UO_1103 (O_1103,N_9816,N_9318);
nor UO_1104 (O_1104,N_8312,N_8472);
or UO_1105 (O_1105,N_9796,N_8642);
and UO_1106 (O_1106,N_9295,N_9815);
and UO_1107 (O_1107,N_8723,N_9575);
xnor UO_1108 (O_1108,N_8351,N_8679);
and UO_1109 (O_1109,N_9406,N_8173);
nor UO_1110 (O_1110,N_8985,N_9355);
nand UO_1111 (O_1111,N_9942,N_9661);
or UO_1112 (O_1112,N_9590,N_9115);
nand UO_1113 (O_1113,N_9464,N_8618);
or UO_1114 (O_1114,N_9363,N_8467);
and UO_1115 (O_1115,N_8416,N_9116);
and UO_1116 (O_1116,N_9313,N_9711);
nor UO_1117 (O_1117,N_8915,N_9139);
nand UO_1118 (O_1118,N_9167,N_9516);
and UO_1119 (O_1119,N_8319,N_9046);
xor UO_1120 (O_1120,N_8937,N_8962);
nor UO_1121 (O_1121,N_9525,N_8795);
nor UO_1122 (O_1122,N_9519,N_8458);
nor UO_1123 (O_1123,N_9762,N_8443);
and UO_1124 (O_1124,N_9657,N_9261);
xnor UO_1125 (O_1125,N_8358,N_9767);
xnor UO_1126 (O_1126,N_8502,N_8699);
nand UO_1127 (O_1127,N_9009,N_8390);
and UO_1128 (O_1128,N_8547,N_9285);
and UO_1129 (O_1129,N_9960,N_9117);
nor UO_1130 (O_1130,N_8101,N_9343);
xnor UO_1131 (O_1131,N_9425,N_9309);
and UO_1132 (O_1132,N_9415,N_8047);
and UO_1133 (O_1133,N_9074,N_9427);
xnor UO_1134 (O_1134,N_9832,N_8121);
and UO_1135 (O_1135,N_8187,N_9077);
xnor UO_1136 (O_1136,N_9563,N_9606);
nor UO_1137 (O_1137,N_8865,N_8772);
xor UO_1138 (O_1138,N_8441,N_9818);
nand UO_1139 (O_1139,N_9468,N_9373);
nor UO_1140 (O_1140,N_8848,N_8320);
and UO_1141 (O_1141,N_8407,N_9793);
or UO_1142 (O_1142,N_9362,N_9352);
and UO_1143 (O_1143,N_8352,N_8414);
or UO_1144 (O_1144,N_8739,N_9360);
and UO_1145 (O_1145,N_8541,N_8002);
or UO_1146 (O_1146,N_9302,N_9901);
nor UO_1147 (O_1147,N_9857,N_9690);
or UO_1148 (O_1148,N_8988,N_8363);
and UO_1149 (O_1149,N_9384,N_9893);
or UO_1150 (O_1150,N_8601,N_9827);
nor UO_1151 (O_1151,N_8400,N_9570);
and UO_1152 (O_1152,N_8329,N_9640);
or UO_1153 (O_1153,N_9561,N_8893);
nand UO_1154 (O_1154,N_8933,N_9817);
or UO_1155 (O_1155,N_8247,N_9270);
and UO_1156 (O_1156,N_9609,N_9728);
xnor UO_1157 (O_1157,N_9930,N_8696);
xor UO_1158 (O_1158,N_9779,N_8426);
or UO_1159 (O_1159,N_9150,N_9110);
xnor UO_1160 (O_1160,N_8574,N_9120);
or UO_1161 (O_1161,N_8512,N_8841);
xnor UO_1162 (O_1162,N_9536,N_8815);
xnor UO_1163 (O_1163,N_9503,N_8271);
xnor UO_1164 (O_1164,N_9150,N_9642);
and UO_1165 (O_1165,N_8364,N_8397);
xnor UO_1166 (O_1166,N_8462,N_8501);
xor UO_1167 (O_1167,N_8581,N_9306);
xnor UO_1168 (O_1168,N_9430,N_8995);
xnor UO_1169 (O_1169,N_8257,N_8757);
xor UO_1170 (O_1170,N_9148,N_8048);
and UO_1171 (O_1171,N_9821,N_9786);
or UO_1172 (O_1172,N_8926,N_9777);
nor UO_1173 (O_1173,N_8664,N_8763);
or UO_1174 (O_1174,N_9323,N_9642);
nand UO_1175 (O_1175,N_8394,N_8854);
xnor UO_1176 (O_1176,N_9611,N_8529);
nand UO_1177 (O_1177,N_9560,N_9196);
and UO_1178 (O_1178,N_9914,N_8145);
nand UO_1179 (O_1179,N_8580,N_9397);
or UO_1180 (O_1180,N_9571,N_8410);
or UO_1181 (O_1181,N_9859,N_8080);
xnor UO_1182 (O_1182,N_9988,N_8273);
nand UO_1183 (O_1183,N_8858,N_9788);
nor UO_1184 (O_1184,N_9073,N_8248);
nand UO_1185 (O_1185,N_8997,N_9909);
or UO_1186 (O_1186,N_9387,N_9501);
nor UO_1187 (O_1187,N_8061,N_8856);
nand UO_1188 (O_1188,N_8944,N_8264);
or UO_1189 (O_1189,N_8361,N_8895);
nand UO_1190 (O_1190,N_8557,N_8652);
or UO_1191 (O_1191,N_9412,N_9929);
or UO_1192 (O_1192,N_9193,N_8554);
or UO_1193 (O_1193,N_8107,N_9403);
nand UO_1194 (O_1194,N_9578,N_9717);
xor UO_1195 (O_1195,N_8881,N_8644);
nand UO_1196 (O_1196,N_8063,N_8179);
nand UO_1197 (O_1197,N_8726,N_9595);
xor UO_1198 (O_1198,N_8813,N_9943);
nor UO_1199 (O_1199,N_9635,N_8087);
or UO_1200 (O_1200,N_8727,N_8217);
and UO_1201 (O_1201,N_8857,N_9440);
and UO_1202 (O_1202,N_9736,N_8051);
nand UO_1203 (O_1203,N_8933,N_8193);
and UO_1204 (O_1204,N_8394,N_8346);
and UO_1205 (O_1205,N_8317,N_8102);
xor UO_1206 (O_1206,N_8654,N_8700);
or UO_1207 (O_1207,N_8239,N_8760);
or UO_1208 (O_1208,N_9871,N_9914);
and UO_1209 (O_1209,N_9089,N_9336);
and UO_1210 (O_1210,N_8493,N_9084);
and UO_1211 (O_1211,N_8413,N_9672);
or UO_1212 (O_1212,N_8096,N_8139);
or UO_1213 (O_1213,N_9487,N_9310);
and UO_1214 (O_1214,N_9946,N_8463);
xnor UO_1215 (O_1215,N_8735,N_8532);
and UO_1216 (O_1216,N_9551,N_9905);
nor UO_1217 (O_1217,N_9452,N_8796);
nand UO_1218 (O_1218,N_9081,N_8198);
xor UO_1219 (O_1219,N_9746,N_8971);
nand UO_1220 (O_1220,N_9722,N_9123);
nand UO_1221 (O_1221,N_8018,N_8587);
xnor UO_1222 (O_1222,N_9335,N_9219);
or UO_1223 (O_1223,N_9369,N_8087);
xor UO_1224 (O_1224,N_9212,N_9596);
and UO_1225 (O_1225,N_9056,N_8953);
nand UO_1226 (O_1226,N_8771,N_8986);
and UO_1227 (O_1227,N_8305,N_8454);
xnor UO_1228 (O_1228,N_9507,N_8731);
and UO_1229 (O_1229,N_8407,N_8182);
nor UO_1230 (O_1230,N_9338,N_9012);
and UO_1231 (O_1231,N_8701,N_8532);
nor UO_1232 (O_1232,N_9368,N_8948);
and UO_1233 (O_1233,N_8028,N_9605);
nor UO_1234 (O_1234,N_9952,N_8442);
xnor UO_1235 (O_1235,N_8632,N_8397);
and UO_1236 (O_1236,N_8667,N_8212);
or UO_1237 (O_1237,N_8755,N_8141);
or UO_1238 (O_1238,N_9279,N_8821);
or UO_1239 (O_1239,N_8511,N_9434);
and UO_1240 (O_1240,N_8178,N_9957);
nand UO_1241 (O_1241,N_9887,N_9862);
and UO_1242 (O_1242,N_9452,N_8110);
nor UO_1243 (O_1243,N_8952,N_9850);
xnor UO_1244 (O_1244,N_9521,N_9769);
or UO_1245 (O_1245,N_8161,N_8816);
or UO_1246 (O_1246,N_8199,N_8392);
xor UO_1247 (O_1247,N_9685,N_8837);
and UO_1248 (O_1248,N_9363,N_8350);
xor UO_1249 (O_1249,N_8695,N_9494);
nand UO_1250 (O_1250,N_8085,N_8331);
or UO_1251 (O_1251,N_8217,N_8791);
nand UO_1252 (O_1252,N_9162,N_9965);
or UO_1253 (O_1253,N_8817,N_9043);
nand UO_1254 (O_1254,N_9912,N_8540);
or UO_1255 (O_1255,N_9780,N_9839);
nor UO_1256 (O_1256,N_9444,N_8384);
xnor UO_1257 (O_1257,N_8559,N_9371);
and UO_1258 (O_1258,N_9358,N_9077);
and UO_1259 (O_1259,N_8973,N_9961);
and UO_1260 (O_1260,N_8102,N_8959);
xnor UO_1261 (O_1261,N_8270,N_9868);
nand UO_1262 (O_1262,N_8665,N_8033);
xnor UO_1263 (O_1263,N_8107,N_9454);
and UO_1264 (O_1264,N_8385,N_8233);
nand UO_1265 (O_1265,N_8956,N_8052);
nand UO_1266 (O_1266,N_9470,N_9039);
or UO_1267 (O_1267,N_9274,N_8809);
nor UO_1268 (O_1268,N_9303,N_9962);
and UO_1269 (O_1269,N_8231,N_9991);
nand UO_1270 (O_1270,N_9712,N_9150);
xor UO_1271 (O_1271,N_8544,N_8270);
nand UO_1272 (O_1272,N_9106,N_8971);
xnor UO_1273 (O_1273,N_8015,N_9008);
nand UO_1274 (O_1274,N_8815,N_9147);
or UO_1275 (O_1275,N_9338,N_9358);
nor UO_1276 (O_1276,N_8815,N_9526);
xor UO_1277 (O_1277,N_8788,N_9687);
and UO_1278 (O_1278,N_8762,N_8459);
or UO_1279 (O_1279,N_8998,N_8253);
and UO_1280 (O_1280,N_8557,N_8899);
nand UO_1281 (O_1281,N_9063,N_9885);
nand UO_1282 (O_1282,N_9157,N_8205);
or UO_1283 (O_1283,N_8055,N_9234);
nor UO_1284 (O_1284,N_8494,N_9968);
and UO_1285 (O_1285,N_8157,N_9680);
or UO_1286 (O_1286,N_8027,N_8829);
nand UO_1287 (O_1287,N_9485,N_8332);
or UO_1288 (O_1288,N_8758,N_9662);
nand UO_1289 (O_1289,N_8238,N_8413);
nand UO_1290 (O_1290,N_8479,N_8593);
nor UO_1291 (O_1291,N_8788,N_8298);
nor UO_1292 (O_1292,N_9419,N_9958);
xnor UO_1293 (O_1293,N_9423,N_8725);
and UO_1294 (O_1294,N_9935,N_8487);
nand UO_1295 (O_1295,N_8046,N_9921);
and UO_1296 (O_1296,N_8837,N_9055);
nor UO_1297 (O_1297,N_8508,N_9165);
or UO_1298 (O_1298,N_8760,N_8874);
xnor UO_1299 (O_1299,N_9182,N_8427);
or UO_1300 (O_1300,N_9195,N_8941);
nand UO_1301 (O_1301,N_9102,N_8132);
nor UO_1302 (O_1302,N_9272,N_8621);
nor UO_1303 (O_1303,N_9424,N_9683);
nand UO_1304 (O_1304,N_9034,N_9556);
or UO_1305 (O_1305,N_9772,N_9555);
or UO_1306 (O_1306,N_8555,N_8684);
xnor UO_1307 (O_1307,N_8382,N_8169);
or UO_1308 (O_1308,N_9607,N_9956);
nand UO_1309 (O_1309,N_9042,N_9374);
and UO_1310 (O_1310,N_8554,N_8079);
nand UO_1311 (O_1311,N_9925,N_9893);
or UO_1312 (O_1312,N_8034,N_8223);
nand UO_1313 (O_1313,N_8712,N_9629);
and UO_1314 (O_1314,N_9214,N_9697);
and UO_1315 (O_1315,N_8199,N_8295);
nand UO_1316 (O_1316,N_9485,N_8488);
xor UO_1317 (O_1317,N_9643,N_8459);
nor UO_1318 (O_1318,N_9112,N_9557);
or UO_1319 (O_1319,N_8282,N_8368);
nand UO_1320 (O_1320,N_9305,N_9229);
and UO_1321 (O_1321,N_9593,N_8822);
nor UO_1322 (O_1322,N_9761,N_9682);
and UO_1323 (O_1323,N_9563,N_9131);
nand UO_1324 (O_1324,N_9858,N_8712);
and UO_1325 (O_1325,N_8052,N_9891);
xor UO_1326 (O_1326,N_8806,N_8721);
or UO_1327 (O_1327,N_9924,N_8816);
or UO_1328 (O_1328,N_8563,N_8808);
or UO_1329 (O_1329,N_8188,N_9065);
nand UO_1330 (O_1330,N_9442,N_9259);
and UO_1331 (O_1331,N_9601,N_9746);
and UO_1332 (O_1332,N_8425,N_8484);
xnor UO_1333 (O_1333,N_8263,N_8076);
or UO_1334 (O_1334,N_9384,N_8493);
xor UO_1335 (O_1335,N_9658,N_9392);
or UO_1336 (O_1336,N_8406,N_9711);
or UO_1337 (O_1337,N_8662,N_9064);
nand UO_1338 (O_1338,N_9726,N_9312);
and UO_1339 (O_1339,N_8135,N_9484);
nand UO_1340 (O_1340,N_9769,N_9850);
xor UO_1341 (O_1341,N_8659,N_8952);
nor UO_1342 (O_1342,N_8735,N_9171);
and UO_1343 (O_1343,N_8154,N_8060);
nor UO_1344 (O_1344,N_9345,N_8655);
or UO_1345 (O_1345,N_9691,N_8691);
xor UO_1346 (O_1346,N_8547,N_8160);
xnor UO_1347 (O_1347,N_8852,N_9304);
xor UO_1348 (O_1348,N_9379,N_9413);
nand UO_1349 (O_1349,N_8569,N_9298);
xor UO_1350 (O_1350,N_9420,N_9934);
nand UO_1351 (O_1351,N_9350,N_9000);
nand UO_1352 (O_1352,N_8216,N_9547);
and UO_1353 (O_1353,N_8860,N_8197);
nor UO_1354 (O_1354,N_8756,N_8996);
and UO_1355 (O_1355,N_8941,N_9474);
or UO_1356 (O_1356,N_9638,N_8997);
nor UO_1357 (O_1357,N_9647,N_9962);
nor UO_1358 (O_1358,N_9151,N_9173);
and UO_1359 (O_1359,N_9990,N_9912);
nand UO_1360 (O_1360,N_8457,N_8565);
nor UO_1361 (O_1361,N_9985,N_9322);
and UO_1362 (O_1362,N_9695,N_9746);
nand UO_1363 (O_1363,N_8065,N_8658);
nand UO_1364 (O_1364,N_9105,N_8116);
and UO_1365 (O_1365,N_9349,N_8432);
nand UO_1366 (O_1366,N_8555,N_9656);
or UO_1367 (O_1367,N_9109,N_8714);
nor UO_1368 (O_1368,N_9812,N_8865);
nand UO_1369 (O_1369,N_9132,N_8911);
nand UO_1370 (O_1370,N_8697,N_9195);
and UO_1371 (O_1371,N_8160,N_9914);
xor UO_1372 (O_1372,N_8261,N_9411);
nand UO_1373 (O_1373,N_8781,N_8749);
and UO_1374 (O_1374,N_8660,N_9074);
nand UO_1375 (O_1375,N_9316,N_9326);
or UO_1376 (O_1376,N_8307,N_8775);
and UO_1377 (O_1377,N_9356,N_9373);
and UO_1378 (O_1378,N_9136,N_8691);
nand UO_1379 (O_1379,N_9726,N_9816);
nor UO_1380 (O_1380,N_8784,N_8691);
nor UO_1381 (O_1381,N_9133,N_8443);
nor UO_1382 (O_1382,N_8762,N_9626);
or UO_1383 (O_1383,N_8778,N_8112);
nor UO_1384 (O_1384,N_9755,N_8136);
nor UO_1385 (O_1385,N_8787,N_9854);
nor UO_1386 (O_1386,N_9920,N_9853);
xor UO_1387 (O_1387,N_9118,N_8957);
or UO_1388 (O_1388,N_8708,N_8338);
or UO_1389 (O_1389,N_8910,N_8488);
or UO_1390 (O_1390,N_9553,N_9896);
nand UO_1391 (O_1391,N_8135,N_8429);
nor UO_1392 (O_1392,N_8534,N_9323);
or UO_1393 (O_1393,N_9044,N_9950);
nand UO_1394 (O_1394,N_8791,N_8609);
xnor UO_1395 (O_1395,N_8812,N_9480);
or UO_1396 (O_1396,N_9807,N_9383);
nor UO_1397 (O_1397,N_8228,N_8634);
and UO_1398 (O_1398,N_9850,N_8656);
nor UO_1399 (O_1399,N_9465,N_8262);
xnor UO_1400 (O_1400,N_9161,N_9865);
xor UO_1401 (O_1401,N_8315,N_9687);
nor UO_1402 (O_1402,N_9848,N_8676);
xor UO_1403 (O_1403,N_9234,N_9901);
and UO_1404 (O_1404,N_8736,N_8575);
xnor UO_1405 (O_1405,N_8568,N_9694);
and UO_1406 (O_1406,N_9802,N_8946);
nor UO_1407 (O_1407,N_8677,N_9615);
xnor UO_1408 (O_1408,N_9451,N_8864);
nand UO_1409 (O_1409,N_8034,N_8326);
nand UO_1410 (O_1410,N_9307,N_8258);
xor UO_1411 (O_1411,N_8422,N_9296);
nand UO_1412 (O_1412,N_8619,N_8665);
nor UO_1413 (O_1413,N_8204,N_8405);
or UO_1414 (O_1414,N_9188,N_8808);
xor UO_1415 (O_1415,N_9970,N_9675);
nand UO_1416 (O_1416,N_9568,N_9048);
nand UO_1417 (O_1417,N_8235,N_8374);
xnor UO_1418 (O_1418,N_8730,N_9036);
and UO_1419 (O_1419,N_9626,N_8767);
and UO_1420 (O_1420,N_8971,N_8768);
or UO_1421 (O_1421,N_9043,N_8649);
xor UO_1422 (O_1422,N_9338,N_8793);
or UO_1423 (O_1423,N_9704,N_9938);
or UO_1424 (O_1424,N_8886,N_8781);
or UO_1425 (O_1425,N_9573,N_9029);
and UO_1426 (O_1426,N_8489,N_8574);
and UO_1427 (O_1427,N_8281,N_9919);
nand UO_1428 (O_1428,N_8301,N_9071);
xor UO_1429 (O_1429,N_9440,N_8964);
or UO_1430 (O_1430,N_9043,N_8687);
or UO_1431 (O_1431,N_9407,N_9261);
xor UO_1432 (O_1432,N_9855,N_9620);
nand UO_1433 (O_1433,N_9692,N_8652);
xnor UO_1434 (O_1434,N_9958,N_9464);
nor UO_1435 (O_1435,N_8526,N_8542);
nor UO_1436 (O_1436,N_9458,N_9220);
xor UO_1437 (O_1437,N_8008,N_9688);
or UO_1438 (O_1438,N_8872,N_9816);
or UO_1439 (O_1439,N_9752,N_8589);
and UO_1440 (O_1440,N_9303,N_9797);
nor UO_1441 (O_1441,N_8688,N_9833);
nor UO_1442 (O_1442,N_8558,N_9644);
nor UO_1443 (O_1443,N_8094,N_9606);
or UO_1444 (O_1444,N_9328,N_8124);
nand UO_1445 (O_1445,N_9332,N_8319);
xnor UO_1446 (O_1446,N_9484,N_9997);
and UO_1447 (O_1447,N_9478,N_8159);
nor UO_1448 (O_1448,N_8548,N_8504);
and UO_1449 (O_1449,N_8232,N_8723);
nand UO_1450 (O_1450,N_9211,N_8756);
or UO_1451 (O_1451,N_8677,N_9582);
or UO_1452 (O_1452,N_8485,N_8134);
nand UO_1453 (O_1453,N_9751,N_9612);
nor UO_1454 (O_1454,N_9178,N_9276);
xor UO_1455 (O_1455,N_8114,N_9050);
xor UO_1456 (O_1456,N_9256,N_9784);
nand UO_1457 (O_1457,N_9618,N_9627);
nor UO_1458 (O_1458,N_8119,N_8334);
nand UO_1459 (O_1459,N_9964,N_8028);
or UO_1460 (O_1460,N_9679,N_9121);
and UO_1461 (O_1461,N_9771,N_9815);
and UO_1462 (O_1462,N_8804,N_8612);
nor UO_1463 (O_1463,N_9298,N_9345);
nand UO_1464 (O_1464,N_8324,N_8687);
or UO_1465 (O_1465,N_9317,N_8556);
xnor UO_1466 (O_1466,N_8757,N_9804);
nor UO_1467 (O_1467,N_9798,N_9506);
nand UO_1468 (O_1468,N_8683,N_9509);
nand UO_1469 (O_1469,N_8302,N_8536);
xor UO_1470 (O_1470,N_9299,N_9226);
nand UO_1471 (O_1471,N_8938,N_9924);
xor UO_1472 (O_1472,N_9834,N_9733);
xnor UO_1473 (O_1473,N_9703,N_8414);
xnor UO_1474 (O_1474,N_9525,N_9010);
xnor UO_1475 (O_1475,N_9941,N_9550);
xor UO_1476 (O_1476,N_9073,N_8007);
and UO_1477 (O_1477,N_9922,N_8224);
xor UO_1478 (O_1478,N_8792,N_9485);
or UO_1479 (O_1479,N_9612,N_8985);
nor UO_1480 (O_1480,N_8500,N_8845);
nor UO_1481 (O_1481,N_9339,N_9101);
nor UO_1482 (O_1482,N_8814,N_9012);
and UO_1483 (O_1483,N_9984,N_9998);
nor UO_1484 (O_1484,N_8433,N_9955);
or UO_1485 (O_1485,N_9800,N_9652);
nand UO_1486 (O_1486,N_9072,N_9296);
nor UO_1487 (O_1487,N_9693,N_9999);
and UO_1488 (O_1488,N_9978,N_8164);
nand UO_1489 (O_1489,N_9794,N_9722);
nor UO_1490 (O_1490,N_9071,N_9575);
or UO_1491 (O_1491,N_9533,N_9252);
nor UO_1492 (O_1492,N_9083,N_9289);
nand UO_1493 (O_1493,N_8737,N_9784);
and UO_1494 (O_1494,N_8779,N_8657);
nor UO_1495 (O_1495,N_8897,N_9603);
nor UO_1496 (O_1496,N_9460,N_9022);
xnor UO_1497 (O_1497,N_8342,N_9622);
nand UO_1498 (O_1498,N_8505,N_8904);
or UO_1499 (O_1499,N_8932,N_9962);
endmodule