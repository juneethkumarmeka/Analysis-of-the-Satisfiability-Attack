module basic_2000_20000_2500_125_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xor U0 (N_0,In_38,In_1842);
nor U1 (N_1,In_573,In_1140);
nand U2 (N_2,In_1633,In_1394);
xnor U3 (N_3,In_1660,In_170);
and U4 (N_4,In_293,In_1426);
or U5 (N_5,In_1212,In_425);
nand U6 (N_6,In_1762,In_897);
xor U7 (N_7,In_1466,In_511);
nand U8 (N_8,In_212,In_1843);
or U9 (N_9,In_201,In_297);
xor U10 (N_10,In_801,In_1854);
or U11 (N_11,In_888,In_448);
nor U12 (N_12,In_386,In_1853);
or U13 (N_13,In_1628,In_1113);
and U14 (N_14,In_1339,In_1338);
nor U15 (N_15,In_110,In_413);
nor U16 (N_16,In_1138,In_662);
nor U17 (N_17,In_1003,In_850);
nand U18 (N_18,In_1320,In_1952);
nand U19 (N_19,In_1543,In_751);
xnor U20 (N_20,In_762,In_1174);
or U21 (N_21,In_924,In_1624);
and U22 (N_22,In_1258,In_518);
and U23 (N_23,In_1354,In_1719);
or U24 (N_24,In_1645,In_1746);
xnor U25 (N_25,In_47,In_1159);
nand U26 (N_26,In_161,In_1246);
nor U27 (N_27,In_97,In_177);
nand U28 (N_28,In_280,In_527);
or U29 (N_29,In_1502,In_257);
xor U30 (N_30,In_183,In_1401);
nor U31 (N_31,In_1035,In_1717);
nor U32 (N_32,In_228,In_1880);
and U33 (N_33,In_968,In_1532);
xor U34 (N_34,In_661,In_1089);
nand U35 (N_35,In_842,In_782);
and U36 (N_36,In_1263,In_1770);
or U37 (N_37,In_11,In_725);
xor U38 (N_38,In_697,In_1464);
or U39 (N_39,In_1487,In_1877);
or U40 (N_40,In_195,In_1795);
or U41 (N_41,In_532,In_1350);
xnor U42 (N_42,In_982,In_1016);
or U43 (N_43,In_1910,In_829);
xor U44 (N_44,In_375,In_1833);
xor U45 (N_45,In_17,In_790);
or U46 (N_46,In_395,In_1907);
and U47 (N_47,In_152,In_1447);
nor U48 (N_48,In_251,In_876);
and U49 (N_49,In_946,In_649);
and U50 (N_50,In_823,In_1839);
nor U51 (N_51,In_1038,In_760);
nor U52 (N_52,In_932,In_1358);
nand U53 (N_53,In_355,In_1085);
and U54 (N_54,In_1310,In_1826);
or U55 (N_55,In_1033,In_306);
nand U56 (N_56,In_95,In_963);
nand U57 (N_57,In_1531,In_336);
nand U58 (N_58,In_190,In_1824);
nor U59 (N_59,In_1469,In_1793);
nor U60 (N_60,In_365,In_1386);
nor U61 (N_61,In_44,In_241);
nor U62 (N_62,In_1534,In_1345);
and U63 (N_63,In_1385,In_1661);
and U64 (N_64,In_114,In_1555);
nand U65 (N_65,In_1699,In_639);
xnor U66 (N_66,In_1074,In_490);
nand U67 (N_67,In_1922,In_174);
or U68 (N_68,In_929,In_1275);
nor U69 (N_69,In_873,In_1110);
nand U70 (N_70,In_721,In_1070);
nor U71 (N_71,In_545,In_1317);
nor U72 (N_72,In_1481,In_1837);
and U73 (N_73,In_1966,In_574);
and U74 (N_74,In_1973,In_703);
xor U75 (N_75,In_1149,In_1112);
xnor U76 (N_76,In_149,In_1820);
nand U77 (N_77,In_1891,In_1856);
xor U78 (N_78,In_1445,In_1048);
nand U79 (N_79,In_337,In_965);
and U80 (N_80,In_715,In_1219);
and U81 (N_81,In_1707,In_1809);
and U82 (N_82,In_821,In_1941);
and U83 (N_83,In_294,In_1143);
nand U84 (N_84,In_643,In_60);
nand U85 (N_85,In_1790,In_481);
nand U86 (N_86,In_726,In_187);
xnor U87 (N_87,In_235,In_1247);
nor U88 (N_88,In_1117,In_636);
xnor U89 (N_89,In_642,In_1363);
nand U90 (N_90,In_1817,In_1865);
or U91 (N_91,In_1313,In_353);
nor U92 (N_92,In_1946,In_1504);
or U93 (N_93,In_1640,In_1101);
and U94 (N_94,In_1539,In_411);
or U95 (N_95,In_889,In_1751);
and U96 (N_96,In_299,In_261);
xor U97 (N_97,In_1256,In_131);
and U98 (N_98,In_880,In_1103);
xnor U99 (N_99,In_1676,In_571);
nor U100 (N_100,In_470,In_409);
nor U101 (N_101,In_1977,In_1899);
or U102 (N_102,In_867,In_1230);
xnor U103 (N_103,In_397,In_287);
nand U104 (N_104,In_668,In_284);
xor U105 (N_105,In_129,In_1193);
xnor U106 (N_106,In_833,In_633);
nor U107 (N_107,In_812,In_273);
nor U108 (N_108,In_1129,In_1478);
xor U109 (N_109,In_817,In_435);
and U110 (N_110,In_1146,In_391);
and U111 (N_111,In_500,In_1606);
nand U112 (N_112,In_1347,In_1359);
or U113 (N_113,In_449,In_1967);
xor U114 (N_114,In_1620,In_1357);
xor U115 (N_115,In_959,In_1254);
xor U116 (N_116,In_1584,In_750);
or U117 (N_117,In_621,In_1871);
nand U118 (N_118,In_1238,In_341);
or U119 (N_119,In_1370,In_1763);
nand U120 (N_120,In_1902,In_587);
and U121 (N_121,In_1834,In_1988);
or U122 (N_122,In_810,In_164);
nor U123 (N_123,In_1080,In_727);
nor U124 (N_124,In_1395,In_1269);
and U125 (N_125,In_1540,In_1411);
nor U126 (N_126,In_1610,In_533);
nor U127 (N_127,In_1314,In_663);
nand U128 (N_128,In_415,In_848);
nand U129 (N_129,In_1602,In_647);
xor U130 (N_130,In_795,In_342);
and U131 (N_131,In_196,In_1167);
and U132 (N_132,In_485,In_84);
and U133 (N_133,In_1490,In_1928);
and U134 (N_134,In_1692,In_247);
and U135 (N_135,In_430,In_591);
and U136 (N_136,In_981,In_599);
and U137 (N_137,In_298,In_1419);
nand U138 (N_138,In_1991,In_1831);
xor U139 (N_139,In_624,In_180);
nand U140 (N_140,In_75,In_296);
or U141 (N_141,In_1944,In_1202);
nand U142 (N_142,In_349,In_1403);
nand U143 (N_143,In_1563,In_1135);
or U144 (N_144,In_214,In_1960);
nor U145 (N_145,In_389,In_1601);
nand U146 (N_146,In_1327,In_665);
xnor U147 (N_147,In_1201,In_382);
nor U148 (N_148,In_1787,In_1326);
xnor U149 (N_149,In_868,In_1923);
xnor U150 (N_150,In_1734,In_1878);
xnor U151 (N_151,In_1558,In_1);
and U152 (N_152,In_31,In_874);
xor U153 (N_153,In_834,In_454);
or U154 (N_154,In_595,In_901);
or U155 (N_155,In_1852,In_1393);
and U156 (N_156,In_69,In_106);
nor U157 (N_157,In_1816,In_484);
or U158 (N_158,In_575,In_1012);
xnor U159 (N_159,In_410,In_534);
nor U160 (N_160,In_1200,In_285);
or U161 (N_161,In_1162,In_91);
nand U162 (N_162,In_758,N_92);
and U163 (N_163,In_986,In_1303);
nor U164 (N_164,In_1718,In_1547);
nand U165 (N_165,In_1511,In_1832);
nand U166 (N_166,In_1082,In_39);
nand U167 (N_167,In_335,N_133);
nand U168 (N_168,In_846,In_539);
or U169 (N_169,In_869,In_137);
xnor U170 (N_170,In_453,N_156);
nand U171 (N_171,In_1905,In_1776);
nor U172 (N_172,In_1272,N_77);
or U173 (N_173,In_1114,In_1881);
nor U174 (N_174,In_1528,In_1835);
nor U175 (N_175,In_1722,In_597);
xnor U176 (N_176,In_209,In_80);
xnor U177 (N_177,In_111,In_863);
or U178 (N_178,In_517,In_1111);
nor U179 (N_179,In_999,In_1471);
nor U180 (N_180,In_1150,In_1329);
xnor U181 (N_181,In_1716,In_1291);
nand U182 (N_182,In_434,In_1051);
nand U183 (N_183,In_789,In_418);
and U184 (N_184,In_523,N_6);
and U185 (N_185,In_1587,N_130);
nor U186 (N_186,In_1245,In_1997);
nor U187 (N_187,In_1428,In_958);
or U188 (N_188,In_1221,In_1575);
and U189 (N_189,In_1761,In_1286);
or U190 (N_190,In_13,In_947);
or U191 (N_191,N_0,N_157);
nand U192 (N_192,In_1451,N_26);
xnor U193 (N_193,In_879,In_757);
xor U194 (N_194,In_788,In_837);
or U195 (N_195,In_502,In_1622);
nand U196 (N_196,In_358,In_978);
or U197 (N_197,In_992,In_627);
xor U198 (N_198,In_250,In_1232);
nand U199 (N_199,In_676,In_941);
nor U200 (N_200,In_1581,In_1011);
xnor U201 (N_201,In_248,In_471);
nor U202 (N_202,In_1289,In_1192);
and U203 (N_203,In_79,In_1959);
or U204 (N_204,In_1679,In_1690);
and U205 (N_205,In_1672,In_1348);
nor U206 (N_206,In_1203,In_1371);
nor U207 (N_207,In_1706,In_1641);
and U208 (N_208,In_1182,In_680);
or U209 (N_209,In_2,In_1595);
nor U210 (N_210,In_1299,N_95);
nor U211 (N_211,In_1251,In_670);
xor U212 (N_212,In_210,In_1460);
or U213 (N_213,N_22,In_1233);
xor U214 (N_214,In_1594,In_264);
nor U215 (N_215,In_678,In_799);
and U216 (N_216,In_1548,N_110);
or U217 (N_217,In_1281,In_1996);
nand U218 (N_218,In_316,In_1573);
and U219 (N_219,In_1505,N_28);
nor U220 (N_220,In_611,In_230);
nor U221 (N_221,In_1911,In_1674);
xnor U222 (N_222,In_188,In_421);
nand U223 (N_223,In_1368,In_1343);
or U224 (N_224,In_742,In_1639);
or U225 (N_225,In_1943,In_1053);
or U226 (N_226,N_21,In_872);
nor U227 (N_227,N_100,In_1389);
and U228 (N_228,In_267,In_438);
xor U229 (N_229,In_1963,In_974);
nand U230 (N_230,In_383,N_79);
or U231 (N_231,In_260,In_1158);
nand U232 (N_232,In_1413,In_240);
nor U233 (N_233,In_332,In_1607);
nand U234 (N_234,In_1971,In_1227);
nand U235 (N_235,In_844,N_102);
or U236 (N_236,In_1749,In_1638);
or U237 (N_237,In_1778,In_1168);
nor U238 (N_238,In_1183,In_1515);
or U239 (N_239,In_371,In_328);
and U240 (N_240,In_818,In_584);
or U241 (N_241,N_16,In_1617);
xnor U242 (N_242,In_1093,In_900);
or U243 (N_243,In_955,In_761);
or U244 (N_244,In_361,In_1588);
xnor U245 (N_245,In_1470,In_178);
nand U246 (N_246,In_1418,In_52);
and U247 (N_247,In_1637,N_124);
nor U248 (N_248,In_427,In_515);
nor U249 (N_249,In_836,In_985);
nand U250 (N_250,In_891,In_1092);
nand U251 (N_251,In_1260,In_1086);
xor U252 (N_252,N_62,In_1791);
nand U253 (N_253,In_694,In_1955);
and U254 (N_254,In_1866,In_222);
or U255 (N_255,In_1542,In_354);
or U256 (N_256,In_1962,In_274);
nand U257 (N_257,In_559,In_1364);
nor U258 (N_258,In_289,In_1675);
nand U259 (N_259,In_1295,In_1130);
nor U260 (N_260,In_1727,In_603);
and U261 (N_261,In_1204,In_1982);
nand U262 (N_262,In_1618,In_1597);
nor U263 (N_263,In_1328,N_111);
or U264 (N_264,In_579,In_689);
nand U265 (N_265,In_917,In_51);
or U266 (N_266,In_1536,In_1229);
and U267 (N_267,In_333,In_424);
and U268 (N_268,In_1496,In_1404);
and U269 (N_269,N_149,In_105);
nor U270 (N_270,In_550,In_1585);
nor U271 (N_271,In_1644,N_150);
and U272 (N_272,In_1572,In_708);
nor U273 (N_273,In_1990,In_785);
and U274 (N_274,In_1252,In_1745);
xnor U275 (N_275,In_1331,In_994);
xnor U276 (N_276,In_107,In_962);
nor U277 (N_277,N_59,In_1777);
or U278 (N_278,In_1882,In_1268);
xor U279 (N_279,In_1431,N_99);
or U280 (N_280,N_154,In_1147);
nand U281 (N_281,N_144,In_589);
and U282 (N_282,In_1104,In_563);
and U283 (N_283,N_40,In_857);
nand U284 (N_284,In_572,In_1214);
xnor U285 (N_285,In_711,In_89);
or U286 (N_286,In_1467,In_551);
or U287 (N_287,In_1173,In_540);
xor U288 (N_288,In_1398,In_566);
nor U289 (N_289,In_856,N_159);
or U290 (N_290,N_67,In_360);
nor U291 (N_291,N_25,In_1334);
and U292 (N_292,In_1935,In_1965);
and U293 (N_293,In_1579,In_1261);
xor U294 (N_294,In_675,In_847);
nand U295 (N_295,In_5,In_154);
nor U296 (N_296,In_893,In_1811);
or U297 (N_297,In_1121,In_1613);
and U298 (N_298,In_1739,In_1609);
nand U299 (N_299,In_367,In_121);
or U300 (N_300,In_1066,N_83);
nand U301 (N_301,In_265,N_74);
or U302 (N_302,N_23,In_1134);
nand U303 (N_303,In_1836,N_88);
nor U304 (N_304,N_2,In_1686);
or U305 (N_305,In_717,In_1559);
nor U306 (N_306,In_269,In_1851);
and U307 (N_307,In_1237,In_989);
and U308 (N_308,In_184,In_1069);
nand U309 (N_309,N_66,In_457);
nor U310 (N_310,In_23,In_814);
nand U311 (N_311,In_775,In_295);
nand U312 (N_312,In_1591,In_1264);
xnor U313 (N_313,In_1550,In_815);
nor U314 (N_314,In_216,In_1766);
or U315 (N_315,In_552,In_1312);
and U316 (N_316,In_472,In_822);
and U317 (N_317,In_1813,In_998);
and U318 (N_318,In_1476,In_1583);
nand U319 (N_319,In_1760,In_150);
and U320 (N_320,In_1500,In_1125);
xor U321 (N_321,In_1535,In_1887);
nor U322 (N_322,In_745,In_1665);
nand U323 (N_323,In_1994,In_1488);
or U324 (N_324,In_570,In_175);
nand U325 (N_325,In_952,In_1729);
xnor U326 (N_326,In_43,N_51);
nor U327 (N_327,In_1044,In_124);
nor U328 (N_328,In_28,In_414);
and U329 (N_329,In_1896,In_1262);
and U330 (N_330,In_112,In_1600);
nand U331 (N_331,In_699,In_218);
or U332 (N_332,N_278,In_1450);
xnor U333 (N_333,In_996,N_318);
and U334 (N_334,In_1294,In_1377);
nand U335 (N_335,In_1556,In_565);
or U336 (N_336,In_1772,In_310);
nand U337 (N_337,N_257,N_120);
or U338 (N_338,N_91,In_381);
and U339 (N_339,In_286,In_226);
xnor U340 (N_340,In_315,In_255);
and U341 (N_341,N_223,In_1266);
xnor U342 (N_342,In_505,In_1844);
and U343 (N_343,In_864,In_786);
xor U344 (N_344,N_211,In_77);
or U345 (N_345,In_322,N_60);
or U346 (N_346,In_1480,In_1666);
or U347 (N_347,In_640,In_1397);
nor U348 (N_348,In_1000,In_1355);
nand U349 (N_349,In_1822,In_100);
xnor U350 (N_350,In_1987,In_1634);
nor U351 (N_351,In_637,In_1062);
or U352 (N_352,N_52,In_899);
and U353 (N_353,N_267,In_707);
xor U354 (N_354,In_508,In_1517);
nand U355 (N_355,In_776,In_909);
nand U356 (N_356,In_548,In_1410);
or U357 (N_357,In_657,In_1325);
nand U358 (N_358,N_199,In_652);
nor U359 (N_359,In_1094,In_811);
xnor U360 (N_360,In_86,In_98);
nand U361 (N_361,In_1346,N_214);
and U362 (N_362,In_1732,In_57);
or U363 (N_363,In_519,In_308);
nor U364 (N_364,In_1870,In_1424);
nand U365 (N_365,In_768,In_1925);
nor U366 (N_366,In_1152,In_743);
or U367 (N_367,In_1443,In_1455);
nand U368 (N_368,In_1222,N_68);
and U369 (N_369,N_166,N_277);
or U370 (N_370,In_1297,In_1166);
nor U371 (N_371,N_76,In_1611);
or U372 (N_372,In_229,In_93);
nand U373 (N_373,In_19,N_262);
xnor U374 (N_374,In_921,In_70);
nand U375 (N_375,N_94,In_223);
or U376 (N_376,In_1280,In_1305);
xnor U377 (N_377,In_234,In_890);
xnor U378 (N_378,In_63,N_30);
or U379 (N_379,In_1034,In_1537);
nand U380 (N_380,In_1097,N_236);
nor U381 (N_381,In_462,N_314);
xnor U382 (N_382,In_231,In_705);
xnor U383 (N_383,In_498,In_1697);
nand U384 (N_384,In_233,In_1118);
nor U385 (N_385,In_733,In_1735);
nand U386 (N_386,In_1945,In_1917);
or U387 (N_387,In_720,In_292);
nand U388 (N_388,In_1438,N_104);
nand U389 (N_389,In_1574,In_1914);
or U390 (N_390,In_1934,N_84);
nand U391 (N_391,In_82,In_1105);
nand U392 (N_392,In_807,In_1884);
or U393 (N_393,N_19,In_1412);
nor U394 (N_394,In_141,In_253);
nand U395 (N_395,In_27,In_1191);
xor U396 (N_396,In_1646,In_1840);
xnor U397 (N_397,In_674,In_1196);
nand U398 (N_398,In_1850,In_46);
or U399 (N_399,In_773,N_134);
xor U400 (N_400,In_1224,In_276);
or U401 (N_401,In_25,In_466);
or U402 (N_402,In_1198,In_1892);
or U403 (N_403,In_1919,In_72);
or U404 (N_404,N_163,In_1803);
or U405 (N_405,N_114,In_1384);
and U406 (N_406,N_237,In_507);
nor U407 (N_407,In_860,In_1789);
nand U408 (N_408,N_316,In_135);
nand U409 (N_409,In_1938,N_197);
nand U410 (N_410,N_127,In_653);
and U411 (N_411,N_41,In_553);
xor U412 (N_412,In_94,In_585);
nand U413 (N_413,In_852,In_92);
xnor U414 (N_414,In_58,N_106);
nor U415 (N_415,In_442,N_220);
xnor U416 (N_416,In_1593,In_1590);
xor U417 (N_417,In_957,In_1197);
nand U418 (N_418,In_1071,In_136);
nor U419 (N_419,In_1099,In_1972);
xor U420 (N_420,N_215,In_1562);
or U421 (N_421,In_1172,In_827);
xor U422 (N_422,In_1715,In_35);
or U423 (N_423,N_238,In_1440);
nor U424 (N_424,In_1700,N_273);
or U425 (N_425,N_245,In_1045);
nor U426 (N_426,In_194,In_1818);
and U427 (N_427,In_1879,N_300);
and U428 (N_428,N_80,In_1360);
or U429 (N_429,In_325,In_1796);
or U430 (N_430,In_496,In_309);
and U431 (N_431,N_303,In_684);
nor U432 (N_432,In_1042,N_293);
or U433 (N_433,In_1171,In_718);
nor U434 (N_434,In_991,In_1804);
xnor U435 (N_435,In_156,In_1926);
nand U436 (N_436,In_582,In_1545);
nor U437 (N_437,In_1376,In_878);
and U438 (N_438,In_1217,In_347);
xnor U439 (N_439,In_1475,In_330);
and U440 (N_440,In_666,In_1889);
and U441 (N_441,N_239,In_1259);
nand U442 (N_442,In_1136,In_221);
and U443 (N_443,In_1039,In_1847);
xnor U444 (N_444,In_918,In_747);
nand U445 (N_445,In_464,In_1499);
xor U446 (N_446,N_263,N_295);
nand U447 (N_447,In_997,In_282);
or U448 (N_448,In_133,In_580);
or U449 (N_449,In_1372,In_1554);
and U450 (N_450,In_147,In_1319);
and U451 (N_451,N_232,In_76);
or U452 (N_452,In_1119,In_1170);
nor U453 (N_453,In_1378,In_1151);
or U454 (N_454,N_45,In_344);
or U455 (N_455,N_319,In_1181);
xnor U456 (N_456,In_1736,In_1888);
nand U457 (N_457,In_1387,In_1560);
nand U458 (N_458,In_1797,In_1332);
nor U459 (N_459,In_1037,N_259);
xnor U460 (N_460,N_275,In_96);
xor U461 (N_461,In_1724,N_308);
and U462 (N_462,N_170,N_141);
or U463 (N_463,In_1434,In_117);
xor U464 (N_464,In_1383,In_1065);
xor U465 (N_465,In_1703,In_1514);
nand U466 (N_466,In_1489,In_1022);
nor U467 (N_467,N_285,In_1408);
xnor U468 (N_468,N_158,In_1276);
xnor U469 (N_469,In_146,In_56);
xor U470 (N_470,In_1670,N_235);
nand U471 (N_471,In_1862,In_151);
and U472 (N_472,In_1165,In_528);
or U473 (N_473,In_1195,In_1465);
nand U474 (N_474,In_513,In_970);
nand U475 (N_475,In_641,In_854);
or U476 (N_476,N_195,In_1918);
nand U477 (N_477,In_1282,In_1626);
and U478 (N_478,In_167,In_408);
nor U479 (N_479,In_1421,In_1041);
xor U480 (N_480,In_1462,In_1702);
or U481 (N_481,N_233,In_631);
nor U482 (N_482,N_93,In_975);
and U483 (N_483,In_1758,In_906);
or U484 (N_484,In_443,In_926);
nor U485 (N_485,N_403,In_1740);
nand U486 (N_486,In_1895,In_351);
nand U487 (N_487,In_1253,In_625);
nor U488 (N_488,N_177,In_499);
xor U489 (N_489,In_682,In_1605);
xor U490 (N_490,In_1897,N_396);
and U491 (N_491,In_783,In_215);
and U492 (N_492,N_37,In_979);
xor U493 (N_493,N_430,N_392);
nor U494 (N_494,N_473,In_1614);
nor U495 (N_495,In_62,In_366);
or U496 (N_496,In_1783,In_1569);
or U497 (N_497,In_1767,N_87);
xnor U498 (N_498,In_509,In_1933);
nor U499 (N_499,In_1890,In_537);
nand U500 (N_500,In_1544,In_1341);
nand U501 (N_501,N_153,In_1240);
and U502 (N_502,N_375,In_1362);
nor U503 (N_503,In_1283,In_1961);
or U504 (N_504,In_1784,In_1599);
nand U505 (N_505,In_774,In_486);
nand U506 (N_506,N_82,In_208);
nand U507 (N_507,N_345,In_1425);
and U508 (N_508,N_286,In_1430);
or U509 (N_509,N_382,N_377);
and U510 (N_510,In_904,In_1029);
nand U511 (N_511,In_961,N_39);
nor U512 (N_512,In_895,In_1860);
xnor U513 (N_513,In_1709,N_422);
or U514 (N_514,In_1728,In_168);
xnor U515 (N_515,In_74,N_174);
xnor U516 (N_516,In_103,In_1306);
nand U517 (N_517,In_547,N_188);
nor U518 (N_518,In_1091,In_1047);
or U519 (N_519,In_207,N_65);
or U520 (N_520,N_454,In_1388);
or U521 (N_521,N_390,In_567);
nor U522 (N_522,N_255,N_90);
or U523 (N_523,In_1983,N_397);
and U524 (N_524,In_1508,In_936);
and U525 (N_525,In_1519,In_1442);
nor U526 (N_526,N_331,In_224);
nor U527 (N_527,N_12,N_89);
and U528 (N_528,In_907,In_609);
xor U529 (N_529,In_514,N_347);
xnor U530 (N_530,In_1586,In_1512);
or U531 (N_531,N_289,In_16);
nor U532 (N_532,N_205,In_1141);
and U533 (N_533,In_387,In_504);
xor U534 (N_534,In_767,In_185);
xor U535 (N_535,In_808,In_1493);
xor U536 (N_536,N_187,In_350);
or U537 (N_537,In_278,In_569);
nor U538 (N_538,In_1215,N_394);
xor U539 (N_539,N_47,N_186);
xnor U540 (N_540,In_938,In_1279);
nand U541 (N_541,In_12,In_816);
nor U542 (N_542,In_108,In_1498);
xor U543 (N_543,N_410,In_348);
nor U544 (N_544,In_1330,In_598);
and U545 (N_545,In_1714,N_43);
and U546 (N_546,In_1001,N_132);
and U547 (N_547,N_409,In_1366);
or U548 (N_548,In_883,In_1453);
and U549 (N_549,In_1503,N_20);
and U550 (N_550,N_117,In_1900);
nand U551 (N_551,In_728,N_441);
and U552 (N_552,In_21,N_406);
or U553 (N_553,N_368,In_393);
nor U554 (N_554,N_85,In_538);
xnor U555 (N_555,N_426,N_281);
or U556 (N_556,In_1073,In_1969);
or U557 (N_557,In_554,In_1226);
xor U558 (N_558,In_1405,N_477);
and U559 (N_559,In_139,N_306);
nor U560 (N_560,In_263,In_1570);
or U561 (N_561,In_1307,In_1659);
and U562 (N_562,In_143,N_13);
nor U563 (N_563,In_1932,N_475);
or U564 (N_564,In_142,In_193);
nand U565 (N_565,In_1416,In_1005);
nor U566 (N_566,In_612,N_175);
and U567 (N_567,In_1270,In_1211);
or U568 (N_568,In_1250,In_586);
and U569 (N_569,In_696,In_18);
nand U570 (N_570,In_1652,N_399);
nand U571 (N_571,In_1979,In_380);
nor U572 (N_572,N_208,In_1433);
or U573 (N_573,In_50,In_695);
nor U574 (N_574,In_832,In_927);
and U575 (N_575,N_387,In_1949);
or U576 (N_576,In_1904,In_971);
or U577 (N_577,In_1603,N_328);
or U578 (N_578,In_1807,In_236);
nand U579 (N_579,N_408,In_118);
and U580 (N_580,In_1235,In_1825);
xnor U581 (N_581,In_1023,In_1993);
or U582 (N_582,In_1989,In_1571);
and U583 (N_583,In_331,In_1218);
or U584 (N_584,In_1974,In_1523);
and U585 (N_585,In_1507,In_719);
and U586 (N_586,In_851,In_1695);
nand U587 (N_587,In_390,In_990);
nand U588 (N_588,N_414,In_125);
or U589 (N_589,In_1998,In_1509);
nor U590 (N_590,In_701,N_361);
xor U591 (N_591,In_1802,N_456);
or U592 (N_592,In_480,N_270);
xnor U593 (N_593,In_1849,N_416);
nor U594 (N_594,In_497,In_1648);
and U595 (N_595,In_179,In_610);
nand U596 (N_596,N_189,In_1190);
nand U597 (N_597,In_1948,In_734);
and U598 (N_598,In_1608,In_969);
xor U599 (N_599,In_802,N_251);
and U600 (N_600,N_317,In_1582);
or U601 (N_601,N_449,N_269);
and U602 (N_602,In_1635,In_1698);
xnor U603 (N_603,In_321,In_1333);
xor U604 (N_604,In_450,In_651);
nand U605 (N_605,N_115,In_1055);
and U606 (N_606,In_805,In_618);
or U607 (N_607,In_1392,In_1604);
and U608 (N_608,N_17,In_1164);
nand U609 (N_609,N_284,In_1194);
or U610 (N_610,In_792,In_885);
nand U611 (N_611,In_1527,N_453);
or U612 (N_612,In_271,N_322);
xor U613 (N_613,N_228,In_1576);
xnor U614 (N_614,In_949,In_845);
nand U615 (N_615,In_1186,In_1311);
nand U616 (N_616,In_602,In_1682);
or U617 (N_617,In_495,In_1738);
or U618 (N_618,In_487,In_1936);
or U619 (N_619,In_712,In_1274);
nand U620 (N_620,In_1792,In_1768);
nor U621 (N_621,N_138,In_20);
or U622 (N_622,N_450,In_1771);
nor U623 (N_623,In_428,In_831);
and U624 (N_624,In_1506,In_1859);
nand U625 (N_625,In_288,In_493);
xor U626 (N_626,In_771,In_1457);
and U627 (N_627,In_272,In_1551);
xor U628 (N_628,In_419,In_1422);
or U629 (N_629,In_1940,In_473);
or U630 (N_630,In_755,In_1701);
or U631 (N_631,In_564,In_677);
nor U632 (N_632,In_281,In_866);
nand U633 (N_633,In_892,N_151);
nor U634 (N_634,In_1957,In_238);
nand U635 (N_635,In_1510,In_385);
xnor U636 (N_636,In_1209,In_1942);
or U637 (N_637,N_167,N_434);
nor U638 (N_638,In_173,In_345);
and U639 (N_639,In_36,In_593);
xor U640 (N_640,In_1309,In_320);
nor U641 (N_641,In_420,N_3);
xnor U642 (N_642,N_471,In_809);
nor U643 (N_643,In_1720,In_1516);
xor U644 (N_644,In_1231,In_1557);
xor U645 (N_645,In_664,In_1801);
nor U646 (N_646,N_507,N_231);
nor U647 (N_647,N_260,In_290);
nand U648 (N_648,In_1036,N_570);
or U649 (N_649,In_916,In_176);
or U650 (N_650,In_628,In_882);
nand U651 (N_651,N_592,N_612);
nand U652 (N_652,In_83,In_739);
xnor U653 (N_653,N_604,N_461);
nand U654 (N_654,In_15,In_544);
and U655 (N_655,N_446,In_1142);
or U656 (N_656,In_1636,In_561);
nand U657 (N_657,In_1207,N_557);
xor U658 (N_658,In_744,In_126);
or U659 (N_659,In_1684,In_1342);
xnor U660 (N_660,In_803,N_563);
nand U661 (N_661,N_234,In_398);
nand U662 (N_662,N_439,In_1349);
xnor U663 (N_663,N_352,In_1883);
or U664 (N_664,In_1951,N_423);
nand U665 (N_665,N_591,In_1894);
and U666 (N_666,N_323,In_1427);
and U667 (N_667,In_536,In_1980);
or U668 (N_668,N_311,N_622);
nor U669 (N_669,In_459,In_1014);
or U670 (N_670,In_1485,N_488);
nand U671 (N_671,In_1521,In_865);
nand U672 (N_672,N_624,In_1316);
nor U673 (N_673,N_487,In_444);
xor U674 (N_674,In_644,In_429);
nand U675 (N_675,In_4,N_298);
and U676 (N_676,In_446,In_1064);
nor U677 (N_677,In_1667,In_300);
nor U678 (N_678,In_1673,In_417);
nand U679 (N_679,N_586,In_1271);
nand U680 (N_680,N_627,N_324);
and U681 (N_681,In_153,In_613);
nand U682 (N_682,In_993,In_779);
and U683 (N_683,N_571,N_596);
or U684 (N_684,In_1857,N_18);
nand U685 (N_685,In_191,In_1819);
or U686 (N_686,In_1446,N_344);
xnor U687 (N_687,N_46,N_54);
or U688 (N_688,In_64,In_145);
xnor U689 (N_689,In_1156,In_3);
or U690 (N_690,In_227,In_102);
or U691 (N_691,In_467,In_828);
or U692 (N_692,In_113,In_1930);
nor U693 (N_693,N_244,In_549);
nand U694 (N_694,N_31,In_312);
or U695 (N_695,N_179,In_370);
or U696 (N_696,In_1127,N_330);
and U697 (N_697,N_218,In_138);
nor U698 (N_698,N_265,In_1391);
or U699 (N_699,In_1913,In_1009);
xor U700 (N_700,N_605,N_210);
or U701 (N_701,In_157,In_1019);
or U702 (N_702,In_884,In_160);
or U703 (N_703,In_148,In_1322);
or U704 (N_704,In_714,N_630);
and U705 (N_705,N_492,In_90);
or U706 (N_706,In_1072,In_686);
nand U707 (N_707,In_706,In_1375);
xnor U708 (N_708,In_1058,In_1920);
and U709 (N_709,In_219,N_183);
nor U710 (N_710,In_202,In_1721);
xor U711 (N_711,N_384,In_1629);
xor U712 (N_712,In_960,In_531);
nand U713 (N_713,In_54,In_1437);
nor U714 (N_714,In_59,N_548);
and U715 (N_715,N_33,N_336);
nand U716 (N_716,N_516,In_1642);
and U717 (N_717,In_578,In_692);
nor U718 (N_718,In_158,In_1567);
and U719 (N_719,In_1417,In_1956);
or U720 (N_720,In_384,N_447);
and U721 (N_721,N_63,In_1292);
xor U722 (N_722,In_134,N_398);
or U723 (N_723,In_1999,In_492);
or U724 (N_724,In_416,In_1087);
or U725 (N_725,In_501,In_1175);
nor U726 (N_726,In_913,In_422);
and U727 (N_727,In_1439,In_1863);
or U728 (N_728,In_752,N_626);
and U729 (N_729,N_638,N_198);
and U730 (N_730,In_1906,N_628);
nand U731 (N_731,In_859,In_483);
or U732 (N_732,In_1903,N_116);
nor U733 (N_733,In_920,In_951);
nand U734 (N_734,In_1621,N_168);
xor U735 (N_735,In_1180,In_1861);
nand U736 (N_736,N_178,In_630);
nor U737 (N_737,In_1169,In_806);
or U738 (N_738,N_160,In_1188);
xnor U739 (N_739,N_472,In_769);
xor U740 (N_740,In_1630,N_249);
xnor U741 (N_741,In_1708,N_530);
xor U742 (N_742,N_497,N_247);
xnor U743 (N_743,N_600,In_503);
xnor U744 (N_744,N_369,In_568);
and U745 (N_745,N_505,N_221);
nand U746 (N_746,In_716,N_343);
or U747 (N_747,In_115,In_1223);
and U748 (N_748,In_645,In_616);
xor U749 (N_749,In_203,N_512);
or U750 (N_750,In_915,In_1612);
xnor U751 (N_751,N_196,In_1241);
and U752 (N_752,N_405,N_121);
nor U753 (N_753,N_313,N_617);
xnor U754 (N_754,In_1337,In_700);
and U755 (N_755,N_629,In_323);
and U756 (N_756,In_363,N_553);
nor U757 (N_757,In_1220,N_32);
or U758 (N_758,N_534,In_660);
xor U759 (N_759,N_86,In_1937);
nand U760 (N_760,In_313,In_1561);
and U761 (N_761,In_339,N_565);
nand U762 (N_762,N_602,In_671);
and U763 (N_763,N_561,In_607);
or U764 (N_764,In_488,N_365);
nor U765 (N_765,In_650,N_9);
nand U766 (N_766,In_1525,In_1486);
and U767 (N_767,N_385,In_600);
xor U768 (N_768,In_26,N_501);
and U769 (N_769,In_1318,In_482);
or U770 (N_770,In_307,N_383);
or U771 (N_771,In_1678,In_144);
and U772 (N_772,N_229,In_546);
xnor U773 (N_773,In_953,In_1315);
xor U774 (N_774,N_142,In_283);
or U775 (N_775,In_973,N_618);
nand U776 (N_776,In_681,N_162);
nor U777 (N_777,In_1855,In_1052);
nand U778 (N_778,In_311,In_781);
xnor U779 (N_779,N_484,In_1079);
and U780 (N_780,In_1623,N_107);
and U781 (N_781,In_945,In_1799);
xor U782 (N_782,In_524,In_373);
xor U783 (N_783,In_1027,In_1096);
nor U784 (N_784,In_1098,In_838);
or U785 (N_785,In_1553,In_1876);
and U786 (N_786,In_629,N_44);
xnor U787 (N_787,N_268,In_691);
nor U788 (N_788,In_1725,N_126);
nand U789 (N_789,In_359,In_601);
nor U790 (N_790,In_270,In_562);
and U791 (N_791,N_579,In_1078);
nand U792 (N_792,N_140,N_435);
and U793 (N_793,In_1381,N_415);
nor U794 (N_794,In_1351,N_555);
xor U795 (N_795,In_1407,In_352);
nand U796 (N_796,In_1773,In_1908);
or U797 (N_797,In_445,In_244);
nand U798 (N_798,In_688,In_948);
and U799 (N_799,In_1664,In_1454);
nand U800 (N_800,In_1361,In_535);
nand U801 (N_801,In_1985,N_536);
xnor U802 (N_802,N_659,In_1828);
or U803 (N_803,In_1015,In_1102);
or U804 (N_804,N_274,N_332);
and U805 (N_805,N_712,N_583);
xnor U806 (N_806,In_935,In_232);
and U807 (N_807,In_556,N_688);
nor U808 (N_808,In_655,In_394);
or U809 (N_809,In_1248,In_1176);
or U810 (N_810,In_1976,N_350);
and U811 (N_811,N_452,In_710);
nand U812 (N_812,N_676,In_1800);
or U813 (N_813,In_1909,N_702);
nand U814 (N_814,N_769,In_1806);
nor U815 (N_815,In_905,In_1302);
and U816 (N_816,N_225,N_357);
or U817 (N_817,In_1461,In_1473);
nor U818 (N_818,In_887,N_620);
xor U819 (N_819,In_1781,N_593);
or U820 (N_820,N_476,In_1075);
and U821 (N_821,In_1981,In_1669);
xnor U822 (N_822,In_843,N_706);
or U823 (N_823,N_202,N_610);
and U824 (N_824,In_1759,In_356);
nor U825 (N_825,In_279,N_1);
xor U826 (N_826,N_176,In_1578);
nor U827 (N_827,N_674,N_474);
nor U828 (N_828,In_24,In_954);
nand U829 (N_829,In_494,In_291);
and U830 (N_830,In_338,In_1290);
or U831 (N_831,N_524,In_912);
and U832 (N_832,N_680,In_452);
nand U833 (N_833,In_1077,In_1046);
xor U834 (N_834,N_272,In_376);
nand U835 (N_835,In_1694,In_1137);
nor U836 (N_836,N_460,In_784);
or U837 (N_837,In_48,In_377);
and U838 (N_838,In_702,N_217);
or U839 (N_839,In_673,In_1010);
xnor U840 (N_840,In_1680,In_617);
or U841 (N_841,In_976,In_200);
nand U842 (N_842,In_778,In_577);
nand U843 (N_843,N_129,In_1810);
xnor U844 (N_844,N_81,N_573);
nor U845 (N_845,In_871,N_432);
or U846 (N_846,N_528,N_282);
or U847 (N_847,In_1677,In_626);
or U848 (N_848,In_1838,N_296);
nand U849 (N_849,N_580,N_486);
and U850 (N_850,In_1300,N_625);
nand U851 (N_851,N_651,In_1927);
or U852 (N_852,In_262,In_1647);
xor U853 (N_853,N_496,In_875);
or U854 (N_854,In_980,In_1288);
and U855 (N_855,N_219,N_458);
nand U856 (N_856,In_30,In_378);
and U857 (N_857,N_5,In_1912);
nor U858 (N_858,N_669,In_305);
or U859 (N_859,In_685,N_572);
xnor U860 (N_860,N_118,In_506);
and U861 (N_861,N_668,In_9);
or U862 (N_862,In_423,In_1533);
nor U863 (N_863,N_64,N_564);
nor U864 (N_864,N_71,N_725);
xor U865 (N_865,In_1655,N_291);
and U866 (N_866,N_788,In_956);
xnor U867 (N_867,In_748,In_127);
nor U868 (N_868,In_1013,N_551);
nand U869 (N_869,In_619,In_245);
nor U870 (N_870,N_784,N_180);
nor U871 (N_871,In_1161,N_748);
or U872 (N_872,N_443,In_654);
and U873 (N_873,In_67,N_635);
nor U874 (N_874,In_1522,N_310);
nand U875 (N_875,N_354,N_672);
xor U876 (N_876,N_351,In_605);
nand U877 (N_877,In_1369,In_877);
and U878 (N_878,In_314,N_616);
nor U879 (N_879,N_733,N_283);
and U880 (N_880,N_606,In_1255);
nor U881 (N_881,N_226,N_537);
and U882 (N_882,N_436,In_1798);
xor U883 (N_883,N_288,In_1456);
or U884 (N_884,N_619,N_707);
nand U885 (N_885,N_632,In_1964);
and U886 (N_886,N_584,N_613);
or U887 (N_887,In_1177,N_401);
and U888 (N_888,In_923,In_372);
or U889 (N_889,N_667,N_798);
or U890 (N_890,In_362,N_342);
nand U891 (N_891,N_276,N_412);
xor U892 (N_892,In_242,In_1468);
nand U893 (N_893,In_1494,N_506);
xor U894 (N_894,N_391,N_400);
and U895 (N_895,In_171,In_400);
xor U896 (N_896,In_615,In_1380);
xor U897 (N_897,In_1139,In_1748);
and U898 (N_898,N_206,N_614);
nand U899 (N_899,In_1336,N_508);
nand U900 (N_900,In_753,N_749);
or U901 (N_901,N_777,In_606);
nor U902 (N_902,In_1841,N_424);
and U903 (N_903,N_790,In_984);
nand U904 (N_904,N_57,N_608);
nand U905 (N_905,N_768,N_184);
nand U906 (N_906,N_653,In_919);
or U907 (N_907,N_601,N_695);
xor U908 (N_908,N_243,In_474);
xor U909 (N_909,N_690,N_660);
and U910 (N_910,In_1444,In_1228);
nor U911 (N_911,In_1953,N_594);
nand U912 (N_912,In_608,In_709);
xnor U913 (N_913,In_1580,In_1484);
nand U914 (N_914,In_862,N_531);
nor U915 (N_915,In_1875,N_779);
nand U916 (N_916,In_399,In_690);
nor U917 (N_917,In_460,In_88);
and U918 (N_918,N_681,N_732);
nor U919 (N_919,N_647,N_27);
nor U920 (N_920,In_1225,In_729);
xnor U921 (N_921,In_163,N_139);
xnor U922 (N_922,In_1713,N_438);
xor U923 (N_923,In_407,N_719);
and U924 (N_924,N_711,In_1115);
and U925 (N_925,N_147,N_722);
nand U926 (N_926,In_166,N_746);
xnor U927 (N_927,N_459,N_366);
xor U928 (N_928,In_1869,N_717);
xnor U929 (N_929,In_1805,N_562);
nor U930 (N_930,In_1757,In_259);
nand U931 (N_931,In_1858,N_726);
or U932 (N_932,In_1452,N_685);
and U933 (N_933,In_1872,In_1868);
or U934 (N_934,In_1324,N_417);
and U935 (N_935,In_1685,In_192);
or U936 (N_936,N_7,N_774);
or U937 (N_937,N_339,N_250);
or U938 (N_938,N_348,In_1821);
or U939 (N_939,In_252,In_510);
nand U940 (N_940,N_56,N_8);
and U941 (N_941,N_201,N_666);
and U942 (N_942,In_1367,In_277);
nor U943 (N_943,In_950,N_216);
or U944 (N_944,In_1132,N_775);
or U945 (N_945,In_1598,In_1415);
xnor U946 (N_946,N_137,N_358);
or U947 (N_947,In_576,In_1992);
nor U948 (N_948,In_1435,N_455);
and U949 (N_949,N_24,In_967);
nand U950 (N_950,In_1423,N_181);
xor U951 (N_951,In_1002,N_294);
nor U952 (N_952,N_302,In_512);
nand U953 (N_953,In_1107,N_662);
or U954 (N_954,N_445,In_246);
and U955 (N_955,N_527,In_469);
nand U956 (N_956,N_763,In_1353);
xnor U957 (N_957,In_1020,In_780);
xor U958 (N_958,N_780,N_587);
xnor U959 (N_959,In_172,N_327);
nor U960 (N_960,N_465,In_1273);
xnor U961 (N_961,In_1340,In_8);
xor U962 (N_962,N_890,In_1124);
nor U963 (N_963,N_655,N_607);
nor U964 (N_964,In_303,N_305);
nand U965 (N_965,In_839,N_145);
and U966 (N_966,In_1662,In_1631);
or U967 (N_967,N_811,N_663);
xnor U968 (N_968,N_190,In_620);
or U969 (N_969,N_597,N_479);
or U970 (N_970,N_312,In_1615);
and U971 (N_971,In_1030,N_892);
nor U972 (N_972,In_800,In_1774);
and U973 (N_973,In_40,In_765);
nand U974 (N_974,In_754,In_1374);
xor U975 (N_975,N_914,In_468);
and U976 (N_976,In_1287,N_480);
nand U977 (N_977,In_1323,In_243);
and U978 (N_978,N_736,N_917);
nor U979 (N_979,N_785,In_318);
or U980 (N_980,In_186,In_1929);
and U981 (N_981,In_1524,N_549);
and U982 (N_982,In_357,In_1566);
nor U983 (N_983,In_1779,In_165);
nor U984 (N_984,In_7,N_934);
nor U985 (N_985,In_604,In_1068);
nor U986 (N_986,N_38,In_475);
nand U987 (N_987,N_710,In_896);
or U988 (N_988,N_922,N_908);
xnor U989 (N_989,N_713,N_822);
nand U990 (N_990,N_849,N_833);
or U991 (N_991,In_1007,In_1491);
nand U992 (N_992,N_585,In_304);
and U993 (N_993,In_1726,In_1786);
and U994 (N_994,In_1400,In_206);
and U995 (N_995,In_855,In_1278);
nand U996 (N_996,In_756,N_776);
xor U997 (N_997,N_812,In_1744);
nor U998 (N_998,N_402,N_395);
or U999 (N_999,In_340,N_113);
xnor U1000 (N_1000,In_436,N_529);
or U1001 (N_1001,N_898,In_1742);
nor U1002 (N_1002,N_590,N_743);
nand U1003 (N_1003,In_1402,In_964);
or U1004 (N_1004,N_692,In_763);
and U1005 (N_1005,N_797,In_594);
or U1006 (N_1006,N_419,N_173);
and U1007 (N_1007,In_746,In_204);
nor U1008 (N_1008,N_885,In_1145);
and U1009 (N_1009,N_428,In_1061);
and U1010 (N_1010,In_672,N_671);
xnor U1011 (N_1011,N_912,In_1154);
xor U1012 (N_1012,N_14,N_538);
nand U1013 (N_1013,In_396,In_1552);
and U1014 (N_1014,N_792,In_189);
nand U1015 (N_1015,N_489,In_1382);
or U1016 (N_1016,N_705,In_1365);
or U1017 (N_1017,In_1024,In_368);
nand U1018 (N_1018,N_913,N_376);
nor U1019 (N_1019,N_902,In_1090);
nand U1020 (N_1020,N_230,In_1184);
and U1021 (N_1021,N_927,In_1782);
xor U1022 (N_1022,In_1691,N_878);
xnor U1023 (N_1023,In_1864,N_337);
nor U1024 (N_1024,N_684,In_723);
nor U1025 (N_1025,N_261,In_1472);
nand U1026 (N_1026,N_844,In_1441);
and U1027 (N_1027,In_326,In_1808);
or U1028 (N_1028,N_910,In_53);
and U1029 (N_1029,N_222,N_661);
or U1030 (N_1030,N_915,N_621);
and U1031 (N_1031,N_541,N_363);
nor U1032 (N_1032,N_742,In_1178);
xor U1033 (N_1033,N_520,In_198);
and U1034 (N_1034,N_789,N_509);
nand U1035 (N_1035,N_654,N_727);
and U1036 (N_1036,In_329,N_491);
xor U1037 (N_1037,N_700,In_764);
nand U1038 (N_1038,In_791,In_543);
and U1039 (N_1039,In_522,N_290);
nand U1040 (N_1040,In_42,N_864);
nor U1041 (N_1041,In_529,N_325);
nor U1042 (N_1042,In_766,N_253);
nor U1043 (N_1043,In_1163,N_832);
xor U1044 (N_1044,In_737,In_1755);
and U1045 (N_1045,In_455,N_865);
and U1046 (N_1046,N_916,In_794);
xnor U1047 (N_1047,In_256,N_919);
xor U1048 (N_1048,In_1296,N_714);
and U1049 (N_1049,In_1043,N_96);
nand U1050 (N_1050,In_841,In_1497);
nand U1051 (N_1051,N_297,N_411);
or U1052 (N_1052,In_477,N_716);
nor U1053 (N_1053,N_522,N_388);
nand U1054 (N_1054,N_697,N_945);
xor U1055 (N_1055,In_853,In_1131);
and U1056 (N_1056,N_879,In_1589);
or U1057 (N_1057,In_1153,In_1308);
xor U1058 (N_1058,N_427,N_128);
nor U1059 (N_1059,In_1788,In_123);
nand U1060 (N_1060,In_1432,N_904);
nand U1061 (N_1061,In_211,N_599);
and U1062 (N_1062,In_71,In_592);
and U1063 (N_1063,In_1984,N_341);
or U1064 (N_1064,In_736,In_588);
xor U1065 (N_1065,N_69,N_643);
or U1066 (N_1066,In_922,In_433);
nor U1067 (N_1067,N_374,In_476);
or U1068 (N_1068,In_1650,In_1546);
or U1069 (N_1069,In_169,In_33);
or U1070 (N_1070,In_1654,In_1213);
and U1071 (N_1071,N_734,In_379);
xor U1072 (N_1072,N_36,N_457);
and U1073 (N_1073,N_485,In_1513);
xnor U1074 (N_1074,N_837,In_516);
nor U1075 (N_1075,N_918,In_1063);
and U1076 (N_1076,In_596,In_911);
and U1077 (N_1077,N_109,In_738);
nand U1078 (N_1078,N_928,In_1095);
or U1079 (N_1079,In_249,N_440);
nand U1080 (N_1080,N_568,In_1975);
xor U1081 (N_1081,In_1954,In_1040);
nand U1082 (N_1082,N_61,N_193);
or U1083 (N_1083,In_456,N_871);
xor U1084 (N_1084,In_1122,In_940);
and U1085 (N_1085,N_581,In_1463);
and U1086 (N_1086,N_333,N_519);
nand U1087 (N_1087,N_648,In_104);
nor U1088 (N_1088,N_539,In_1492);
nand U1089 (N_1089,In_669,N_778);
or U1090 (N_1090,N_821,N_731);
nor U1091 (N_1091,In_412,N_633);
and U1092 (N_1092,N_739,N_828);
xnor U1093 (N_1093,N_634,In_858);
nand U1094 (N_1094,In_1750,In_6);
and U1095 (N_1095,In_1148,N_224);
nor U1096 (N_1096,In_634,N_279);
nand U1097 (N_1097,In_119,N_773);
nand U1098 (N_1098,N_481,N_463);
xor U1099 (N_1099,N_874,In_820);
or U1100 (N_1100,In_939,In_930);
xnor U1101 (N_1101,N_11,N_362);
nand U1102 (N_1102,In_894,In_489);
or U1103 (N_1103,In_942,In_793);
nor U1104 (N_1104,N_958,In_122);
xnor U1105 (N_1105,In_825,N_574);
and U1106 (N_1106,In_667,N_378);
xnor U1107 (N_1107,N_136,In_1747);
or U1108 (N_1108,N_148,In_1705);
xnor U1109 (N_1109,In_944,In_1257);
and U1110 (N_1110,In_182,N_698);
or U1111 (N_1111,N_741,In_1683);
xnor U1112 (N_1112,In_1657,N_786);
nand U1113 (N_1113,N_595,N_125);
nor U1114 (N_1114,N_155,In_1916);
xnor U1115 (N_1115,In_1482,N_386);
nand U1116 (N_1116,N_266,N_326);
or U1117 (N_1117,In_1109,In_1057);
and U1118 (N_1118,In_458,In_1123);
nor U1119 (N_1119,N_642,N_433);
nand U1120 (N_1120,N_609,N_696);
or U1121 (N_1121,N_191,In_835);
and U1122 (N_1122,N_469,N_360);
or U1123 (N_1123,N_728,In_1088);
or U1124 (N_1124,In_99,N_1119);
and U1125 (N_1125,In_275,In_1373);
nor U1126 (N_1126,In_1100,N_823);
or U1127 (N_1127,N_1090,N_765);
nand U1128 (N_1128,N_1017,N_280);
or U1129 (N_1129,In_1265,In_1128);
nand U1130 (N_1130,N_806,N_729);
and U1131 (N_1131,N_192,N_1051);
xor U1132 (N_1132,N_379,In_1429);
xnor U1133 (N_1133,In_693,N_500);
or U1134 (N_1134,N_598,N_464);
nor U1135 (N_1135,N_1097,N_511);
xnor U1136 (N_1136,In_1668,In_181);
or U1137 (N_1137,In_85,In_1120);
nand U1138 (N_1138,In_886,N_999);
nand U1139 (N_1139,N_1109,N_271);
nand U1140 (N_1140,N_953,In_1284);
nor U1141 (N_1141,In_1915,In_925);
xnor U1142 (N_1142,In_220,In_1155);
nor U1143 (N_1143,N_751,N_544);
nor U1144 (N_1144,In_327,N_356);
nor U1145 (N_1145,N_816,N_862);
nor U1146 (N_1146,In_555,N_747);
nor U1147 (N_1147,N_756,In_1688);
or U1148 (N_1148,N_1038,N_854);
xor U1149 (N_1149,N_29,In_319);
and U1150 (N_1150,N_523,N_542);
and U1151 (N_1151,In_1564,N_996);
and U1152 (N_1152,N_442,In_1304);
nor U1153 (N_1153,N_1094,N_545);
nand U1154 (N_1154,In_590,N_985);
xnor U1155 (N_1155,N_830,In_1627);
nor U1156 (N_1156,N_820,N_373);
xor U1157 (N_1157,N_1050,In_1236);
xor U1158 (N_1158,In_759,In_1848);
and U1159 (N_1159,N_850,In_1199);
nor U1160 (N_1160,In_1017,N_502);
and U1161 (N_1161,N_930,N_204);
xnor U1162 (N_1162,In_1242,In_41);
nand U1163 (N_1163,In_656,In_937);
and U1164 (N_1164,N_421,In_558);
xor U1165 (N_1165,N_693,In_987);
and U1166 (N_1166,N_526,N_924);
and U1167 (N_1167,N_611,N_495);
nor U1168 (N_1168,In_749,In_977);
or U1169 (N_1169,In_1711,N_558);
nand U1170 (N_1170,In_1815,N_973);
nor U1171 (N_1171,In_162,N_657);
nand U1172 (N_1172,N_577,N_359);
and U1173 (N_1173,N_1002,N_1070);
or U1174 (N_1174,N_894,In_1032);
and U1175 (N_1175,In_1765,N_744);
nand U1176 (N_1176,In_301,N_703);
nor U1177 (N_1177,N_78,N_842);
and U1178 (N_1178,N_860,In_797);
and U1179 (N_1179,N_925,In_1208);
xnor U1180 (N_1180,N_493,N_540);
xnor U1181 (N_1181,N_73,In_1737);
or U1182 (N_1182,N_1067,N_735);
nor U1183 (N_1183,In_1301,N_525);
nor U1184 (N_1184,N_772,In_1769);
or U1185 (N_1185,In_648,N_767);
or U1186 (N_1186,N_944,N_977);
nor U1187 (N_1187,N_567,In_1893);
and U1188 (N_1188,N_701,N_1058);
and U1189 (N_1189,In_130,N_1001);
nand U1190 (N_1190,N_75,In_461);
and U1191 (N_1191,N_1096,In_1873);
or U1192 (N_1192,In_1931,N_498);
and U1193 (N_1193,In_302,N_550);
or U1194 (N_1194,N_227,In_81);
nand U1195 (N_1195,N_974,N_787);
and U1196 (N_1196,N_877,N_900);
and U1197 (N_1197,N_380,N_761);
xnor U1198 (N_1198,In_1006,In_266);
or U1199 (N_1199,In_1986,In_1743);
and U1200 (N_1200,In_1687,N_636);
nand U1201 (N_1201,In_1681,N_431);
or U1202 (N_1202,In_61,N_886);
or U1203 (N_1203,N_292,N_838);
nor U1204 (N_1204,In_1731,N_940);
nand U1205 (N_1205,In_1206,N_315);
nand U1206 (N_1206,N_839,N_929);
nor U1207 (N_1207,In_1321,N_355);
nand U1208 (N_1208,N_883,N_757);
xor U1209 (N_1209,In_1663,N_1069);
nor U1210 (N_1210,N_704,N_760);
or U1211 (N_1211,N_880,N_950);
xnor U1212 (N_1212,In_881,N_578);
or U1213 (N_1213,N_1031,N_738);
nand U1214 (N_1214,N_42,In_439);
and U1215 (N_1215,In_109,N_510);
nor U1216 (N_1216,N_1106,In_659);
or U1217 (N_1217,N_978,N_656);
nand U1218 (N_1218,In_1846,In_1775);
or U1219 (N_1219,In_804,N_943);
and U1220 (N_1220,N_889,N_407);
xnor U1221 (N_1221,In_1898,N_346);
nand U1222 (N_1222,In_1067,N_855);
nor U1223 (N_1223,N_972,In_1356);
or U1224 (N_1224,N_623,In_581);
xnor U1225 (N_1225,N_947,In_1874);
nor U1226 (N_1226,In_1028,In_1116);
nand U1227 (N_1227,N_482,N_652);
and U1228 (N_1228,N_1039,N_242);
nand U1229 (N_1229,N_299,In_1733);
nand U1230 (N_1230,In_638,In_542);
xor U1231 (N_1231,In_1785,N_691);
nand U1232 (N_1232,N_825,N_956);
nor U1233 (N_1233,In_1619,In_698);
and U1234 (N_1234,N_1007,In_1479);
xor U1235 (N_1235,In_426,N_895);
xor U1236 (N_1236,In_1704,In_861);
nor U1237 (N_1237,In_623,N_1100);
xnor U1238 (N_1238,N_1110,N_1101);
nand U1239 (N_1239,N_213,In_451);
or U1240 (N_1240,N_252,N_887);
and U1241 (N_1241,N_1071,N_1092);
nand U1242 (N_1242,In_520,In_1658);
nand U1243 (N_1243,In_1958,N_905);
xor U1244 (N_1244,In_140,In_1277);
and U1245 (N_1245,In_1160,In_1671);
or U1246 (N_1246,N_961,N_589);
nor U1247 (N_1247,N_1009,In_1549);
or U1248 (N_1248,N_1105,N_831);
xor U1249 (N_1249,N_962,In_1059);
nand U1250 (N_1250,In_972,In_1414);
or U1251 (N_1251,N_888,N_989);
and U1252 (N_1252,In_521,In_870);
nand U1253 (N_1253,In_120,In_988);
nand U1254 (N_1254,N_923,In_78);
nor U1255 (N_1255,N_840,N_771);
nand U1256 (N_1256,N_35,N_334);
xor U1257 (N_1257,N_131,N_1045);
xnor U1258 (N_1258,N_1010,N_34);
nand U1259 (N_1259,N_1068,N_770);
and U1260 (N_1260,In_155,N_1086);
or U1261 (N_1261,N_875,In_254);
xor U1262 (N_1262,N_800,N_826);
and U1263 (N_1263,N_984,In_1249);
or U1264 (N_1264,In_557,N_301);
or U1265 (N_1265,N_212,In_1794);
nand U1266 (N_1266,In_777,N_1065);
or U1267 (N_1267,N_1046,In_1335);
and U1268 (N_1268,N_1028,N_50);
and U1269 (N_1269,N_58,N_164);
and U1270 (N_1270,N_108,N_194);
nand U1271 (N_1271,N_105,N_1014);
nor U1272 (N_1272,N_979,N_1057);
and U1273 (N_1273,N_853,In_1625);
nor U1274 (N_1274,In_1352,In_1712);
nand U1275 (N_1275,N_437,N_576);
xnor U1276 (N_1276,N_404,In_128);
and U1277 (N_1277,In_560,N_320);
xor U1278 (N_1278,N_1042,In_1592);
nor U1279 (N_1279,N_810,N_813);
or U1280 (N_1280,N_55,N_4);
or U1281 (N_1281,N_935,N_851);
nor U1282 (N_1282,N_1161,N_1238);
nand U1283 (N_1283,N_1080,N_329);
nor U1284 (N_1284,N_1198,N_1208);
and U1285 (N_1285,In_402,N_1202);
xnor U1286 (N_1286,N_413,N_1267);
and U1287 (N_1287,In_1520,N_1081);
nor U1288 (N_1288,N_1089,N_1183);
xor U1289 (N_1289,N_1091,N_1074);
nand U1290 (N_1290,N_1254,N_876);
nor U1291 (N_1291,N_1193,In_324);
nand U1292 (N_1292,N_451,N_1118);
and U1293 (N_1293,N_665,N_1279);
or U1294 (N_1294,N_899,In_1049);
or U1295 (N_1295,N_675,N_720);
nand U1296 (N_1296,N_1248,N_980);
or U1297 (N_1297,In_1483,N_1251);
and U1298 (N_1298,In_491,In_787);
xnor U1299 (N_1299,N_639,N_1011);
or U1300 (N_1300,N_881,In_1406);
xor U1301 (N_1301,N_1229,N_1205);
nor U1302 (N_1302,N_782,In_632);
or U1303 (N_1303,N_1240,N_1224);
xnor U1304 (N_1304,N_1213,In_197);
or U1305 (N_1305,N_1196,In_1133);
nor U1306 (N_1306,In_1643,N_998);
and U1307 (N_1307,N_1135,N_1177);
xnor U1308 (N_1308,N_1232,N_53);
nand U1309 (N_1309,N_1197,In_463);
xnor U1310 (N_1310,N_1079,N_1130);
nand U1311 (N_1311,N_644,In_995);
nor U1312 (N_1312,N_799,In_258);
nand U1313 (N_1313,N_10,N_1150);
or U1314 (N_1314,N_841,In_440);
nor U1315 (N_1315,In_614,N_1114);
nor U1316 (N_1316,N_1163,In_1947);
nor U1317 (N_1317,N_939,N_1040);
and U1318 (N_1318,N_1262,N_1125);
xor U1319 (N_1319,In_1939,N_112);
nand U1320 (N_1320,N_1060,In_432);
or U1321 (N_1321,N_687,N_1021);
nor U1322 (N_1322,N_781,N_1148);
or U1323 (N_1323,In_1696,N_1004);
and U1324 (N_1324,N_209,N_1066);
or U1325 (N_1325,N_686,In_819);
nand U1326 (N_1326,In_405,In_343);
nand U1327 (N_1327,N_1128,N_560);
nand U1328 (N_1328,N_1049,In_1885);
nor U1329 (N_1329,In_334,In_1458);
and U1330 (N_1330,In_1632,N_920);
xor U1331 (N_1331,N_682,N_835);
nand U1332 (N_1332,N_903,N_827);
nor U1333 (N_1333,N_1250,In_1031);
or U1334 (N_1334,N_952,N_1180);
and U1335 (N_1335,N_468,N_836);
and U1336 (N_1336,In_1436,N_1054);
or U1337 (N_1337,N_1030,N_70);
nand U1338 (N_1338,N_466,In_772);
nor U1339 (N_1339,In_431,N_287);
nor U1340 (N_1340,N_1273,N_1003);
xor U1341 (N_1341,N_679,N_946);
and U1342 (N_1342,N_970,N_650);
or U1343 (N_1343,N_1024,N_1033);
or U1344 (N_1344,N_1237,N_1036);
xor U1345 (N_1345,N_335,N_852);
nand U1346 (N_1346,N_808,N_1158);
or U1347 (N_1347,In_646,N_976);
xnor U1348 (N_1348,N_448,N_1129);
nor U1349 (N_1349,N_1176,N_814);
or U1350 (N_1350,In_704,N_848);
and U1351 (N_1351,N_1020,In_1390);
nand U1352 (N_1352,N_1152,In_1126);
nor U1353 (N_1353,In_1812,N_1195);
and U1354 (N_1354,N_1063,N_1173);
and U1355 (N_1355,In_478,In_1021);
and U1356 (N_1356,N_1243,N_1244);
or U1357 (N_1357,N_1027,In_735);
nand U1358 (N_1358,N_483,In_1596);
nor U1359 (N_1359,N_794,N_699);
nor U1360 (N_1360,N_1225,N_1189);
nor U1361 (N_1361,N_1055,N_256);
nor U1362 (N_1362,In_983,N_1276);
or U1363 (N_1363,In_1538,In_1216);
and U1364 (N_1364,In_1144,In_101);
nor U1365 (N_1365,In_403,N_1137);
or U1366 (N_1366,N_1082,N_1235);
nand U1367 (N_1367,N_1192,N_951);
and U1368 (N_1368,N_882,In_849);
and U1369 (N_1369,N_949,N_631);
xor U1370 (N_1370,In_1568,In_199);
xnor U1371 (N_1371,N_907,N_1005);
nor U1372 (N_1372,In_364,N_1167);
or U1373 (N_1373,In_1577,N_740);
nand U1374 (N_1374,N_891,N_207);
or U1375 (N_1375,In_1653,N_1190);
xor U1376 (N_1376,N_169,In_1616);
and U1377 (N_1377,N_490,N_1034);
nor U1378 (N_1378,In_1752,In_1814);
or U1379 (N_1379,N_165,N_393);
and U1380 (N_1380,N_1120,N_1000);
nand U1381 (N_1381,In_14,N_152);
nand U1382 (N_1382,N_1154,N_101);
nor U1383 (N_1383,N_1093,N_1239);
xnor U1384 (N_1384,N_1241,In_1921);
and U1385 (N_1385,N_957,N_646);
nor U1386 (N_1386,N_1187,N_1217);
nand U1387 (N_1387,N_1052,N_869);
nand U1388 (N_1388,N_677,In_826);
xor U1389 (N_1389,N_103,N_1061);
nor U1390 (N_1390,N_805,N_1191);
and U1391 (N_1391,N_863,N_1278);
xor U1392 (N_1392,N_1157,N_494);
or U1393 (N_1393,In_1081,N_834);
and U1394 (N_1394,N_370,In_1060);
xnor U1395 (N_1395,N_246,N_559);
nand U1396 (N_1396,N_575,N_1162);
or U1397 (N_1397,N_1168,N_119);
or U1398 (N_1398,In_374,In_1901);
nand U1399 (N_1399,In_796,N_694);
or U1400 (N_1400,N_1008,In_1234);
or U1401 (N_1401,In_1924,N_1136);
xor U1402 (N_1402,N_1149,N_1041);
xor U1403 (N_1403,N_97,N_1221);
and U1404 (N_1404,N_1134,N_1083);
nor U1405 (N_1405,N_802,N_1078);
and U1406 (N_1406,N_783,In_530);
and U1407 (N_1407,N_425,In_1829);
or U1408 (N_1408,N_983,N_868);
nor U1409 (N_1409,N_1223,N_678);
or U1410 (N_1410,N_603,N_1006);
nand U1411 (N_1411,N_755,In_824);
xor U1412 (N_1412,N_1246,In_116);
and U1413 (N_1413,In_943,N_843);
and U1414 (N_1414,In_914,In_87);
or U1415 (N_1415,N_543,N_340);
nor U1416 (N_1416,N_911,In_401);
or U1417 (N_1417,N_1104,N_1077);
or U1418 (N_1418,In_0,N_909);
xnor U1419 (N_1419,N_803,N_938);
and U1420 (N_1420,In_479,N_1132);
or U1421 (N_1421,N_758,In_1076);
xor U1422 (N_1422,N_515,N_959);
xor U1423 (N_1423,N_248,N_960);
nor U1424 (N_1424,N_745,N_637);
xnor U1425 (N_1425,In_34,N_1085);
or U1426 (N_1426,N_967,N_1220);
nor U1427 (N_1427,N_1037,N_937);
nor U1428 (N_1428,In_205,N_1075);
xor U1429 (N_1429,N_1147,In_1004);
or U1430 (N_1430,N_546,N_1143);
nor U1431 (N_1431,In_225,In_1244);
and U1432 (N_1432,In_317,N_1088);
nor U1433 (N_1433,N_1206,N_870);
or U1434 (N_1434,N_1146,N_364);
or U1435 (N_1435,N_965,N_649);
and U1436 (N_1436,N_1259,N_1214);
nor U1437 (N_1437,In_1754,In_65);
xnor U1438 (N_1438,N_15,In_1239);
and U1439 (N_1439,N_200,N_122);
nor U1440 (N_1440,N_1122,N_1292);
or U1441 (N_1441,In_441,N_673);
or U1442 (N_1442,N_1102,N_367);
or U1443 (N_1443,N_98,N_1338);
nor U1444 (N_1444,N_664,N_1347);
xnor U1445 (N_1445,N_1431,N_1419);
nand U1446 (N_1446,N_906,In_1018);
or U1447 (N_1447,N_1164,N_72);
nor U1448 (N_1448,N_1182,N_1399);
or U1449 (N_1449,In_1420,N_658);
and U1450 (N_1450,N_764,N_1062);
nor U1451 (N_1451,N_1178,N_371);
nand U1452 (N_1452,N_1266,N_1286);
or U1453 (N_1453,N_1326,In_1968);
nor U1454 (N_1454,N_1282,N_49);
xnor U1455 (N_1455,In_32,In_813);
nand U1456 (N_1456,N_1207,In_159);
and U1457 (N_1457,N_1159,N_1295);
xor U1458 (N_1458,In_732,N_1321);
xor U1459 (N_1459,N_754,N_1123);
nand U1460 (N_1460,N_645,In_1530);
xor U1461 (N_1461,N_1421,N_1059);
nand U1462 (N_1462,In_66,In_369);
or U1463 (N_1463,N_535,In_713);
or U1464 (N_1464,In_1756,N_1376);
or U1465 (N_1465,N_670,N_1290);
or U1466 (N_1466,N_514,N_1412);
xor U1467 (N_1467,In_1656,In_898);
or U1468 (N_1468,N_1218,In_1108);
nor U1469 (N_1469,N_859,N_796);
or U1470 (N_1470,N_873,N_1381);
nor U1471 (N_1471,N_321,N_1437);
or U1472 (N_1472,N_721,N_1255);
or U1473 (N_1473,N_809,In_1409);
xnor U1474 (N_1474,N_1349,N_1404);
nand U1475 (N_1475,N_1138,N_1379);
or U1476 (N_1476,N_552,N_1160);
nand U1477 (N_1477,N_135,N_1098);
nand U1478 (N_1478,N_1409,N_964);
and U1479 (N_1479,In_1243,N_1099);
nor U1480 (N_1480,N_240,In_1689);
and U1481 (N_1481,N_954,N_182);
nor U1482 (N_1482,N_1116,N_123);
nor U1483 (N_1483,N_1056,N_304);
nor U1484 (N_1484,In_966,N_1258);
xnor U1485 (N_1485,N_1289,N_1139);
nand U1486 (N_1486,N_941,N_1185);
xor U1487 (N_1487,N_615,In_1298);
and U1488 (N_1488,N_708,N_1043);
or U1489 (N_1489,In_1185,N_1407);
or U1490 (N_1490,N_1300,In_931);
xor U1491 (N_1491,N_1212,N_1385);
nand U1492 (N_1492,N_478,N_1414);
nand U1493 (N_1493,In_1026,N_418);
xnor U1494 (N_1494,In_1541,N_1126);
nor U1495 (N_1495,N_1253,N_1332);
xnor U1496 (N_1496,In_687,N_1417);
nand U1497 (N_1497,In_1285,N_1144);
nor U1498 (N_1498,N_1352,N_1336);
or U1499 (N_1499,N_750,N_1303);
xor U1500 (N_1500,In_1054,N_752);
nand U1501 (N_1501,N_1402,N_521);
or U1502 (N_1502,N_1319,In_910);
or U1503 (N_1503,N_1272,N_171);
and U1504 (N_1504,In_1399,N_1174);
nor U1505 (N_1505,N_1142,N_1287);
xor U1506 (N_1506,In_1344,N_1277);
xor U1507 (N_1507,N_1400,N_1307);
or U1508 (N_1508,N_429,In_1830);
xor U1509 (N_1509,N_1423,N_1297);
and U1510 (N_1510,N_1335,N_582);
xnor U1511 (N_1511,N_1345,In_1501);
and U1512 (N_1512,In_1179,N_981);
or U1513 (N_1513,N_975,N_1181);
and U1514 (N_1514,N_815,N_1401);
nand U1515 (N_1515,N_1231,N_715);
and U1516 (N_1516,N_1166,N_1264);
or U1517 (N_1517,N_689,N_389);
or U1518 (N_1518,N_381,In_217);
xnor U1519 (N_1519,N_1302,N_1023);
xnor U1520 (N_1520,N_1179,N_254);
xor U1521 (N_1521,N_1438,In_526);
nor U1522 (N_1522,N_467,N_641);
or U1523 (N_1523,N_1245,N_1234);
nand U1524 (N_1524,N_1354,N_997);
or U1525 (N_1525,N_1357,In_1886);
nand U1526 (N_1526,N_804,In_722);
nand U1527 (N_1527,N_1350,N_753);
or U1528 (N_1528,N_1200,N_1124);
nor U1529 (N_1529,In_1477,N_1382);
xnor U1530 (N_1530,N_1351,N_1151);
or U1531 (N_1531,In_1764,In_1693);
nand U1532 (N_1532,N_1029,N_723);
or U1533 (N_1533,N_1084,N_1340);
and U1534 (N_1534,In_1995,N_1211);
or U1535 (N_1535,N_1170,N_1247);
and U1536 (N_1536,N_1439,In_45);
nor U1537 (N_1537,N_791,N_1342);
or U1538 (N_1538,N_1209,N_884);
nand U1539 (N_1539,N_1064,N_896);
xnor U1540 (N_1540,N_1398,In_1649);
nand U1541 (N_1541,N_1425,N_462);
xor U1542 (N_1542,N_817,N_866);
or U1543 (N_1543,N_991,N_987);
nor U1544 (N_1544,N_1230,N_982);
nand U1545 (N_1545,In_1526,N_1366);
nand U1546 (N_1546,N_1271,N_1107);
nand U1547 (N_1547,N_1432,N_901);
or U1548 (N_1548,In_541,N_1219);
nor U1549 (N_1549,N_1044,N_1330);
and U1550 (N_1550,N_1072,N_1328);
nor U1551 (N_1551,N_1265,N_1397);
or U1552 (N_1552,N_824,N_1314);
xor U1553 (N_1553,N_1344,In_928);
xor U1554 (N_1554,N_1194,In_1293);
and U1555 (N_1555,N_1018,N_1308);
nor U1556 (N_1556,In_213,In_406);
xnor U1557 (N_1557,N_420,N_307);
nand U1558 (N_1558,N_819,N_1296);
or U1559 (N_1559,In_1710,N_172);
and U1560 (N_1560,In_902,N_1413);
xnor U1561 (N_1561,N_795,In_731);
nor U1562 (N_1562,N_1053,In_1845);
nor U1563 (N_1563,N_513,N_1315);
xnor U1564 (N_1564,N_737,N_1012);
or U1565 (N_1565,N_857,N_1371);
nand U1566 (N_1566,N_1184,N_1370);
nand U1567 (N_1567,In_658,In_1474);
and U1568 (N_1568,N_1121,N_1233);
nand U1569 (N_1569,In_1157,N_1216);
or U1570 (N_1570,N_1171,In_683);
xor U1571 (N_1571,In_1379,In_1396);
xnor U1572 (N_1572,N_766,N_48);
or U1573 (N_1573,N_1141,N_1016);
xnor U1574 (N_1574,In_68,N_569);
and U1575 (N_1575,In_1459,In_1189);
nand U1576 (N_1576,In_934,In_1780);
and U1577 (N_1577,N_793,In_1867);
nor U1578 (N_1578,N_203,N_1406);
or U1579 (N_1579,In_1651,N_1426);
or U1580 (N_1580,N_807,N_353);
and U1581 (N_1581,N_1363,N_1257);
nor U1582 (N_1582,N_1383,N_372);
nand U1583 (N_1583,N_1334,N_143);
and U1584 (N_1584,N_1108,In_1210);
xnor U1585 (N_1585,N_932,In_1008);
nand U1586 (N_1586,N_518,N_1390);
nor U1587 (N_1587,N_995,N_1204);
and U1588 (N_1588,N_988,N_1372);
xor U1589 (N_1589,In_1050,N_1384);
nor U1590 (N_1590,N_1429,N_1377);
or U1591 (N_1591,N_846,In_1083);
nor U1592 (N_1592,In_679,N_1133);
xnor U1593 (N_1593,N_1320,N_1285);
or U1594 (N_1594,N_1396,N_1284);
and U1595 (N_1595,N_1387,N_1201);
nand U1596 (N_1596,N_1294,N_858);
or U1597 (N_1597,N_1269,N_470);
and U1598 (N_1598,N_1117,N_861);
or U1599 (N_1599,N_1435,N_829);
or U1600 (N_1600,N_1153,N_1252);
or U1601 (N_1601,In_1978,N_1445);
nand U1602 (N_1602,N_801,N_1508);
nand U1603 (N_1603,N_1015,N_1567);
xnor U1604 (N_1604,N_309,N_1562);
xor U1605 (N_1605,N_1365,N_1403);
nor U1606 (N_1606,N_1422,N_1480);
nand U1607 (N_1607,In_770,N_1323);
nand U1608 (N_1608,In_55,N_931);
or U1609 (N_1609,In_29,N_1468);
or U1610 (N_1610,N_1156,N_1581);
xor U1611 (N_1611,N_1364,In_132);
nand U1612 (N_1612,N_1465,In_1448);
nand U1613 (N_1613,N_1293,In_1730);
nand U1614 (N_1614,N_1509,N_1518);
nand U1615 (N_1615,N_1550,N_1496);
nor U1616 (N_1616,N_994,N_1433);
xor U1617 (N_1617,N_1593,N_942);
nor U1618 (N_1618,N_1561,N_1578);
xnor U1619 (N_1619,In_1025,N_1448);
and U1620 (N_1620,N_1533,N_1270);
and U1621 (N_1621,N_1543,N_1458);
or U1622 (N_1622,N_992,N_1513);
nand U1623 (N_1623,N_1467,N_1275);
or U1624 (N_1624,N_845,N_1405);
and U1625 (N_1625,N_1501,N_1327);
nor U1626 (N_1626,N_185,N_1488);
and U1627 (N_1627,N_1486,N_1483);
xor U1628 (N_1628,N_1579,N_1484);
or U1629 (N_1629,N_1476,N_1242);
xnor U1630 (N_1630,N_1316,N_1313);
xor U1631 (N_1631,N_1510,N_1298);
xnor U1632 (N_1632,N_1460,In_622);
xnor U1633 (N_1633,In_1495,N_1362);
or U1634 (N_1634,N_1443,N_1359);
nand U1635 (N_1635,N_444,N_1353);
nand U1636 (N_1636,N_1280,N_1495);
nand U1637 (N_1637,N_1536,N_241);
and U1638 (N_1638,N_1115,N_1199);
and U1639 (N_1639,N_1544,N_1459);
nand U1640 (N_1640,N_1331,N_872);
nor U1641 (N_1641,N_1268,N_1474);
nand U1642 (N_1642,N_1203,N_1585);
nor U1643 (N_1643,In_933,N_1022);
nand U1644 (N_1644,N_1457,N_1595);
and U1645 (N_1645,N_1369,In_392);
nand U1646 (N_1646,N_1535,In_1267);
or U1647 (N_1647,In_1970,N_1519);
xor U1648 (N_1648,N_1380,N_503);
nand U1649 (N_1649,N_1591,N_1337);
and U1650 (N_1650,In_49,In_1084);
nand U1651 (N_1651,N_1583,N_161);
or U1652 (N_1652,N_1322,N_1317);
nor U1653 (N_1653,N_1343,N_1589);
or U1654 (N_1654,N_926,N_532);
or U1655 (N_1655,N_1261,In_724);
and U1656 (N_1656,In_73,N_762);
xor U1657 (N_1657,N_1538,N_1512);
xnor U1658 (N_1658,N_724,N_1442);
or U1659 (N_1659,N_1288,N_1594);
nor U1660 (N_1660,N_966,In_268);
nor U1661 (N_1661,N_554,N_1073);
or U1662 (N_1662,N_1545,N_1348);
xor U1663 (N_1663,In_583,N_1528);
nor U1664 (N_1664,N_971,In_239);
or U1665 (N_1665,N_1392,N_1227);
xor U1666 (N_1666,N_1569,N_1524);
nor U1667 (N_1667,N_1522,N_1568);
xnor U1668 (N_1668,N_1339,In_1827);
and U1669 (N_1669,N_1514,N_1103);
xor U1670 (N_1670,N_1358,In_1529);
and U1671 (N_1671,N_1534,N_1582);
or U1672 (N_1672,N_1441,N_1304);
nor U1673 (N_1673,N_1140,N_1440);
nor U1674 (N_1674,N_1175,N_1580);
nand U1675 (N_1675,N_1222,N_1450);
and U1676 (N_1676,N_1573,N_1575);
xor U1677 (N_1677,N_1471,N_1549);
xor U1678 (N_1678,N_1333,N_1375);
xnor U1679 (N_1679,N_1542,N_1418);
nor U1680 (N_1680,In_830,N_1479);
or U1681 (N_1681,N_1517,In_437);
or U1682 (N_1682,N_847,N_1490);
nor U1683 (N_1683,N_1539,N_1145);
and U1684 (N_1684,N_1299,N_1306);
or U1685 (N_1685,N_588,N_1572);
nand U1686 (N_1686,N_1494,N_517);
or U1687 (N_1687,N_897,N_1599);
nand U1688 (N_1688,In_10,N_1449);
xnor U1689 (N_1689,In_37,In_635);
or U1690 (N_1690,N_1428,N_1032);
and U1691 (N_1691,N_718,N_1415);
and U1692 (N_1692,N_1493,In_840);
nor U1693 (N_1693,N_1368,In_1753);
xnor U1694 (N_1694,N_1455,N_1311);
xor U1695 (N_1695,N_1360,N_146);
nor U1696 (N_1696,N_1047,N_893);
xnor U1697 (N_1697,N_1527,N_1525);
nand U1698 (N_1698,N_1447,N_1095);
nor U1699 (N_1699,N_1558,N_1436);
nand U1700 (N_1700,In_1741,In_1723);
nand U1701 (N_1701,N_1236,In_741);
nor U1702 (N_1702,In_1950,N_1389);
nor U1703 (N_1703,N_1587,N_1420);
xnor U1704 (N_1704,N_1408,N_1111);
nor U1705 (N_1705,N_1546,N_1453);
nor U1706 (N_1706,In_1518,N_1013);
or U1707 (N_1707,N_1552,N_1592);
and U1708 (N_1708,N_1215,N_1274);
xor U1709 (N_1709,N_1391,N_1019);
nand U1710 (N_1710,N_1557,N_1491);
nand U1711 (N_1711,N_1410,N_1521);
nor U1712 (N_1712,N_1256,N_1131);
nor U1713 (N_1713,N_1388,N_1025);
xor U1714 (N_1714,N_1548,N_1035);
or U1715 (N_1715,N_1565,N_1260);
nand U1716 (N_1716,N_1547,N_1263);
nor U1717 (N_1717,N_1464,N_1394);
and U1718 (N_1718,N_1374,N_1430);
xnor U1719 (N_1719,N_1540,N_969);
nand U1720 (N_1720,N_968,N_1511);
nand U1721 (N_1721,N_1596,In_903);
nor U1722 (N_1722,In_1565,N_1165);
nor U1723 (N_1723,N_1588,N_1411);
nand U1724 (N_1724,N_1466,N_1434);
xnor U1725 (N_1725,N_1507,N_1461);
nand U1726 (N_1726,In_237,N_1470);
xnor U1727 (N_1727,N_1598,N_1427);
xor U1728 (N_1728,N_1487,N_533);
or U1729 (N_1729,N_1566,In_908);
and U1730 (N_1730,N_1577,N_1462);
xor U1731 (N_1731,In_1823,N_264);
xor U1732 (N_1732,N_1532,N_1463);
nand U1733 (N_1733,N_1186,N_1324);
or U1734 (N_1734,N_1169,N_1473);
and U1735 (N_1735,In_730,N_1472);
and U1736 (N_1736,N_1386,N_338);
and U1737 (N_1737,N_1451,N_1485);
nor U1738 (N_1738,N_504,N_1452);
nor U1739 (N_1739,In_1106,N_1502);
xnor U1740 (N_1740,N_1341,N_1393);
or U1741 (N_1741,N_1556,N_1444);
and U1742 (N_1742,N_1481,N_1226);
nand U1743 (N_1743,N_1560,N_1482);
nor U1744 (N_1744,N_1559,In_1205);
xnor U1745 (N_1745,N_1492,N_948);
nor U1746 (N_1746,N_963,N_993);
xnor U1747 (N_1747,N_955,N_1515);
and U1748 (N_1748,N_1489,N_730);
or U1749 (N_1749,N_1499,N_986);
nand U1750 (N_1750,N_1475,N_1318);
nand U1751 (N_1751,N_1361,N_1570);
nand U1752 (N_1752,N_1597,N_1586);
nand U1753 (N_1753,N_1541,N_1188);
nor U1754 (N_1754,N_349,N_990);
nor U1755 (N_1755,N_1503,In_22);
nor U1756 (N_1756,N_818,N_1574);
nor U1757 (N_1757,N_1564,N_1530);
nor U1758 (N_1758,N_1505,N_1172);
xnor U1759 (N_1759,N_1249,N_1500);
or U1760 (N_1760,N_1639,N_1701);
xor U1761 (N_1761,N_1623,In_346);
nor U1762 (N_1762,N_1714,N_1661);
and U1763 (N_1763,N_258,N_921);
or U1764 (N_1764,N_1529,N_1076);
nand U1765 (N_1765,N_1621,N_1506);
or U1766 (N_1766,N_1715,N_1367);
or U1767 (N_1767,N_1692,N_1708);
xnor U1768 (N_1768,N_1355,N_1378);
or U1769 (N_1769,N_1728,N_1590);
nand U1770 (N_1770,N_1609,N_1456);
or U1771 (N_1771,N_683,In_388);
and U1772 (N_1772,N_1716,N_936);
nand U1773 (N_1773,N_1753,N_1671);
or U1774 (N_1774,N_1697,N_1283);
nor U1775 (N_1775,N_1659,N_1622);
or U1776 (N_1776,N_1416,N_1497);
and U1777 (N_1777,N_1696,N_1633);
or U1778 (N_1778,N_1676,N_1624);
nor U1779 (N_1779,N_856,N_1691);
xnor U1780 (N_1780,N_1758,N_1618);
xnor U1781 (N_1781,N_1674,N_1210);
nor U1782 (N_1782,N_1611,N_1744);
nor U1783 (N_1783,N_1739,N_1601);
and U1784 (N_1784,N_1640,N_1608);
nor U1785 (N_1785,N_1720,In_525);
xnor U1786 (N_1786,N_1722,N_1632);
nand U1787 (N_1787,N_1638,In_740);
and U1788 (N_1788,N_640,N_1710);
nand U1789 (N_1789,N_1698,N_1620);
or U1790 (N_1790,N_1757,N_1755);
xor U1791 (N_1791,N_1685,N_1663);
xor U1792 (N_1792,In_1056,N_1395);
or U1793 (N_1793,N_1660,N_1733);
nor U1794 (N_1794,N_1329,N_1662);
nand U1795 (N_1795,N_1651,N_1026);
or U1796 (N_1796,N_1713,N_1644);
nor U1797 (N_1797,N_1703,N_1686);
and U1798 (N_1798,N_1738,N_1325);
or U1799 (N_1799,N_1615,N_709);
nand U1800 (N_1800,N_1523,N_1649);
and U1801 (N_1801,N_1643,N_1673);
and U1802 (N_1802,N_1301,N_566);
nor U1803 (N_1803,N_1571,N_1127);
nand U1804 (N_1804,N_1756,N_1048);
nor U1805 (N_1805,N_1725,N_1747);
and U1806 (N_1806,N_1666,N_1576);
and U1807 (N_1807,N_1682,N_1610);
nand U1808 (N_1808,N_1678,N_1498);
and U1809 (N_1809,N_1729,N_1356);
and U1810 (N_1810,N_499,N_1625);
xor U1811 (N_1811,N_1469,N_1658);
nor U1812 (N_1812,N_1600,N_1746);
nor U1813 (N_1813,N_1631,N_1630);
or U1814 (N_1814,N_1749,N_1635);
and U1815 (N_1815,N_1113,N_1646);
or U1816 (N_1816,N_1687,N_1705);
or U1817 (N_1817,N_1668,N_1641);
and U1818 (N_1818,N_1653,In_1449);
nor U1819 (N_1819,N_1626,N_1684);
nand U1820 (N_1820,N_1604,N_1712);
or U1821 (N_1821,N_1584,N_1667);
or U1822 (N_1822,N_1657,N_1717);
nand U1823 (N_1823,N_1735,N_1748);
or U1824 (N_1824,N_1637,N_1677);
xor U1825 (N_1825,N_1628,N_1726);
nor U1826 (N_1826,N_1634,N_1740);
nor U1827 (N_1827,N_1724,N_1612);
nor U1828 (N_1828,N_1723,N_1614);
nor U1829 (N_1829,N_1695,N_1478);
or U1830 (N_1830,N_1754,In_465);
nor U1831 (N_1831,N_1424,N_1636);
xor U1832 (N_1832,N_1629,N_1605);
nor U1833 (N_1833,N_1616,N_1537);
nor U1834 (N_1834,N_1750,N_1759);
and U1835 (N_1835,N_1656,N_1155);
nor U1836 (N_1836,N_1718,N_1732);
xnor U1837 (N_1837,N_1642,N_1690);
nor U1838 (N_1838,N_1606,N_1309);
xor U1839 (N_1839,N_1617,N_547);
nand U1840 (N_1840,N_1680,N_1373);
nor U1841 (N_1841,N_1291,N_1699);
or U1842 (N_1842,N_1709,N_1702);
nor U1843 (N_1843,N_1688,N_1719);
and U1844 (N_1844,N_1664,N_1520);
or U1845 (N_1845,In_798,N_1737);
nor U1846 (N_1846,N_1669,N_1689);
xnor U1847 (N_1847,N_1553,N_1736);
and U1848 (N_1848,N_1446,N_1312);
and U1849 (N_1849,N_1087,N_1281);
xor U1850 (N_1850,N_1310,N_1454);
nand U1851 (N_1851,N_1675,N_1665);
nor U1852 (N_1852,N_1652,N_1711);
and U1853 (N_1853,N_1504,N_933);
and U1854 (N_1854,N_1693,N_1516);
xor U1855 (N_1855,N_1305,N_1707);
xor U1856 (N_1856,N_1563,In_447);
nand U1857 (N_1857,N_1602,N_1645);
or U1858 (N_1858,N_1551,N_1477);
nor U1859 (N_1859,N_1679,N_1554);
xor U1860 (N_1860,N_1706,N_1742);
nand U1861 (N_1861,N_1613,N_1655);
nand U1862 (N_1862,N_1730,N_1727);
nor U1863 (N_1863,N_1741,N_556);
nand U1864 (N_1864,N_1731,N_1721);
or U1865 (N_1865,N_1603,N_1751);
xor U1866 (N_1866,N_1700,N_1648);
nand U1867 (N_1867,N_1112,N_1734);
nand U1868 (N_1868,N_1526,N_1672);
or U1869 (N_1869,N_1681,N_1650);
and U1870 (N_1870,N_1745,N_1683);
nand U1871 (N_1871,N_1619,N_1752);
nand U1872 (N_1872,In_404,N_759);
nor U1873 (N_1873,N_1704,N_867);
or U1874 (N_1874,N_1627,N_1607);
or U1875 (N_1875,N_1346,N_1228);
or U1876 (N_1876,N_1694,N_1647);
xor U1877 (N_1877,N_1531,N_1743);
nor U1878 (N_1878,N_1654,N_1670);
nand U1879 (N_1879,In_1187,N_1555);
or U1880 (N_1880,N_1750,N_1699);
or U1881 (N_1881,N_1726,N_1724);
or U1882 (N_1882,N_867,N_1737);
or U1883 (N_1883,N_921,N_1684);
nand U1884 (N_1884,N_1720,N_1711);
and U1885 (N_1885,N_1738,N_1603);
nand U1886 (N_1886,N_1702,N_1736);
xor U1887 (N_1887,N_640,N_1704);
and U1888 (N_1888,N_1620,N_1730);
and U1889 (N_1889,N_1662,N_1751);
nand U1890 (N_1890,N_1454,N_1571);
nor U1891 (N_1891,N_1690,N_1655);
or U1892 (N_1892,N_1611,N_1614);
xor U1893 (N_1893,N_1721,N_1291);
nor U1894 (N_1894,N_1694,In_447);
nand U1895 (N_1895,N_1087,N_1642);
and U1896 (N_1896,N_1646,N_1708);
or U1897 (N_1897,N_1309,N_1620);
xnor U1898 (N_1898,N_1754,N_1692);
nand U1899 (N_1899,N_1757,N_1669);
xnor U1900 (N_1900,N_1625,N_1626);
or U1901 (N_1901,N_1696,N_1681);
xnor U1902 (N_1902,N_1613,In_798);
nor U1903 (N_1903,N_1614,N_1755);
nor U1904 (N_1904,N_1416,N_1756);
nand U1905 (N_1905,N_683,N_1650);
xor U1906 (N_1906,N_566,N_1706);
nor U1907 (N_1907,N_1416,N_1621);
and U1908 (N_1908,N_1424,N_1687);
and U1909 (N_1909,N_1633,N_1683);
or U1910 (N_1910,N_1755,N_1749);
nor U1911 (N_1911,N_1689,N_1667);
or U1912 (N_1912,N_1731,N_1647);
nor U1913 (N_1913,N_1703,N_566);
nor U1914 (N_1914,N_1705,N_1609);
or U1915 (N_1915,N_1723,In_404);
nand U1916 (N_1916,N_1424,N_1656);
or U1917 (N_1917,N_1684,N_1687);
xnor U1918 (N_1918,N_1291,N_1677);
xnor U1919 (N_1919,N_258,N_640);
nand U1920 (N_1920,N_1893,N_1811);
xnor U1921 (N_1921,N_1854,N_1883);
nor U1922 (N_1922,N_1888,N_1886);
and U1923 (N_1923,N_1802,N_1859);
and U1924 (N_1924,N_1774,N_1798);
or U1925 (N_1925,N_1837,N_1917);
nor U1926 (N_1926,N_1861,N_1875);
nand U1927 (N_1927,N_1773,N_1817);
nand U1928 (N_1928,N_1789,N_1918);
nand U1929 (N_1929,N_1842,N_1795);
xor U1930 (N_1930,N_1783,N_1806);
nor U1931 (N_1931,N_1819,N_1770);
nand U1932 (N_1932,N_1782,N_1838);
nor U1933 (N_1933,N_1906,N_1820);
or U1934 (N_1934,N_1829,N_1801);
and U1935 (N_1935,N_1902,N_1821);
nor U1936 (N_1936,N_1777,N_1912);
and U1937 (N_1937,N_1824,N_1813);
or U1938 (N_1938,N_1788,N_1855);
nor U1939 (N_1939,N_1803,N_1775);
xor U1940 (N_1940,N_1852,N_1863);
nand U1941 (N_1941,N_1841,N_1907);
or U1942 (N_1942,N_1772,N_1884);
nand U1943 (N_1943,N_1786,N_1908);
nand U1944 (N_1944,N_1849,N_1816);
nor U1945 (N_1945,N_1919,N_1810);
and U1946 (N_1946,N_1878,N_1891);
xnor U1947 (N_1947,N_1840,N_1911);
and U1948 (N_1948,N_1763,N_1784);
nand U1949 (N_1949,N_1880,N_1808);
nand U1950 (N_1950,N_1851,N_1887);
or U1951 (N_1951,N_1885,N_1792);
and U1952 (N_1952,N_1867,N_1881);
and U1953 (N_1953,N_1853,N_1876);
nor U1954 (N_1954,N_1901,N_1909);
or U1955 (N_1955,N_1903,N_1780);
xor U1956 (N_1956,N_1761,N_1866);
or U1957 (N_1957,N_1825,N_1769);
nand U1958 (N_1958,N_1896,N_1860);
and U1959 (N_1959,N_1843,N_1815);
or U1960 (N_1960,N_1895,N_1762);
nand U1961 (N_1961,N_1828,N_1915);
nand U1962 (N_1962,N_1832,N_1799);
or U1963 (N_1963,N_1862,N_1882);
or U1964 (N_1964,N_1847,N_1812);
and U1965 (N_1965,N_1776,N_1796);
nand U1966 (N_1966,N_1794,N_1916);
or U1967 (N_1967,N_1899,N_1823);
and U1968 (N_1968,N_1864,N_1913);
nand U1969 (N_1969,N_1850,N_1848);
or U1970 (N_1970,N_1904,N_1768);
xnor U1971 (N_1971,N_1897,N_1830);
or U1972 (N_1972,N_1809,N_1834);
nand U1973 (N_1973,N_1839,N_1800);
and U1974 (N_1974,N_1857,N_1833);
xor U1975 (N_1975,N_1890,N_1807);
or U1976 (N_1976,N_1845,N_1791);
and U1977 (N_1977,N_1826,N_1804);
nor U1978 (N_1978,N_1785,N_1892);
nand U1979 (N_1979,N_1844,N_1835);
nor U1980 (N_1980,N_1778,N_1831);
nor U1981 (N_1981,N_1894,N_1879);
nand U1982 (N_1982,N_1900,N_1873);
xor U1983 (N_1983,N_1781,N_1771);
or U1984 (N_1984,N_1797,N_1805);
or U1985 (N_1985,N_1793,N_1872);
nor U1986 (N_1986,N_1874,N_1818);
xor U1987 (N_1987,N_1814,N_1870);
or U1988 (N_1988,N_1767,N_1869);
and U1989 (N_1989,N_1836,N_1905);
and U1990 (N_1990,N_1790,N_1846);
or U1991 (N_1991,N_1764,N_1822);
or U1992 (N_1992,N_1865,N_1858);
or U1993 (N_1993,N_1856,N_1910);
or U1994 (N_1994,N_1765,N_1779);
nand U1995 (N_1995,N_1787,N_1766);
nand U1996 (N_1996,N_1868,N_1898);
nand U1997 (N_1997,N_1889,N_1760);
xnor U1998 (N_1998,N_1914,N_1871);
and U1999 (N_1999,N_1877,N_1827);
xor U2000 (N_2000,N_1877,N_1795);
nand U2001 (N_2001,N_1761,N_1850);
nor U2002 (N_2002,N_1882,N_1878);
nand U2003 (N_2003,N_1849,N_1785);
nand U2004 (N_2004,N_1841,N_1772);
or U2005 (N_2005,N_1824,N_1919);
xor U2006 (N_2006,N_1826,N_1763);
xnor U2007 (N_2007,N_1791,N_1868);
xor U2008 (N_2008,N_1800,N_1763);
xnor U2009 (N_2009,N_1875,N_1839);
xor U2010 (N_2010,N_1836,N_1879);
or U2011 (N_2011,N_1841,N_1823);
nand U2012 (N_2012,N_1819,N_1905);
xnor U2013 (N_2013,N_1893,N_1803);
nand U2014 (N_2014,N_1803,N_1844);
nand U2015 (N_2015,N_1903,N_1835);
nor U2016 (N_2016,N_1802,N_1769);
nand U2017 (N_2017,N_1816,N_1916);
and U2018 (N_2018,N_1830,N_1892);
xnor U2019 (N_2019,N_1812,N_1867);
or U2020 (N_2020,N_1768,N_1918);
nor U2021 (N_2021,N_1909,N_1794);
nand U2022 (N_2022,N_1857,N_1881);
nand U2023 (N_2023,N_1770,N_1864);
or U2024 (N_2024,N_1845,N_1916);
xnor U2025 (N_2025,N_1822,N_1762);
or U2026 (N_2026,N_1786,N_1864);
nor U2027 (N_2027,N_1807,N_1798);
and U2028 (N_2028,N_1872,N_1779);
or U2029 (N_2029,N_1763,N_1906);
xnor U2030 (N_2030,N_1783,N_1804);
nor U2031 (N_2031,N_1903,N_1789);
xor U2032 (N_2032,N_1794,N_1883);
nand U2033 (N_2033,N_1793,N_1783);
and U2034 (N_2034,N_1784,N_1828);
xor U2035 (N_2035,N_1902,N_1901);
nor U2036 (N_2036,N_1847,N_1856);
nand U2037 (N_2037,N_1799,N_1827);
or U2038 (N_2038,N_1767,N_1855);
xnor U2039 (N_2039,N_1839,N_1780);
xor U2040 (N_2040,N_1884,N_1764);
nor U2041 (N_2041,N_1839,N_1887);
or U2042 (N_2042,N_1862,N_1766);
nor U2043 (N_2043,N_1781,N_1832);
nand U2044 (N_2044,N_1839,N_1905);
nor U2045 (N_2045,N_1761,N_1841);
nand U2046 (N_2046,N_1804,N_1825);
or U2047 (N_2047,N_1761,N_1868);
nand U2048 (N_2048,N_1843,N_1862);
xor U2049 (N_2049,N_1793,N_1789);
and U2050 (N_2050,N_1884,N_1818);
and U2051 (N_2051,N_1852,N_1847);
and U2052 (N_2052,N_1815,N_1818);
xor U2053 (N_2053,N_1841,N_1844);
xnor U2054 (N_2054,N_1893,N_1791);
xor U2055 (N_2055,N_1783,N_1791);
xnor U2056 (N_2056,N_1914,N_1894);
xor U2057 (N_2057,N_1779,N_1858);
and U2058 (N_2058,N_1826,N_1778);
nor U2059 (N_2059,N_1762,N_1870);
nor U2060 (N_2060,N_1814,N_1767);
or U2061 (N_2061,N_1825,N_1812);
or U2062 (N_2062,N_1888,N_1892);
nor U2063 (N_2063,N_1796,N_1896);
or U2064 (N_2064,N_1804,N_1801);
and U2065 (N_2065,N_1879,N_1797);
nor U2066 (N_2066,N_1866,N_1843);
or U2067 (N_2067,N_1813,N_1841);
nand U2068 (N_2068,N_1871,N_1897);
or U2069 (N_2069,N_1853,N_1796);
and U2070 (N_2070,N_1913,N_1879);
xor U2071 (N_2071,N_1800,N_1774);
nand U2072 (N_2072,N_1892,N_1848);
nand U2073 (N_2073,N_1826,N_1792);
nor U2074 (N_2074,N_1912,N_1869);
xor U2075 (N_2075,N_1840,N_1784);
nor U2076 (N_2076,N_1791,N_1778);
and U2077 (N_2077,N_1762,N_1912);
nand U2078 (N_2078,N_1771,N_1778);
xnor U2079 (N_2079,N_1831,N_1841);
xnor U2080 (N_2080,N_2027,N_2047);
xor U2081 (N_2081,N_2035,N_1927);
and U2082 (N_2082,N_1988,N_1938);
nor U2083 (N_2083,N_1923,N_1920);
nor U2084 (N_2084,N_1926,N_2066);
nand U2085 (N_2085,N_1959,N_2025);
or U2086 (N_2086,N_2071,N_1940);
nor U2087 (N_2087,N_2021,N_2008);
xnor U2088 (N_2088,N_2051,N_2073);
nand U2089 (N_2089,N_2067,N_2009);
and U2090 (N_2090,N_2006,N_1961);
nand U2091 (N_2091,N_1962,N_1969);
and U2092 (N_2092,N_2003,N_1954);
nor U2093 (N_2093,N_2039,N_1939);
and U2094 (N_2094,N_1978,N_2043);
or U2095 (N_2095,N_2011,N_1946);
nor U2096 (N_2096,N_2049,N_2062);
nor U2097 (N_2097,N_2077,N_2028);
xnor U2098 (N_2098,N_2017,N_2002);
or U2099 (N_2099,N_2001,N_2057);
and U2100 (N_2100,N_2068,N_2020);
and U2101 (N_2101,N_1932,N_2034);
nand U2102 (N_2102,N_1950,N_1925);
nand U2103 (N_2103,N_1922,N_2014);
nand U2104 (N_2104,N_1955,N_1973);
xnor U2105 (N_2105,N_2069,N_2063);
nand U2106 (N_2106,N_1945,N_2030);
xnor U2107 (N_2107,N_2050,N_2076);
nor U2108 (N_2108,N_2053,N_2056);
and U2109 (N_2109,N_2072,N_2012);
or U2110 (N_2110,N_2042,N_2064);
nand U2111 (N_2111,N_2061,N_2023);
nor U2112 (N_2112,N_1958,N_1951);
and U2113 (N_2113,N_2007,N_1936);
nand U2114 (N_2114,N_2044,N_2018);
xor U2115 (N_2115,N_1931,N_2022);
and U2116 (N_2116,N_2046,N_2037);
and U2117 (N_2117,N_2054,N_1965);
and U2118 (N_2118,N_1997,N_1921);
nor U2119 (N_2119,N_2045,N_1993);
xnor U2120 (N_2120,N_1928,N_1963);
nor U2121 (N_2121,N_2010,N_1980);
and U2122 (N_2122,N_2058,N_1970);
and U2123 (N_2123,N_1983,N_1935);
or U2124 (N_2124,N_2060,N_1995);
or U2125 (N_2125,N_1986,N_2040);
or U2126 (N_2126,N_1957,N_2031);
nand U2127 (N_2127,N_1953,N_1942);
and U2128 (N_2128,N_1998,N_2016);
and U2129 (N_2129,N_2005,N_1999);
or U2130 (N_2130,N_1982,N_2033);
xnor U2131 (N_2131,N_1979,N_2041);
and U2132 (N_2132,N_2024,N_1981);
or U2133 (N_2133,N_2029,N_2000);
nand U2134 (N_2134,N_1992,N_1972);
xnor U2135 (N_2135,N_1975,N_1934);
or U2136 (N_2136,N_1971,N_2015);
or U2137 (N_2137,N_2013,N_2038);
nand U2138 (N_2138,N_1976,N_2004);
nand U2139 (N_2139,N_2079,N_2059);
or U2140 (N_2140,N_2048,N_1930);
nand U2141 (N_2141,N_2065,N_1943);
or U2142 (N_2142,N_1989,N_1947);
xor U2143 (N_2143,N_2078,N_1960);
nor U2144 (N_2144,N_1964,N_1929);
and U2145 (N_2145,N_1937,N_1991);
xnor U2146 (N_2146,N_1985,N_1974);
xor U2147 (N_2147,N_2074,N_2019);
and U2148 (N_2148,N_2026,N_2052);
and U2149 (N_2149,N_1994,N_1949);
nor U2150 (N_2150,N_1966,N_1956);
nand U2151 (N_2151,N_1990,N_1941);
xnor U2152 (N_2152,N_1933,N_1987);
nor U2153 (N_2153,N_1967,N_2070);
nand U2154 (N_2154,N_1968,N_1924);
and U2155 (N_2155,N_2032,N_1944);
nand U2156 (N_2156,N_2036,N_1977);
or U2157 (N_2157,N_1996,N_1984);
xor U2158 (N_2158,N_1948,N_1952);
xnor U2159 (N_2159,N_2055,N_2075);
and U2160 (N_2160,N_1972,N_2057);
and U2161 (N_2161,N_1962,N_2059);
nand U2162 (N_2162,N_2001,N_1943);
and U2163 (N_2163,N_2035,N_1976);
or U2164 (N_2164,N_1993,N_2051);
xnor U2165 (N_2165,N_1972,N_2029);
nand U2166 (N_2166,N_1999,N_1983);
xor U2167 (N_2167,N_2058,N_1929);
and U2168 (N_2168,N_1964,N_2001);
nand U2169 (N_2169,N_2071,N_2030);
nand U2170 (N_2170,N_1997,N_2041);
nand U2171 (N_2171,N_1987,N_2064);
nand U2172 (N_2172,N_2028,N_2018);
or U2173 (N_2173,N_2004,N_1982);
nand U2174 (N_2174,N_1990,N_1930);
nor U2175 (N_2175,N_2077,N_1939);
or U2176 (N_2176,N_1993,N_1931);
nand U2177 (N_2177,N_1990,N_1977);
or U2178 (N_2178,N_1938,N_2016);
nand U2179 (N_2179,N_1925,N_2070);
xnor U2180 (N_2180,N_1982,N_1988);
nor U2181 (N_2181,N_1961,N_2049);
nor U2182 (N_2182,N_2011,N_1994);
nor U2183 (N_2183,N_2038,N_1997);
xor U2184 (N_2184,N_1998,N_1960);
nand U2185 (N_2185,N_2076,N_2045);
nand U2186 (N_2186,N_1954,N_1992);
nor U2187 (N_2187,N_2046,N_1958);
nor U2188 (N_2188,N_2073,N_2071);
nor U2189 (N_2189,N_2036,N_2047);
or U2190 (N_2190,N_1998,N_1985);
or U2191 (N_2191,N_2079,N_1948);
and U2192 (N_2192,N_1968,N_1983);
and U2193 (N_2193,N_2017,N_2074);
xnor U2194 (N_2194,N_2027,N_2069);
or U2195 (N_2195,N_1941,N_2073);
xnor U2196 (N_2196,N_1956,N_2003);
xor U2197 (N_2197,N_1920,N_2072);
or U2198 (N_2198,N_2024,N_1995);
nand U2199 (N_2199,N_1953,N_2000);
nor U2200 (N_2200,N_1928,N_2033);
nand U2201 (N_2201,N_1943,N_1947);
and U2202 (N_2202,N_1996,N_1995);
nor U2203 (N_2203,N_2037,N_2009);
nand U2204 (N_2204,N_2046,N_2074);
xor U2205 (N_2205,N_1977,N_1969);
nor U2206 (N_2206,N_1989,N_2028);
nor U2207 (N_2207,N_1942,N_1947);
xnor U2208 (N_2208,N_1983,N_1984);
nor U2209 (N_2209,N_2029,N_1927);
nand U2210 (N_2210,N_2016,N_2051);
or U2211 (N_2211,N_2075,N_2071);
nand U2212 (N_2212,N_1981,N_1926);
or U2213 (N_2213,N_1969,N_1938);
and U2214 (N_2214,N_2026,N_1962);
xnor U2215 (N_2215,N_1952,N_2042);
xnor U2216 (N_2216,N_1978,N_2077);
or U2217 (N_2217,N_1925,N_1965);
nor U2218 (N_2218,N_2063,N_1992);
nor U2219 (N_2219,N_2055,N_2004);
nor U2220 (N_2220,N_2036,N_1944);
nor U2221 (N_2221,N_2047,N_1979);
nand U2222 (N_2222,N_1929,N_1946);
xor U2223 (N_2223,N_1925,N_2051);
or U2224 (N_2224,N_2055,N_1959);
nand U2225 (N_2225,N_1952,N_2077);
xnor U2226 (N_2226,N_1967,N_1939);
nand U2227 (N_2227,N_2011,N_2033);
or U2228 (N_2228,N_2023,N_1961);
nor U2229 (N_2229,N_1944,N_1964);
nor U2230 (N_2230,N_1984,N_1950);
or U2231 (N_2231,N_2047,N_1953);
nor U2232 (N_2232,N_1942,N_1968);
and U2233 (N_2233,N_1991,N_2018);
nand U2234 (N_2234,N_2036,N_2073);
xnor U2235 (N_2235,N_1944,N_2005);
nor U2236 (N_2236,N_2026,N_1987);
xor U2237 (N_2237,N_1974,N_1941);
nand U2238 (N_2238,N_2022,N_2011);
xnor U2239 (N_2239,N_2036,N_2005);
and U2240 (N_2240,N_2195,N_2092);
or U2241 (N_2241,N_2208,N_2084);
xnor U2242 (N_2242,N_2115,N_2151);
nand U2243 (N_2243,N_2100,N_2197);
nand U2244 (N_2244,N_2209,N_2202);
or U2245 (N_2245,N_2160,N_2238);
nor U2246 (N_2246,N_2112,N_2130);
xnor U2247 (N_2247,N_2085,N_2237);
nor U2248 (N_2248,N_2186,N_2143);
or U2249 (N_2249,N_2146,N_2175);
nor U2250 (N_2250,N_2181,N_2118);
or U2251 (N_2251,N_2194,N_2217);
or U2252 (N_2252,N_2179,N_2207);
or U2253 (N_2253,N_2124,N_2223);
or U2254 (N_2254,N_2236,N_2239);
nand U2255 (N_2255,N_2180,N_2110);
nor U2256 (N_2256,N_2184,N_2164);
nand U2257 (N_2257,N_2083,N_2128);
nor U2258 (N_2258,N_2171,N_2159);
nand U2259 (N_2259,N_2107,N_2101);
or U2260 (N_2260,N_2196,N_2129);
or U2261 (N_2261,N_2225,N_2133);
or U2262 (N_2262,N_2188,N_2087);
xor U2263 (N_2263,N_2139,N_2229);
nor U2264 (N_2264,N_2104,N_2154);
xnor U2265 (N_2265,N_2105,N_2114);
nand U2266 (N_2266,N_2169,N_2199);
xnor U2267 (N_2267,N_2149,N_2190);
nor U2268 (N_2268,N_2155,N_2233);
or U2269 (N_2269,N_2132,N_2235);
nand U2270 (N_2270,N_2117,N_2113);
and U2271 (N_2271,N_2156,N_2141);
and U2272 (N_2272,N_2150,N_2173);
xnor U2273 (N_2273,N_2096,N_2123);
nor U2274 (N_2274,N_2178,N_2191);
and U2275 (N_2275,N_2203,N_2089);
and U2276 (N_2276,N_2142,N_2152);
nor U2277 (N_2277,N_2095,N_2106);
xor U2278 (N_2278,N_2200,N_2140);
or U2279 (N_2279,N_2214,N_2116);
xnor U2280 (N_2280,N_2182,N_2111);
nor U2281 (N_2281,N_2082,N_2192);
nor U2282 (N_2282,N_2131,N_2187);
or U2283 (N_2283,N_2090,N_2094);
or U2284 (N_2284,N_2163,N_2127);
xor U2285 (N_2285,N_2162,N_2088);
nand U2286 (N_2286,N_2204,N_2174);
or U2287 (N_2287,N_2153,N_2224);
and U2288 (N_2288,N_2125,N_2138);
and U2289 (N_2289,N_2103,N_2157);
xor U2290 (N_2290,N_2212,N_2185);
nor U2291 (N_2291,N_2231,N_2218);
nand U2292 (N_2292,N_2098,N_2222);
nor U2293 (N_2293,N_2126,N_2215);
and U2294 (N_2294,N_2161,N_2172);
and U2295 (N_2295,N_2136,N_2122);
nand U2296 (N_2296,N_2220,N_2099);
or U2297 (N_2297,N_2165,N_2091);
nor U2298 (N_2298,N_2093,N_2216);
or U2299 (N_2299,N_2213,N_2234);
nand U2300 (N_2300,N_2145,N_2228);
xnor U2301 (N_2301,N_2137,N_2206);
or U2302 (N_2302,N_2168,N_2176);
nand U2303 (N_2303,N_2205,N_2144);
or U2304 (N_2304,N_2193,N_2120);
xnor U2305 (N_2305,N_2097,N_2226);
xnor U2306 (N_2306,N_2211,N_2148);
nand U2307 (N_2307,N_2177,N_2189);
nand U2308 (N_2308,N_2210,N_2158);
and U2309 (N_2309,N_2119,N_2221);
xnor U2310 (N_2310,N_2230,N_2198);
nor U2311 (N_2311,N_2108,N_2081);
nor U2312 (N_2312,N_2121,N_2227);
and U2313 (N_2313,N_2219,N_2183);
nor U2314 (N_2314,N_2167,N_2109);
xnor U2315 (N_2315,N_2102,N_2147);
and U2316 (N_2316,N_2201,N_2086);
or U2317 (N_2317,N_2166,N_2170);
nand U2318 (N_2318,N_2134,N_2080);
nor U2319 (N_2319,N_2232,N_2135);
nand U2320 (N_2320,N_2092,N_2139);
and U2321 (N_2321,N_2116,N_2216);
nor U2322 (N_2322,N_2107,N_2160);
xnor U2323 (N_2323,N_2218,N_2159);
nor U2324 (N_2324,N_2160,N_2146);
nor U2325 (N_2325,N_2133,N_2228);
or U2326 (N_2326,N_2119,N_2143);
nor U2327 (N_2327,N_2189,N_2149);
xnor U2328 (N_2328,N_2123,N_2179);
or U2329 (N_2329,N_2199,N_2148);
nand U2330 (N_2330,N_2173,N_2096);
nor U2331 (N_2331,N_2201,N_2092);
nor U2332 (N_2332,N_2083,N_2159);
nand U2333 (N_2333,N_2239,N_2100);
or U2334 (N_2334,N_2119,N_2223);
nor U2335 (N_2335,N_2084,N_2140);
and U2336 (N_2336,N_2218,N_2134);
and U2337 (N_2337,N_2087,N_2107);
or U2338 (N_2338,N_2169,N_2103);
or U2339 (N_2339,N_2154,N_2203);
and U2340 (N_2340,N_2215,N_2113);
nor U2341 (N_2341,N_2187,N_2118);
and U2342 (N_2342,N_2173,N_2228);
nand U2343 (N_2343,N_2153,N_2217);
xor U2344 (N_2344,N_2234,N_2156);
and U2345 (N_2345,N_2167,N_2210);
or U2346 (N_2346,N_2221,N_2160);
xnor U2347 (N_2347,N_2219,N_2084);
xnor U2348 (N_2348,N_2222,N_2167);
and U2349 (N_2349,N_2140,N_2212);
nand U2350 (N_2350,N_2126,N_2144);
nor U2351 (N_2351,N_2196,N_2161);
nand U2352 (N_2352,N_2112,N_2142);
and U2353 (N_2353,N_2192,N_2121);
xor U2354 (N_2354,N_2152,N_2133);
nand U2355 (N_2355,N_2097,N_2187);
nor U2356 (N_2356,N_2208,N_2163);
and U2357 (N_2357,N_2096,N_2212);
or U2358 (N_2358,N_2231,N_2136);
xnor U2359 (N_2359,N_2215,N_2151);
nand U2360 (N_2360,N_2185,N_2092);
nand U2361 (N_2361,N_2131,N_2146);
xnor U2362 (N_2362,N_2230,N_2135);
nand U2363 (N_2363,N_2215,N_2115);
or U2364 (N_2364,N_2116,N_2091);
nand U2365 (N_2365,N_2238,N_2145);
and U2366 (N_2366,N_2121,N_2197);
nor U2367 (N_2367,N_2105,N_2106);
xor U2368 (N_2368,N_2129,N_2219);
and U2369 (N_2369,N_2092,N_2203);
nor U2370 (N_2370,N_2092,N_2158);
nor U2371 (N_2371,N_2118,N_2106);
or U2372 (N_2372,N_2086,N_2231);
and U2373 (N_2373,N_2096,N_2149);
nor U2374 (N_2374,N_2199,N_2112);
nor U2375 (N_2375,N_2129,N_2092);
xnor U2376 (N_2376,N_2239,N_2146);
or U2377 (N_2377,N_2167,N_2206);
xor U2378 (N_2378,N_2089,N_2123);
nand U2379 (N_2379,N_2215,N_2191);
xor U2380 (N_2380,N_2202,N_2218);
nand U2381 (N_2381,N_2237,N_2086);
and U2382 (N_2382,N_2238,N_2117);
nor U2383 (N_2383,N_2119,N_2231);
and U2384 (N_2384,N_2217,N_2129);
xnor U2385 (N_2385,N_2233,N_2205);
and U2386 (N_2386,N_2165,N_2100);
and U2387 (N_2387,N_2092,N_2216);
nand U2388 (N_2388,N_2209,N_2183);
or U2389 (N_2389,N_2152,N_2125);
or U2390 (N_2390,N_2128,N_2206);
nor U2391 (N_2391,N_2205,N_2161);
nand U2392 (N_2392,N_2225,N_2151);
nor U2393 (N_2393,N_2167,N_2106);
xnor U2394 (N_2394,N_2189,N_2237);
and U2395 (N_2395,N_2129,N_2149);
nor U2396 (N_2396,N_2132,N_2091);
and U2397 (N_2397,N_2168,N_2210);
nor U2398 (N_2398,N_2214,N_2157);
or U2399 (N_2399,N_2193,N_2176);
xor U2400 (N_2400,N_2395,N_2255);
nand U2401 (N_2401,N_2376,N_2315);
nor U2402 (N_2402,N_2289,N_2385);
and U2403 (N_2403,N_2354,N_2311);
xnor U2404 (N_2404,N_2269,N_2291);
or U2405 (N_2405,N_2375,N_2275);
nor U2406 (N_2406,N_2303,N_2391);
and U2407 (N_2407,N_2325,N_2253);
or U2408 (N_2408,N_2397,N_2295);
nor U2409 (N_2409,N_2280,N_2331);
xnor U2410 (N_2410,N_2353,N_2358);
and U2411 (N_2411,N_2265,N_2324);
and U2412 (N_2412,N_2254,N_2258);
nand U2413 (N_2413,N_2259,N_2349);
nor U2414 (N_2414,N_2297,N_2389);
and U2415 (N_2415,N_2316,N_2320);
nand U2416 (N_2416,N_2330,N_2342);
nor U2417 (N_2417,N_2362,N_2244);
xnor U2418 (N_2418,N_2347,N_2266);
nand U2419 (N_2419,N_2336,N_2261);
or U2420 (N_2420,N_2248,N_2398);
xor U2421 (N_2421,N_2262,N_2240);
nand U2422 (N_2422,N_2250,N_2283);
or U2423 (N_2423,N_2293,N_2251);
nand U2424 (N_2424,N_2267,N_2318);
nor U2425 (N_2425,N_2360,N_2359);
xnor U2426 (N_2426,N_2386,N_2279);
and U2427 (N_2427,N_2392,N_2271);
xnor U2428 (N_2428,N_2356,N_2334);
nor U2429 (N_2429,N_2305,N_2317);
or U2430 (N_2430,N_2340,N_2301);
or U2431 (N_2431,N_2270,N_2309);
and U2432 (N_2432,N_2304,N_2390);
xnor U2433 (N_2433,N_2241,N_2296);
or U2434 (N_2434,N_2257,N_2346);
or U2435 (N_2435,N_2322,N_2287);
nor U2436 (N_2436,N_2246,N_2285);
xor U2437 (N_2437,N_2380,N_2276);
nand U2438 (N_2438,N_2307,N_2326);
or U2439 (N_2439,N_2278,N_2306);
or U2440 (N_2440,N_2374,N_2286);
nor U2441 (N_2441,N_2284,N_2387);
nor U2442 (N_2442,N_2394,N_2335);
xnor U2443 (N_2443,N_2345,N_2399);
or U2444 (N_2444,N_2256,N_2328);
nor U2445 (N_2445,N_2366,N_2355);
nor U2446 (N_2446,N_2370,N_2393);
nand U2447 (N_2447,N_2351,N_2302);
nor U2448 (N_2448,N_2298,N_2282);
or U2449 (N_2449,N_2323,N_2382);
and U2450 (N_2450,N_2350,N_2357);
nor U2451 (N_2451,N_2364,N_2365);
xor U2452 (N_2452,N_2319,N_2272);
xor U2453 (N_2453,N_2273,N_2245);
or U2454 (N_2454,N_2333,N_2383);
xnor U2455 (N_2455,N_2344,N_2367);
nand U2456 (N_2456,N_2348,N_2388);
xor U2457 (N_2457,N_2252,N_2381);
and U2458 (N_2458,N_2292,N_2314);
or U2459 (N_2459,N_2379,N_2290);
xor U2460 (N_2460,N_2332,N_2341);
nand U2461 (N_2461,N_2260,N_2361);
nand U2462 (N_2462,N_2243,N_2338);
nor U2463 (N_2463,N_2329,N_2321);
nand U2464 (N_2464,N_2310,N_2369);
and U2465 (N_2465,N_2277,N_2249);
nand U2466 (N_2466,N_2372,N_2242);
and U2467 (N_2467,N_2371,N_2396);
nand U2468 (N_2468,N_2343,N_2288);
or U2469 (N_2469,N_2247,N_2268);
and U2470 (N_2470,N_2308,N_2312);
and U2471 (N_2471,N_2352,N_2378);
or U2472 (N_2472,N_2313,N_2300);
nor U2473 (N_2473,N_2263,N_2264);
nand U2474 (N_2474,N_2274,N_2337);
and U2475 (N_2475,N_2327,N_2377);
or U2476 (N_2476,N_2373,N_2281);
nand U2477 (N_2477,N_2299,N_2363);
nand U2478 (N_2478,N_2384,N_2294);
and U2479 (N_2479,N_2339,N_2368);
xnor U2480 (N_2480,N_2353,N_2371);
nand U2481 (N_2481,N_2330,N_2286);
nor U2482 (N_2482,N_2302,N_2256);
nor U2483 (N_2483,N_2254,N_2335);
and U2484 (N_2484,N_2354,N_2264);
and U2485 (N_2485,N_2331,N_2376);
or U2486 (N_2486,N_2269,N_2355);
nor U2487 (N_2487,N_2273,N_2300);
nand U2488 (N_2488,N_2387,N_2249);
nand U2489 (N_2489,N_2244,N_2297);
nor U2490 (N_2490,N_2295,N_2386);
and U2491 (N_2491,N_2332,N_2280);
and U2492 (N_2492,N_2389,N_2312);
nand U2493 (N_2493,N_2273,N_2333);
and U2494 (N_2494,N_2348,N_2393);
xnor U2495 (N_2495,N_2350,N_2338);
and U2496 (N_2496,N_2256,N_2305);
and U2497 (N_2497,N_2358,N_2316);
xor U2498 (N_2498,N_2296,N_2249);
or U2499 (N_2499,N_2329,N_2290);
or U2500 (N_2500,N_2396,N_2342);
nor U2501 (N_2501,N_2379,N_2275);
and U2502 (N_2502,N_2294,N_2281);
xor U2503 (N_2503,N_2340,N_2241);
nor U2504 (N_2504,N_2303,N_2241);
and U2505 (N_2505,N_2306,N_2281);
xor U2506 (N_2506,N_2315,N_2348);
xnor U2507 (N_2507,N_2253,N_2304);
nand U2508 (N_2508,N_2357,N_2259);
nor U2509 (N_2509,N_2372,N_2256);
nand U2510 (N_2510,N_2283,N_2356);
and U2511 (N_2511,N_2276,N_2399);
nor U2512 (N_2512,N_2344,N_2329);
xnor U2513 (N_2513,N_2324,N_2313);
or U2514 (N_2514,N_2361,N_2348);
xnor U2515 (N_2515,N_2283,N_2304);
nor U2516 (N_2516,N_2338,N_2394);
nor U2517 (N_2517,N_2318,N_2284);
and U2518 (N_2518,N_2346,N_2291);
nor U2519 (N_2519,N_2260,N_2391);
or U2520 (N_2520,N_2341,N_2327);
or U2521 (N_2521,N_2397,N_2275);
nand U2522 (N_2522,N_2266,N_2334);
and U2523 (N_2523,N_2261,N_2366);
nor U2524 (N_2524,N_2251,N_2333);
nor U2525 (N_2525,N_2322,N_2266);
nor U2526 (N_2526,N_2396,N_2377);
nor U2527 (N_2527,N_2393,N_2394);
and U2528 (N_2528,N_2317,N_2288);
and U2529 (N_2529,N_2327,N_2289);
xor U2530 (N_2530,N_2253,N_2252);
or U2531 (N_2531,N_2301,N_2272);
nand U2532 (N_2532,N_2281,N_2305);
nand U2533 (N_2533,N_2389,N_2336);
nor U2534 (N_2534,N_2270,N_2329);
nand U2535 (N_2535,N_2373,N_2258);
nor U2536 (N_2536,N_2399,N_2395);
or U2537 (N_2537,N_2368,N_2348);
or U2538 (N_2538,N_2379,N_2293);
nand U2539 (N_2539,N_2269,N_2337);
nor U2540 (N_2540,N_2246,N_2387);
and U2541 (N_2541,N_2320,N_2291);
nand U2542 (N_2542,N_2368,N_2260);
nor U2543 (N_2543,N_2367,N_2330);
or U2544 (N_2544,N_2339,N_2291);
nor U2545 (N_2545,N_2330,N_2394);
nor U2546 (N_2546,N_2307,N_2374);
xnor U2547 (N_2547,N_2335,N_2323);
nor U2548 (N_2548,N_2313,N_2311);
nor U2549 (N_2549,N_2284,N_2386);
xor U2550 (N_2550,N_2299,N_2322);
nand U2551 (N_2551,N_2310,N_2247);
xor U2552 (N_2552,N_2349,N_2380);
or U2553 (N_2553,N_2281,N_2329);
and U2554 (N_2554,N_2375,N_2348);
xnor U2555 (N_2555,N_2283,N_2338);
nand U2556 (N_2556,N_2353,N_2285);
nor U2557 (N_2557,N_2241,N_2373);
or U2558 (N_2558,N_2311,N_2287);
nand U2559 (N_2559,N_2394,N_2392);
nand U2560 (N_2560,N_2516,N_2403);
xor U2561 (N_2561,N_2435,N_2417);
nand U2562 (N_2562,N_2532,N_2511);
and U2563 (N_2563,N_2542,N_2484);
nor U2564 (N_2564,N_2528,N_2538);
nor U2565 (N_2565,N_2420,N_2544);
or U2566 (N_2566,N_2414,N_2457);
nor U2567 (N_2567,N_2413,N_2526);
nor U2568 (N_2568,N_2551,N_2423);
nand U2569 (N_2569,N_2469,N_2454);
nand U2570 (N_2570,N_2477,N_2547);
nand U2571 (N_2571,N_2410,N_2549);
or U2572 (N_2572,N_2529,N_2557);
nand U2573 (N_2573,N_2452,N_2463);
xnor U2574 (N_2574,N_2491,N_2422);
or U2575 (N_2575,N_2558,N_2552);
or U2576 (N_2576,N_2508,N_2426);
nor U2577 (N_2577,N_2522,N_2464);
nor U2578 (N_2578,N_2418,N_2424);
or U2579 (N_2579,N_2407,N_2539);
nand U2580 (N_2580,N_2408,N_2404);
xor U2581 (N_2581,N_2536,N_2482);
or U2582 (N_2582,N_2523,N_2412);
xnor U2583 (N_2583,N_2546,N_2447);
xnor U2584 (N_2584,N_2441,N_2541);
nor U2585 (N_2585,N_2489,N_2462);
or U2586 (N_2586,N_2493,N_2535);
nor U2587 (N_2587,N_2531,N_2442);
nor U2588 (N_2588,N_2451,N_2554);
nand U2589 (N_2589,N_2445,N_2470);
and U2590 (N_2590,N_2439,N_2505);
or U2591 (N_2591,N_2425,N_2460);
nor U2592 (N_2592,N_2517,N_2510);
and U2593 (N_2593,N_2540,N_2409);
nor U2594 (N_2594,N_2416,N_2525);
or U2595 (N_2595,N_2448,N_2427);
and U2596 (N_2596,N_2437,N_2483);
nand U2597 (N_2597,N_2429,N_2436);
or U2598 (N_2598,N_2475,N_2518);
xnor U2599 (N_2599,N_2485,N_2455);
nand U2600 (N_2600,N_2497,N_2486);
nand U2601 (N_2601,N_2471,N_2548);
nor U2602 (N_2602,N_2472,N_2402);
nand U2603 (N_2603,N_2405,N_2465);
nor U2604 (N_2604,N_2456,N_2432);
and U2605 (N_2605,N_2507,N_2433);
xor U2606 (N_2606,N_2496,N_2492);
or U2607 (N_2607,N_2476,N_2478);
or U2608 (N_2608,N_2503,N_2506);
nand U2609 (N_2609,N_2556,N_2501);
or U2610 (N_2610,N_2499,N_2512);
or U2611 (N_2611,N_2480,N_2530);
nor U2612 (N_2612,N_2490,N_2509);
and U2613 (N_2613,N_2521,N_2553);
xnor U2614 (N_2614,N_2487,N_2550);
xor U2615 (N_2615,N_2449,N_2520);
and U2616 (N_2616,N_2504,N_2500);
or U2617 (N_2617,N_2559,N_2400);
nor U2618 (N_2618,N_2431,N_2440);
nor U2619 (N_2619,N_2438,N_2494);
nor U2620 (N_2620,N_2415,N_2545);
and U2621 (N_2621,N_2466,N_2481);
nor U2622 (N_2622,N_2419,N_2519);
nand U2623 (N_2623,N_2458,N_2524);
nor U2624 (N_2624,N_2446,N_2428);
and U2625 (N_2625,N_2461,N_2498);
nor U2626 (N_2626,N_2401,N_2434);
and U2627 (N_2627,N_2513,N_2453);
nand U2628 (N_2628,N_2473,N_2495);
xor U2629 (N_2629,N_2543,N_2555);
xnor U2630 (N_2630,N_2459,N_2502);
nor U2631 (N_2631,N_2450,N_2488);
xnor U2632 (N_2632,N_2527,N_2515);
and U2633 (N_2633,N_2444,N_2514);
nand U2634 (N_2634,N_2468,N_2533);
nand U2635 (N_2635,N_2474,N_2479);
and U2636 (N_2636,N_2537,N_2467);
xor U2637 (N_2637,N_2406,N_2421);
nand U2638 (N_2638,N_2411,N_2534);
and U2639 (N_2639,N_2430,N_2443);
xor U2640 (N_2640,N_2431,N_2492);
and U2641 (N_2641,N_2433,N_2531);
xor U2642 (N_2642,N_2466,N_2504);
nor U2643 (N_2643,N_2420,N_2455);
or U2644 (N_2644,N_2421,N_2452);
xor U2645 (N_2645,N_2520,N_2552);
xnor U2646 (N_2646,N_2450,N_2510);
or U2647 (N_2647,N_2483,N_2538);
xor U2648 (N_2648,N_2549,N_2489);
xor U2649 (N_2649,N_2535,N_2526);
xnor U2650 (N_2650,N_2411,N_2526);
nor U2651 (N_2651,N_2504,N_2539);
xor U2652 (N_2652,N_2487,N_2512);
nand U2653 (N_2653,N_2531,N_2457);
or U2654 (N_2654,N_2498,N_2516);
and U2655 (N_2655,N_2486,N_2559);
or U2656 (N_2656,N_2543,N_2538);
or U2657 (N_2657,N_2540,N_2459);
and U2658 (N_2658,N_2474,N_2482);
and U2659 (N_2659,N_2492,N_2515);
nand U2660 (N_2660,N_2468,N_2412);
or U2661 (N_2661,N_2500,N_2515);
xor U2662 (N_2662,N_2538,N_2450);
xnor U2663 (N_2663,N_2408,N_2417);
nor U2664 (N_2664,N_2546,N_2450);
xnor U2665 (N_2665,N_2552,N_2542);
nand U2666 (N_2666,N_2489,N_2425);
nor U2667 (N_2667,N_2427,N_2468);
or U2668 (N_2668,N_2486,N_2443);
and U2669 (N_2669,N_2491,N_2523);
and U2670 (N_2670,N_2454,N_2453);
and U2671 (N_2671,N_2410,N_2440);
and U2672 (N_2672,N_2440,N_2452);
xor U2673 (N_2673,N_2471,N_2421);
nand U2674 (N_2674,N_2495,N_2549);
nand U2675 (N_2675,N_2457,N_2516);
and U2676 (N_2676,N_2442,N_2471);
nor U2677 (N_2677,N_2446,N_2467);
xnor U2678 (N_2678,N_2555,N_2547);
xnor U2679 (N_2679,N_2456,N_2495);
or U2680 (N_2680,N_2458,N_2503);
nand U2681 (N_2681,N_2523,N_2405);
or U2682 (N_2682,N_2540,N_2521);
nand U2683 (N_2683,N_2503,N_2476);
nand U2684 (N_2684,N_2506,N_2420);
xor U2685 (N_2685,N_2479,N_2549);
nand U2686 (N_2686,N_2505,N_2529);
nor U2687 (N_2687,N_2419,N_2471);
nor U2688 (N_2688,N_2423,N_2507);
and U2689 (N_2689,N_2527,N_2440);
nor U2690 (N_2690,N_2464,N_2555);
nand U2691 (N_2691,N_2492,N_2501);
nand U2692 (N_2692,N_2535,N_2418);
xor U2693 (N_2693,N_2435,N_2421);
xnor U2694 (N_2694,N_2426,N_2467);
nand U2695 (N_2695,N_2467,N_2401);
nor U2696 (N_2696,N_2515,N_2524);
nand U2697 (N_2697,N_2513,N_2471);
or U2698 (N_2698,N_2512,N_2485);
xnor U2699 (N_2699,N_2439,N_2434);
xnor U2700 (N_2700,N_2536,N_2519);
xnor U2701 (N_2701,N_2457,N_2542);
and U2702 (N_2702,N_2440,N_2435);
nor U2703 (N_2703,N_2543,N_2528);
and U2704 (N_2704,N_2558,N_2469);
xor U2705 (N_2705,N_2544,N_2414);
and U2706 (N_2706,N_2494,N_2471);
xor U2707 (N_2707,N_2417,N_2455);
and U2708 (N_2708,N_2421,N_2423);
or U2709 (N_2709,N_2458,N_2508);
or U2710 (N_2710,N_2441,N_2474);
nand U2711 (N_2711,N_2411,N_2539);
and U2712 (N_2712,N_2558,N_2556);
or U2713 (N_2713,N_2533,N_2469);
nand U2714 (N_2714,N_2413,N_2448);
and U2715 (N_2715,N_2482,N_2456);
or U2716 (N_2716,N_2428,N_2471);
or U2717 (N_2717,N_2460,N_2463);
or U2718 (N_2718,N_2485,N_2451);
xnor U2719 (N_2719,N_2541,N_2525);
xor U2720 (N_2720,N_2677,N_2714);
nand U2721 (N_2721,N_2719,N_2632);
or U2722 (N_2722,N_2614,N_2574);
or U2723 (N_2723,N_2686,N_2671);
nand U2724 (N_2724,N_2585,N_2660);
xor U2725 (N_2725,N_2705,N_2624);
and U2726 (N_2726,N_2664,N_2644);
nor U2727 (N_2727,N_2667,N_2687);
or U2728 (N_2728,N_2608,N_2635);
xor U2729 (N_2729,N_2629,N_2586);
or U2730 (N_2730,N_2665,N_2592);
nand U2731 (N_2731,N_2628,N_2616);
xor U2732 (N_2732,N_2668,N_2692);
and U2733 (N_2733,N_2607,N_2690);
or U2734 (N_2734,N_2681,N_2684);
or U2735 (N_2735,N_2706,N_2653);
xor U2736 (N_2736,N_2560,N_2562);
xor U2737 (N_2737,N_2646,N_2716);
or U2738 (N_2738,N_2656,N_2617);
or U2739 (N_2739,N_2654,N_2642);
or U2740 (N_2740,N_2680,N_2682);
nand U2741 (N_2741,N_2584,N_2701);
xnor U2742 (N_2742,N_2703,N_2566);
and U2743 (N_2743,N_2593,N_2622);
and U2744 (N_2744,N_2702,N_2674);
nand U2745 (N_2745,N_2599,N_2565);
nand U2746 (N_2746,N_2641,N_2619);
nor U2747 (N_2747,N_2672,N_2568);
nor U2748 (N_2748,N_2579,N_2572);
nor U2749 (N_2749,N_2620,N_2655);
xor U2750 (N_2750,N_2673,N_2580);
nor U2751 (N_2751,N_2689,N_2604);
xnor U2752 (N_2752,N_2658,N_2691);
or U2753 (N_2753,N_2577,N_2631);
xor U2754 (N_2754,N_2713,N_2567);
or U2755 (N_2755,N_2563,N_2570);
xnor U2756 (N_2756,N_2670,N_2715);
nor U2757 (N_2757,N_2615,N_2657);
or U2758 (N_2758,N_2602,N_2693);
nor U2759 (N_2759,N_2587,N_2611);
or U2760 (N_2760,N_2700,N_2571);
nand U2761 (N_2761,N_2695,N_2596);
nand U2762 (N_2762,N_2634,N_2613);
nand U2763 (N_2763,N_2662,N_2609);
or U2764 (N_2764,N_2650,N_2603);
nor U2765 (N_2765,N_2645,N_2589);
xor U2766 (N_2766,N_2709,N_2661);
nand U2767 (N_2767,N_2649,N_2712);
and U2768 (N_2768,N_2694,N_2651);
nand U2769 (N_2769,N_2663,N_2626);
xnor U2770 (N_2770,N_2711,N_2679);
and U2771 (N_2771,N_2643,N_2697);
nand U2772 (N_2772,N_2704,N_2647);
or U2773 (N_2773,N_2588,N_2618);
or U2774 (N_2774,N_2582,N_2698);
xor U2775 (N_2775,N_2666,N_2576);
nand U2776 (N_2776,N_2605,N_2623);
or U2777 (N_2777,N_2638,N_2600);
and U2778 (N_2778,N_2710,N_2669);
or U2779 (N_2779,N_2606,N_2583);
nor U2780 (N_2780,N_2636,N_2696);
and U2781 (N_2781,N_2569,N_2652);
xor U2782 (N_2782,N_2640,N_2625);
nand U2783 (N_2783,N_2627,N_2639);
xnor U2784 (N_2784,N_2573,N_2678);
nand U2785 (N_2785,N_2594,N_2708);
nand U2786 (N_2786,N_2718,N_2659);
or U2787 (N_2787,N_2621,N_2630);
nand U2788 (N_2788,N_2685,N_2610);
nor U2789 (N_2789,N_2717,N_2676);
nand U2790 (N_2790,N_2707,N_2595);
xor U2791 (N_2791,N_2699,N_2561);
and U2792 (N_2792,N_2601,N_2648);
and U2793 (N_2793,N_2581,N_2564);
xnor U2794 (N_2794,N_2675,N_2633);
nand U2795 (N_2795,N_2597,N_2683);
nand U2796 (N_2796,N_2591,N_2575);
and U2797 (N_2797,N_2688,N_2578);
xnor U2798 (N_2798,N_2590,N_2637);
nand U2799 (N_2799,N_2598,N_2612);
and U2800 (N_2800,N_2714,N_2607);
and U2801 (N_2801,N_2584,N_2564);
nor U2802 (N_2802,N_2635,N_2606);
nor U2803 (N_2803,N_2621,N_2681);
and U2804 (N_2804,N_2560,N_2588);
or U2805 (N_2805,N_2595,N_2666);
nand U2806 (N_2806,N_2680,N_2645);
xnor U2807 (N_2807,N_2646,N_2575);
or U2808 (N_2808,N_2581,N_2667);
nor U2809 (N_2809,N_2690,N_2579);
nand U2810 (N_2810,N_2657,N_2692);
nor U2811 (N_2811,N_2623,N_2695);
nand U2812 (N_2812,N_2706,N_2635);
nand U2813 (N_2813,N_2700,N_2715);
nor U2814 (N_2814,N_2684,N_2668);
or U2815 (N_2815,N_2638,N_2633);
nor U2816 (N_2816,N_2674,N_2597);
or U2817 (N_2817,N_2562,N_2705);
or U2818 (N_2818,N_2593,N_2652);
and U2819 (N_2819,N_2683,N_2713);
xnor U2820 (N_2820,N_2626,N_2620);
xnor U2821 (N_2821,N_2677,N_2648);
and U2822 (N_2822,N_2656,N_2625);
nor U2823 (N_2823,N_2629,N_2605);
xor U2824 (N_2824,N_2691,N_2711);
nor U2825 (N_2825,N_2637,N_2610);
nand U2826 (N_2826,N_2565,N_2714);
nand U2827 (N_2827,N_2617,N_2639);
nand U2828 (N_2828,N_2568,N_2645);
or U2829 (N_2829,N_2561,N_2565);
or U2830 (N_2830,N_2568,N_2692);
nand U2831 (N_2831,N_2583,N_2711);
nand U2832 (N_2832,N_2672,N_2619);
nand U2833 (N_2833,N_2688,N_2634);
and U2834 (N_2834,N_2606,N_2611);
or U2835 (N_2835,N_2663,N_2659);
or U2836 (N_2836,N_2579,N_2619);
nand U2837 (N_2837,N_2596,N_2632);
and U2838 (N_2838,N_2618,N_2626);
xor U2839 (N_2839,N_2642,N_2656);
and U2840 (N_2840,N_2709,N_2696);
nand U2841 (N_2841,N_2651,N_2709);
and U2842 (N_2842,N_2561,N_2569);
or U2843 (N_2843,N_2631,N_2608);
nor U2844 (N_2844,N_2641,N_2674);
and U2845 (N_2845,N_2700,N_2614);
and U2846 (N_2846,N_2664,N_2600);
nand U2847 (N_2847,N_2666,N_2640);
or U2848 (N_2848,N_2566,N_2682);
or U2849 (N_2849,N_2676,N_2561);
nand U2850 (N_2850,N_2598,N_2652);
or U2851 (N_2851,N_2599,N_2579);
nor U2852 (N_2852,N_2572,N_2633);
xor U2853 (N_2853,N_2576,N_2645);
nand U2854 (N_2854,N_2628,N_2623);
nor U2855 (N_2855,N_2620,N_2688);
nor U2856 (N_2856,N_2620,N_2665);
nand U2857 (N_2857,N_2645,N_2606);
or U2858 (N_2858,N_2651,N_2706);
and U2859 (N_2859,N_2570,N_2634);
or U2860 (N_2860,N_2597,N_2593);
xor U2861 (N_2861,N_2662,N_2615);
xor U2862 (N_2862,N_2712,N_2579);
nor U2863 (N_2863,N_2586,N_2695);
nor U2864 (N_2864,N_2645,N_2693);
and U2865 (N_2865,N_2588,N_2595);
nand U2866 (N_2866,N_2635,N_2579);
and U2867 (N_2867,N_2632,N_2618);
nand U2868 (N_2868,N_2671,N_2571);
nand U2869 (N_2869,N_2625,N_2677);
nor U2870 (N_2870,N_2642,N_2684);
xor U2871 (N_2871,N_2583,N_2682);
nand U2872 (N_2872,N_2700,N_2699);
nand U2873 (N_2873,N_2574,N_2596);
and U2874 (N_2874,N_2651,N_2662);
nand U2875 (N_2875,N_2687,N_2571);
xor U2876 (N_2876,N_2620,N_2647);
nand U2877 (N_2877,N_2715,N_2685);
and U2878 (N_2878,N_2602,N_2699);
nor U2879 (N_2879,N_2588,N_2673);
nand U2880 (N_2880,N_2804,N_2801);
nor U2881 (N_2881,N_2724,N_2822);
xor U2882 (N_2882,N_2872,N_2798);
nand U2883 (N_2883,N_2863,N_2784);
xnor U2884 (N_2884,N_2857,N_2855);
nand U2885 (N_2885,N_2749,N_2738);
nand U2886 (N_2886,N_2764,N_2809);
xnor U2887 (N_2887,N_2788,N_2879);
nand U2888 (N_2888,N_2769,N_2736);
and U2889 (N_2889,N_2779,N_2852);
or U2890 (N_2890,N_2806,N_2866);
xor U2891 (N_2891,N_2861,N_2792);
xnor U2892 (N_2892,N_2723,N_2790);
nor U2893 (N_2893,N_2754,N_2878);
nor U2894 (N_2894,N_2793,N_2766);
and U2895 (N_2895,N_2753,N_2858);
xor U2896 (N_2896,N_2759,N_2831);
nor U2897 (N_2897,N_2745,N_2829);
or U2898 (N_2898,N_2851,N_2826);
or U2899 (N_2899,N_2803,N_2744);
nor U2900 (N_2900,N_2808,N_2807);
and U2901 (N_2901,N_2842,N_2867);
xor U2902 (N_2902,N_2871,N_2802);
nand U2903 (N_2903,N_2735,N_2805);
or U2904 (N_2904,N_2833,N_2785);
and U2905 (N_2905,N_2873,N_2752);
nand U2906 (N_2906,N_2875,N_2787);
and U2907 (N_2907,N_2732,N_2786);
and U2908 (N_2908,N_2824,N_2874);
or U2909 (N_2909,N_2853,N_2728);
xor U2910 (N_2910,N_2854,N_2725);
and U2911 (N_2911,N_2812,N_2856);
nand U2912 (N_2912,N_2835,N_2832);
and U2913 (N_2913,N_2747,N_2839);
and U2914 (N_2914,N_2814,N_2734);
nor U2915 (N_2915,N_2750,N_2763);
xnor U2916 (N_2916,N_2834,N_2840);
and U2917 (N_2917,N_2870,N_2774);
or U2918 (N_2918,N_2865,N_2755);
xnor U2919 (N_2919,N_2844,N_2848);
and U2920 (N_2920,N_2761,N_2841);
nor U2921 (N_2921,N_2776,N_2799);
and U2922 (N_2922,N_2756,N_2862);
nor U2923 (N_2923,N_2739,N_2817);
xor U2924 (N_2924,N_2827,N_2860);
and U2925 (N_2925,N_2737,N_2820);
nor U2926 (N_2926,N_2777,N_2795);
nand U2927 (N_2927,N_2876,N_2746);
nor U2928 (N_2928,N_2741,N_2772);
or U2929 (N_2929,N_2730,N_2836);
or U2930 (N_2930,N_2760,N_2810);
and U2931 (N_2931,N_2846,N_2849);
nand U2932 (N_2932,N_2773,N_2778);
and U2933 (N_2933,N_2765,N_2775);
xnor U2934 (N_2934,N_2823,N_2722);
xor U2935 (N_2935,N_2830,N_2850);
xor U2936 (N_2936,N_2800,N_2859);
and U2937 (N_2937,N_2758,N_2762);
nor U2938 (N_2938,N_2843,N_2733);
nand U2939 (N_2939,N_2748,N_2726);
or U2940 (N_2940,N_2821,N_2813);
nor U2941 (N_2941,N_2782,N_2811);
xor U2942 (N_2942,N_2794,N_2868);
and U2943 (N_2943,N_2721,N_2847);
xnor U2944 (N_2944,N_2740,N_2742);
and U2945 (N_2945,N_2789,N_2757);
and U2946 (N_2946,N_2791,N_2767);
nand U2947 (N_2947,N_2828,N_2731);
xor U2948 (N_2948,N_2877,N_2838);
nor U2949 (N_2949,N_2727,N_2819);
or U2950 (N_2950,N_2825,N_2720);
nand U2951 (N_2951,N_2743,N_2751);
nand U2952 (N_2952,N_2837,N_2729);
xor U2953 (N_2953,N_2770,N_2818);
or U2954 (N_2954,N_2869,N_2816);
nor U2955 (N_2955,N_2768,N_2864);
nand U2956 (N_2956,N_2783,N_2796);
nor U2957 (N_2957,N_2845,N_2781);
xnor U2958 (N_2958,N_2780,N_2797);
or U2959 (N_2959,N_2815,N_2771);
nand U2960 (N_2960,N_2875,N_2760);
nand U2961 (N_2961,N_2854,N_2779);
nand U2962 (N_2962,N_2824,N_2813);
or U2963 (N_2963,N_2720,N_2862);
and U2964 (N_2964,N_2839,N_2766);
xor U2965 (N_2965,N_2809,N_2851);
nor U2966 (N_2966,N_2771,N_2877);
nand U2967 (N_2967,N_2769,N_2837);
and U2968 (N_2968,N_2737,N_2822);
or U2969 (N_2969,N_2850,N_2849);
or U2970 (N_2970,N_2739,N_2876);
nor U2971 (N_2971,N_2726,N_2801);
nor U2972 (N_2972,N_2814,N_2843);
or U2973 (N_2973,N_2778,N_2800);
nor U2974 (N_2974,N_2727,N_2768);
nand U2975 (N_2975,N_2725,N_2812);
nand U2976 (N_2976,N_2853,N_2740);
xnor U2977 (N_2977,N_2799,N_2748);
xnor U2978 (N_2978,N_2775,N_2801);
nor U2979 (N_2979,N_2761,N_2820);
nand U2980 (N_2980,N_2837,N_2834);
nand U2981 (N_2981,N_2807,N_2762);
and U2982 (N_2982,N_2841,N_2821);
nand U2983 (N_2983,N_2819,N_2729);
nor U2984 (N_2984,N_2832,N_2874);
nand U2985 (N_2985,N_2757,N_2838);
nand U2986 (N_2986,N_2877,N_2793);
or U2987 (N_2987,N_2802,N_2778);
or U2988 (N_2988,N_2728,N_2779);
nand U2989 (N_2989,N_2732,N_2858);
nor U2990 (N_2990,N_2814,N_2869);
nand U2991 (N_2991,N_2870,N_2722);
xor U2992 (N_2992,N_2793,N_2804);
or U2993 (N_2993,N_2759,N_2791);
nor U2994 (N_2994,N_2775,N_2878);
nor U2995 (N_2995,N_2764,N_2772);
or U2996 (N_2996,N_2819,N_2853);
or U2997 (N_2997,N_2798,N_2879);
nand U2998 (N_2998,N_2813,N_2726);
nand U2999 (N_2999,N_2838,N_2805);
nand U3000 (N_3000,N_2786,N_2821);
and U3001 (N_3001,N_2770,N_2871);
and U3002 (N_3002,N_2812,N_2762);
or U3003 (N_3003,N_2740,N_2793);
or U3004 (N_3004,N_2809,N_2834);
or U3005 (N_3005,N_2878,N_2873);
and U3006 (N_3006,N_2814,N_2771);
nor U3007 (N_3007,N_2752,N_2827);
xnor U3008 (N_3008,N_2729,N_2870);
or U3009 (N_3009,N_2875,N_2837);
or U3010 (N_3010,N_2801,N_2866);
and U3011 (N_3011,N_2786,N_2772);
or U3012 (N_3012,N_2848,N_2797);
nor U3013 (N_3013,N_2835,N_2773);
and U3014 (N_3014,N_2781,N_2756);
and U3015 (N_3015,N_2817,N_2801);
nor U3016 (N_3016,N_2770,N_2801);
xnor U3017 (N_3017,N_2839,N_2876);
nand U3018 (N_3018,N_2772,N_2756);
xnor U3019 (N_3019,N_2837,N_2757);
xor U3020 (N_3020,N_2837,N_2826);
nand U3021 (N_3021,N_2804,N_2843);
or U3022 (N_3022,N_2774,N_2761);
and U3023 (N_3023,N_2774,N_2820);
nor U3024 (N_3024,N_2876,N_2795);
nor U3025 (N_3025,N_2766,N_2782);
nand U3026 (N_3026,N_2740,N_2876);
and U3027 (N_3027,N_2738,N_2864);
xnor U3028 (N_3028,N_2875,N_2871);
or U3029 (N_3029,N_2859,N_2866);
nor U3030 (N_3030,N_2755,N_2756);
nand U3031 (N_3031,N_2757,N_2797);
nand U3032 (N_3032,N_2819,N_2736);
or U3033 (N_3033,N_2818,N_2760);
xor U3034 (N_3034,N_2817,N_2777);
nor U3035 (N_3035,N_2809,N_2833);
or U3036 (N_3036,N_2746,N_2756);
xor U3037 (N_3037,N_2828,N_2720);
nand U3038 (N_3038,N_2808,N_2834);
or U3039 (N_3039,N_2862,N_2773);
nor U3040 (N_3040,N_2932,N_2928);
and U3041 (N_3041,N_3013,N_2925);
or U3042 (N_3042,N_2948,N_3026);
nor U3043 (N_3043,N_2902,N_3020);
or U3044 (N_3044,N_2908,N_3006);
xnor U3045 (N_3045,N_2979,N_2963);
nand U3046 (N_3046,N_2880,N_3035);
or U3047 (N_3047,N_2969,N_2938);
and U3048 (N_3048,N_2915,N_3009);
and U3049 (N_3049,N_2968,N_3008);
nor U3050 (N_3050,N_2929,N_2895);
or U3051 (N_3051,N_2951,N_2980);
nand U3052 (N_3052,N_2947,N_3011);
and U3053 (N_3053,N_2972,N_3027);
or U3054 (N_3054,N_2894,N_2921);
and U3055 (N_3055,N_3010,N_3021);
and U3056 (N_3056,N_2960,N_2967);
xnor U3057 (N_3057,N_3037,N_2961);
and U3058 (N_3058,N_2996,N_2907);
nand U3059 (N_3059,N_2887,N_3028);
or U3060 (N_3060,N_3005,N_2909);
and U3061 (N_3061,N_3019,N_2978);
xnor U3062 (N_3062,N_2949,N_2985);
nor U3063 (N_3063,N_3015,N_2953);
nand U3064 (N_3064,N_2919,N_2910);
nor U3065 (N_3065,N_2924,N_2883);
nand U3066 (N_3066,N_2935,N_2882);
nand U3067 (N_3067,N_3025,N_3022);
xnor U3068 (N_3068,N_2990,N_2981);
nand U3069 (N_3069,N_3016,N_2999);
nand U3070 (N_3070,N_2957,N_3023);
nor U3071 (N_3071,N_2946,N_2931);
and U3072 (N_3072,N_2916,N_2993);
nor U3073 (N_3073,N_2898,N_3031);
nand U3074 (N_3074,N_2889,N_2998);
xor U3075 (N_3075,N_2984,N_2965);
nand U3076 (N_3076,N_2950,N_2930);
or U3077 (N_3077,N_2896,N_2973);
xor U3078 (N_3078,N_3030,N_2913);
xor U3079 (N_3079,N_2987,N_3007);
nor U3080 (N_3080,N_2891,N_2892);
xor U3081 (N_3081,N_2970,N_2983);
nand U3082 (N_3082,N_2986,N_3039);
nand U3083 (N_3083,N_3036,N_2955);
nor U3084 (N_3084,N_2994,N_3018);
and U3085 (N_3085,N_2927,N_3014);
xnor U3086 (N_3086,N_2936,N_2899);
nor U3087 (N_3087,N_2958,N_3001);
nor U3088 (N_3088,N_2939,N_2975);
nand U3089 (N_3089,N_2901,N_2988);
or U3090 (N_3090,N_2942,N_2923);
and U3091 (N_3091,N_2962,N_2897);
nand U3092 (N_3092,N_3002,N_2922);
or U3093 (N_3093,N_2971,N_2995);
nand U3094 (N_3094,N_3003,N_2933);
or U3095 (N_3095,N_2954,N_2884);
nand U3096 (N_3096,N_3032,N_2934);
and U3097 (N_3097,N_2945,N_2881);
or U3098 (N_3098,N_2952,N_3029);
nor U3099 (N_3099,N_3017,N_2918);
or U3100 (N_3100,N_2900,N_3033);
xor U3101 (N_3101,N_2966,N_2976);
and U3102 (N_3102,N_2917,N_2885);
and U3103 (N_3103,N_2905,N_2991);
nor U3104 (N_3104,N_2959,N_2912);
nand U3105 (N_3105,N_2893,N_2997);
nor U3106 (N_3106,N_2977,N_2940);
and U3107 (N_3107,N_2890,N_2920);
and U3108 (N_3108,N_3034,N_2888);
and U3109 (N_3109,N_2937,N_3024);
nor U3110 (N_3110,N_2941,N_2911);
or U3111 (N_3111,N_2982,N_3038);
xor U3112 (N_3112,N_2914,N_2956);
and U3113 (N_3113,N_2989,N_2943);
nand U3114 (N_3114,N_2944,N_2906);
and U3115 (N_3115,N_2903,N_3012);
nand U3116 (N_3116,N_2926,N_3000);
and U3117 (N_3117,N_2886,N_2904);
or U3118 (N_3118,N_3004,N_2974);
nor U3119 (N_3119,N_2964,N_2992);
or U3120 (N_3120,N_2987,N_3037);
and U3121 (N_3121,N_2990,N_3001);
xor U3122 (N_3122,N_3031,N_2886);
nor U3123 (N_3123,N_3026,N_2972);
or U3124 (N_3124,N_3034,N_2946);
nand U3125 (N_3125,N_3024,N_3011);
or U3126 (N_3126,N_3011,N_2908);
or U3127 (N_3127,N_2969,N_2966);
nand U3128 (N_3128,N_2939,N_2976);
xor U3129 (N_3129,N_3004,N_3030);
or U3130 (N_3130,N_3000,N_2952);
nand U3131 (N_3131,N_3016,N_3021);
nor U3132 (N_3132,N_3009,N_3017);
xnor U3133 (N_3133,N_2910,N_2889);
or U3134 (N_3134,N_2893,N_3018);
or U3135 (N_3135,N_2897,N_2895);
nor U3136 (N_3136,N_3013,N_3021);
or U3137 (N_3137,N_2976,N_3007);
or U3138 (N_3138,N_2924,N_2965);
and U3139 (N_3139,N_2979,N_2923);
and U3140 (N_3140,N_2960,N_2905);
xor U3141 (N_3141,N_2940,N_2905);
nand U3142 (N_3142,N_3009,N_2925);
xnor U3143 (N_3143,N_2926,N_2949);
nand U3144 (N_3144,N_2929,N_2961);
or U3145 (N_3145,N_2952,N_2881);
or U3146 (N_3146,N_2985,N_2973);
nand U3147 (N_3147,N_2995,N_2889);
nor U3148 (N_3148,N_2957,N_2914);
xor U3149 (N_3149,N_3013,N_2965);
xor U3150 (N_3150,N_3030,N_2998);
nor U3151 (N_3151,N_2999,N_3033);
nand U3152 (N_3152,N_2938,N_3039);
or U3153 (N_3153,N_2961,N_2909);
and U3154 (N_3154,N_2967,N_2890);
xor U3155 (N_3155,N_2979,N_2992);
nor U3156 (N_3156,N_2883,N_2929);
nor U3157 (N_3157,N_2995,N_2937);
or U3158 (N_3158,N_2986,N_2936);
and U3159 (N_3159,N_2901,N_2927);
or U3160 (N_3160,N_3027,N_3030);
xor U3161 (N_3161,N_2880,N_2934);
or U3162 (N_3162,N_2937,N_2885);
or U3163 (N_3163,N_2901,N_3003);
or U3164 (N_3164,N_2889,N_2962);
xnor U3165 (N_3165,N_2947,N_2923);
or U3166 (N_3166,N_2955,N_2930);
nor U3167 (N_3167,N_2941,N_2899);
nand U3168 (N_3168,N_3038,N_2911);
xnor U3169 (N_3169,N_2888,N_3028);
nor U3170 (N_3170,N_2905,N_3027);
nand U3171 (N_3171,N_2900,N_2924);
nand U3172 (N_3172,N_2912,N_2960);
or U3173 (N_3173,N_2949,N_2934);
nor U3174 (N_3174,N_3003,N_3024);
nand U3175 (N_3175,N_2912,N_2921);
or U3176 (N_3176,N_2959,N_2910);
or U3177 (N_3177,N_2901,N_2957);
or U3178 (N_3178,N_2888,N_2919);
nor U3179 (N_3179,N_2929,N_2966);
nor U3180 (N_3180,N_2932,N_2961);
nand U3181 (N_3181,N_3026,N_2903);
xnor U3182 (N_3182,N_2995,N_2936);
nand U3183 (N_3183,N_2962,N_2902);
or U3184 (N_3184,N_2953,N_2914);
nand U3185 (N_3185,N_3032,N_2988);
nor U3186 (N_3186,N_2928,N_2982);
nand U3187 (N_3187,N_2982,N_3007);
or U3188 (N_3188,N_3027,N_2998);
and U3189 (N_3189,N_2972,N_2984);
and U3190 (N_3190,N_2939,N_2986);
xor U3191 (N_3191,N_3014,N_2945);
nor U3192 (N_3192,N_2929,N_2916);
xor U3193 (N_3193,N_2883,N_2923);
and U3194 (N_3194,N_2993,N_2912);
xnor U3195 (N_3195,N_2910,N_2955);
nand U3196 (N_3196,N_2941,N_2902);
nor U3197 (N_3197,N_2910,N_2900);
or U3198 (N_3198,N_3031,N_2908);
or U3199 (N_3199,N_2949,N_2897);
and U3200 (N_3200,N_3093,N_3192);
nor U3201 (N_3201,N_3062,N_3199);
nor U3202 (N_3202,N_3165,N_3123);
and U3203 (N_3203,N_3127,N_3098);
and U3204 (N_3204,N_3063,N_3190);
and U3205 (N_3205,N_3166,N_3099);
and U3206 (N_3206,N_3147,N_3115);
or U3207 (N_3207,N_3044,N_3110);
nor U3208 (N_3208,N_3103,N_3089);
xnor U3209 (N_3209,N_3171,N_3073);
or U3210 (N_3210,N_3104,N_3059);
xor U3211 (N_3211,N_3079,N_3094);
nand U3212 (N_3212,N_3120,N_3184);
and U3213 (N_3213,N_3135,N_3131);
nand U3214 (N_3214,N_3149,N_3130);
and U3215 (N_3215,N_3183,N_3067);
and U3216 (N_3216,N_3168,N_3145);
and U3217 (N_3217,N_3185,N_3197);
nand U3218 (N_3218,N_3071,N_3117);
nor U3219 (N_3219,N_3143,N_3161);
and U3220 (N_3220,N_3174,N_3179);
xor U3221 (N_3221,N_3153,N_3097);
and U3222 (N_3222,N_3084,N_3111);
xnor U3223 (N_3223,N_3081,N_3181);
xnor U3224 (N_3224,N_3072,N_3055);
xor U3225 (N_3225,N_3057,N_3060);
nor U3226 (N_3226,N_3090,N_3085);
and U3227 (N_3227,N_3066,N_3116);
and U3228 (N_3228,N_3163,N_3188);
xor U3229 (N_3229,N_3195,N_3102);
xor U3230 (N_3230,N_3113,N_3096);
nor U3231 (N_3231,N_3041,N_3042);
xnor U3232 (N_3232,N_3162,N_3140);
xnor U3233 (N_3233,N_3069,N_3124);
nor U3234 (N_3234,N_3114,N_3178);
nor U3235 (N_3235,N_3164,N_3095);
xnor U3236 (N_3236,N_3076,N_3138);
xnor U3237 (N_3237,N_3158,N_3061);
nand U3238 (N_3238,N_3048,N_3086);
nand U3239 (N_3239,N_3170,N_3133);
nor U3240 (N_3240,N_3101,N_3121);
and U3241 (N_3241,N_3125,N_3045);
nor U3242 (N_3242,N_3100,N_3077);
xor U3243 (N_3243,N_3106,N_3068);
nand U3244 (N_3244,N_3191,N_3180);
nand U3245 (N_3245,N_3107,N_3128);
and U3246 (N_3246,N_3047,N_3075);
xor U3247 (N_3247,N_3169,N_3186);
or U3248 (N_3248,N_3088,N_3142);
and U3249 (N_3249,N_3046,N_3155);
xnor U3250 (N_3250,N_3141,N_3160);
nand U3251 (N_3251,N_3156,N_3052);
xor U3252 (N_3252,N_3056,N_3126);
or U3253 (N_3253,N_3118,N_3187);
nand U3254 (N_3254,N_3083,N_3176);
xnor U3255 (N_3255,N_3144,N_3196);
or U3256 (N_3256,N_3050,N_3119);
nor U3257 (N_3257,N_3177,N_3112);
and U3258 (N_3258,N_3122,N_3108);
nand U3259 (N_3259,N_3132,N_3080);
xnor U3260 (N_3260,N_3129,N_3198);
xnor U3261 (N_3261,N_3058,N_3078);
nor U3262 (N_3262,N_3148,N_3070);
nor U3263 (N_3263,N_3193,N_3139);
xnor U3264 (N_3264,N_3087,N_3040);
or U3265 (N_3265,N_3064,N_3189);
and U3266 (N_3266,N_3043,N_3151);
and U3267 (N_3267,N_3172,N_3173);
or U3268 (N_3268,N_3167,N_3105);
and U3269 (N_3269,N_3175,N_3154);
and U3270 (N_3270,N_3137,N_3053);
and U3271 (N_3271,N_3157,N_3049);
nor U3272 (N_3272,N_3065,N_3051);
or U3273 (N_3273,N_3194,N_3159);
and U3274 (N_3274,N_3091,N_3134);
nand U3275 (N_3275,N_3082,N_3146);
nor U3276 (N_3276,N_3182,N_3092);
or U3277 (N_3277,N_3150,N_3109);
and U3278 (N_3278,N_3136,N_3054);
xnor U3279 (N_3279,N_3152,N_3074);
and U3280 (N_3280,N_3119,N_3081);
xor U3281 (N_3281,N_3100,N_3090);
and U3282 (N_3282,N_3114,N_3143);
or U3283 (N_3283,N_3104,N_3188);
or U3284 (N_3284,N_3170,N_3119);
nor U3285 (N_3285,N_3161,N_3047);
xor U3286 (N_3286,N_3197,N_3048);
and U3287 (N_3287,N_3054,N_3195);
xor U3288 (N_3288,N_3073,N_3103);
xnor U3289 (N_3289,N_3199,N_3188);
and U3290 (N_3290,N_3106,N_3074);
nand U3291 (N_3291,N_3089,N_3170);
and U3292 (N_3292,N_3095,N_3122);
xnor U3293 (N_3293,N_3097,N_3113);
or U3294 (N_3294,N_3172,N_3144);
nand U3295 (N_3295,N_3128,N_3073);
nor U3296 (N_3296,N_3088,N_3160);
nand U3297 (N_3297,N_3193,N_3072);
nand U3298 (N_3298,N_3082,N_3168);
or U3299 (N_3299,N_3157,N_3191);
nand U3300 (N_3300,N_3142,N_3138);
nand U3301 (N_3301,N_3192,N_3077);
or U3302 (N_3302,N_3099,N_3108);
or U3303 (N_3303,N_3125,N_3041);
and U3304 (N_3304,N_3134,N_3045);
xor U3305 (N_3305,N_3125,N_3065);
xnor U3306 (N_3306,N_3123,N_3093);
or U3307 (N_3307,N_3168,N_3092);
nor U3308 (N_3308,N_3054,N_3122);
nor U3309 (N_3309,N_3082,N_3053);
and U3310 (N_3310,N_3135,N_3101);
xnor U3311 (N_3311,N_3134,N_3177);
xnor U3312 (N_3312,N_3077,N_3062);
nand U3313 (N_3313,N_3167,N_3143);
or U3314 (N_3314,N_3074,N_3121);
and U3315 (N_3315,N_3125,N_3103);
or U3316 (N_3316,N_3041,N_3108);
nor U3317 (N_3317,N_3188,N_3040);
xor U3318 (N_3318,N_3114,N_3186);
and U3319 (N_3319,N_3086,N_3155);
nor U3320 (N_3320,N_3086,N_3148);
and U3321 (N_3321,N_3062,N_3086);
nor U3322 (N_3322,N_3077,N_3160);
and U3323 (N_3323,N_3049,N_3198);
and U3324 (N_3324,N_3077,N_3093);
and U3325 (N_3325,N_3179,N_3176);
nor U3326 (N_3326,N_3193,N_3050);
and U3327 (N_3327,N_3119,N_3132);
xor U3328 (N_3328,N_3172,N_3198);
and U3329 (N_3329,N_3153,N_3116);
nand U3330 (N_3330,N_3163,N_3103);
xor U3331 (N_3331,N_3152,N_3070);
nand U3332 (N_3332,N_3072,N_3177);
or U3333 (N_3333,N_3131,N_3095);
or U3334 (N_3334,N_3112,N_3136);
nor U3335 (N_3335,N_3192,N_3137);
or U3336 (N_3336,N_3166,N_3110);
nor U3337 (N_3337,N_3096,N_3060);
and U3338 (N_3338,N_3114,N_3166);
and U3339 (N_3339,N_3126,N_3095);
nor U3340 (N_3340,N_3146,N_3197);
or U3341 (N_3341,N_3097,N_3176);
nor U3342 (N_3342,N_3101,N_3158);
nand U3343 (N_3343,N_3194,N_3077);
or U3344 (N_3344,N_3040,N_3069);
xnor U3345 (N_3345,N_3059,N_3108);
or U3346 (N_3346,N_3169,N_3128);
nand U3347 (N_3347,N_3194,N_3198);
nor U3348 (N_3348,N_3183,N_3162);
nor U3349 (N_3349,N_3071,N_3182);
and U3350 (N_3350,N_3198,N_3147);
xor U3351 (N_3351,N_3161,N_3157);
xnor U3352 (N_3352,N_3151,N_3075);
or U3353 (N_3353,N_3077,N_3061);
nand U3354 (N_3354,N_3197,N_3139);
nor U3355 (N_3355,N_3191,N_3057);
or U3356 (N_3356,N_3140,N_3199);
nand U3357 (N_3357,N_3092,N_3091);
and U3358 (N_3358,N_3117,N_3180);
nand U3359 (N_3359,N_3170,N_3064);
nand U3360 (N_3360,N_3219,N_3276);
xor U3361 (N_3361,N_3342,N_3306);
and U3362 (N_3362,N_3348,N_3319);
or U3363 (N_3363,N_3334,N_3290);
or U3364 (N_3364,N_3208,N_3269);
nor U3365 (N_3365,N_3346,N_3321);
nand U3366 (N_3366,N_3256,N_3252);
or U3367 (N_3367,N_3280,N_3325);
and U3368 (N_3368,N_3258,N_3358);
and U3369 (N_3369,N_3273,N_3215);
nand U3370 (N_3370,N_3201,N_3270);
nor U3371 (N_3371,N_3309,N_3304);
nand U3372 (N_3372,N_3209,N_3329);
nand U3373 (N_3373,N_3274,N_3217);
nand U3374 (N_3374,N_3243,N_3301);
and U3375 (N_3375,N_3331,N_3293);
nor U3376 (N_3376,N_3231,N_3356);
or U3377 (N_3377,N_3259,N_3235);
xor U3378 (N_3378,N_3339,N_3347);
and U3379 (N_3379,N_3204,N_3350);
nor U3380 (N_3380,N_3324,N_3253);
nor U3381 (N_3381,N_3246,N_3267);
or U3382 (N_3382,N_3299,N_3357);
and U3383 (N_3383,N_3330,N_3249);
nand U3384 (N_3384,N_3220,N_3233);
nand U3385 (N_3385,N_3335,N_3326);
or U3386 (N_3386,N_3203,N_3320);
and U3387 (N_3387,N_3300,N_3302);
nor U3388 (N_3388,N_3266,N_3359);
nand U3389 (N_3389,N_3238,N_3344);
xor U3390 (N_3390,N_3232,N_3323);
xnor U3391 (N_3391,N_3277,N_3336);
nor U3392 (N_3392,N_3227,N_3250);
and U3393 (N_3393,N_3272,N_3279);
or U3394 (N_3394,N_3212,N_3285);
or U3395 (N_3395,N_3353,N_3295);
or U3396 (N_3396,N_3244,N_3206);
or U3397 (N_3397,N_3332,N_3303);
nand U3398 (N_3398,N_3223,N_3247);
nor U3399 (N_3399,N_3322,N_3224);
nor U3400 (N_3400,N_3265,N_3207);
nand U3401 (N_3401,N_3355,N_3287);
nor U3402 (N_3402,N_3318,N_3283);
nor U3403 (N_3403,N_3281,N_3349);
nand U3404 (N_3404,N_3257,N_3205);
or U3405 (N_3405,N_3316,N_3288);
or U3406 (N_3406,N_3333,N_3228);
or U3407 (N_3407,N_3222,N_3340);
or U3408 (N_3408,N_3352,N_3234);
xor U3409 (N_3409,N_3292,N_3278);
nand U3410 (N_3410,N_3341,N_3296);
nor U3411 (N_3411,N_3310,N_3328);
and U3412 (N_3412,N_3307,N_3343);
and U3413 (N_3413,N_3245,N_3236);
or U3414 (N_3414,N_3241,N_3314);
or U3415 (N_3415,N_3251,N_3214);
and U3416 (N_3416,N_3275,N_3327);
or U3417 (N_3417,N_3239,N_3337);
or U3418 (N_3418,N_3262,N_3268);
and U3419 (N_3419,N_3291,N_3221);
or U3420 (N_3420,N_3213,N_3254);
nand U3421 (N_3421,N_3216,N_3230);
and U3422 (N_3422,N_3226,N_3294);
nor U3423 (N_3423,N_3264,N_3313);
nand U3424 (N_3424,N_3286,N_3242);
nand U3425 (N_3425,N_3354,N_3282);
nor U3426 (N_3426,N_3312,N_3345);
xor U3427 (N_3427,N_3211,N_3218);
xor U3428 (N_3428,N_3225,N_3284);
nor U3429 (N_3429,N_3263,N_3248);
nand U3430 (N_3430,N_3202,N_3315);
or U3431 (N_3431,N_3311,N_3298);
or U3432 (N_3432,N_3338,N_3210);
nor U3433 (N_3433,N_3229,N_3305);
nand U3434 (N_3434,N_3271,N_3317);
nand U3435 (N_3435,N_3297,N_3261);
nor U3436 (N_3436,N_3289,N_3260);
nor U3437 (N_3437,N_3240,N_3308);
nor U3438 (N_3438,N_3255,N_3351);
or U3439 (N_3439,N_3200,N_3237);
or U3440 (N_3440,N_3277,N_3358);
nand U3441 (N_3441,N_3317,N_3233);
or U3442 (N_3442,N_3337,N_3278);
or U3443 (N_3443,N_3328,N_3263);
nand U3444 (N_3444,N_3229,N_3205);
nor U3445 (N_3445,N_3330,N_3288);
nor U3446 (N_3446,N_3272,N_3314);
nor U3447 (N_3447,N_3285,N_3227);
and U3448 (N_3448,N_3208,N_3202);
nor U3449 (N_3449,N_3258,N_3237);
or U3450 (N_3450,N_3281,N_3212);
nor U3451 (N_3451,N_3314,N_3337);
and U3452 (N_3452,N_3217,N_3208);
nand U3453 (N_3453,N_3327,N_3300);
nand U3454 (N_3454,N_3352,N_3243);
nor U3455 (N_3455,N_3213,N_3296);
xor U3456 (N_3456,N_3279,N_3290);
nor U3457 (N_3457,N_3207,N_3308);
and U3458 (N_3458,N_3200,N_3309);
or U3459 (N_3459,N_3222,N_3328);
xnor U3460 (N_3460,N_3303,N_3295);
xnor U3461 (N_3461,N_3329,N_3286);
xnor U3462 (N_3462,N_3342,N_3248);
or U3463 (N_3463,N_3233,N_3232);
and U3464 (N_3464,N_3286,N_3235);
or U3465 (N_3465,N_3265,N_3295);
nor U3466 (N_3466,N_3313,N_3338);
and U3467 (N_3467,N_3228,N_3252);
and U3468 (N_3468,N_3253,N_3295);
and U3469 (N_3469,N_3314,N_3208);
or U3470 (N_3470,N_3296,N_3332);
nor U3471 (N_3471,N_3288,N_3244);
and U3472 (N_3472,N_3217,N_3319);
and U3473 (N_3473,N_3207,N_3250);
and U3474 (N_3474,N_3335,N_3221);
nand U3475 (N_3475,N_3327,N_3352);
nor U3476 (N_3476,N_3266,N_3299);
xor U3477 (N_3477,N_3228,N_3348);
and U3478 (N_3478,N_3352,N_3222);
xor U3479 (N_3479,N_3287,N_3235);
or U3480 (N_3480,N_3325,N_3242);
xor U3481 (N_3481,N_3353,N_3215);
nor U3482 (N_3482,N_3325,N_3276);
nor U3483 (N_3483,N_3287,N_3301);
xor U3484 (N_3484,N_3357,N_3224);
nand U3485 (N_3485,N_3290,N_3212);
xnor U3486 (N_3486,N_3335,N_3260);
or U3487 (N_3487,N_3242,N_3266);
xnor U3488 (N_3488,N_3218,N_3343);
nand U3489 (N_3489,N_3288,N_3221);
or U3490 (N_3490,N_3230,N_3226);
or U3491 (N_3491,N_3205,N_3247);
and U3492 (N_3492,N_3322,N_3250);
nand U3493 (N_3493,N_3231,N_3224);
nand U3494 (N_3494,N_3227,N_3347);
and U3495 (N_3495,N_3321,N_3240);
or U3496 (N_3496,N_3236,N_3331);
nand U3497 (N_3497,N_3307,N_3354);
xnor U3498 (N_3498,N_3271,N_3245);
nand U3499 (N_3499,N_3250,N_3285);
or U3500 (N_3500,N_3354,N_3245);
or U3501 (N_3501,N_3243,N_3215);
nor U3502 (N_3502,N_3267,N_3268);
nor U3503 (N_3503,N_3259,N_3344);
nor U3504 (N_3504,N_3226,N_3224);
nor U3505 (N_3505,N_3355,N_3238);
xnor U3506 (N_3506,N_3304,N_3278);
and U3507 (N_3507,N_3216,N_3239);
nand U3508 (N_3508,N_3261,N_3301);
nor U3509 (N_3509,N_3353,N_3278);
and U3510 (N_3510,N_3247,N_3300);
nand U3511 (N_3511,N_3287,N_3267);
and U3512 (N_3512,N_3215,N_3213);
or U3513 (N_3513,N_3276,N_3251);
or U3514 (N_3514,N_3236,N_3297);
nor U3515 (N_3515,N_3211,N_3323);
nor U3516 (N_3516,N_3304,N_3344);
xnor U3517 (N_3517,N_3297,N_3207);
nand U3518 (N_3518,N_3214,N_3356);
nor U3519 (N_3519,N_3321,N_3299);
or U3520 (N_3520,N_3466,N_3363);
xor U3521 (N_3521,N_3465,N_3391);
nand U3522 (N_3522,N_3386,N_3468);
nand U3523 (N_3523,N_3410,N_3360);
nor U3524 (N_3524,N_3500,N_3473);
nand U3525 (N_3525,N_3477,N_3372);
and U3526 (N_3526,N_3417,N_3446);
xor U3527 (N_3527,N_3416,N_3368);
nor U3528 (N_3528,N_3402,N_3380);
xor U3529 (N_3529,N_3451,N_3482);
xor U3530 (N_3530,N_3361,N_3415);
nor U3531 (N_3531,N_3432,N_3405);
or U3532 (N_3532,N_3491,N_3404);
or U3533 (N_3533,N_3429,N_3454);
nand U3534 (N_3534,N_3371,N_3367);
nand U3535 (N_3535,N_3495,N_3407);
nand U3536 (N_3536,N_3448,N_3467);
or U3537 (N_3537,N_3397,N_3508);
nor U3538 (N_3538,N_3369,N_3438);
xor U3539 (N_3539,N_3471,N_3479);
or U3540 (N_3540,N_3437,N_3506);
nand U3541 (N_3541,N_3488,N_3374);
xor U3542 (N_3542,N_3449,N_3444);
nand U3543 (N_3543,N_3411,N_3489);
nand U3544 (N_3544,N_3445,N_3392);
xnor U3545 (N_3545,N_3375,N_3514);
or U3546 (N_3546,N_3396,N_3409);
or U3547 (N_3547,N_3431,N_3439);
nand U3548 (N_3548,N_3426,N_3510);
xnor U3549 (N_3549,N_3377,N_3502);
nor U3550 (N_3550,N_3399,N_3455);
nand U3551 (N_3551,N_3378,N_3494);
and U3552 (N_3552,N_3475,N_3383);
or U3553 (N_3553,N_3370,N_3428);
nand U3554 (N_3554,N_3458,N_3453);
or U3555 (N_3555,N_3464,N_3517);
and U3556 (N_3556,N_3513,N_3456);
or U3557 (N_3557,N_3503,N_3376);
nand U3558 (N_3558,N_3390,N_3447);
or U3559 (N_3559,N_3459,N_3476);
nor U3560 (N_3560,N_3393,N_3486);
xnor U3561 (N_3561,N_3507,N_3373);
xnor U3562 (N_3562,N_3496,N_3450);
nand U3563 (N_3563,N_3457,N_3501);
nand U3564 (N_3564,N_3497,N_3434);
and U3565 (N_3565,N_3519,N_3385);
nor U3566 (N_3566,N_3420,N_3460);
or U3567 (N_3567,N_3505,N_3483);
xnor U3568 (N_3568,N_3461,N_3427);
nor U3569 (N_3569,N_3425,N_3487);
and U3570 (N_3570,N_3480,N_3462);
xnor U3571 (N_3571,N_3436,N_3400);
and U3572 (N_3572,N_3443,N_3413);
nor U3573 (N_3573,N_3463,N_3504);
nor U3574 (N_3574,N_3384,N_3511);
nor U3575 (N_3575,N_3516,N_3469);
or U3576 (N_3576,N_3419,N_3493);
and U3577 (N_3577,N_3435,N_3379);
nor U3578 (N_3578,N_3509,N_3498);
nand U3579 (N_3579,N_3403,N_3470);
nor U3580 (N_3580,N_3387,N_3422);
xor U3581 (N_3581,N_3364,N_3366);
nand U3582 (N_3582,N_3414,N_3382);
xor U3583 (N_3583,N_3484,N_3430);
xor U3584 (N_3584,N_3472,N_3492);
or U3585 (N_3585,N_3398,N_3395);
nor U3586 (N_3586,N_3452,N_3442);
xnor U3587 (N_3587,N_3418,N_3515);
or U3588 (N_3588,N_3440,N_3362);
and U3589 (N_3589,N_3394,N_3441);
xor U3590 (N_3590,N_3424,N_3499);
and U3591 (N_3591,N_3412,N_3481);
xor U3592 (N_3592,N_3423,N_3518);
nand U3593 (N_3593,N_3381,N_3401);
nand U3594 (N_3594,N_3388,N_3490);
nor U3595 (N_3595,N_3421,N_3365);
nand U3596 (N_3596,N_3512,N_3433);
nand U3597 (N_3597,N_3406,N_3408);
and U3598 (N_3598,N_3478,N_3474);
nor U3599 (N_3599,N_3389,N_3485);
or U3600 (N_3600,N_3408,N_3385);
nor U3601 (N_3601,N_3478,N_3378);
xor U3602 (N_3602,N_3496,N_3414);
or U3603 (N_3603,N_3487,N_3415);
or U3604 (N_3604,N_3375,N_3414);
nor U3605 (N_3605,N_3363,N_3416);
nand U3606 (N_3606,N_3449,N_3496);
or U3607 (N_3607,N_3413,N_3427);
nor U3608 (N_3608,N_3428,N_3498);
xnor U3609 (N_3609,N_3504,N_3506);
and U3610 (N_3610,N_3478,N_3407);
xor U3611 (N_3611,N_3455,N_3373);
nor U3612 (N_3612,N_3409,N_3478);
nand U3613 (N_3613,N_3404,N_3394);
nor U3614 (N_3614,N_3481,N_3479);
nor U3615 (N_3615,N_3406,N_3385);
nand U3616 (N_3616,N_3409,N_3388);
nand U3617 (N_3617,N_3490,N_3360);
nor U3618 (N_3618,N_3380,N_3516);
nor U3619 (N_3619,N_3519,N_3438);
xnor U3620 (N_3620,N_3444,N_3447);
nand U3621 (N_3621,N_3463,N_3515);
nand U3622 (N_3622,N_3425,N_3446);
or U3623 (N_3623,N_3435,N_3462);
and U3624 (N_3624,N_3452,N_3408);
nor U3625 (N_3625,N_3505,N_3423);
or U3626 (N_3626,N_3447,N_3506);
nor U3627 (N_3627,N_3373,N_3426);
xor U3628 (N_3628,N_3402,N_3395);
nor U3629 (N_3629,N_3477,N_3486);
xnor U3630 (N_3630,N_3388,N_3421);
xor U3631 (N_3631,N_3371,N_3361);
xnor U3632 (N_3632,N_3466,N_3455);
and U3633 (N_3633,N_3499,N_3459);
nand U3634 (N_3634,N_3477,N_3472);
nor U3635 (N_3635,N_3518,N_3453);
xnor U3636 (N_3636,N_3395,N_3485);
and U3637 (N_3637,N_3508,N_3453);
or U3638 (N_3638,N_3399,N_3479);
and U3639 (N_3639,N_3442,N_3481);
xnor U3640 (N_3640,N_3475,N_3420);
or U3641 (N_3641,N_3376,N_3360);
nor U3642 (N_3642,N_3389,N_3493);
and U3643 (N_3643,N_3443,N_3464);
nand U3644 (N_3644,N_3430,N_3409);
nand U3645 (N_3645,N_3466,N_3378);
or U3646 (N_3646,N_3480,N_3390);
or U3647 (N_3647,N_3380,N_3360);
or U3648 (N_3648,N_3406,N_3490);
and U3649 (N_3649,N_3510,N_3518);
and U3650 (N_3650,N_3500,N_3426);
nand U3651 (N_3651,N_3446,N_3458);
nor U3652 (N_3652,N_3383,N_3390);
or U3653 (N_3653,N_3495,N_3454);
or U3654 (N_3654,N_3493,N_3426);
nor U3655 (N_3655,N_3499,N_3471);
nor U3656 (N_3656,N_3415,N_3479);
nor U3657 (N_3657,N_3362,N_3450);
nor U3658 (N_3658,N_3503,N_3409);
or U3659 (N_3659,N_3399,N_3431);
nor U3660 (N_3660,N_3364,N_3439);
and U3661 (N_3661,N_3499,N_3503);
nand U3662 (N_3662,N_3407,N_3493);
and U3663 (N_3663,N_3456,N_3493);
nand U3664 (N_3664,N_3438,N_3444);
or U3665 (N_3665,N_3484,N_3373);
xnor U3666 (N_3666,N_3397,N_3401);
nor U3667 (N_3667,N_3463,N_3364);
or U3668 (N_3668,N_3409,N_3473);
or U3669 (N_3669,N_3472,N_3460);
and U3670 (N_3670,N_3411,N_3479);
xnor U3671 (N_3671,N_3516,N_3430);
nor U3672 (N_3672,N_3478,N_3369);
and U3673 (N_3673,N_3479,N_3398);
xor U3674 (N_3674,N_3420,N_3446);
and U3675 (N_3675,N_3450,N_3431);
nand U3676 (N_3676,N_3517,N_3442);
or U3677 (N_3677,N_3413,N_3498);
and U3678 (N_3678,N_3480,N_3393);
xor U3679 (N_3679,N_3493,N_3483);
and U3680 (N_3680,N_3638,N_3559);
nor U3681 (N_3681,N_3612,N_3616);
nand U3682 (N_3682,N_3552,N_3597);
and U3683 (N_3683,N_3540,N_3579);
and U3684 (N_3684,N_3541,N_3549);
or U3685 (N_3685,N_3642,N_3520);
nor U3686 (N_3686,N_3652,N_3627);
nand U3687 (N_3687,N_3610,N_3626);
nor U3688 (N_3688,N_3600,N_3560);
or U3689 (N_3689,N_3528,N_3548);
or U3690 (N_3690,N_3584,N_3524);
nor U3691 (N_3691,N_3654,N_3662);
or U3692 (N_3692,N_3608,N_3580);
nor U3693 (N_3693,N_3525,N_3550);
xnor U3694 (N_3694,N_3633,N_3635);
xnor U3695 (N_3695,N_3545,N_3583);
or U3696 (N_3696,N_3533,N_3565);
nand U3697 (N_3697,N_3667,N_3581);
or U3698 (N_3698,N_3615,N_3531);
or U3699 (N_3699,N_3539,N_3669);
nor U3700 (N_3700,N_3598,N_3561);
nor U3701 (N_3701,N_3587,N_3521);
nand U3702 (N_3702,N_3606,N_3529);
nor U3703 (N_3703,N_3641,N_3535);
nor U3704 (N_3704,N_3611,N_3653);
nand U3705 (N_3705,N_3640,N_3673);
or U3706 (N_3706,N_3630,N_3646);
or U3707 (N_3707,N_3596,N_3574);
nor U3708 (N_3708,N_3647,N_3607);
xnor U3709 (N_3709,N_3601,N_3672);
nor U3710 (N_3710,N_3563,N_3588);
and U3711 (N_3711,N_3621,N_3553);
and U3712 (N_3712,N_3655,N_3522);
and U3713 (N_3713,N_3547,N_3567);
xnor U3714 (N_3714,N_3677,N_3542);
nand U3715 (N_3715,N_3523,N_3644);
nor U3716 (N_3716,N_3544,N_3631);
and U3717 (N_3717,N_3656,N_3634);
and U3718 (N_3718,N_3557,N_3603);
and U3719 (N_3719,N_3623,N_3632);
nand U3720 (N_3720,N_3532,N_3613);
or U3721 (N_3721,N_3594,N_3566);
nor U3722 (N_3722,N_3671,N_3675);
nand U3723 (N_3723,N_3617,N_3593);
nor U3724 (N_3724,N_3624,N_3658);
xnor U3725 (N_3725,N_3551,N_3649);
and U3726 (N_3726,N_3629,N_3537);
nand U3727 (N_3727,N_3605,N_3586);
and U3728 (N_3728,N_3538,N_3674);
nor U3729 (N_3729,N_3555,N_3679);
nor U3730 (N_3730,N_3534,N_3546);
xnor U3731 (N_3731,N_3657,N_3558);
nor U3732 (N_3732,N_3628,N_3576);
and U3733 (N_3733,N_3573,N_3575);
or U3734 (N_3734,N_3591,N_3651);
and U3735 (N_3735,N_3637,N_3636);
nand U3736 (N_3736,N_3670,N_3582);
nor U3737 (N_3737,N_3570,N_3625);
or U3738 (N_3738,N_3664,N_3622);
and U3739 (N_3739,N_3556,N_3543);
and U3740 (N_3740,N_3645,N_3530);
and U3741 (N_3741,N_3578,N_3668);
and U3742 (N_3742,N_3663,N_3659);
xnor U3743 (N_3743,N_3585,N_3660);
and U3744 (N_3744,N_3618,N_3595);
or U3745 (N_3745,N_3536,N_3648);
or U3746 (N_3746,N_3562,N_3602);
xor U3747 (N_3747,N_3572,N_3650);
xnor U3748 (N_3748,N_3527,N_3620);
xnor U3749 (N_3749,N_3589,N_3665);
nor U3750 (N_3750,N_3577,N_3526);
nor U3751 (N_3751,N_3678,N_3661);
nand U3752 (N_3752,N_3609,N_3639);
nor U3753 (N_3753,N_3590,N_3614);
and U3754 (N_3754,N_3554,N_3564);
or U3755 (N_3755,N_3619,N_3571);
or U3756 (N_3756,N_3643,N_3568);
xnor U3757 (N_3757,N_3666,N_3569);
or U3758 (N_3758,N_3604,N_3599);
xnor U3759 (N_3759,N_3592,N_3676);
xor U3760 (N_3760,N_3582,N_3645);
xor U3761 (N_3761,N_3657,N_3543);
nor U3762 (N_3762,N_3603,N_3591);
xor U3763 (N_3763,N_3588,N_3543);
or U3764 (N_3764,N_3555,N_3576);
xnor U3765 (N_3765,N_3525,N_3538);
nand U3766 (N_3766,N_3537,N_3677);
or U3767 (N_3767,N_3617,N_3532);
xnor U3768 (N_3768,N_3550,N_3574);
nand U3769 (N_3769,N_3671,N_3640);
nor U3770 (N_3770,N_3564,N_3584);
nand U3771 (N_3771,N_3534,N_3574);
or U3772 (N_3772,N_3577,N_3640);
nand U3773 (N_3773,N_3538,N_3676);
nand U3774 (N_3774,N_3653,N_3549);
nand U3775 (N_3775,N_3531,N_3596);
and U3776 (N_3776,N_3639,N_3520);
or U3777 (N_3777,N_3636,N_3559);
and U3778 (N_3778,N_3550,N_3598);
nor U3779 (N_3779,N_3595,N_3614);
nor U3780 (N_3780,N_3531,N_3631);
and U3781 (N_3781,N_3635,N_3571);
or U3782 (N_3782,N_3526,N_3542);
and U3783 (N_3783,N_3522,N_3611);
xnor U3784 (N_3784,N_3622,N_3528);
nor U3785 (N_3785,N_3540,N_3527);
or U3786 (N_3786,N_3623,N_3555);
and U3787 (N_3787,N_3656,N_3530);
xnor U3788 (N_3788,N_3571,N_3582);
xor U3789 (N_3789,N_3634,N_3599);
xnor U3790 (N_3790,N_3543,N_3612);
xnor U3791 (N_3791,N_3524,N_3540);
xor U3792 (N_3792,N_3678,N_3535);
nor U3793 (N_3793,N_3676,N_3525);
xor U3794 (N_3794,N_3654,N_3561);
and U3795 (N_3795,N_3674,N_3534);
nand U3796 (N_3796,N_3537,N_3651);
or U3797 (N_3797,N_3630,N_3579);
nor U3798 (N_3798,N_3615,N_3671);
nor U3799 (N_3799,N_3573,N_3558);
and U3800 (N_3800,N_3638,N_3535);
or U3801 (N_3801,N_3633,N_3589);
or U3802 (N_3802,N_3655,N_3529);
nand U3803 (N_3803,N_3581,N_3642);
and U3804 (N_3804,N_3584,N_3672);
nand U3805 (N_3805,N_3617,N_3636);
xor U3806 (N_3806,N_3662,N_3656);
nor U3807 (N_3807,N_3593,N_3538);
or U3808 (N_3808,N_3609,N_3585);
nand U3809 (N_3809,N_3608,N_3630);
and U3810 (N_3810,N_3550,N_3541);
xnor U3811 (N_3811,N_3626,N_3584);
xor U3812 (N_3812,N_3622,N_3577);
or U3813 (N_3813,N_3555,N_3672);
nor U3814 (N_3814,N_3541,N_3646);
nor U3815 (N_3815,N_3677,N_3670);
nor U3816 (N_3816,N_3548,N_3664);
and U3817 (N_3817,N_3624,N_3559);
nand U3818 (N_3818,N_3535,N_3589);
and U3819 (N_3819,N_3546,N_3637);
nor U3820 (N_3820,N_3642,N_3671);
xnor U3821 (N_3821,N_3652,N_3663);
and U3822 (N_3822,N_3635,N_3600);
nor U3823 (N_3823,N_3604,N_3650);
nor U3824 (N_3824,N_3573,N_3560);
or U3825 (N_3825,N_3671,N_3529);
and U3826 (N_3826,N_3561,N_3551);
and U3827 (N_3827,N_3566,N_3637);
and U3828 (N_3828,N_3595,N_3607);
or U3829 (N_3829,N_3572,N_3604);
nor U3830 (N_3830,N_3587,N_3580);
nor U3831 (N_3831,N_3556,N_3562);
and U3832 (N_3832,N_3549,N_3584);
or U3833 (N_3833,N_3658,N_3583);
nor U3834 (N_3834,N_3606,N_3679);
or U3835 (N_3835,N_3594,N_3553);
and U3836 (N_3836,N_3661,N_3613);
nand U3837 (N_3837,N_3646,N_3647);
nand U3838 (N_3838,N_3631,N_3660);
nor U3839 (N_3839,N_3585,N_3616);
nand U3840 (N_3840,N_3739,N_3777);
nand U3841 (N_3841,N_3826,N_3808);
nand U3842 (N_3842,N_3695,N_3815);
nand U3843 (N_3843,N_3834,N_3697);
or U3844 (N_3844,N_3779,N_3776);
nand U3845 (N_3845,N_3820,N_3747);
nor U3846 (N_3846,N_3713,N_3728);
or U3847 (N_3847,N_3734,N_3833);
or U3848 (N_3848,N_3788,N_3839);
nand U3849 (N_3849,N_3759,N_3832);
nor U3850 (N_3850,N_3787,N_3763);
and U3851 (N_3851,N_3757,N_3723);
nor U3852 (N_3852,N_3748,N_3824);
nor U3853 (N_3853,N_3708,N_3794);
nand U3854 (N_3854,N_3680,N_3838);
nand U3855 (N_3855,N_3692,N_3689);
and U3856 (N_3856,N_3827,N_3807);
and U3857 (N_3857,N_3720,N_3732);
nand U3858 (N_3858,N_3740,N_3704);
nor U3859 (N_3859,N_3780,N_3684);
nor U3860 (N_3860,N_3831,N_3786);
xnor U3861 (N_3861,N_3690,N_3691);
and U3862 (N_3862,N_3836,N_3792);
or U3863 (N_3863,N_3770,N_3712);
nand U3864 (N_3864,N_3778,N_3722);
nor U3865 (N_3865,N_3781,N_3715);
nor U3866 (N_3866,N_3765,N_3819);
xor U3867 (N_3867,N_3764,N_3750);
and U3868 (N_3868,N_3731,N_3791);
xnor U3869 (N_3869,N_3823,N_3798);
and U3870 (N_3870,N_3774,N_3802);
nor U3871 (N_3871,N_3800,N_3804);
nand U3872 (N_3872,N_3741,N_3737);
nor U3873 (N_3873,N_3688,N_3789);
or U3874 (N_3874,N_3809,N_3822);
nand U3875 (N_3875,N_3761,N_3727);
nand U3876 (N_3876,N_3711,N_3771);
and U3877 (N_3877,N_3795,N_3736);
nand U3878 (N_3878,N_3810,N_3726);
and U3879 (N_3879,N_3801,N_3714);
xor U3880 (N_3880,N_3694,N_3796);
xor U3881 (N_3881,N_3706,N_3814);
or U3882 (N_3882,N_3783,N_3830);
nand U3883 (N_3883,N_3721,N_3698);
nand U3884 (N_3884,N_3835,N_3773);
xnor U3885 (N_3885,N_3805,N_3710);
nand U3886 (N_3886,N_3701,N_3735);
nor U3887 (N_3887,N_3828,N_3754);
xnor U3888 (N_3888,N_3769,N_3816);
nor U3889 (N_3889,N_3725,N_3719);
or U3890 (N_3890,N_3745,N_3752);
and U3891 (N_3891,N_3782,N_3790);
and U3892 (N_3892,N_3775,N_3813);
and U3893 (N_3893,N_3756,N_3829);
and U3894 (N_3894,N_3716,N_3811);
and U3895 (N_3895,N_3793,N_3705);
nor U3896 (N_3896,N_3803,N_3733);
and U3897 (N_3897,N_3766,N_3785);
nand U3898 (N_3898,N_3758,N_3742);
nor U3899 (N_3899,N_3753,N_3784);
nor U3900 (N_3900,N_3700,N_3709);
and U3901 (N_3901,N_3738,N_3696);
xnor U3902 (N_3902,N_3730,N_3703);
or U3903 (N_3903,N_3825,N_3812);
nand U3904 (N_3904,N_3767,N_3686);
xor U3905 (N_3905,N_3682,N_3718);
nand U3906 (N_3906,N_3751,N_3729);
nor U3907 (N_3907,N_3685,N_3702);
or U3908 (N_3908,N_3724,N_3693);
nor U3909 (N_3909,N_3749,N_3699);
or U3910 (N_3910,N_3821,N_3760);
nand U3911 (N_3911,N_3799,N_3772);
xnor U3912 (N_3912,N_3707,N_3717);
nor U3913 (N_3913,N_3837,N_3806);
nand U3914 (N_3914,N_3818,N_3797);
or U3915 (N_3915,N_3762,N_3683);
and U3916 (N_3916,N_3744,N_3817);
nor U3917 (N_3917,N_3768,N_3746);
nand U3918 (N_3918,N_3687,N_3743);
nand U3919 (N_3919,N_3681,N_3755);
nor U3920 (N_3920,N_3810,N_3706);
nor U3921 (N_3921,N_3700,N_3698);
nand U3922 (N_3922,N_3805,N_3764);
nor U3923 (N_3923,N_3685,N_3726);
nand U3924 (N_3924,N_3810,N_3762);
nor U3925 (N_3925,N_3771,N_3784);
xnor U3926 (N_3926,N_3705,N_3753);
nand U3927 (N_3927,N_3731,N_3801);
and U3928 (N_3928,N_3732,N_3711);
xnor U3929 (N_3929,N_3777,N_3831);
and U3930 (N_3930,N_3698,N_3815);
nor U3931 (N_3931,N_3803,N_3696);
nor U3932 (N_3932,N_3752,N_3808);
or U3933 (N_3933,N_3793,N_3776);
and U3934 (N_3934,N_3773,N_3782);
and U3935 (N_3935,N_3789,N_3724);
nand U3936 (N_3936,N_3837,N_3748);
or U3937 (N_3937,N_3723,N_3754);
or U3938 (N_3938,N_3814,N_3821);
and U3939 (N_3939,N_3683,N_3786);
xor U3940 (N_3940,N_3721,N_3717);
nor U3941 (N_3941,N_3714,N_3823);
and U3942 (N_3942,N_3699,N_3713);
nand U3943 (N_3943,N_3757,N_3783);
and U3944 (N_3944,N_3709,N_3838);
xnor U3945 (N_3945,N_3788,N_3686);
nor U3946 (N_3946,N_3737,N_3798);
nand U3947 (N_3947,N_3689,N_3746);
or U3948 (N_3948,N_3700,N_3699);
or U3949 (N_3949,N_3764,N_3752);
nor U3950 (N_3950,N_3730,N_3833);
nor U3951 (N_3951,N_3821,N_3724);
nor U3952 (N_3952,N_3696,N_3839);
or U3953 (N_3953,N_3720,N_3771);
nand U3954 (N_3954,N_3692,N_3814);
nand U3955 (N_3955,N_3756,N_3741);
and U3956 (N_3956,N_3706,N_3807);
xnor U3957 (N_3957,N_3685,N_3696);
xnor U3958 (N_3958,N_3765,N_3731);
nand U3959 (N_3959,N_3748,N_3702);
and U3960 (N_3960,N_3726,N_3710);
and U3961 (N_3961,N_3750,N_3780);
and U3962 (N_3962,N_3710,N_3713);
nand U3963 (N_3963,N_3816,N_3753);
and U3964 (N_3964,N_3725,N_3716);
nand U3965 (N_3965,N_3793,N_3722);
xnor U3966 (N_3966,N_3816,N_3754);
and U3967 (N_3967,N_3752,N_3741);
and U3968 (N_3968,N_3737,N_3758);
nor U3969 (N_3969,N_3750,N_3823);
or U3970 (N_3970,N_3710,N_3753);
nor U3971 (N_3971,N_3769,N_3830);
nor U3972 (N_3972,N_3832,N_3804);
nor U3973 (N_3973,N_3695,N_3682);
xor U3974 (N_3974,N_3726,N_3714);
nand U3975 (N_3975,N_3829,N_3696);
nand U3976 (N_3976,N_3780,N_3710);
xor U3977 (N_3977,N_3778,N_3835);
nor U3978 (N_3978,N_3756,N_3806);
xnor U3979 (N_3979,N_3787,N_3772);
nor U3980 (N_3980,N_3818,N_3798);
xor U3981 (N_3981,N_3784,N_3713);
xnor U3982 (N_3982,N_3760,N_3750);
nand U3983 (N_3983,N_3699,N_3711);
and U3984 (N_3984,N_3728,N_3818);
nor U3985 (N_3985,N_3785,N_3798);
xnor U3986 (N_3986,N_3735,N_3739);
nand U3987 (N_3987,N_3721,N_3827);
xnor U3988 (N_3988,N_3756,N_3766);
or U3989 (N_3989,N_3751,N_3773);
and U3990 (N_3990,N_3717,N_3749);
nand U3991 (N_3991,N_3796,N_3700);
xor U3992 (N_3992,N_3729,N_3808);
and U3993 (N_3993,N_3766,N_3800);
nor U3994 (N_3994,N_3718,N_3824);
nand U3995 (N_3995,N_3716,N_3741);
or U3996 (N_3996,N_3738,N_3785);
nand U3997 (N_3997,N_3774,N_3825);
nand U3998 (N_3998,N_3705,N_3803);
or U3999 (N_3999,N_3749,N_3789);
nor U4000 (N_4000,N_3996,N_3884);
and U4001 (N_4001,N_3912,N_3991);
nand U4002 (N_4002,N_3863,N_3989);
nand U4003 (N_4003,N_3887,N_3964);
or U4004 (N_4004,N_3979,N_3876);
nand U4005 (N_4005,N_3971,N_3921);
or U4006 (N_4006,N_3847,N_3853);
or U4007 (N_4007,N_3990,N_3875);
xor U4008 (N_4008,N_3981,N_3942);
nor U4009 (N_4009,N_3848,N_3877);
nand U4010 (N_4010,N_3856,N_3886);
or U4011 (N_4011,N_3901,N_3963);
xnor U4012 (N_4012,N_3986,N_3854);
or U4013 (N_4013,N_3920,N_3915);
and U4014 (N_4014,N_3843,N_3992);
nor U4015 (N_4015,N_3926,N_3943);
nor U4016 (N_4016,N_3902,N_3850);
or U4017 (N_4017,N_3894,N_3871);
or U4018 (N_4018,N_3851,N_3952);
nor U4019 (N_4019,N_3862,N_3881);
nand U4020 (N_4020,N_3883,N_3983);
nand U4021 (N_4021,N_3978,N_3977);
and U4022 (N_4022,N_3919,N_3914);
or U4023 (N_4023,N_3845,N_3932);
or U4024 (N_4024,N_3903,N_3842);
xnor U4025 (N_4025,N_3951,N_3997);
or U4026 (N_4026,N_3947,N_3861);
nor U4027 (N_4027,N_3878,N_3959);
nor U4028 (N_4028,N_3999,N_3998);
and U4029 (N_4029,N_3950,N_3905);
xnor U4030 (N_4030,N_3893,N_3958);
xor U4031 (N_4031,N_3962,N_3873);
nand U4032 (N_4032,N_3841,N_3867);
nand U4033 (N_4033,N_3872,N_3895);
and U4034 (N_4034,N_3885,N_3944);
xor U4035 (N_4035,N_3890,N_3935);
nor U4036 (N_4036,N_3972,N_3868);
nand U4037 (N_4037,N_3953,N_3938);
or U4038 (N_4038,N_3975,N_3954);
nand U4039 (N_4039,N_3858,N_3968);
xnor U4040 (N_4040,N_3846,N_3980);
nand U4041 (N_4041,N_3866,N_3945);
and U4042 (N_4042,N_3922,N_3948);
nand U4043 (N_4043,N_3987,N_3900);
and U4044 (N_4044,N_3949,N_3988);
or U4045 (N_4045,N_3936,N_3995);
nand U4046 (N_4046,N_3940,N_3907);
nor U4047 (N_4047,N_3882,N_3870);
nand U4048 (N_4048,N_3840,N_3925);
nor U4049 (N_4049,N_3984,N_3974);
and U4050 (N_4050,N_3865,N_3928);
xor U4051 (N_4051,N_3898,N_3916);
xnor U4052 (N_4052,N_3946,N_3906);
and U4053 (N_4053,N_3879,N_3924);
nor U4054 (N_4054,N_3930,N_3957);
nand U4055 (N_4055,N_3860,N_3880);
and U4056 (N_4056,N_3888,N_3970);
nand U4057 (N_4057,N_3955,N_3909);
and U4058 (N_4058,N_3849,N_3956);
and U4059 (N_4059,N_3966,N_3982);
xnor U4060 (N_4060,N_3976,N_3859);
nor U4061 (N_4061,N_3904,N_3985);
nand U4062 (N_4062,N_3913,N_3933);
nor U4063 (N_4063,N_3896,N_3960);
or U4064 (N_4064,N_3891,N_3973);
nor U4065 (N_4065,N_3939,N_3937);
or U4066 (N_4066,N_3929,N_3993);
xor U4067 (N_4067,N_3918,N_3889);
nand U4068 (N_4068,N_3844,N_3899);
nand U4069 (N_4069,N_3857,N_3961);
nor U4070 (N_4070,N_3931,N_3994);
nor U4071 (N_4071,N_3941,N_3917);
or U4072 (N_4072,N_3855,N_3874);
or U4073 (N_4073,N_3892,N_3965);
nor U4074 (N_4074,N_3908,N_3852);
or U4075 (N_4075,N_3927,N_3910);
nand U4076 (N_4076,N_3934,N_3864);
xnor U4077 (N_4077,N_3923,N_3897);
nand U4078 (N_4078,N_3869,N_3967);
xnor U4079 (N_4079,N_3911,N_3969);
nor U4080 (N_4080,N_3944,N_3866);
nor U4081 (N_4081,N_3851,N_3937);
or U4082 (N_4082,N_3957,N_3872);
nand U4083 (N_4083,N_3988,N_3922);
and U4084 (N_4084,N_3844,N_3984);
nand U4085 (N_4085,N_3866,N_3931);
nor U4086 (N_4086,N_3875,N_3976);
nor U4087 (N_4087,N_3949,N_3924);
nand U4088 (N_4088,N_3929,N_3941);
or U4089 (N_4089,N_3928,N_3965);
xnor U4090 (N_4090,N_3879,N_3996);
nand U4091 (N_4091,N_3987,N_3903);
and U4092 (N_4092,N_3891,N_3994);
or U4093 (N_4093,N_3946,N_3993);
and U4094 (N_4094,N_3984,N_3895);
nand U4095 (N_4095,N_3840,N_3993);
nand U4096 (N_4096,N_3999,N_3936);
xnor U4097 (N_4097,N_3999,N_3971);
or U4098 (N_4098,N_3971,N_3919);
nor U4099 (N_4099,N_3907,N_3934);
nand U4100 (N_4100,N_3866,N_3971);
or U4101 (N_4101,N_3910,N_3867);
nand U4102 (N_4102,N_3924,N_3982);
nand U4103 (N_4103,N_3854,N_3968);
and U4104 (N_4104,N_3853,N_3991);
nand U4105 (N_4105,N_3853,N_3972);
xnor U4106 (N_4106,N_3877,N_3875);
and U4107 (N_4107,N_3908,N_3939);
or U4108 (N_4108,N_3852,N_3891);
nor U4109 (N_4109,N_3927,N_3860);
and U4110 (N_4110,N_3937,N_3980);
and U4111 (N_4111,N_3875,N_3893);
xnor U4112 (N_4112,N_3934,N_3997);
and U4113 (N_4113,N_3911,N_3856);
xnor U4114 (N_4114,N_3959,N_3939);
and U4115 (N_4115,N_3898,N_3891);
or U4116 (N_4116,N_3894,N_3903);
nand U4117 (N_4117,N_3855,N_3977);
nand U4118 (N_4118,N_3861,N_3989);
or U4119 (N_4119,N_3969,N_3848);
or U4120 (N_4120,N_3948,N_3853);
nand U4121 (N_4121,N_3907,N_3880);
or U4122 (N_4122,N_3923,N_3919);
nand U4123 (N_4123,N_3876,N_3924);
nor U4124 (N_4124,N_3909,N_3929);
nand U4125 (N_4125,N_3879,N_3925);
nor U4126 (N_4126,N_3928,N_3873);
xnor U4127 (N_4127,N_3960,N_3953);
and U4128 (N_4128,N_3860,N_3980);
nor U4129 (N_4129,N_3963,N_3993);
xnor U4130 (N_4130,N_3953,N_3915);
and U4131 (N_4131,N_3988,N_3916);
or U4132 (N_4132,N_3873,N_3965);
nand U4133 (N_4133,N_3941,N_3973);
nor U4134 (N_4134,N_3849,N_3843);
nor U4135 (N_4135,N_3966,N_3905);
xor U4136 (N_4136,N_3906,N_3866);
or U4137 (N_4137,N_3987,N_3930);
or U4138 (N_4138,N_3921,N_3962);
and U4139 (N_4139,N_3902,N_3905);
nor U4140 (N_4140,N_3848,N_3855);
nand U4141 (N_4141,N_3901,N_3941);
xor U4142 (N_4142,N_3889,N_3938);
nor U4143 (N_4143,N_3979,N_3956);
nor U4144 (N_4144,N_3871,N_3951);
nand U4145 (N_4145,N_3957,N_3934);
nand U4146 (N_4146,N_3926,N_3997);
xor U4147 (N_4147,N_3956,N_3843);
or U4148 (N_4148,N_3863,N_3900);
and U4149 (N_4149,N_3910,N_3946);
nor U4150 (N_4150,N_3974,N_3988);
and U4151 (N_4151,N_3877,N_3969);
nand U4152 (N_4152,N_3923,N_3925);
or U4153 (N_4153,N_3999,N_3876);
or U4154 (N_4154,N_3951,N_3987);
or U4155 (N_4155,N_3938,N_3959);
nand U4156 (N_4156,N_3871,N_3937);
or U4157 (N_4157,N_3861,N_3844);
xor U4158 (N_4158,N_3957,N_3881);
xor U4159 (N_4159,N_3911,N_3956);
xor U4160 (N_4160,N_4088,N_4019);
and U4161 (N_4161,N_4128,N_4090);
and U4162 (N_4162,N_4077,N_4076);
nand U4163 (N_4163,N_4105,N_4124);
nand U4164 (N_4164,N_4007,N_4002);
xnor U4165 (N_4165,N_4149,N_4006);
or U4166 (N_4166,N_4009,N_4156);
and U4167 (N_4167,N_4049,N_4152);
xor U4168 (N_4168,N_4089,N_4092);
and U4169 (N_4169,N_4091,N_4146);
and U4170 (N_4170,N_4079,N_4022);
or U4171 (N_4171,N_4071,N_4108);
or U4172 (N_4172,N_4129,N_4078);
and U4173 (N_4173,N_4042,N_4011);
nor U4174 (N_4174,N_4017,N_4093);
nand U4175 (N_4175,N_4046,N_4066);
or U4176 (N_4176,N_4104,N_4056);
xor U4177 (N_4177,N_4125,N_4106);
nand U4178 (N_4178,N_4113,N_4060);
or U4179 (N_4179,N_4097,N_4121);
and U4180 (N_4180,N_4098,N_4032);
nor U4181 (N_4181,N_4118,N_4094);
nor U4182 (N_4182,N_4100,N_4029);
or U4183 (N_4183,N_4087,N_4127);
or U4184 (N_4184,N_4159,N_4158);
nand U4185 (N_4185,N_4034,N_4138);
and U4186 (N_4186,N_4052,N_4116);
xnor U4187 (N_4187,N_4024,N_4144);
xor U4188 (N_4188,N_4039,N_4120);
xor U4189 (N_4189,N_4036,N_4123);
or U4190 (N_4190,N_4148,N_4048);
xnor U4191 (N_4191,N_4139,N_4016);
xor U4192 (N_4192,N_4145,N_4083);
nand U4193 (N_4193,N_4101,N_4154);
xor U4194 (N_4194,N_4081,N_4050);
and U4195 (N_4195,N_4054,N_4045);
xnor U4196 (N_4196,N_4119,N_4080);
nor U4197 (N_4197,N_4133,N_4044);
and U4198 (N_4198,N_4131,N_4020);
or U4199 (N_4199,N_4137,N_4059);
nor U4200 (N_4200,N_4040,N_4103);
nand U4201 (N_4201,N_4150,N_4115);
nand U4202 (N_4202,N_4063,N_4099);
or U4203 (N_4203,N_4065,N_4111);
nand U4204 (N_4204,N_4010,N_4110);
xor U4205 (N_4205,N_4140,N_4025);
xor U4206 (N_4206,N_4096,N_4068);
xnor U4207 (N_4207,N_4155,N_4073);
and U4208 (N_4208,N_4109,N_4122);
xor U4209 (N_4209,N_4082,N_4058);
nand U4210 (N_4210,N_4041,N_4037);
or U4211 (N_4211,N_4153,N_4107);
xor U4212 (N_4212,N_4134,N_4057);
and U4213 (N_4213,N_4033,N_4067);
xor U4214 (N_4214,N_4051,N_4136);
or U4215 (N_4215,N_4074,N_4014);
nor U4216 (N_4216,N_4126,N_4013);
and U4217 (N_4217,N_4043,N_4064);
xnor U4218 (N_4218,N_4028,N_4004);
nand U4219 (N_4219,N_4085,N_4142);
nor U4220 (N_4220,N_4070,N_4021);
nand U4221 (N_4221,N_4069,N_4157);
and U4222 (N_4222,N_4143,N_4023);
xnor U4223 (N_4223,N_4095,N_4027);
nor U4224 (N_4224,N_4005,N_4001);
and U4225 (N_4225,N_4062,N_4047);
or U4226 (N_4226,N_4000,N_4075);
or U4227 (N_4227,N_4130,N_4061);
and U4228 (N_4228,N_4026,N_4084);
nor U4229 (N_4229,N_4117,N_4147);
xnor U4230 (N_4230,N_4141,N_4102);
nand U4231 (N_4231,N_4031,N_4030);
nand U4232 (N_4232,N_4035,N_4055);
or U4233 (N_4233,N_4053,N_4018);
nand U4234 (N_4234,N_4114,N_4003);
nand U4235 (N_4235,N_4072,N_4015);
and U4236 (N_4236,N_4135,N_4151);
xor U4237 (N_4237,N_4008,N_4112);
or U4238 (N_4238,N_4086,N_4132);
nand U4239 (N_4239,N_4012,N_4038);
nor U4240 (N_4240,N_4109,N_4105);
or U4241 (N_4241,N_4009,N_4074);
nand U4242 (N_4242,N_4071,N_4091);
xnor U4243 (N_4243,N_4038,N_4122);
nand U4244 (N_4244,N_4044,N_4057);
and U4245 (N_4245,N_4115,N_4071);
nand U4246 (N_4246,N_4141,N_4099);
xor U4247 (N_4247,N_4142,N_4132);
nand U4248 (N_4248,N_4141,N_4144);
and U4249 (N_4249,N_4099,N_4014);
nor U4250 (N_4250,N_4125,N_4094);
or U4251 (N_4251,N_4012,N_4152);
xor U4252 (N_4252,N_4093,N_4005);
nor U4253 (N_4253,N_4013,N_4082);
and U4254 (N_4254,N_4034,N_4067);
nand U4255 (N_4255,N_4135,N_4143);
xnor U4256 (N_4256,N_4034,N_4066);
and U4257 (N_4257,N_4016,N_4010);
or U4258 (N_4258,N_4003,N_4010);
or U4259 (N_4259,N_4103,N_4061);
and U4260 (N_4260,N_4015,N_4030);
and U4261 (N_4261,N_4028,N_4145);
and U4262 (N_4262,N_4088,N_4117);
xnor U4263 (N_4263,N_4104,N_4071);
and U4264 (N_4264,N_4059,N_4016);
and U4265 (N_4265,N_4145,N_4146);
or U4266 (N_4266,N_4156,N_4029);
or U4267 (N_4267,N_4155,N_4014);
xnor U4268 (N_4268,N_4132,N_4064);
or U4269 (N_4269,N_4034,N_4030);
and U4270 (N_4270,N_4050,N_4052);
and U4271 (N_4271,N_4017,N_4044);
nor U4272 (N_4272,N_4045,N_4099);
nor U4273 (N_4273,N_4158,N_4123);
nor U4274 (N_4274,N_4120,N_4109);
and U4275 (N_4275,N_4137,N_4072);
or U4276 (N_4276,N_4037,N_4064);
nor U4277 (N_4277,N_4079,N_4032);
xor U4278 (N_4278,N_4069,N_4093);
xor U4279 (N_4279,N_4010,N_4149);
xor U4280 (N_4280,N_4070,N_4113);
and U4281 (N_4281,N_4085,N_4077);
nor U4282 (N_4282,N_4086,N_4075);
or U4283 (N_4283,N_4100,N_4112);
or U4284 (N_4284,N_4076,N_4088);
nand U4285 (N_4285,N_4086,N_4100);
xor U4286 (N_4286,N_4031,N_4015);
and U4287 (N_4287,N_4135,N_4025);
or U4288 (N_4288,N_4083,N_4044);
or U4289 (N_4289,N_4097,N_4014);
xnor U4290 (N_4290,N_4044,N_4153);
and U4291 (N_4291,N_4139,N_4109);
or U4292 (N_4292,N_4090,N_4141);
xor U4293 (N_4293,N_4016,N_4137);
or U4294 (N_4294,N_4117,N_4142);
or U4295 (N_4295,N_4080,N_4113);
xnor U4296 (N_4296,N_4120,N_4084);
or U4297 (N_4297,N_4076,N_4082);
or U4298 (N_4298,N_4066,N_4068);
or U4299 (N_4299,N_4086,N_4078);
nand U4300 (N_4300,N_4159,N_4041);
nor U4301 (N_4301,N_4017,N_4154);
nor U4302 (N_4302,N_4051,N_4052);
or U4303 (N_4303,N_4031,N_4140);
or U4304 (N_4304,N_4041,N_4122);
xor U4305 (N_4305,N_4057,N_4005);
and U4306 (N_4306,N_4154,N_4087);
nand U4307 (N_4307,N_4081,N_4106);
and U4308 (N_4308,N_4150,N_4060);
xor U4309 (N_4309,N_4109,N_4099);
or U4310 (N_4310,N_4145,N_4131);
xor U4311 (N_4311,N_4084,N_4052);
or U4312 (N_4312,N_4048,N_4017);
xnor U4313 (N_4313,N_4087,N_4137);
or U4314 (N_4314,N_4016,N_4058);
nor U4315 (N_4315,N_4008,N_4152);
xor U4316 (N_4316,N_4092,N_4062);
nor U4317 (N_4317,N_4025,N_4152);
nor U4318 (N_4318,N_4089,N_4029);
or U4319 (N_4319,N_4111,N_4064);
nand U4320 (N_4320,N_4198,N_4256);
nand U4321 (N_4321,N_4222,N_4261);
and U4322 (N_4322,N_4253,N_4281);
nand U4323 (N_4323,N_4263,N_4269);
and U4324 (N_4324,N_4296,N_4235);
nor U4325 (N_4325,N_4208,N_4203);
or U4326 (N_4326,N_4291,N_4178);
xor U4327 (N_4327,N_4249,N_4276);
and U4328 (N_4328,N_4277,N_4307);
nor U4329 (N_4329,N_4248,N_4262);
or U4330 (N_4330,N_4241,N_4271);
nor U4331 (N_4331,N_4184,N_4251);
nand U4332 (N_4332,N_4314,N_4227);
xor U4333 (N_4333,N_4200,N_4225);
nand U4334 (N_4334,N_4245,N_4266);
or U4335 (N_4335,N_4302,N_4246);
nand U4336 (N_4336,N_4259,N_4176);
nand U4337 (N_4337,N_4247,N_4220);
nand U4338 (N_4338,N_4183,N_4228);
xor U4339 (N_4339,N_4181,N_4286);
nor U4340 (N_4340,N_4289,N_4257);
or U4341 (N_4341,N_4308,N_4299);
xnor U4342 (N_4342,N_4219,N_4311);
or U4343 (N_4343,N_4309,N_4167);
or U4344 (N_4344,N_4194,N_4306);
or U4345 (N_4345,N_4190,N_4215);
nand U4346 (N_4346,N_4317,N_4162);
or U4347 (N_4347,N_4265,N_4292);
or U4348 (N_4348,N_4172,N_4285);
nand U4349 (N_4349,N_4210,N_4230);
xor U4350 (N_4350,N_4312,N_4244);
or U4351 (N_4351,N_4211,N_4279);
nor U4352 (N_4352,N_4187,N_4221);
nor U4353 (N_4353,N_4218,N_4171);
nor U4354 (N_4354,N_4204,N_4165);
and U4355 (N_4355,N_4193,N_4315);
xnor U4356 (N_4356,N_4169,N_4258);
and U4357 (N_4357,N_4295,N_4170);
xnor U4358 (N_4358,N_4216,N_4229);
nand U4359 (N_4359,N_4264,N_4318);
and U4360 (N_4360,N_4267,N_4166);
and U4361 (N_4361,N_4182,N_4283);
xor U4362 (N_4362,N_4243,N_4260);
and U4363 (N_4363,N_4237,N_4214);
and U4364 (N_4364,N_4310,N_4206);
nor U4365 (N_4365,N_4313,N_4189);
xor U4366 (N_4366,N_4254,N_4305);
nor U4367 (N_4367,N_4233,N_4185);
or U4368 (N_4368,N_4290,N_4252);
and U4369 (N_4369,N_4234,N_4192);
and U4370 (N_4370,N_4304,N_4188);
and U4371 (N_4371,N_4199,N_4196);
xor U4372 (N_4372,N_4212,N_4161);
nor U4373 (N_4373,N_4207,N_4236);
xor U4374 (N_4374,N_4278,N_4280);
and U4375 (N_4375,N_4273,N_4272);
xnor U4376 (N_4376,N_4179,N_4239);
nor U4377 (N_4377,N_4191,N_4270);
xnor U4378 (N_4378,N_4319,N_4282);
or U4379 (N_4379,N_4275,N_4160);
or U4380 (N_4380,N_4301,N_4186);
nand U4381 (N_4381,N_4174,N_4177);
xor U4382 (N_4382,N_4180,N_4268);
xor U4383 (N_4383,N_4175,N_4298);
nand U4384 (N_4384,N_4300,N_4231);
nor U4385 (N_4385,N_4238,N_4217);
or U4386 (N_4386,N_4205,N_4240);
nor U4387 (N_4387,N_4201,N_4274);
nor U4388 (N_4388,N_4213,N_4284);
xnor U4389 (N_4389,N_4224,N_4288);
xor U4390 (N_4390,N_4255,N_4294);
nor U4391 (N_4391,N_4293,N_4197);
nand U4392 (N_4392,N_4226,N_4297);
xnor U4393 (N_4393,N_4250,N_4195);
xnor U4394 (N_4394,N_4316,N_4242);
nor U4395 (N_4395,N_4163,N_4232);
and U4396 (N_4396,N_4202,N_4223);
or U4397 (N_4397,N_4164,N_4168);
and U4398 (N_4398,N_4173,N_4287);
or U4399 (N_4399,N_4209,N_4303);
nor U4400 (N_4400,N_4197,N_4226);
or U4401 (N_4401,N_4223,N_4243);
nor U4402 (N_4402,N_4316,N_4246);
nand U4403 (N_4403,N_4204,N_4162);
xnor U4404 (N_4404,N_4277,N_4233);
and U4405 (N_4405,N_4168,N_4191);
nor U4406 (N_4406,N_4175,N_4265);
or U4407 (N_4407,N_4266,N_4217);
nand U4408 (N_4408,N_4261,N_4181);
nor U4409 (N_4409,N_4311,N_4187);
or U4410 (N_4410,N_4292,N_4196);
or U4411 (N_4411,N_4251,N_4230);
xor U4412 (N_4412,N_4161,N_4230);
and U4413 (N_4413,N_4317,N_4222);
xnor U4414 (N_4414,N_4277,N_4285);
and U4415 (N_4415,N_4256,N_4229);
xor U4416 (N_4416,N_4169,N_4291);
xnor U4417 (N_4417,N_4182,N_4180);
xor U4418 (N_4418,N_4269,N_4259);
or U4419 (N_4419,N_4255,N_4162);
xor U4420 (N_4420,N_4239,N_4297);
xnor U4421 (N_4421,N_4215,N_4225);
and U4422 (N_4422,N_4290,N_4205);
nand U4423 (N_4423,N_4197,N_4261);
or U4424 (N_4424,N_4275,N_4176);
nand U4425 (N_4425,N_4170,N_4312);
and U4426 (N_4426,N_4187,N_4209);
or U4427 (N_4427,N_4179,N_4282);
nand U4428 (N_4428,N_4306,N_4178);
or U4429 (N_4429,N_4299,N_4293);
nand U4430 (N_4430,N_4286,N_4242);
and U4431 (N_4431,N_4229,N_4311);
and U4432 (N_4432,N_4191,N_4257);
nor U4433 (N_4433,N_4299,N_4317);
or U4434 (N_4434,N_4278,N_4187);
nand U4435 (N_4435,N_4278,N_4303);
nor U4436 (N_4436,N_4277,N_4167);
nor U4437 (N_4437,N_4247,N_4312);
xor U4438 (N_4438,N_4218,N_4224);
or U4439 (N_4439,N_4179,N_4308);
and U4440 (N_4440,N_4182,N_4256);
nand U4441 (N_4441,N_4275,N_4265);
and U4442 (N_4442,N_4296,N_4236);
nor U4443 (N_4443,N_4281,N_4318);
and U4444 (N_4444,N_4275,N_4245);
or U4445 (N_4445,N_4181,N_4267);
or U4446 (N_4446,N_4166,N_4307);
nor U4447 (N_4447,N_4258,N_4253);
nand U4448 (N_4448,N_4317,N_4245);
nor U4449 (N_4449,N_4302,N_4215);
nand U4450 (N_4450,N_4242,N_4218);
nor U4451 (N_4451,N_4222,N_4281);
xnor U4452 (N_4452,N_4246,N_4238);
and U4453 (N_4453,N_4288,N_4311);
nor U4454 (N_4454,N_4270,N_4291);
xor U4455 (N_4455,N_4260,N_4232);
and U4456 (N_4456,N_4163,N_4178);
nor U4457 (N_4457,N_4317,N_4318);
nor U4458 (N_4458,N_4301,N_4294);
nor U4459 (N_4459,N_4296,N_4182);
xor U4460 (N_4460,N_4205,N_4232);
xor U4461 (N_4461,N_4194,N_4231);
nand U4462 (N_4462,N_4222,N_4229);
nor U4463 (N_4463,N_4211,N_4238);
xor U4464 (N_4464,N_4196,N_4235);
or U4465 (N_4465,N_4273,N_4261);
xor U4466 (N_4466,N_4264,N_4286);
xor U4467 (N_4467,N_4299,N_4309);
xor U4468 (N_4468,N_4227,N_4166);
and U4469 (N_4469,N_4170,N_4227);
nor U4470 (N_4470,N_4198,N_4240);
or U4471 (N_4471,N_4276,N_4235);
or U4472 (N_4472,N_4245,N_4243);
xor U4473 (N_4473,N_4290,N_4197);
nor U4474 (N_4474,N_4240,N_4318);
nand U4475 (N_4475,N_4235,N_4240);
xnor U4476 (N_4476,N_4176,N_4181);
xnor U4477 (N_4477,N_4290,N_4298);
nor U4478 (N_4478,N_4198,N_4292);
nand U4479 (N_4479,N_4253,N_4268);
and U4480 (N_4480,N_4436,N_4343);
xnor U4481 (N_4481,N_4327,N_4468);
xor U4482 (N_4482,N_4370,N_4361);
and U4483 (N_4483,N_4409,N_4342);
nand U4484 (N_4484,N_4366,N_4472);
nor U4485 (N_4485,N_4330,N_4404);
nand U4486 (N_4486,N_4416,N_4438);
or U4487 (N_4487,N_4332,N_4453);
xnor U4488 (N_4488,N_4395,N_4458);
and U4489 (N_4489,N_4364,N_4393);
nand U4490 (N_4490,N_4392,N_4406);
xor U4491 (N_4491,N_4403,N_4389);
or U4492 (N_4492,N_4352,N_4459);
or U4493 (N_4493,N_4339,N_4323);
nor U4494 (N_4494,N_4450,N_4381);
nor U4495 (N_4495,N_4391,N_4382);
nor U4496 (N_4496,N_4440,N_4449);
xor U4497 (N_4497,N_4375,N_4470);
and U4498 (N_4498,N_4463,N_4347);
nand U4499 (N_4499,N_4385,N_4451);
xor U4500 (N_4500,N_4325,N_4348);
nor U4501 (N_4501,N_4429,N_4402);
nor U4502 (N_4502,N_4349,N_4419);
or U4503 (N_4503,N_4473,N_4322);
nor U4504 (N_4504,N_4418,N_4407);
or U4505 (N_4505,N_4466,N_4390);
xnor U4506 (N_4506,N_4377,N_4456);
xor U4507 (N_4507,N_4360,N_4460);
nand U4508 (N_4508,N_4431,N_4452);
and U4509 (N_4509,N_4413,N_4426);
or U4510 (N_4510,N_4331,N_4379);
nor U4511 (N_4511,N_4457,N_4367);
nand U4512 (N_4512,N_4401,N_4405);
nor U4513 (N_4513,N_4462,N_4356);
nand U4514 (N_4514,N_4424,N_4464);
nand U4515 (N_4515,N_4444,N_4357);
nor U4516 (N_4516,N_4376,N_4400);
nor U4517 (N_4517,N_4467,N_4420);
and U4518 (N_4518,N_4411,N_4439);
nand U4519 (N_4519,N_4469,N_4371);
nor U4520 (N_4520,N_4320,N_4386);
nor U4521 (N_4521,N_4394,N_4479);
nand U4522 (N_4522,N_4410,N_4399);
nand U4523 (N_4523,N_4355,N_4372);
xnor U4524 (N_4524,N_4447,N_4368);
xor U4525 (N_4525,N_4324,N_4337);
nand U4526 (N_4526,N_4471,N_4358);
xnor U4527 (N_4527,N_4414,N_4383);
xor U4528 (N_4528,N_4445,N_4387);
nor U4529 (N_4529,N_4334,N_4345);
and U4530 (N_4530,N_4474,N_4398);
and U4531 (N_4531,N_4422,N_4423);
and U4532 (N_4532,N_4374,N_4461);
and U4533 (N_4533,N_4321,N_4359);
xor U4534 (N_4534,N_4415,N_4441);
xor U4535 (N_4535,N_4454,N_4408);
or U4536 (N_4536,N_4437,N_4388);
or U4537 (N_4537,N_4378,N_4373);
nor U4538 (N_4538,N_4435,N_4351);
or U4539 (N_4539,N_4427,N_4328);
and U4540 (N_4540,N_4448,N_4354);
or U4541 (N_4541,N_4336,N_4335);
or U4542 (N_4542,N_4442,N_4428);
nand U4543 (N_4543,N_4475,N_4434);
and U4544 (N_4544,N_4465,N_4455);
xnor U4545 (N_4545,N_4412,N_4340);
nor U4546 (N_4546,N_4344,N_4333);
xor U4547 (N_4547,N_4443,N_4430);
and U4548 (N_4548,N_4397,N_4365);
or U4549 (N_4549,N_4369,N_4417);
nand U4550 (N_4550,N_4350,N_4338);
nor U4551 (N_4551,N_4425,N_4346);
and U4552 (N_4552,N_4363,N_4446);
xor U4553 (N_4553,N_4477,N_4326);
xnor U4554 (N_4554,N_4384,N_4353);
or U4555 (N_4555,N_4329,N_4380);
or U4556 (N_4556,N_4433,N_4476);
nand U4557 (N_4557,N_4362,N_4396);
or U4558 (N_4558,N_4421,N_4341);
or U4559 (N_4559,N_4432,N_4478);
and U4560 (N_4560,N_4409,N_4418);
and U4561 (N_4561,N_4474,N_4424);
or U4562 (N_4562,N_4398,N_4382);
nand U4563 (N_4563,N_4428,N_4377);
nand U4564 (N_4564,N_4428,N_4340);
or U4565 (N_4565,N_4456,N_4415);
xor U4566 (N_4566,N_4380,N_4455);
xor U4567 (N_4567,N_4345,N_4355);
and U4568 (N_4568,N_4423,N_4458);
and U4569 (N_4569,N_4414,N_4477);
nor U4570 (N_4570,N_4437,N_4383);
xnor U4571 (N_4571,N_4440,N_4370);
nor U4572 (N_4572,N_4446,N_4375);
and U4573 (N_4573,N_4327,N_4375);
and U4574 (N_4574,N_4332,N_4474);
nor U4575 (N_4575,N_4409,N_4336);
nor U4576 (N_4576,N_4452,N_4389);
and U4577 (N_4577,N_4373,N_4465);
nand U4578 (N_4578,N_4383,N_4446);
nor U4579 (N_4579,N_4383,N_4344);
nor U4580 (N_4580,N_4411,N_4322);
nand U4581 (N_4581,N_4387,N_4389);
xor U4582 (N_4582,N_4445,N_4432);
nand U4583 (N_4583,N_4337,N_4370);
nand U4584 (N_4584,N_4406,N_4357);
nand U4585 (N_4585,N_4353,N_4393);
nor U4586 (N_4586,N_4434,N_4436);
or U4587 (N_4587,N_4344,N_4433);
or U4588 (N_4588,N_4467,N_4459);
nand U4589 (N_4589,N_4432,N_4328);
or U4590 (N_4590,N_4359,N_4430);
or U4591 (N_4591,N_4411,N_4370);
xor U4592 (N_4592,N_4404,N_4466);
nor U4593 (N_4593,N_4328,N_4475);
or U4594 (N_4594,N_4472,N_4468);
nor U4595 (N_4595,N_4385,N_4339);
or U4596 (N_4596,N_4470,N_4333);
or U4597 (N_4597,N_4458,N_4475);
nand U4598 (N_4598,N_4367,N_4399);
or U4599 (N_4599,N_4325,N_4426);
nand U4600 (N_4600,N_4322,N_4399);
xnor U4601 (N_4601,N_4435,N_4407);
nand U4602 (N_4602,N_4355,N_4329);
or U4603 (N_4603,N_4407,N_4441);
or U4604 (N_4604,N_4392,N_4431);
and U4605 (N_4605,N_4476,N_4329);
or U4606 (N_4606,N_4322,N_4437);
or U4607 (N_4607,N_4322,N_4468);
nand U4608 (N_4608,N_4400,N_4378);
and U4609 (N_4609,N_4341,N_4433);
nand U4610 (N_4610,N_4328,N_4356);
and U4611 (N_4611,N_4379,N_4338);
xnor U4612 (N_4612,N_4433,N_4383);
nor U4613 (N_4613,N_4439,N_4383);
or U4614 (N_4614,N_4339,N_4404);
xnor U4615 (N_4615,N_4474,N_4350);
or U4616 (N_4616,N_4439,N_4434);
nor U4617 (N_4617,N_4379,N_4368);
xor U4618 (N_4618,N_4451,N_4421);
nand U4619 (N_4619,N_4359,N_4467);
and U4620 (N_4620,N_4378,N_4454);
and U4621 (N_4621,N_4374,N_4449);
nand U4622 (N_4622,N_4337,N_4334);
nand U4623 (N_4623,N_4363,N_4436);
or U4624 (N_4624,N_4450,N_4456);
nand U4625 (N_4625,N_4367,N_4406);
or U4626 (N_4626,N_4414,N_4476);
and U4627 (N_4627,N_4321,N_4478);
nand U4628 (N_4628,N_4359,N_4376);
xor U4629 (N_4629,N_4426,N_4422);
and U4630 (N_4630,N_4468,N_4385);
and U4631 (N_4631,N_4456,N_4402);
nand U4632 (N_4632,N_4460,N_4467);
or U4633 (N_4633,N_4445,N_4363);
or U4634 (N_4634,N_4347,N_4427);
and U4635 (N_4635,N_4395,N_4477);
nor U4636 (N_4636,N_4452,N_4395);
nor U4637 (N_4637,N_4442,N_4361);
nand U4638 (N_4638,N_4337,N_4377);
or U4639 (N_4639,N_4336,N_4470);
and U4640 (N_4640,N_4534,N_4612);
nand U4641 (N_4641,N_4608,N_4598);
or U4642 (N_4642,N_4495,N_4563);
and U4643 (N_4643,N_4507,N_4535);
nor U4644 (N_4644,N_4617,N_4490);
xnor U4645 (N_4645,N_4581,N_4508);
nor U4646 (N_4646,N_4550,N_4591);
or U4647 (N_4647,N_4638,N_4515);
nor U4648 (N_4648,N_4639,N_4599);
xor U4649 (N_4649,N_4526,N_4564);
nor U4650 (N_4650,N_4540,N_4580);
and U4651 (N_4651,N_4592,N_4492);
nand U4652 (N_4652,N_4603,N_4551);
nand U4653 (N_4653,N_4505,N_4630);
xnor U4654 (N_4654,N_4514,N_4568);
xnor U4655 (N_4655,N_4579,N_4528);
nor U4656 (N_4656,N_4511,N_4622);
nand U4657 (N_4657,N_4553,N_4525);
nand U4658 (N_4658,N_4596,N_4493);
nand U4659 (N_4659,N_4618,N_4619);
xor U4660 (N_4660,N_4633,N_4572);
nand U4661 (N_4661,N_4506,N_4588);
or U4662 (N_4662,N_4518,N_4593);
xnor U4663 (N_4663,N_4554,N_4635);
nor U4664 (N_4664,N_4586,N_4561);
nor U4665 (N_4665,N_4602,N_4556);
or U4666 (N_4666,N_4611,N_4589);
and U4667 (N_4667,N_4557,N_4530);
xor U4668 (N_4668,N_4627,N_4637);
nor U4669 (N_4669,N_4629,N_4516);
and U4670 (N_4670,N_4547,N_4524);
nand U4671 (N_4671,N_4536,N_4546);
or U4672 (N_4672,N_4520,N_4610);
nand U4673 (N_4673,N_4494,N_4616);
or U4674 (N_4674,N_4539,N_4570);
or U4675 (N_4675,N_4573,N_4583);
nand U4676 (N_4676,N_4480,N_4527);
or U4677 (N_4677,N_4585,N_4487);
or U4678 (N_4678,N_4489,N_4571);
or U4679 (N_4679,N_4614,N_4574);
and U4680 (N_4680,N_4632,N_4523);
nand U4681 (N_4681,N_4538,N_4541);
nand U4682 (N_4682,N_4620,N_4482);
and U4683 (N_4683,N_4595,N_4509);
nor U4684 (N_4684,N_4631,N_4519);
and U4685 (N_4685,N_4569,N_4483);
or U4686 (N_4686,N_4628,N_4513);
xnor U4687 (N_4687,N_4576,N_4559);
nand U4688 (N_4688,N_4594,N_4634);
and U4689 (N_4689,N_4517,N_4607);
xnor U4690 (N_4690,N_4496,N_4500);
xor U4691 (N_4691,N_4504,N_4481);
xnor U4692 (N_4692,N_4488,N_4625);
nand U4693 (N_4693,N_4510,N_4548);
xnor U4694 (N_4694,N_4584,N_4578);
or U4695 (N_4695,N_4545,N_4562);
xor U4696 (N_4696,N_4542,N_4497);
nand U4697 (N_4697,N_4609,N_4531);
nand U4698 (N_4698,N_4624,N_4636);
and U4699 (N_4699,N_4575,N_4486);
nand U4700 (N_4700,N_4587,N_4501);
and U4701 (N_4701,N_4626,N_4543);
nand U4702 (N_4702,N_4605,N_4537);
nor U4703 (N_4703,N_4544,N_4521);
xor U4704 (N_4704,N_4503,N_4498);
xnor U4705 (N_4705,N_4533,N_4577);
nand U4706 (N_4706,N_4615,N_4600);
xnor U4707 (N_4707,N_4555,N_4522);
xnor U4708 (N_4708,N_4552,N_4485);
xor U4709 (N_4709,N_4491,N_4604);
nor U4710 (N_4710,N_4590,N_4597);
nor U4711 (N_4711,N_4549,N_4512);
and U4712 (N_4712,N_4567,N_4582);
or U4713 (N_4713,N_4613,N_4623);
nand U4714 (N_4714,N_4560,N_4565);
or U4715 (N_4715,N_4621,N_4499);
nor U4716 (N_4716,N_4601,N_4502);
xor U4717 (N_4717,N_4606,N_4558);
and U4718 (N_4718,N_4532,N_4566);
nor U4719 (N_4719,N_4529,N_4484);
nor U4720 (N_4720,N_4491,N_4489);
nand U4721 (N_4721,N_4592,N_4505);
nor U4722 (N_4722,N_4561,N_4584);
nand U4723 (N_4723,N_4536,N_4618);
xor U4724 (N_4724,N_4578,N_4490);
and U4725 (N_4725,N_4507,N_4527);
and U4726 (N_4726,N_4552,N_4503);
xnor U4727 (N_4727,N_4620,N_4539);
xor U4728 (N_4728,N_4556,N_4574);
and U4729 (N_4729,N_4480,N_4621);
and U4730 (N_4730,N_4541,N_4625);
or U4731 (N_4731,N_4591,N_4612);
nand U4732 (N_4732,N_4547,N_4571);
or U4733 (N_4733,N_4492,N_4513);
xor U4734 (N_4734,N_4578,N_4512);
xnor U4735 (N_4735,N_4559,N_4482);
and U4736 (N_4736,N_4563,N_4521);
nor U4737 (N_4737,N_4594,N_4602);
xnor U4738 (N_4738,N_4489,N_4513);
nand U4739 (N_4739,N_4547,N_4565);
xor U4740 (N_4740,N_4617,N_4606);
nand U4741 (N_4741,N_4508,N_4502);
and U4742 (N_4742,N_4530,N_4618);
nor U4743 (N_4743,N_4576,N_4589);
nand U4744 (N_4744,N_4601,N_4533);
xnor U4745 (N_4745,N_4638,N_4635);
nand U4746 (N_4746,N_4559,N_4637);
and U4747 (N_4747,N_4582,N_4526);
or U4748 (N_4748,N_4519,N_4520);
and U4749 (N_4749,N_4518,N_4523);
or U4750 (N_4750,N_4497,N_4587);
nand U4751 (N_4751,N_4594,N_4493);
and U4752 (N_4752,N_4494,N_4550);
nor U4753 (N_4753,N_4498,N_4543);
or U4754 (N_4754,N_4568,N_4524);
and U4755 (N_4755,N_4636,N_4599);
or U4756 (N_4756,N_4556,N_4607);
and U4757 (N_4757,N_4559,N_4606);
xor U4758 (N_4758,N_4634,N_4566);
and U4759 (N_4759,N_4575,N_4613);
xnor U4760 (N_4760,N_4546,N_4613);
nor U4761 (N_4761,N_4592,N_4591);
nor U4762 (N_4762,N_4544,N_4537);
nor U4763 (N_4763,N_4487,N_4496);
or U4764 (N_4764,N_4522,N_4569);
xor U4765 (N_4765,N_4487,N_4532);
or U4766 (N_4766,N_4513,N_4484);
xor U4767 (N_4767,N_4534,N_4507);
and U4768 (N_4768,N_4595,N_4627);
nand U4769 (N_4769,N_4601,N_4483);
and U4770 (N_4770,N_4622,N_4528);
nor U4771 (N_4771,N_4534,N_4584);
nor U4772 (N_4772,N_4627,N_4560);
xor U4773 (N_4773,N_4639,N_4636);
and U4774 (N_4774,N_4628,N_4610);
xnor U4775 (N_4775,N_4521,N_4575);
nand U4776 (N_4776,N_4621,N_4599);
and U4777 (N_4777,N_4609,N_4629);
xnor U4778 (N_4778,N_4595,N_4638);
nor U4779 (N_4779,N_4487,N_4632);
xor U4780 (N_4780,N_4574,N_4639);
or U4781 (N_4781,N_4570,N_4604);
xnor U4782 (N_4782,N_4618,N_4639);
xor U4783 (N_4783,N_4586,N_4486);
nand U4784 (N_4784,N_4598,N_4562);
and U4785 (N_4785,N_4525,N_4500);
or U4786 (N_4786,N_4551,N_4504);
nand U4787 (N_4787,N_4537,N_4519);
nor U4788 (N_4788,N_4631,N_4635);
nand U4789 (N_4789,N_4525,N_4575);
xnor U4790 (N_4790,N_4494,N_4486);
xor U4791 (N_4791,N_4548,N_4527);
nor U4792 (N_4792,N_4502,N_4600);
or U4793 (N_4793,N_4594,N_4593);
or U4794 (N_4794,N_4571,N_4560);
or U4795 (N_4795,N_4529,N_4526);
or U4796 (N_4796,N_4611,N_4509);
and U4797 (N_4797,N_4539,N_4519);
nand U4798 (N_4798,N_4526,N_4506);
xnor U4799 (N_4799,N_4510,N_4525);
xnor U4800 (N_4800,N_4774,N_4750);
or U4801 (N_4801,N_4790,N_4715);
and U4802 (N_4802,N_4783,N_4709);
nor U4803 (N_4803,N_4699,N_4723);
or U4804 (N_4804,N_4720,N_4760);
nand U4805 (N_4805,N_4736,N_4640);
nand U4806 (N_4806,N_4717,N_4671);
xnor U4807 (N_4807,N_4719,N_4652);
nand U4808 (N_4808,N_4748,N_4672);
and U4809 (N_4809,N_4757,N_4673);
and U4810 (N_4810,N_4680,N_4799);
or U4811 (N_4811,N_4716,N_4698);
nor U4812 (N_4812,N_4666,N_4686);
and U4813 (N_4813,N_4741,N_4758);
xor U4814 (N_4814,N_4688,N_4775);
and U4815 (N_4815,N_4789,N_4773);
nand U4816 (N_4816,N_4645,N_4728);
xor U4817 (N_4817,N_4661,N_4689);
and U4818 (N_4818,N_4786,N_4745);
nor U4819 (N_4819,N_4793,N_4743);
or U4820 (N_4820,N_4795,N_4687);
nand U4821 (N_4821,N_4667,N_4788);
nor U4822 (N_4822,N_4655,N_4762);
xnor U4823 (N_4823,N_4718,N_4796);
xor U4824 (N_4824,N_4659,N_4650);
and U4825 (N_4825,N_4776,N_4792);
or U4826 (N_4826,N_4646,N_4765);
nor U4827 (N_4827,N_4681,N_4654);
or U4828 (N_4828,N_4791,N_4772);
and U4829 (N_4829,N_4653,N_4764);
nand U4830 (N_4830,N_4771,N_4710);
or U4831 (N_4831,N_4664,N_4756);
or U4832 (N_4832,N_4701,N_4683);
nand U4833 (N_4833,N_4733,N_4721);
or U4834 (N_4834,N_4735,N_4727);
nand U4835 (N_4835,N_4676,N_4729);
and U4836 (N_4836,N_4660,N_4724);
nand U4837 (N_4837,N_4693,N_4755);
and U4838 (N_4838,N_4782,N_4781);
and U4839 (N_4839,N_4794,N_4752);
nor U4840 (N_4840,N_4731,N_4641);
nor U4841 (N_4841,N_4700,N_4777);
and U4842 (N_4842,N_4695,N_4679);
or U4843 (N_4843,N_4778,N_4647);
xnor U4844 (N_4844,N_4726,N_4669);
xnor U4845 (N_4845,N_4751,N_4770);
or U4846 (N_4846,N_4712,N_4670);
and U4847 (N_4847,N_4649,N_4656);
nand U4848 (N_4848,N_4759,N_4707);
nand U4849 (N_4849,N_4668,N_4749);
xnor U4850 (N_4850,N_4754,N_4785);
xor U4851 (N_4851,N_4704,N_4768);
xnor U4852 (N_4852,N_4730,N_4753);
or U4853 (N_4853,N_4696,N_4746);
and U4854 (N_4854,N_4761,N_4739);
nor U4855 (N_4855,N_4797,N_4779);
nand U4856 (N_4856,N_4713,N_4702);
and U4857 (N_4857,N_4651,N_4662);
nand U4858 (N_4858,N_4703,N_4737);
xnor U4859 (N_4859,N_4722,N_4747);
or U4860 (N_4860,N_4690,N_4705);
xor U4861 (N_4861,N_4742,N_4663);
and U4862 (N_4862,N_4769,N_4734);
nor U4863 (N_4863,N_4648,N_4711);
or U4864 (N_4864,N_4740,N_4766);
nor U4865 (N_4865,N_4675,N_4763);
or U4866 (N_4866,N_4643,N_4706);
nor U4867 (N_4867,N_4692,N_4685);
nand U4868 (N_4868,N_4697,N_4738);
or U4869 (N_4869,N_4725,N_4678);
or U4870 (N_4870,N_4714,N_4665);
and U4871 (N_4871,N_4657,N_4744);
or U4872 (N_4872,N_4682,N_4732);
and U4873 (N_4873,N_4674,N_4677);
xnor U4874 (N_4874,N_4684,N_4708);
and U4875 (N_4875,N_4798,N_4787);
and U4876 (N_4876,N_4644,N_4694);
nand U4877 (N_4877,N_4691,N_4780);
and U4878 (N_4878,N_4658,N_4767);
and U4879 (N_4879,N_4784,N_4642);
nand U4880 (N_4880,N_4779,N_4647);
xnor U4881 (N_4881,N_4754,N_4742);
nor U4882 (N_4882,N_4673,N_4728);
nor U4883 (N_4883,N_4743,N_4659);
xor U4884 (N_4884,N_4747,N_4710);
nor U4885 (N_4885,N_4794,N_4663);
and U4886 (N_4886,N_4765,N_4641);
and U4887 (N_4887,N_4716,N_4788);
nor U4888 (N_4888,N_4644,N_4792);
xnor U4889 (N_4889,N_4734,N_4719);
nor U4890 (N_4890,N_4746,N_4728);
xor U4891 (N_4891,N_4799,N_4657);
nand U4892 (N_4892,N_4745,N_4654);
or U4893 (N_4893,N_4790,N_4668);
nor U4894 (N_4894,N_4682,N_4725);
or U4895 (N_4895,N_4794,N_4770);
nand U4896 (N_4896,N_4771,N_4722);
nor U4897 (N_4897,N_4756,N_4768);
or U4898 (N_4898,N_4792,N_4744);
or U4899 (N_4899,N_4650,N_4670);
or U4900 (N_4900,N_4686,N_4757);
xnor U4901 (N_4901,N_4692,N_4769);
xor U4902 (N_4902,N_4693,N_4736);
xor U4903 (N_4903,N_4696,N_4794);
xnor U4904 (N_4904,N_4719,N_4685);
nand U4905 (N_4905,N_4677,N_4698);
or U4906 (N_4906,N_4795,N_4781);
and U4907 (N_4907,N_4785,N_4706);
or U4908 (N_4908,N_4759,N_4767);
nand U4909 (N_4909,N_4759,N_4769);
or U4910 (N_4910,N_4674,N_4659);
nor U4911 (N_4911,N_4708,N_4698);
or U4912 (N_4912,N_4776,N_4769);
and U4913 (N_4913,N_4660,N_4736);
and U4914 (N_4914,N_4658,N_4771);
xnor U4915 (N_4915,N_4750,N_4681);
xnor U4916 (N_4916,N_4742,N_4705);
or U4917 (N_4917,N_4751,N_4689);
and U4918 (N_4918,N_4709,N_4739);
nand U4919 (N_4919,N_4725,N_4723);
nor U4920 (N_4920,N_4712,N_4782);
nor U4921 (N_4921,N_4797,N_4688);
xor U4922 (N_4922,N_4766,N_4700);
xor U4923 (N_4923,N_4709,N_4661);
and U4924 (N_4924,N_4671,N_4709);
nor U4925 (N_4925,N_4773,N_4644);
nand U4926 (N_4926,N_4645,N_4655);
nor U4927 (N_4927,N_4729,N_4652);
or U4928 (N_4928,N_4703,N_4738);
nor U4929 (N_4929,N_4748,N_4719);
nor U4930 (N_4930,N_4744,N_4674);
or U4931 (N_4931,N_4698,N_4655);
xor U4932 (N_4932,N_4765,N_4775);
or U4933 (N_4933,N_4650,N_4787);
and U4934 (N_4934,N_4644,N_4736);
xor U4935 (N_4935,N_4642,N_4759);
nand U4936 (N_4936,N_4704,N_4711);
nor U4937 (N_4937,N_4675,N_4686);
or U4938 (N_4938,N_4723,N_4763);
nand U4939 (N_4939,N_4785,N_4752);
xnor U4940 (N_4940,N_4765,N_4660);
xor U4941 (N_4941,N_4671,N_4762);
and U4942 (N_4942,N_4748,N_4735);
and U4943 (N_4943,N_4737,N_4690);
xor U4944 (N_4944,N_4664,N_4675);
nor U4945 (N_4945,N_4746,N_4662);
xor U4946 (N_4946,N_4764,N_4674);
nor U4947 (N_4947,N_4659,N_4759);
and U4948 (N_4948,N_4657,N_4715);
and U4949 (N_4949,N_4724,N_4790);
nand U4950 (N_4950,N_4781,N_4793);
nor U4951 (N_4951,N_4657,N_4756);
nand U4952 (N_4952,N_4684,N_4656);
or U4953 (N_4953,N_4757,N_4676);
and U4954 (N_4954,N_4732,N_4762);
or U4955 (N_4955,N_4710,N_4741);
xnor U4956 (N_4956,N_4728,N_4684);
nand U4957 (N_4957,N_4733,N_4737);
nor U4958 (N_4958,N_4644,N_4793);
or U4959 (N_4959,N_4675,N_4644);
or U4960 (N_4960,N_4927,N_4955);
xnor U4961 (N_4961,N_4869,N_4843);
and U4962 (N_4962,N_4953,N_4828);
nor U4963 (N_4963,N_4868,N_4809);
nand U4964 (N_4964,N_4951,N_4924);
xor U4965 (N_4965,N_4889,N_4884);
xnor U4966 (N_4966,N_4818,N_4856);
nand U4967 (N_4967,N_4958,N_4886);
nand U4968 (N_4968,N_4820,N_4875);
nand U4969 (N_4969,N_4907,N_4812);
and U4970 (N_4970,N_4878,N_4861);
and U4971 (N_4971,N_4939,N_4943);
and U4972 (N_4972,N_4805,N_4913);
or U4973 (N_4973,N_4823,N_4804);
nor U4974 (N_4974,N_4853,N_4948);
xor U4975 (N_4975,N_4942,N_4959);
xnor U4976 (N_4976,N_4956,N_4867);
or U4977 (N_4977,N_4883,N_4814);
nand U4978 (N_4978,N_4895,N_4802);
xor U4979 (N_4979,N_4826,N_4892);
nand U4980 (N_4980,N_4935,N_4844);
or U4981 (N_4981,N_4899,N_4834);
xnor U4982 (N_4982,N_4932,N_4877);
nand U4983 (N_4983,N_4946,N_4950);
xor U4984 (N_4984,N_4837,N_4842);
nor U4985 (N_4985,N_4825,N_4905);
and U4986 (N_4986,N_4819,N_4839);
nor U4987 (N_4987,N_4903,N_4830);
nand U4988 (N_4988,N_4841,N_4938);
nand U4989 (N_4989,N_4929,N_4850);
and U4990 (N_4990,N_4816,N_4919);
xnor U4991 (N_4991,N_4925,N_4847);
and U4992 (N_4992,N_4945,N_4858);
and U4993 (N_4993,N_4926,N_4901);
xor U4994 (N_4994,N_4846,N_4915);
nor U4995 (N_4995,N_4917,N_4888);
nor U4996 (N_4996,N_4934,N_4952);
xnor U4997 (N_4997,N_4872,N_4936);
nand U4998 (N_4998,N_4876,N_4920);
nor U4999 (N_4999,N_4957,N_4849);
nor U5000 (N_5000,N_4949,N_4824);
or U5001 (N_5001,N_4882,N_4801);
nor U5002 (N_5002,N_4918,N_4864);
or U5003 (N_5003,N_4885,N_4833);
or U5004 (N_5004,N_4848,N_4887);
nand U5005 (N_5005,N_4822,N_4813);
nand U5006 (N_5006,N_4898,N_4912);
xnor U5007 (N_5007,N_4896,N_4923);
xor U5008 (N_5008,N_4921,N_4863);
xnor U5009 (N_5009,N_4928,N_4832);
xnor U5010 (N_5010,N_4803,N_4831);
xnor U5011 (N_5011,N_4893,N_4810);
xor U5012 (N_5012,N_4811,N_4922);
or U5013 (N_5013,N_4827,N_4859);
or U5014 (N_5014,N_4947,N_4890);
xnor U5015 (N_5015,N_4906,N_4891);
nand U5016 (N_5016,N_4931,N_4808);
nor U5017 (N_5017,N_4866,N_4851);
nor U5018 (N_5018,N_4930,N_4916);
xor U5019 (N_5019,N_4910,N_4835);
and U5020 (N_5020,N_4902,N_4829);
nand U5021 (N_5021,N_4865,N_4852);
or U5022 (N_5022,N_4880,N_4817);
xnor U5023 (N_5023,N_4904,N_4840);
and U5024 (N_5024,N_4954,N_4914);
nor U5025 (N_5025,N_4838,N_4881);
or U5026 (N_5026,N_4933,N_4944);
nor U5027 (N_5027,N_4815,N_4807);
and U5028 (N_5028,N_4821,N_4873);
xor U5029 (N_5029,N_4806,N_4940);
nor U5030 (N_5030,N_4874,N_4836);
and U5031 (N_5031,N_4860,N_4879);
nor U5032 (N_5032,N_4909,N_4941);
xnor U5033 (N_5033,N_4897,N_4871);
nor U5034 (N_5034,N_4894,N_4937);
and U5035 (N_5035,N_4900,N_4862);
or U5036 (N_5036,N_4854,N_4855);
nor U5037 (N_5037,N_4857,N_4845);
or U5038 (N_5038,N_4870,N_4911);
nor U5039 (N_5039,N_4908,N_4800);
and U5040 (N_5040,N_4813,N_4865);
nor U5041 (N_5041,N_4950,N_4874);
and U5042 (N_5042,N_4949,N_4808);
xnor U5043 (N_5043,N_4843,N_4959);
nor U5044 (N_5044,N_4870,N_4841);
xor U5045 (N_5045,N_4860,N_4831);
or U5046 (N_5046,N_4867,N_4827);
nor U5047 (N_5047,N_4839,N_4936);
nor U5048 (N_5048,N_4875,N_4945);
nor U5049 (N_5049,N_4955,N_4959);
xnor U5050 (N_5050,N_4930,N_4811);
nor U5051 (N_5051,N_4894,N_4946);
nor U5052 (N_5052,N_4853,N_4949);
xnor U5053 (N_5053,N_4854,N_4816);
nor U5054 (N_5054,N_4894,N_4883);
xor U5055 (N_5055,N_4873,N_4916);
xnor U5056 (N_5056,N_4879,N_4835);
and U5057 (N_5057,N_4830,N_4812);
nor U5058 (N_5058,N_4852,N_4907);
nor U5059 (N_5059,N_4920,N_4858);
and U5060 (N_5060,N_4855,N_4826);
nand U5061 (N_5061,N_4958,N_4808);
xnor U5062 (N_5062,N_4926,N_4824);
xor U5063 (N_5063,N_4914,N_4803);
xnor U5064 (N_5064,N_4910,N_4872);
nor U5065 (N_5065,N_4811,N_4921);
nand U5066 (N_5066,N_4928,N_4880);
nor U5067 (N_5067,N_4954,N_4945);
xnor U5068 (N_5068,N_4945,N_4910);
and U5069 (N_5069,N_4944,N_4864);
nand U5070 (N_5070,N_4944,N_4825);
xnor U5071 (N_5071,N_4916,N_4881);
and U5072 (N_5072,N_4931,N_4896);
or U5073 (N_5073,N_4828,N_4898);
xor U5074 (N_5074,N_4906,N_4808);
and U5075 (N_5075,N_4938,N_4909);
xor U5076 (N_5076,N_4880,N_4870);
and U5077 (N_5077,N_4854,N_4911);
nand U5078 (N_5078,N_4917,N_4815);
xor U5079 (N_5079,N_4896,N_4821);
or U5080 (N_5080,N_4935,N_4939);
nand U5081 (N_5081,N_4857,N_4878);
or U5082 (N_5082,N_4888,N_4878);
nor U5083 (N_5083,N_4875,N_4851);
nor U5084 (N_5084,N_4870,N_4919);
or U5085 (N_5085,N_4852,N_4940);
xor U5086 (N_5086,N_4811,N_4931);
and U5087 (N_5087,N_4834,N_4936);
or U5088 (N_5088,N_4949,N_4866);
nor U5089 (N_5089,N_4847,N_4891);
nor U5090 (N_5090,N_4808,N_4822);
nor U5091 (N_5091,N_4853,N_4910);
or U5092 (N_5092,N_4921,N_4825);
nor U5093 (N_5093,N_4937,N_4867);
nand U5094 (N_5094,N_4957,N_4850);
nor U5095 (N_5095,N_4826,N_4927);
nand U5096 (N_5096,N_4935,N_4877);
nor U5097 (N_5097,N_4811,N_4846);
nand U5098 (N_5098,N_4910,N_4812);
xor U5099 (N_5099,N_4930,N_4828);
nand U5100 (N_5100,N_4803,N_4920);
and U5101 (N_5101,N_4876,N_4958);
or U5102 (N_5102,N_4916,N_4842);
nand U5103 (N_5103,N_4827,N_4886);
and U5104 (N_5104,N_4921,N_4892);
and U5105 (N_5105,N_4873,N_4958);
xor U5106 (N_5106,N_4832,N_4937);
nand U5107 (N_5107,N_4931,N_4852);
nor U5108 (N_5108,N_4806,N_4933);
nor U5109 (N_5109,N_4847,N_4839);
xor U5110 (N_5110,N_4884,N_4954);
xnor U5111 (N_5111,N_4847,N_4929);
xnor U5112 (N_5112,N_4812,N_4851);
xor U5113 (N_5113,N_4925,N_4869);
xor U5114 (N_5114,N_4841,N_4813);
and U5115 (N_5115,N_4893,N_4867);
or U5116 (N_5116,N_4904,N_4874);
xnor U5117 (N_5117,N_4886,N_4879);
and U5118 (N_5118,N_4815,N_4908);
xor U5119 (N_5119,N_4958,N_4956);
xnor U5120 (N_5120,N_5071,N_5019);
nand U5121 (N_5121,N_5027,N_5025);
nand U5122 (N_5122,N_5016,N_5045);
and U5123 (N_5123,N_4968,N_5086);
or U5124 (N_5124,N_5040,N_5073);
or U5125 (N_5125,N_5030,N_5098);
nand U5126 (N_5126,N_5107,N_5056);
nand U5127 (N_5127,N_5119,N_5028);
nor U5128 (N_5128,N_5072,N_4997);
xor U5129 (N_5129,N_4975,N_4969);
nor U5130 (N_5130,N_4989,N_5088);
or U5131 (N_5131,N_5109,N_4999);
nor U5132 (N_5132,N_5042,N_5101);
xnor U5133 (N_5133,N_5106,N_4967);
nand U5134 (N_5134,N_4974,N_5022);
xnor U5135 (N_5135,N_5012,N_5113);
and U5136 (N_5136,N_5116,N_5058);
nor U5137 (N_5137,N_5067,N_5021);
and U5138 (N_5138,N_4962,N_5105);
xnor U5139 (N_5139,N_5080,N_5061);
nor U5140 (N_5140,N_5082,N_5000);
or U5141 (N_5141,N_4984,N_5038);
xnor U5142 (N_5142,N_4990,N_5094);
or U5143 (N_5143,N_4986,N_5029);
xor U5144 (N_5144,N_5005,N_5010);
xnor U5145 (N_5145,N_5104,N_5114);
and U5146 (N_5146,N_5066,N_4970);
xnor U5147 (N_5147,N_5091,N_5002);
and U5148 (N_5148,N_4996,N_5014);
nand U5149 (N_5149,N_5011,N_5070);
nand U5150 (N_5150,N_5095,N_5099);
nand U5151 (N_5151,N_5090,N_5069);
or U5152 (N_5152,N_5075,N_5003);
nor U5153 (N_5153,N_5064,N_4977);
nand U5154 (N_5154,N_5103,N_4991);
or U5155 (N_5155,N_5039,N_5063);
or U5156 (N_5156,N_5115,N_5048);
and U5157 (N_5157,N_5052,N_5087);
nand U5158 (N_5158,N_4971,N_4972);
and U5159 (N_5159,N_4979,N_4994);
and U5160 (N_5160,N_5015,N_5089);
nand U5161 (N_5161,N_5044,N_5023);
or U5162 (N_5162,N_5043,N_5057);
nand U5163 (N_5163,N_5111,N_5033);
or U5164 (N_5164,N_4982,N_4988);
and U5165 (N_5165,N_4985,N_5081);
or U5166 (N_5166,N_4966,N_5026);
and U5167 (N_5167,N_5096,N_5031);
nand U5168 (N_5168,N_5112,N_5110);
nor U5169 (N_5169,N_4980,N_5051);
nor U5170 (N_5170,N_4981,N_5001);
xor U5171 (N_5171,N_5085,N_5074);
xnor U5172 (N_5172,N_4973,N_5083);
or U5173 (N_5173,N_4987,N_5008);
and U5174 (N_5174,N_5092,N_5036);
nor U5175 (N_5175,N_4992,N_5035);
nor U5176 (N_5176,N_5100,N_4983);
or U5177 (N_5177,N_5076,N_5013);
or U5178 (N_5178,N_5017,N_5053);
or U5179 (N_5179,N_5037,N_5117);
xnor U5180 (N_5180,N_4960,N_5050);
and U5181 (N_5181,N_5004,N_5009);
and U5182 (N_5182,N_5078,N_5007);
or U5183 (N_5183,N_4998,N_5108);
or U5184 (N_5184,N_5060,N_5034);
or U5185 (N_5185,N_5049,N_5079);
nand U5186 (N_5186,N_5055,N_5006);
nand U5187 (N_5187,N_4995,N_4965);
or U5188 (N_5188,N_5047,N_4993);
nand U5189 (N_5189,N_5054,N_4963);
nand U5190 (N_5190,N_5046,N_4964);
xnor U5191 (N_5191,N_5018,N_5097);
xnor U5192 (N_5192,N_4978,N_5024);
nor U5193 (N_5193,N_5041,N_5068);
and U5194 (N_5194,N_4961,N_4976);
nand U5195 (N_5195,N_5118,N_5059);
or U5196 (N_5196,N_5062,N_5020);
and U5197 (N_5197,N_5093,N_5065);
and U5198 (N_5198,N_5084,N_5032);
xor U5199 (N_5199,N_5077,N_5102);
nand U5200 (N_5200,N_4999,N_4997);
and U5201 (N_5201,N_4973,N_5060);
nor U5202 (N_5202,N_4994,N_5089);
and U5203 (N_5203,N_5041,N_5006);
and U5204 (N_5204,N_5071,N_4998);
or U5205 (N_5205,N_5021,N_4993);
or U5206 (N_5206,N_5086,N_5003);
or U5207 (N_5207,N_5031,N_5018);
nand U5208 (N_5208,N_5103,N_5019);
xnor U5209 (N_5209,N_4995,N_5115);
nor U5210 (N_5210,N_5004,N_5040);
xnor U5211 (N_5211,N_4996,N_4972);
xor U5212 (N_5212,N_5001,N_5067);
nor U5213 (N_5213,N_5094,N_5012);
or U5214 (N_5214,N_4987,N_5110);
xnor U5215 (N_5215,N_5066,N_5027);
nor U5216 (N_5216,N_5059,N_4971);
and U5217 (N_5217,N_5027,N_5096);
and U5218 (N_5218,N_4969,N_4974);
xor U5219 (N_5219,N_5091,N_5078);
or U5220 (N_5220,N_4967,N_5012);
and U5221 (N_5221,N_5012,N_5103);
nand U5222 (N_5222,N_5060,N_5050);
or U5223 (N_5223,N_4992,N_4977);
nor U5224 (N_5224,N_4968,N_4982);
and U5225 (N_5225,N_5039,N_4974);
and U5226 (N_5226,N_4991,N_5058);
and U5227 (N_5227,N_5075,N_5074);
nor U5228 (N_5228,N_4973,N_4963);
xnor U5229 (N_5229,N_5064,N_5083);
nand U5230 (N_5230,N_5068,N_5031);
xnor U5231 (N_5231,N_5081,N_5116);
xnor U5232 (N_5232,N_5038,N_4982);
or U5233 (N_5233,N_5098,N_4981);
xor U5234 (N_5234,N_5094,N_5050);
and U5235 (N_5235,N_5007,N_5077);
xor U5236 (N_5236,N_4985,N_5096);
nor U5237 (N_5237,N_5040,N_5064);
or U5238 (N_5238,N_5081,N_5079);
or U5239 (N_5239,N_5090,N_4970);
xnor U5240 (N_5240,N_5058,N_4996);
nor U5241 (N_5241,N_4985,N_5043);
or U5242 (N_5242,N_5045,N_4981);
or U5243 (N_5243,N_5093,N_4979);
nor U5244 (N_5244,N_5098,N_5051);
xor U5245 (N_5245,N_5016,N_5077);
xnor U5246 (N_5246,N_5028,N_5118);
and U5247 (N_5247,N_5067,N_5104);
xnor U5248 (N_5248,N_5115,N_5029);
nor U5249 (N_5249,N_4979,N_4965);
xor U5250 (N_5250,N_5038,N_4988);
xnor U5251 (N_5251,N_5075,N_4978);
or U5252 (N_5252,N_5063,N_5075);
nand U5253 (N_5253,N_5032,N_5005);
nor U5254 (N_5254,N_5052,N_5022);
nand U5255 (N_5255,N_5099,N_5060);
or U5256 (N_5256,N_5087,N_5099);
xnor U5257 (N_5257,N_5023,N_5066);
xnor U5258 (N_5258,N_5050,N_4970);
xnor U5259 (N_5259,N_5118,N_5021);
xnor U5260 (N_5260,N_4972,N_5095);
nor U5261 (N_5261,N_5039,N_5102);
nor U5262 (N_5262,N_5000,N_5099);
or U5263 (N_5263,N_5085,N_5049);
or U5264 (N_5264,N_4964,N_4965);
nor U5265 (N_5265,N_5030,N_5065);
nor U5266 (N_5266,N_4979,N_4976);
nand U5267 (N_5267,N_5046,N_5004);
nand U5268 (N_5268,N_5110,N_4982);
nor U5269 (N_5269,N_5027,N_5088);
or U5270 (N_5270,N_5021,N_5109);
and U5271 (N_5271,N_5099,N_5045);
and U5272 (N_5272,N_5058,N_5110);
and U5273 (N_5273,N_5072,N_5039);
nand U5274 (N_5274,N_5085,N_5099);
and U5275 (N_5275,N_5070,N_5119);
nor U5276 (N_5276,N_5098,N_4966);
nor U5277 (N_5277,N_5116,N_5037);
nand U5278 (N_5278,N_4965,N_5092);
or U5279 (N_5279,N_5043,N_4990);
nand U5280 (N_5280,N_5262,N_5207);
nand U5281 (N_5281,N_5199,N_5212);
nand U5282 (N_5282,N_5268,N_5228);
nor U5283 (N_5283,N_5139,N_5197);
xnor U5284 (N_5284,N_5180,N_5184);
nand U5285 (N_5285,N_5128,N_5146);
nor U5286 (N_5286,N_5269,N_5270);
nand U5287 (N_5287,N_5263,N_5179);
and U5288 (N_5288,N_5177,N_5126);
xor U5289 (N_5289,N_5244,N_5222);
nor U5290 (N_5290,N_5196,N_5232);
or U5291 (N_5291,N_5276,N_5264);
or U5292 (N_5292,N_5208,N_5153);
or U5293 (N_5293,N_5145,N_5242);
nand U5294 (N_5294,N_5188,N_5267);
xnor U5295 (N_5295,N_5175,N_5141);
xnor U5296 (N_5296,N_5246,N_5178);
nand U5297 (N_5297,N_5190,N_5174);
and U5298 (N_5298,N_5233,N_5223);
xnor U5299 (N_5299,N_5252,N_5278);
nand U5300 (N_5300,N_5189,N_5200);
and U5301 (N_5301,N_5234,N_5271);
xor U5302 (N_5302,N_5221,N_5193);
nand U5303 (N_5303,N_5220,N_5168);
nand U5304 (N_5304,N_5137,N_5202);
nor U5305 (N_5305,N_5226,N_5261);
and U5306 (N_5306,N_5143,N_5227);
or U5307 (N_5307,N_5127,N_5206);
xnor U5308 (N_5308,N_5237,N_5135);
xor U5309 (N_5309,N_5218,N_5272);
xor U5310 (N_5310,N_5253,N_5257);
nor U5311 (N_5311,N_5159,N_5245);
or U5312 (N_5312,N_5192,N_5260);
nand U5313 (N_5313,N_5195,N_5191);
xor U5314 (N_5314,N_5130,N_5140);
nor U5315 (N_5315,N_5120,N_5172);
xnor U5316 (N_5316,N_5254,N_5170);
nor U5317 (N_5317,N_5256,N_5249);
or U5318 (N_5318,N_5204,N_5229);
nor U5319 (N_5319,N_5219,N_5149);
or U5320 (N_5320,N_5185,N_5147);
and U5321 (N_5321,N_5144,N_5131);
and U5322 (N_5322,N_5166,N_5169);
and U5323 (N_5323,N_5123,N_5214);
and U5324 (N_5324,N_5181,N_5125);
nand U5325 (N_5325,N_5156,N_5194);
nand U5326 (N_5326,N_5163,N_5129);
xnor U5327 (N_5327,N_5230,N_5250);
nor U5328 (N_5328,N_5121,N_5225);
xnor U5329 (N_5329,N_5183,N_5162);
nand U5330 (N_5330,N_5186,N_5251);
or U5331 (N_5331,N_5224,N_5157);
or U5332 (N_5332,N_5164,N_5167);
or U5333 (N_5333,N_5236,N_5133);
xnor U5334 (N_5334,N_5255,N_5205);
or U5335 (N_5335,N_5241,N_5160);
or U5336 (N_5336,N_5266,N_5258);
or U5337 (N_5337,N_5279,N_5134);
xor U5338 (N_5338,N_5217,N_5171);
or U5339 (N_5339,N_5238,N_5124);
and U5340 (N_5340,N_5235,N_5273);
xnor U5341 (N_5341,N_5122,N_5136);
nand U5342 (N_5342,N_5148,N_5138);
nand U5343 (N_5343,N_5176,N_5265);
and U5344 (N_5344,N_5158,N_5216);
or U5345 (N_5345,N_5154,N_5239);
nand U5346 (N_5346,N_5150,N_5161);
and U5347 (N_5347,N_5259,N_5274);
xnor U5348 (N_5348,N_5132,N_5243);
or U5349 (N_5349,N_5155,N_5215);
xor U5350 (N_5350,N_5173,N_5248);
and U5351 (N_5351,N_5165,N_5231);
nor U5352 (N_5352,N_5213,N_5182);
nand U5353 (N_5353,N_5198,N_5209);
or U5354 (N_5354,N_5151,N_5142);
and U5355 (N_5355,N_5187,N_5201);
nor U5356 (N_5356,N_5203,N_5275);
and U5357 (N_5357,N_5240,N_5277);
xnor U5358 (N_5358,N_5211,N_5247);
or U5359 (N_5359,N_5210,N_5152);
nand U5360 (N_5360,N_5173,N_5152);
and U5361 (N_5361,N_5143,N_5229);
xnor U5362 (N_5362,N_5245,N_5227);
nor U5363 (N_5363,N_5272,N_5157);
and U5364 (N_5364,N_5147,N_5151);
nand U5365 (N_5365,N_5278,N_5258);
xnor U5366 (N_5366,N_5272,N_5186);
xnor U5367 (N_5367,N_5215,N_5220);
nor U5368 (N_5368,N_5234,N_5133);
or U5369 (N_5369,N_5220,N_5139);
nand U5370 (N_5370,N_5206,N_5176);
nand U5371 (N_5371,N_5184,N_5155);
nor U5372 (N_5372,N_5276,N_5233);
and U5373 (N_5373,N_5275,N_5237);
nor U5374 (N_5374,N_5262,N_5276);
or U5375 (N_5375,N_5212,N_5129);
nor U5376 (N_5376,N_5236,N_5242);
or U5377 (N_5377,N_5153,N_5256);
nand U5378 (N_5378,N_5246,N_5124);
nor U5379 (N_5379,N_5245,N_5232);
xnor U5380 (N_5380,N_5155,N_5196);
or U5381 (N_5381,N_5181,N_5197);
nor U5382 (N_5382,N_5271,N_5208);
or U5383 (N_5383,N_5205,N_5250);
nand U5384 (N_5384,N_5262,N_5264);
nand U5385 (N_5385,N_5220,N_5239);
nor U5386 (N_5386,N_5197,N_5123);
and U5387 (N_5387,N_5181,N_5216);
nor U5388 (N_5388,N_5120,N_5265);
nor U5389 (N_5389,N_5203,N_5164);
or U5390 (N_5390,N_5245,N_5267);
xnor U5391 (N_5391,N_5217,N_5145);
or U5392 (N_5392,N_5198,N_5167);
nand U5393 (N_5393,N_5195,N_5209);
and U5394 (N_5394,N_5165,N_5166);
nor U5395 (N_5395,N_5122,N_5147);
nand U5396 (N_5396,N_5216,N_5251);
nor U5397 (N_5397,N_5246,N_5270);
nor U5398 (N_5398,N_5189,N_5255);
nand U5399 (N_5399,N_5183,N_5218);
nor U5400 (N_5400,N_5161,N_5121);
xnor U5401 (N_5401,N_5221,N_5279);
xnor U5402 (N_5402,N_5155,N_5211);
nand U5403 (N_5403,N_5181,N_5158);
xnor U5404 (N_5404,N_5241,N_5143);
xor U5405 (N_5405,N_5150,N_5279);
nand U5406 (N_5406,N_5236,N_5156);
or U5407 (N_5407,N_5137,N_5182);
and U5408 (N_5408,N_5240,N_5261);
or U5409 (N_5409,N_5145,N_5129);
xor U5410 (N_5410,N_5233,N_5146);
nand U5411 (N_5411,N_5277,N_5190);
xor U5412 (N_5412,N_5158,N_5187);
nand U5413 (N_5413,N_5192,N_5258);
or U5414 (N_5414,N_5120,N_5248);
or U5415 (N_5415,N_5200,N_5248);
xnor U5416 (N_5416,N_5244,N_5224);
nor U5417 (N_5417,N_5195,N_5197);
nor U5418 (N_5418,N_5221,N_5216);
or U5419 (N_5419,N_5157,N_5256);
and U5420 (N_5420,N_5238,N_5150);
or U5421 (N_5421,N_5130,N_5260);
xnor U5422 (N_5422,N_5279,N_5168);
or U5423 (N_5423,N_5206,N_5168);
nand U5424 (N_5424,N_5209,N_5205);
or U5425 (N_5425,N_5170,N_5127);
xnor U5426 (N_5426,N_5152,N_5233);
or U5427 (N_5427,N_5273,N_5157);
or U5428 (N_5428,N_5167,N_5185);
nand U5429 (N_5429,N_5155,N_5239);
and U5430 (N_5430,N_5202,N_5265);
and U5431 (N_5431,N_5224,N_5188);
xnor U5432 (N_5432,N_5274,N_5269);
xor U5433 (N_5433,N_5213,N_5245);
nand U5434 (N_5434,N_5141,N_5172);
and U5435 (N_5435,N_5191,N_5144);
nand U5436 (N_5436,N_5196,N_5137);
nand U5437 (N_5437,N_5267,N_5211);
nor U5438 (N_5438,N_5128,N_5184);
and U5439 (N_5439,N_5204,N_5183);
or U5440 (N_5440,N_5429,N_5425);
xor U5441 (N_5441,N_5325,N_5369);
xnor U5442 (N_5442,N_5301,N_5405);
nand U5443 (N_5443,N_5391,N_5299);
xnor U5444 (N_5444,N_5416,N_5312);
and U5445 (N_5445,N_5439,N_5414);
and U5446 (N_5446,N_5387,N_5359);
nor U5447 (N_5447,N_5404,N_5373);
nor U5448 (N_5448,N_5345,N_5317);
xnor U5449 (N_5449,N_5284,N_5386);
or U5450 (N_5450,N_5367,N_5356);
and U5451 (N_5451,N_5381,N_5407);
xor U5452 (N_5452,N_5287,N_5360);
nor U5453 (N_5453,N_5349,N_5357);
nand U5454 (N_5454,N_5318,N_5298);
and U5455 (N_5455,N_5435,N_5438);
xor U5456 (N_5456,N_5437,N_5344);
nand U5457 (N_5457,N_5358,N_5342);
xor U5458 (N_5458,N_5306,N_5412);
xnor U5459 (N_5459,N_5285,N_5286);
and U5460 (N_5460,N_5341,N_5374);
nand U5461 (N_5461,N_5346,N_5333);
or U5462 (N_5462,N_5324,N_5400);
or U5463 (N_5463,N_5361,N_5427);
nand U5464 (N_5464,N_5422,N_5331);
nand U5465 (N_5465,N_5314,N_5376);
and U5466 (N_5466,N_5303,N_5355);
xnor U5467 (N_5467,N_5431,N_5434);
xnor U5468 (N_5468,N_5280,N_5430);
nor U5469 (N_5469,N_5281,N_5329);
nand U5470 (N_5470,N_5334,N_5378);
xnor U5471 (N_5471,N_5409,N_5340);
xor U5472 (N_5472,N_5348,N_5418);
nand U5473 (N_5473,N_5370,N_5419);
xnor U5474 (N_5474,N_5377,N_5362);
and U5475 (N_5475,N_5410,N_5297);
and U5476 (N_5476,N_5335,N_5415);
nor U5477 (N_5477,N_5402,N_5296);
or U5478 (N_5478,N_5328,N_5403);
nand U5479 (N_5479,N_5315,N_5321);
and U5480 (N_5480,N_5327,N_5350);
and U5481 (N_5481,N_5379,N_5390);
nor U5482 (N_5482,N_5309,N_5411);
nor U5483 (N_5483,N_5283,N_5320);
or U5484 (N_5484,N_5423,N_5323);
nor U5485 (N_5485,N_5347,N_5282);
and U5486 (N_5486,N_5354,N_5294);
nor U5487 (N_5487,N_5396,N_5308);
xor U5488 (N_5488,N_5424,N_5289);
and U5489 (N_5489,N_5421,N_5385);
nor U5490 (N_5490,N_5338,N_5389);
nand U5491 (N_5491,N_5330,N_5426);
or U5492 (N_5492,N_5295,N_5304);
xor U5493 (N_5493,N_5375,N_5392);
and U5494 (N_5494,N_5319,N_5316);
xnor U5495 (N_5495,N_5313,N_5302);
or U5496 (N_5496,N_5388,N_5332);
xor U5497 (N_5497,N_5326,N_5399);
or U5498 (N_5498,N_5288,N_5292);
nand U5499 (N_5499,N_5366,N_5413);
and U5500 (N_5500,N_5428,N_5408);
xnor U5501 (N_5501,N_5406,N_5351);
or U5502 (N_5502,N_5436,N_5433);
xor U5503 (N_5503,N_5384,N_5365);
and U5504 (N_5504,N_5307,N_5432);
or U5505 (N_5505,N_5291,N_5339);
xor U5506 (N_5506,N_5300,N_5352);
and U5507 (N_5507,N_5310,N_5417);
nor U5508 (N_5508,N_5364,N_5393);
nand U5509 (N_5509,N_5395,N_5337);
or U5510 (N_5510,N_5398,N_5401);
or U5511 (N_5511,N_5353,N_5397);
or U5512 (N_5512,N_5305,N_5371);
or U5513 (N_5513,N_5420,N_5290);
and U5514 (N_5514,N_5394,N_5322);
and U5515 (N_5515,N_5363,N_5368);
nor U5516 (N_5516,N_5380,N_5343);
or U5517 (N_5517,N_5311,N_5336);
nor U5518 (N_5518,N_5293,N_5383);
and U5519 (N_5519,N_5382,N_5372);
and U5520 (N_5520,N_5345,N_5407);
xnor U5521 (N_5521,N_5420,N_5288);
xnor U5522 (N_5522,N_5302,N_5351);
or U5523 (N_5523,N_5427,N_5385);
xnor U5524 (N_5524,N_5304,N_5315);
nor U5525 (N_5525,N_5415,N_5401);
nor U5526 (N_5526,N_5401,N_5285);
nand U5527 (N_5527,N_5340,N_5413);
xnor U5528 (N_5528,N_5388,N_5347);
nand U5529 (N_5529,N_5304,N_5311);
and U5530 (N_5530,N_5305,N_5353);
and U5531 (N_5531,N_5340,N_5291);
or U5532 (N_5532,N_5306,N_5300);
and U5533 (N_5533,N_5401,N_5336);
nand U5534 (N_5534,N_5367,N_5418);
xnor U5535 (N_5535,N_5354,N_5344);
or U5536 (N_5536,N_5409,N_5354);
nand U5537 (N_5537,N_5296,N_5290);
or U5538 (N_5538,N_5366,N_5402);
nor U5539 (N_5539,N_5367,N_5382);
and U5540 (N_5540,N_5388,N_5354);
or U5541 (N_5541,N_5308,N_5342);
xnor U5542 (N_5542,N_5282,N_5319);
xor U5543 (N_5543,N_5344,N_5377);
or U5544 (N_5544,N_5317,N_5408);
nand U5545 (N_5545,N_5285,N_5289);
nor U5546 (N_5546,N_5428,N_5336);
and U5547 (N_5547,N_5384,N_5406);
or U5548 (N_5548,N_5319,N_5435);
nand U5549 (N_5549,N_5410,N_5413);
or U5550 (N_5550,N_5290,N_5292);
or U5551 (N_5551,N_5289,N_5349);
nand U5552 (N_5552,N_5289,N_5306);
xnor U5553 (N_5553,N_5318,N_5376);
nand U5554 (N_5554,N_5297,N_5429);
nor U5555 (N_5555,N_5308,N_5313);
or U5556 (N_5556,N_5345,N_5342);
nor U5557 (N_5557,N_5356,N_5338);
nor U5558 (N_5558,N_5392,N_5290);
nand U5559 (N_5559,N_5337,N_5430);
and U5560 (N_5560,N_5417,N_5326);
nor U5561 (N_5561,N_5424,N_5317);
xnor U5562 (N_5562,N_5401,N_5341);
nand U5563 (N_5563,N_5294,N_5415);
nand U5564 (N_5564,N_5358,N_5408);
nand U5565 (N_5565,N_5434,N_5309);
and U5566 (N_5566,N_5425,N_5294);
nor U5567 (N_5567,N_5290,N_5297);
or U5568 (N_5568,N_5331,N_5344);
and U5569 (N_5569,N_5335,N_5318);
xor U5570 (N_5570,N_5309,N_5345);
nor U5571 (N_5571,N_5341,N_5350);
xor U5572 (N_5572,N_5406,N_5423);
xor U5573 (N_5573,N_5334,N_5288);
nor U5574 (N_5574,N_5430,N_5413);
xor U5575 (N_5575,N_5432,N_5438);
nand U5576 (N_5576,N_5398,N_5337);
nand U5577 (N_5577,N_5285,N_5346);
and U5578 (N_5578,N_5317,N_5342);
xor U5579 (N_5579,N_5297,N_5313);
and U5580 (N_5580,N_5419,N_5355);
nand U5581 (N_5581,N_5345,N_5394);
nor U5582 (N_5582,N_5382,N_5355);
xnor U5583 (N_5583,N_5327,N_5428);
xnor U5584 (N_5584,N_5339,N_5384);
nor U5585 (N_5585,N_5379,N_5317);
nand U5586 (N_5586,N_5373,N_5378);
or U5587 (N_5587,N_5309,N_5286);
and U5588 (N_5588,N_5287,N_5389);
or U5589 (N_5589,N_5386,N_5342);
and U5590 (N_5590,N_5341,N_5421);
and U5591 (N_5591,N_5395,N_5393);
and U5592 (N_5592,N_5302,N_5362);
xor U5593 (N_5593,N_5345,N_5283);
xnor U5594 (N_5594,N_5303,N_5435);
nand U5595 (N_5595,N_5337,N_5386);
xor U5596 (N_5596,N_5381,N_5431);
or U5597 (N_5597,N_5339,N_5335);
xor U5598 (N_5598,N_5301,N_5433);
nand U5599 (N_5599,N_5295,N_5398);
nand U5600 (N_5600,N_5575,N_5581);
nand U5601 (N_5601,N_5565,N_5588);
or U5602 (N_5602,N_5564,N_5510);
nand U5603 (N_5603,N_5506,N_5508);
nor U5604 (N_5604,N_5444,N_5459);
nand U5605 (N_5605,N_5549,N_5519);
nand U5606 (N_5606,N_5532,N_5490);
or U5607 (N_5607,N_5572,N_5596);
or U5608 (N_5608,N_5579,N_5460);
nand U5609 (N_5609,N_5563,N_5523);
and U5610 (N_5610,N_5471,N_5516);
nor U5611 (N_5611,N_5528,N_5480);
or U5612 (N_5612,N_5441,N_5598);
nor U5613 (N_5613,N_5451,N_5538);
nand U5614 (N_5614,N_5507,N_5470);
and U5615 (N_5615,N_5570,N_5560);
and U5616 (N_5616,N_5501,N_5509);
nor U5617 (N_5617,N_5513,N_5592);
nand U5618 (N_5618,N_5478,N_5529);
nor U5619 (N_5619,N_5461,N_5525);
xor U5620 (N_5620,N_5531,N_5553);
xnor U5621 (N_5621,N_5558,N_5540);
xnor U5622 (N_5622,N_5494,N_5554);
xnor U5623 (N_5623,N_5476,N_5517);
xor U5624 (N_5624,N_5449,N_5484);
nand U5625 (N_5625,N_5491,N_5520);
and U5626 (N_5626,N_5534,N_5547);
nor U5627 (N_5627,N_5556,N_5548);
or U5628 (N_5628,N_5530,N_5445);
nor U5629 (N_5629,N_5473,N_5469);
nand U5630 (N_5630,N_5551,N_5504);
nand U5631 (N_5631,N_5442,N_5580);
nor U5632 (N_5632,N_5566,N_5550);
nand U5633 (N_5633,N_5477,N_5489);
xor U5634 (N_5634,N_5485,N_5521);
or U5635 (N_5635,N_5511,N_5535);
and U5636 (N_5636,N_5479,N_5440);
nand U5637 (N_5637,N_5541,N_5487);
nand U5638 (N_5638,N_5464,N_5533);
xor U5639 (N_5639,N_5512,N_5537);
nand U5640 (N_5640,N_5522,N_5542);
and U5641 (N_5641,N_5591,N_5498);
nor U5642 (N_5642,N_5536,N_5552);
or U5643 (N_5643,N_5595,N_5544);
or U5644 (N_5644,N_5545,N_5467);
and U5645 (N_5645,N_5562,N_5455);
and U5646 (N_5646,N_5497,N_5527);
and U5647 (N_5647,N_5447,N_5569);
nor U5648 (N_5648,N_5567,N_5495);
xor U5649 (N_5649,N_5499,N_5446);
and U5650 (N_5650,N_5472,N_5492);
or U5651 (N_5651,N_5597,N_5474);
nand U5652 (N_5652,N_5493,N_5546);
and U5653 (N_5653,N_5524,N_5594);
nand U5654 (N_5654,N_5456,N_5574);
or U5655 (N_5655,N_5568,N_5593);
or U5656 (N_5656,N_5515,N_5454);
nor U5657 (N_5657,N_5584,N_5559);
nand U5658 (N_5658,N_5443,N_5457);
xor U5659 (N_5659,N_5571,N_5573);
xor U5660 (N_5660,N_5483,N_5488);
or U5661 (N_5661,N_5543,N_5496);
nand U5662 (N_5662,N_5578,N_5500);
nand U5663 (N_5663,N_5463,N_5458);
xnor U5664 (N_5664,N_5590,N_5599);
or U5665 (N_5665,N_5586,N_5448);
xnor U5666 (N_5666,N_5468,N_5481);
nand U5667 (N_5667,N_5557,N_5576);
and U5668 (N_5668,N_5502,N_5526);
nand U5669 (N_5669,N_5503,N_5518);
xnor U5670 (N_5670,N_5452,N_5583);
nor U5671 (N_5671,N_5514,N_5587);
nand U5672 (N_5672,N_5505,N_5453);
and U5673 (N_5673,N_5450,N_5466);
xnor U5674 (N_5674,N_5482,N_5539);
and U5675 (N_5675,N_5465,N_5475);
xor U5676 (N_5676,N_5577,N_5555);
and U5677 (N_5677,N_5486,N_5582);
nand U5678 (N_5678,N_5561,N_5462);
and U5679 (N_5679,N_5589,N_5585);
and U5680 (N_5680,N_5474,N_5460);
or U5681 (N_5681,N_5511,N_5569);
or U5682 (N_5682,N_5475,N_5506);
xor U5683 (N_5683,N_5566,N_5528);
and U5684 (N_5684,N_5568,N_5518);
and U5685 (N_5685,N_5445,N_5480);
and U5686 (N_5686,N_5475,N_5504);
or U5687 (N_5687,N_5561,N_5514);
xnor U5688 (N_5688,N_5595,N_5561);
or U5689 (N_5689,N_5451,N_5480);
xor U5690 (N_5690,N_5583,N_5443);
xor U5691 (N_5691,N_5536,N_5590);
xnor U5692 (N_5692,N_5571,N_5456);
or U5693 (N_5693,N_5446,N_5458);
nor U5694 (N_5694,N_5510,N_5443);
nand U5695 (N_5695,N_5458,N_5537);
nor U5696 (N_5696,N_5539,N_5519);
nor U5697 (N_5697,N_5464,N_5591);
nand U5698 (N_5698,N_5558,N_5582);
nand U5699 (N_5699,N_5493,N_5547);
nand U5700 (N_5700,N_5477,N_5509);
xnor U5701 (N_5701,N_5592,N_5471);
nand U5702 (N_5702,N_5530,N_5517);
nor U5703 (N_5703,N_5579,N_5559);
nor U5704 (N_5704,N_5518,N_5570);
nor U5705 (N_5705,N_5457,N_5476);
and U5706 (N_5706,N_5526,N_5443);
xor U5707 (N_5707,N_5525,N_5521);
nor U5708 (N_5708,N_5519,N_5541);
nand U5709 (N_5709,N_5572,N_5500);
xnor U5710 (N_5710,N_5445,N_5577);
or U5711 (N_5711,N_5583,N_5471);
nand U5712 (N_5712,N_5591,N_5478);
nor U5713 (N_5713,N_5532,N_5546);
and U5714 (N_5714,N_5514,N_5543);
xnor U5715 (N_5715,N_5542,N_5478);
and U5716 (N_5716,N_5480,N_5497);
nand U5717 (N_5717,N_5504,N_5510);
nand U5718 (N_5718,N_5494,N_5592);
or U5719 (N_5719,N_5513,N_5499);
xor U5720 (N_5720,N_5509,N_5475);
and U5721 (N_5721,N_5562,N_5516);
nor U5722 (N_5722,N_5487,N_5593);
or U5723 (N_5723,N_5549,N_5477);
xnor U5724 (N_5724,N_5464,N_5498);
nand U5725 (N_5725,N_5596,N_5584);
and U5726 (N_5726,N_5572,N_5508);
xor U5727 (N_5727,N_5475,N_5576);
nand U5728 (N_5728,N_5474,N_5453);
nand U5729 (N_5729,N_5489,N_5595);
or U5730 (N_5730,N_5524,N_5591);
or U5731 (N_5731,N_5555,N_5590);
or U5732 (N_5732,N_5495,N_5534);
nor U5733 (N_5733,N_5560,N_5565);
or U5734 (N_5734,N_5596,N_5533);
and U5735 (N_5735,N_5577,N_5501);
nand U5736 (N_5736,N_5461,N_5456);
and U5737 (N_5737,N_5506,N_5452);
and U5738 (N_5738,N_5467,N_5487);
xnor U5739 (N_5739,N_5514,N_5502);
and U5740 (N_5740,N_5468,N_5447);
and U5741 (N_5741,N_5548,N_5592);
nor U5742 (N_5742,N_5514,N_5598);
xor U5743 (N_5743,N_5473,N_5509);
nand U5744 (N_5744,N_5591,N_5574);
or U5745 (N_5745,N_5561,N_5448);
nor U5746 (N_5746,N_5474,N_5525);
nand U5747 (N_5747,N_5586,N_5506);
and U5748 (N_5748,N_5461,N_5527);
and U5749 (N_5749,N_5581,N_5566);
nand U5750 (N_5750,N_5503,N_5494);
or U5751 (N_5751,N_5539,N_5598);
and U5752 (N_5752,N_5576,N_5593);
nand U5753 (N_5753,N_5583,N_5445);
and U5754 (N_5754,N_5531,N_5530);
or U5755 (N_5755,N_5477,N_5455);
and U5756 (N_5756,N_5487,N_5496);
nand U5757 (N_5757,N_5505,N_5462);
or U5758 (N_5758,N_5483,N_5521);
and U5759 (N_5759,N_5557,N_5475);
xor U5760 (N_5760,N_5664,N_5693);
nor U5761 (N_5761,N_5744,N_5750);
nor U5762 (N_5762,N_5642,N_5681);
and U5763 (N_5763,N_5609,N_5671);
nor U5764 (N_5764,N_5721,N_5648);
nor U5765 (N_5765,N_5646,N_5618);
nor U5766 (N_5766,N_5653,N_5702);
nor U5767 (N_5767,N_5748,N_5705);
xnor U5768 (N_5768,N_5698,N_5651);
and U5769 (N_5769,N_5704,N_5747);
nand U5770 (N_5770,N_5640,N_5746);
or U5771 (N_5771,N_5611,N_5650);
nor U5772 (N_5772,N_5674,N_5645);
xor U5773 (N_5773,N_5628,N_5659);
xor U5774 (N_5774,N_5752,N_5658);
or U5775 (N_5775,N_5652,N_5633);
nor U5776 (N_5776,N_5603,N_5635);
xnor U5777 (N_5777,N_5729,N_5639);
nand U5778 (N_5778,N_5685,N_5662);
and U5779 (N_5779,N_5684,N_5686);
nand U5780 (N_5780,N_5703,N_5757);
nand U5781 (N_5781,N_5696,N_5695);
xnor U5782 (N_5782,N_5690,N_5665);
and U5783 (N_5783,N_5753,N_5682);
nand U5784 (N_5784,N_5656,N_5619);
or U5785 (N_5785,N_5709,N_5631);
or U5786 (N_5786,N_5742,N_5676);
nand U5787 (N_5787,N_5608,N_5740);
nor U5788 (N_5788,N_5636,N_5714);
nand U5789 (N_5789,N_5745,N_5719);
xor U5790 (N_5790,N_5616,N_5623);
nand U5791 (N_5791,N_5755,N_5604);
or U5792 (N_5792,N_5673,N_5624);
and U5793 (N_5793,N_5722,N_5758);
or U5794 (N_5794,N_5672,N_5660);
nand U5795 (N_5795,N_5622,N_5680);
nor U5796 (N_5796,N_5728,N_5675);
nor U5797 (N_5797,N_5710,N_5654);
nor U5798 (N_5798,N_5670,N_5718);
or U5799 (N_5799,N_5661,N_5649);
or U5800 (N_5800,N_5734,N_5739);
nor U5801 (N_5801,N_5699,N_5625);
nand U5802 (N_5802,N_5638,N_5629);
nor U5803 (N_5803,N_5712,N_5706);
nand U5804 (N_5804,N_5663,N_5620);
xnor U5805 (N_5805,N_5741,N_5730);
nand U5806 (N_5806,N_5727,N_5621);
xor U5807 (N_5807,N_5689,N_5708);
or U5808 (N_5808,N_5683,N_5614);
or U5809 (N_5809,N_5617,N_5700);
nor U5810 (N_5810,N_5657,N_5668);
or U5811 (N_5811,N_5627,N_5600);
and U5812 (N_5812,N_5725,N_5759);
nor U5813 (N_5813,N_5641,N_5756);
or U5814 (N_5814,N_5692,N_5688);
xnor U5815 (N_5815,N_5726,N_5711);
and U5816 (N_5816,N_5632,N_5723);
nor U5817 (N_5817,N_5751,N_5601);
xnor U5818 (N_5818,N_5605,N_5738);
or U5819 (N_5819,N_5694,N_5743);
or U5820 (N_5820,N_5717,N_5731);
nor U5821 (N_5821,N_5691,N_5687);
or U5822 (N_5822,N_5630,N_5754);
nand U5823 (N_5823,N_5613,N_5602);
nand U5824 (N_5824,N_5724,N_5607);
or U5825 (N_5825,N_5733,N_5644);
and U5826 (N_5826,N_5677,N_5637);
xor U5827 (N_5827,N_5716,N_5735);
nor U5828 (N_5828,N_5643,N_5610);
and U5829 (N_5829,N_5720,N_5615);
nor U5830 (N_5830,N_5697,N_5655);
nand U5831 (N_5831,N_5626,N_5666);
and U5832 (N_5832,N_5737,N_5749);
xor U5833 (N_5833,N_5713,N_5669);
and U5834 (N_5834,N_5707,N_5634);
nor U5835 (N_5835,N_5701,N_5606);
and U5836 (N_5836,N_5612,N_5736);
or U5837 (N_5837,N_5715,N_5732);
xnor U5838 (N_5838,N_5679,N_5647);
and U5839 (N_5839,N_5667,N_5678);
nand U5840 (N_5840,N_5718,N_5739);
xor U5841 (N_5841,N_5728,N_5749);
and U5842 (N_5842,N_5610,N_5641);
nand U5843 (N_5843,N_5660,N_5729);
xor U5844 (N_5844,N_5618,N_5757);
nor U5845 (N_5845,N_5733,N_5604);
xnor U5846 (N_5846,N_5682,N_5726);
and U5847 (N_5847,N_5747,N_5647);
nand U5848 (N_5848,N_5623,N_5684);
nand U5849 (N_5849,N_5629,N_5675);
and U5850 (N_5850,N_5640,N_5677);
xnor U5851 (N_5851,N_5637,N_5747);
nand U5852 (N_5852,N_5653,N_5663);
and U5853 (N_5853,N_5623,N_5712);
nor U5854 (N_5854,N_5696,N_5759);
nand U5855 (N_5855,N_5726,N_5619);
xnor U5856 (N_5856,N_5679,N_5664);
xnor U5857 (N_5857,N_5713,N_5638);
or U5858 (N_5858,N_5625,N_5663);
and U5859 (N_5859,N_5664,N_5672);
nor U5860 (N_5860,N_5685,N_5749);
xor U5861 (N_5861,N_5636,N_5651);
nor U5862 (N_5862,N_5620,N_5647);
xor U5863 (N_5863,N_5731,N_5675);
nand U5864 (N_5864,N_5748,N_5616);
and U5865 (N_5865,N_5658,N_5640);
xor U5866 (N_5866,N_5742,N_5667);
nand U5867 (N_5867,N_5725,N_5621);
nor U5868 (N_5868,N_5656,N_5749);
or U5869 (N_5869,N_5707,N_5714);
nor U5870 (N_5870,N_5631,N_5608);
and U5871 (N_5871,N_5758,N_5673);
or U5872 (N_5872,N_5736,N_5635);
xor U5873 (N_5873,N_5723,N_5653);
xor U5874 (N_5874,N_5608,N_5687);
xnor U5875 (N_5875,N_5730,N_5615);
xnor U5876 (N_5876,N_5645,N_5751);
xor U5877 (N_5877,N_5618,N_5743);
or U5878 (N_5878,N_5752,N_5709);
xor U5879 (N_5879,N_5677,N_5751);
nor U5880 (N_5880,N_5660,N_5716);
or U5881 (N_5881,N_5669,N_5692);
and U5882 (N_5882,N_5697,N_5724);
nor U5883 (N_5883,N_5726,N_5614);
or U5884 (N_5884,N_5669,N_5675);
or U5885 (N_5885,N_5652,N_5700);
or U5886 (N_5886,N_5735,N_5638);
and U5887 (N_5887,N_5669,N_5664);
nor U5888 (N_5888,N_5738,N_5732);
nand U5889 (N_5889,N_5611,N_5601);
xnor U5890 (N_5890,N_5751,N_5657);
nor U5891 (N_5891,N_5670,N_5698);
xnor U5892 (N_5892,N_5741,N_5617);
and U5893 (N_5893,N_5654,N_5730);
and U5894 (N_5894,N_5683,N_5694);
and U5895 (N_5895,N_5600,N_5654);
or U5896 (N_5896,N_5730,N_5755);
nand U5897 (N_5897,N_5646,N_5663);
or U5898 (N_5898,N_5613,N_5620);
xnor U5899 (N_5899,N_5704,N_5751);
xor U5900 (N_5900,N_5725,N_5664);
nand U5901 (N_5901,N_5613,N_5706);
nor U5902 (N_5902,N_5748,N_5625);
and U5903 (N_5903,N_5606,N_5679);
or U5904 (N_5904,N_5636,N_5722);
nand U5905 (N_5905,N_5686,N_5720);
and U5906 (N_5906,N_5657,N_5670);
nor U5907 (N_5907,N_5605,N_5632);
and U5908 (N_5908,N_5710,N_5711);
xnor U5909 (N_5909,N_5717,N_5677);
and U5910 (N_5910,N_5607,N_5622);
nand U5911 (N_5911,N_5715,N_5627);
nand U5912 (N_5912,N_5681,N_5607);
and U5913 (N_5913,N_5650,N_5737);
nor U5914 (N_5914,N_5702,N_5681);
nand U5915 (N_5915,N_5661,N_5690);
and U5916 (N_5916,N_5643,N_5750);
nand U5917 (N_5917,N_5642,N_5643);
nand U5918 (N_5918,N_5661,N_5716);
nor U5919 (N_5919,N_5628,N_5623);
nor U5920 (N_5920,N_5813,N_5778);
and U5921 (N_5921,N_5860,N_5911);
and U5922 (N_5922,N_5800,N_5843);
nor U5923 (N_5923,N_5831,N_5766);
nor U5924 (N_5924,N_5865,N_5789);
nor U5925 (N_5925,N_5895,N_5799);
nand U5926 (N_5926,N_5822,N_5819);
nor U5927 (N_5927,N_5892,N_5796);
and U5928 (N_5928,N_5883,N_5887);
xnor U5929 (N_5929,N_5891,N_5889);
and U5930 (N_5930,N_5830,N_5797);
xor U5931 (N_5931,N_5795,N_5802);
nand U5932 (N_5932,N_5863,N_5881);
xnor U5933 (N_5933,N_5784,N_5825);
xnor U5934 (N_5934,N_5878,N_5806);
nor U5935 (N_5935,N_5852,N_5905);
and U5936 (N_5936,N_5762,N_5893);
nand U5937 (N_5937,N_5851,N_5815);
or U5938 (N_5938,N_5885,N_5846);
nor U5939 (N_5939,N_5868,N_5782);
xor U5940 (N_5940,N_5788,N_5876);
nand U5941 (N_5941,N_5809,N_5828);
or U5942 (N_5942,N_5760,N_5818);
and U5943 (N_5943,N_5904,N_5888);
nor U5944 (N_5944,N_5859,N_5803);
or U5945 (N_5945,N_5907,N_5875);
nand U5946 (N_5946,N_5804,N_5879);
or U5947 (N_5947,N_5785,N_5835);
nor U5948 (N_5948,N_5764,N_5787);
and U5949 (N_5949,N_5847,N_5770);
nor U5950 (N_5950,N_5914,N_5783);
nand U5951 (N_5951,N_5772,N_5910);
and U5952 (N_5952,N_5861,N_5824);
nor U5953 (N_5953,N_5816,N_5873);
or U5954 (N_5954,N_5842,N_5850);
xor U5955 (N_5955,N_5768,N_5821);
nand U5956 (N_5956,N_5849,N_5886);
nor U5957 (N_5957,N_5794,N_5871);
nand U5958 (N_5958,N_5894,N_5781);
xnor U5959 (N_5959,N_5839,N_5902);
xnor U5960 (N_5960,N_5912,N_5882);
nor U5961 (N_5961,N_5916,N_5771);
xor U5962 (N_5962,N_5792,N_5901);
nor U5963 (N_5963,N_5844,N_5823);
nor U5964 (N_5964,N_5811,N_5864);
nand U5965 (N_5965,N_5870,N_5855);
or U5966 (N_5966,N_5909,N_5791);
and U5967 (N_5967,N_5820,N_5853);
or U5968 (N_5968,N_5856,N_5836);
or U5969 (N_5969,N_5805,N_5918);
nand U5970 (N_5970,N_5906,N_5786);
nand U5971 (N_5971,N_5840,N_5898);
xnor U5972 (N_5972,N_5817,N_5812);
nor U5973 (N_5973,N_5913,N_5777);
xor U5974 (N_5974,N_5845,N_5899);
or U5975 (N_5975,N_5807,N_5769);
nand U5976 (N_5976,N_5874,N_5884);
nand U5977 (N_5977,N_5765,N_5763);
nand U5978 (N_5978,N_5773,N_5775);
nand U5979 (N_5979,N_5779,N_5872);
xnor U5980 (N_5980,N_5767,N_5854);
and U5981 (N_5981,N_5880,N_5867);
and U5982 (N_5982,N_5866,N_5832);
xor U5983 (N_5983,N_5808,N_5917);
nor U5984 (N_5984,N_5838,N_5897);
or U5985 (N_5985,N_5848,N_5908);
nor U5986 (N_5986,N_5810,N_5826);
nand U5987 (N_5987,N_5761,N_5869);
xnor U5988 (N_5988,N_5776,N_5900);
or U5989 (N_5989,N_5857,N_5919);
xnor U5990 (N_5990,N_5858,N_5890);
nand U5991 (N_5991,N_5877,N_5780);
or U5992 (N_5992,N_5827,N_5774);
nand U5993 (N_5993,N_5896,N_5837);
xnor U5994 (N_5994,N_5793,N_5915);
or U5995 (N_5995,N_5798,N_5833);
nand U5996 (N_5996,N_5790,N_5801);
or U5997 (N_5997,N_5862,N_5829);
xnor U5998 (N_5998,N_5903,N_5841);
nand U5999 (N_5999,N_5834,N_5814);
or U6000 (N_6000,N_5887,N_5785);
nand U6001 (N_6001,N_5798,N_5891);
nor U6002 (N_6002,N_5892,N_5791);
xor U6003 (N_6003,N_5784,N_5777);
nand U6004 (N_6004,N_5768,N_5901);
nor U6005 (N_6005,N_5853,N_5810);
or U6006 (N_6006,N_5859,N_5760);
and U6007 (N_6007,N_5913,N_5770);
xnor U6008 (N_6008,N_5833,N_5909);
nor U6009 (N_6009,N_5898,N_5776);
nand U6010 (N_6010,N_5779,N_5890);
xnor U6011 (N_6011,N_5892,N_5899);
nor U6012 (N_6012,N_5845,N_5843);
nor U6013 (N_6013,N_5875,N_5772);
and U6014 (N_6014,N_5830,N_5782);
and U6015 (N_6015,N_5843,N_5809);
nor U6016 (N_6016,N_5866,N_5895);
xnor U6017 (N_6017,N_5867,N_5909);
or U6018 (N_6018,N_5902,N_5802);
xnor U6019 (N_6019,N_5805,N_5862);
nor U6020 (N_6020,N_5874,N_5837);
or U6021 (N_6021,N_5761,N_5810);
xor U6022 (N_6022,N_5874,N_5771);
and U6023 (N_6023,N_5904,N_5918);
nor U6024 (N_6024,N_5825,N_5889);
nor U6025 (N_6025,N_5828,N_5824);
xnor U6026 (N_6026,N_5909,N_5884);
nand U6027 (N_6027,N_5852,N_5859);
nand U6028 (N_6028,N_5830,N_5852);
and U6029 (N_6029,N_5876,N_5835);
nor U6030 (N_6030,N_5778,N_5882);
or U6031 (N_6031,N_5865,N_5854);
nor U6032 (N_6032,N_5781,N_5776);
xnor U6033 (N_6033,N_5790,N_5762);
nand U6034 (N_6034,N_5811,N_5761);
nor U6035 (N_6035,N_5910,N_5795);
or U6036 (N_6036,N_5897,N_5865);
nor U6037 (N_6037,N_5813,N_5809);
and U6038 (N_6038,N_5903,N_5822);
xnor U6039 (N_6039,N_5838,N_5916);
or U6040 (N_6040,N_5814,N_5849);
xor U6041 (N_6041,N_5789,N_5850);
nand U6042 (N_6042,N_5918,N_5898);
or U6043 (N_6043,N_5825,N_5826);
and U6044 (N_6044,N_5847,N_5833);
xor U6045 (N_6045,N_5761,N_5865);
or U6046 (N_6046,N_5804,N_5832);
nand U6047 (N_6047,N_5787,N_5855);
nand U6048 (N_6048,N_5874,N_5861);
nand U6049 (N_6049,N_5806,N_5814);
nand U6050 (N_6050,N_5842,N_5774);
nand U6051 (N_6051,N_5901,N_5817);
nand U6052 (N_6052,N_5899,N_5780);
nor U6053 (N_6053,N_5884,N_5860);
and U6054 (N_6054,N_5770,N_5797);
xor U6055 (N_6055,N_5914,N_5901);
or U6056 (N_6056,N_5794,N_5822);
nand U6057 (N_6057,N_5909,N_5774);
xnor U6058 (N_6058,N_5909,N_5858);
and U6059 (N_6059,N_5842,N_5811);
or U6060 (N_6060,N_5866,N_5794);
and U6061 (N_6061,N_5896,N_5909);
and U6062 (N_6062,N_5877,N_5870);
nand U6063 (N_6063,N_5903,N_5917);
and U6064 (N_6064,N_5906,N_5848);
and U6065 (N_6065,N_5882,N_5859);
and U6066 (N_6066,N_5845,N_5916);
or U6067 (N_6067,N_5775,N_5854);
or U6068 (N_6068,N_5916,N_5867);
xnor U6069 (N_6069,N_5899,N_5884);
or U6070 (N_6070,N_5911,N_5836);
and U6071 (N_6071,N_5803,N_5800);
nor U6072 (N_6072,N_5825,N_5919);
or U6073 (N_6073,N_5895,N_5767);
xnor U6074 (N_6074,N_5788,N_5835);
nor U6075 (N_6075,N_5832,N_5812);
xor U6076 (N_6076,N_5799,N_5892);
or U6077 (N_6077,N_5916,N_5817);
and U6078 (N_6078,N_5833,N_5903);
nor U6079 (N_6079,N_5846,N_5854);
nor U6080 (N_6080,N_5956,N_5986);
nor U6081 (N_6081,N_6058,N_5974);
nand U6082 (N_6082,N_5988,N_6022);
nor U6083 (N_6083,N_5996,N_6019);
and U6084 (N_6084,N_6012,N_5925);
nor U6085 (N_6085,N_5972,N_5934);
nand U6086 (N_6086,N_5955,N_5982);
xor U6087 (N_6087,N_5923,N_5948);
and U6088 (N_6088,N_5951,N_6028);
or U6089 (N_6089,N_6009,N_6056);
or U6090 (N_6090,N_6062,N_6006);
nand U6091 (N_6091,N_6035,N_6011);
xor U6092 (N_6092,N_5924,N_6023);
xnor U6093 (N_6093,N_5940,N_5950);
or U6094 (N_6094,N_6059,N_5946);
or U6095 (N_6095,N_5929,N_6076);
nor U6096 (N_6096,N_5998,N_6048);
nand U6097 (N_6097,N_5999,N_6067);
and U6098 (N_6098,N_5949,N_6003);
nor U6099 (N_6099,N_5971,N_5963);
nor U6100 (N_6100,N_5933,N_6046);
nand U6101 (N_6101,N_6057,N_5975);
nand U6102 (N_6102,N_5927,N_6013);
nor U6103 (N_6103,N_6075,N_5993);
and U6104 (N_6104,N_5990,N_6039);
or U6105 (N_6105,N_5960,N_6029);
nor U6106 (N_6106,N_5964,N_6033);
nand U6107 (N_6107,N_5966,N_5961);
xor U6108 (N_6108,N_6070,N_6038);
nor U6109 (N_6109,N_5939,N_5997);
nor U6110 (N_6110,N_6027,N_6002);
xnor U6111 (N_6111,N_5926,N_5984);
nor U6112 (N_6112,N_5928,N_5991);
nand U6113 (N_6113,N_6040,N_6065);
and U6114 (N_6114,N_5977,N_6015);
xnor U6115 (N_6115,N_6073,N_5957);
nor U6116 (N_6116,N_5969,N_5935);
xnor U6117 (N_6117,N_5994,N_6037);
xnor U6118 (N_6118,N_5947,N_6026);
and U6119 (N_6119,N_5922,N_6021);
and U6120 (N_6120,N_6000,N_6071);
or U6121 (N_6121,N_5941,N_6066);
nor U6122 (N_6122,N_5958,N_5962);
nand U6123 (N_6123,N_6042,N_6079);
and U6124 (N_6124,N_6049,N_5920);
or U6125 (N_6125,N_5973,N_6041);
xor U6126 (N_6126,N_5967,N_6050);
or U6127 (N_6127,N_6034,N_5945);
and U6128 (N_6128,N_5983,N_6055);
or U6129 (N_6129,N_6030,N_5981);
xor U6130 (N_6130,N_6016,N_5989);
xnor U6131 (N_6131,N_6044,N_5979);
nand U6132 (N_6132,N_5976,N_6051);
nor U6133 (N_6133,N_5959,N_5936);
nand U6134 (N_6134,N_6024,N_6032);
or U6135 (N_6135,N_5980,N_6063);
xor U6136 (N_6136,N_6025,N_6064);
nand U6137 (N_6137,N_5970,N_5953);
xor U6138 (N_6138,N_6052,N_6005);
nand U6139 (N_6139,N_6001,N_5944);
and U6140 (N_6140,N_6010,N_5938);
nor U6141 (N_6141,N_5985,N_5995);
and U6142 (N_6142,N_6018,N_5921);
xor U6143 (N_6143,N_6072,N_5987);
nor U6144 (N_6144,N_5965,N_5932);
nand U6145 (N_6145,N_5943,N_5954);
nor U6146 (N_6146,N_6069,N_6014);
nor U6147 (N_6147,N_6068,N_6054);
or U6148 (N_6148,N_6045,N_5937);
nand U6149 (N_6149,N_6008,N_6078);
and U6150 (N_6150,N_6061,N_5952);
or U6151 (N_6151,N_6077,N_5942);
nand U6152 (N_6152,N_6074,N_6007);
xnor U6153 (N_6153,N_5978,N_6036);
and U6154 (N_6154,N_6047,N_6060);
nand U6155 (N_6155,N_6043,N_6020);
nor U6156 (N_6156,N_6004,N_5931);
or U6157 (N_6157,N_6017,N_5968);
nor U6158 (N_6158,N_5930,N_6053);
nor U6159 (N_6159,N_5992,N_6031);
nor U6160 (N_6160,N_5985,N_5990);
or U6161 (N_6161,N_6040,N_5993);
or U6162 (N_6162,N_6023,N_5987);
xor U6163 (N_6163,N_6023,N_5968);
nand U6164 (N_6164,N_6002,N_6057);
nand U6165 (N_6165,N_5978,N_6065);
xnor U6166 (N_6166,N_5945,N_6023);
and U6167 (N_6167,N_6025,N_6022);
and U6168 (N_6168,N_6041,N_5956);
and U6169 (N_6169,N_5957,N_6025);
nand U6170 (N_6170,N_6039,N_5925);
or U6171 (N_6171,N_6060,N_6048);
nor U6172 (N_6172,N_6050,N_6041);
nand U6173 (N_6173,N_5993,N_6030);
nor U6174 (N_6174,N_6015,N_6046);
nor U6175 (N_6175,N_6019,N_6029);
xnor U6176 (N_6176,N_6073,N_6074);
nor U6177 (N_6177,N_5981,N_6069);
nor U6178 (N_6178,N_5965,N_5946);
nor U6179 (N_6179,N_6047,N_6075);
xor U6180 (N_6180,N_6018,N_5927);
xnor U6181 (N_6181,N_6058,N_6053);
and U6182 (N_6182,N_5961,N_5938);
nand U6183 (N_6183,N_5939,N_6053);
or U6184 (N_6184,N_6054,N_6021);
nor U6185 (N_6185,N_6005,N_5923);
and U6186 (N_6186,N_6032,N_5974);
xor U6187 (N_6187,N_5984,N_6029);
xnor U6188 (N_6188,N_6072,N_5979);
nand U6189 (N_6189,N_6055,N_5976);
nand U6190 (N_6190,N_5966,N_5976);
or U6191 (N_6191,N_6009,N_5995);
or U6192 (N_6192,N_6048,N_5982);
nand U6193 (N_6193,N_5965,N_6001);
nor U6194 (N_6194,N_5951,N_5943);
xor U6195 (N_6195,N_5977,N_6057);
xnor U6196 (N_6196,N_5974,N_6076);
xor U6197 (N_6197,N_5966,N_6068);
or U6198 (N_6198,N_6056,N_6057);
xnor U6199 (N_6199,N_6070,N_6045);
xor U6200 (N_6200,N_5988,N_6034);
xor U6201 (N_6201,N_6002,N_6044);
nor U6202 (N_6202,N_6078,N_6000);
xor U6203 (N_6203,N_5990,N_6052);
or U6204 (N_6204,N_6005,N_6008);
nor U6205 (N_6205,N_6033,N_5938);
nor U6206 (N_6206,N_6022,N_6036);
or U6207 (N_6207,N_5957,N_6059);
nor U6208 (N_6208,N_5968,N_5943);
or U6209 (N_6209,N_5921,N_5988);
nand U6210 (N_6210,N_6057,N_5984);
and U6211 (N_6211,N_5946,N_5989);
xor U6212 (N_6212,N_6012,N_6009);
xor U6213 (N_6213,N_5988,N_5942);
nor U6214 (N_6214,N_6078,N_5998);
xor U6215 (N_6215,N_5937,N_5926);
and U6216 (N_6216,N_6042,N_5978);
xnor U6217 (N_6217,N_5933,N_5947);
or U6218 (N_6218,N_6034,N_6037);
or U6219 (N_6219,N_6025,N_6075);
xnor U6220 (N_6220,N_6056,N_6065);
xor U6221 (N_6221,N_6050,N_6051);
xor U6222 (N_6222,N_6003,N_6059);
xor U6223 (N_6223,N_6035,N_5999);
xor U6224 (N_6224,N_5951,N_5993);
nor U6225 (N_6225,N_6029,N_6035);
and U6226 (N_6226,N_5935,N_6046);
nor U6227 (N_6227,N_6025,N_5949);
nand U6228 (N_6228,N_5961,N_6074);
or U6229 (N_6229,N_6072,N_6029);
or U6230 (N_6230,N_6000,N_5986);
nand U6231 (N_6231,N_6072,N_6073);
or U6232 (N_6232,N_5974,N_5960);
and U6233 (N_6233,N_5981,N_5974);
xor U6234 (N_6234,N_5931,N_6071);
or U6235 (N_6235,N_5988,N_5948);
nor U6236 (N_6236,N_5987,N_5958);
nor U6237 (N_6237,N_6017,N_6007);
nand U6238 (N_6238,N_6009,N_6062);
nor U6239 (N_6239,N_5993,N_6068);
xnor U6240 (N_6240,N_6210,N_6126);
xor U6241 (N_6241,N_6208,N_6175);
and U6242 (N_6242,N_6147,N_6109);
nand U6243 (N_6243,N_6094,N_6127);
nor U6244 (N_6244,N_6099,N_6106);
or U6245 (N_6245,N_6098,N_6167);
xnor U6246 (N_6246,N_6237,N_6169);
and U6247 (N_6247,N_6151,N_6107);
xnor U6248 (N_6248,N_6146,N_6081);
xnor U6249 (N_6249,N_6159,N_6201);
nor U6250 (N_6250,N_6233,N_6093);
and U6251 (N_6251,N_6102,N_6224);
xnor U6252 (N_6252,N_6083,N_6212);
or U6253 (N_6253,N_6223,N_6164);
and U6254 (N_6254,N_6217,N_6178);
nand U6255 (N_6255,N_6089,N_6085);
xnor U6256 (N_6256,N_6134,N_6228);
or U6257 (N_6257,N_6189,N_6165);
and U6258 (N_6258,N_6173,N_6234);
and U6259 (N_6259,N_6227,N_6225);
or U6260 (N_6260,N_6101,N_6222);
or U6261 (N_6261,N_6205,N_6095);
nor U6262 (N_6262,N_6176,N_6158);
xor U6263 (N_6263,N_6172,N_6145);
and U6264 (N_6264,N_6181,N_6232);
or U6265 (N_6265,N_6141,N_6136);
or U6266 (N_6266,N_6207,N_6115);
or U6267 (N_6267,N_6137,N_6100);
and U6268 (N_6268,N_6143,N_6196);
nand U6269 (N_6269,N_6156,N_6177);
xor U6270 (N_6270,N_6215,N_6160);
nor U6271 (N_6271,N_6213,N_6219);
nand U6272 (N_6272,N_6186,N_6125);
xnor U6273 (N_6273,N_6216,N_6214);
nor U6274 (N_6274,N_6180,N_6088);
nor U6275 (N_6275,N_6087,N_6197);
xnor U6276 (N_6276,N_6149,N_6105);
xnor U6277 (N_6277,N_6209,N_6163);
nand U6278 (N_6278,N_6211,N_6168);
nor U6279 (N_6279,N_6191,N_6230);
or U6280 (N_6280,N_6157,N_6132);
nand U6281 (N_6281,N_6231,N_6121);
xor U6282 (N_6282,N_6184,N_6204);
or U6283 (N_6283,N_6142,N_6119);
nor U6284 (N_6284,N_6171,N_6080);
or U6285 (N_6285,N_6140,N_6161);
and U6286 (N_6286,N_6104,N_6182);
nor U6287 (N_6287,N_6229,N_6198);
nand U6288 (N_6288,N_6116,N_6091);
nand U6289 (N_6289,N_6084,N_6133);
nor U6290 (N_6290,N_6185,N_6202);
xor U6291 (N_6291,N_6097,N_6110);
nand U6292 (N_6292,N_6113,N_6226);
nand U6293 (N_6293,N_6192,N_6111);
xnor U6294 (N_6294,N_6179,N_6131);
xnor U6295 (N_6295,N_6096,N_6183);
nand U6296 (N_6296,N_6092,N_6139);
nand U6297 (N_6297,N_6162,N_6155);
xor U6298 (N_6298,N_6239,N_6129);
xnor U6299 (N_6299,N_6135,N_6236);
or U6300 (N_6300,N_6170,N_6148);
and U6301 (N_6301,N_6200,N_6190);
or U6302 (N_6302,N_6120,N_6118);
or U6303 (N_6303,N_6194,N_6154);
nand U6304 (N_6304,N_6130,N_6203);
nor U6305 (N_6305,N_6153,N_6090);
nand U6306 (N_6306,N_6124,N_6122);
and U6307 (N_6307,N_6174,N_6150);
nand U6308 (N_6308,N_6114,N_6117);
nand U6309 (N_6309,N_6199,N_6195);
and U6310 (N_6310,N_6166,N_6152);
nand U6311 (N_6311,N_6138,N_6112);
xnor U6312 (N_6312,N_6128,N_6238);
and U6313 (N_6313,N_6103,N_6193);
nand U6314 (N_6314,N_6221,N_6220);
or U6315 (N_6315,N_6206,N_6123);
and U6316 (N_6316,N_6108,N_6082);
nor U6317 (N_6317,N_6144,N_6086);
or U6318 (N_6318,N_6218,N_6188);
and U6319 (N_6319,N_6187,N_6235);
and U6320 (N_6320,N_6213,N_6092);
xor U6321 (N_6321,N_6237,N_6089);
nor U6322 (N_6322,N_6149,N_6089);
and U6323 (N_6323,N_6214,N_6179);
or U6324 (N_6324,N_6197,N_6130);
nor U6325 (N_6325,N_6220,N_6106);
nor U6326 (N_6326,N_6106,N_6154);
nand U6327 (N_6327,N_6105,N_6125);
xnor U6328 (N_6328,N_6122,N_6214);
nand U6329 (N_6329,N_6135,N_6202);
or U6330 (N_6330,N_6181,N_6096);
nor U6331 (N_6331,N_6205,N_6190);
or U6332 (N_6332,N_6131,N_6220);
or U6333 (N_6333,N_6150,N_6181);
or U6334 (N_6334,N_6130,N_6092);
and U6335 (N_6335,N_6144,N_6114);
xnor U6336 (N_6336,N_6139,N_6156);
or U6337 (N_6337,N_6129,N_6114);
nor U6338 (N_6338,N_6156,N_6197);
nand U6339 (N_6339,N_6082,N_6228);
and U6340 (N_6340,N_6112,N_6164);
and U6341 (N_6341,N_6163,N_6198);
nor U6342 (N_6342,N_6150,N_6136);
nor U6343 (N_6343,N_6182,N_6093);
and U6344 (N_6344,N_6203,N_6135);
nand U6345 (N_6345,N_6173,N_6124);
and U6346 (N_6346,N_6185,N_6229);
nand U6347 (N_6347,N_6239,N_6089);
xor U6348 (N_6348,N_6198,N_6231);
nor U6349 (N_6349,N_6229,N_6178);
nand U6350 (N_6350,N_6176,N_6109);
and U6351 (N_6351,N_6098,N_6144);
nor U6352 (N_6352,N_6085,N_6127);
xnor U6353 (N_6353,N_6105,N_6204);
xnor U6354 (N_6354,N_6190,N_6203);
xnor U6355 (N_6355,N_6196,N_6133);
nand U6356 (N_6356,N_6233,N_6202);
and U6357 (N_6357,N_6178,N_6113);
nor U6358 (N_6358,N_6147,N_6228);
nor U6359 (N_6359,N_6146,N_6205);
nor U6360 (N_6360,N_6235,N_6090);
nor U6361 (N_6361,N_6187,N_6101);
and U6362 (N_6362,N_6205,N_6158);
and U6363 (N_6363,N_6095,N_6206);
xnor U6364 (N_6364,N_6138,N_6123);
nand U6365 (N_6365,N_6151,N_6204);
or U6366 (N_6366,N_6170,N_6142);
nor U6367 (N_6367,N_6129,N_6122);
nor U6368 (N_6368,N_6142,N_6183);
nor U6369 (N_6369,N_6237,N_6132);
and U6370 (N_6370,N_6202,N_6096);
or U6371 (N_6371,N_6112,N_6149);
nand U6372 (N_6372,N_6107,N_6086);
or U6373 (N_6373,N_6154,N_6207);
nor U6374 (N_6374,N_6141,N_6119);
and U6375 (N_6375,N_6208,N_6108);
or U6376 (N_6376,N_6190,N_6166);
and U6377 (N_6377,N_6099,N_6113);
and U6378 (N_6378,N_6148,N_6230);
or U6379 (N_6379,N_6139,N_6089);
or U6380 (N_6380,N_6223,N_6092);
and U6381 (N_6381,N_6198,N_6183);
nand U6382 (N_6382,N_6082,N_6105);
nor U6383 (N_6383,N_6148,N_6141);
nand U6384 (N_6384,N_6091,N_6237);
or U6385 (N_6385,N_6132,N_6130);
nor U6386 (N_6386,N_6141,N_6113);
nor U6387 (N_6387,N_6172,N_6221);
nor U6388 (N_6388,N_6101,N_6231);
and U6389 (N_6389,N_6110,N_6198);
and U6390 (N_6390,N_6105,N_6227);
nor U6391 (N_6391,N_6190,N_6215);
and U6392 (N_6392,N_6184,N_6121);
nand U6393 (N_6393,N_6238,N_6151);
nor U6394 (N_6394,N_6115,N_6131);
xnor U6395 (N_6395,N_6183,N_6103);
xor U6396 (N_6396,N_6160,N_6122);
nand U6397 (N_6397,N_6093,N_6159);
nand U6398 (N_6398,N_6147,N_6169);
nand U6399 (N_6399,N_6221,N_6127);
nand U6400 (N_6400,N_6372,N_6308);
and U6401 (N_6401,N_6314,N_6359);
nand U6402 (N_6402,N_6325,N_6381);
and U6403 (N_6403,N_6358,N_6387);
nor U6404 (N_6404,N_6273,N_6365);
xor U6405 (N_6405,N_6317,N_6328);
nand U6406 (N_6406,N_6349,N_6374);
xnor U6407 (N_6407,N_6303,N_6310);
nor U6408 (N_6408,N_6351,N_6391);
and U6409 (N_6409,N_6393,N_6276);
nand U6410 (N_6410,N_6345,N_6338);
or U6411 (N_6411,N_6360,N_6278);
nor U6412 (N_6412,N_6315,N_6257);
and U6413 (N_6413,N_6293,N_6289);
xnor U6414 (N_6414,N_6266,N_6335);
xnor U6415 (N_6415,N_6282,N_6302);
xor U6416 (N_6416,N_6371,N_6390);
nand U6417 (N_6417,N_6250,N_6294);
and U6418 (N_6418,N_6340,N_6313);
nand U6419 (N_6419,N_6274,N_6320);
and U6420 (N_6420,N_6290,N_6251);
xnor U6421 (N_6421,N_6368,N_6243);
xor U6422 (N_6422,N_6279,N_6388);
and U6423 (N_6423,N_6255,N_6307);
or U6424 (N_6424,N_6253,N_6326);
and U6425 (N_6425,N_6248,N_6322);
and U6426 (N_6426,N_6378,N_6382);
nor U6427 (N_6427,N_6342,N_6264);
nand U6428 (N_6428,N_6327,N_6354);
or U6429 (N_6429,N_6269,N_6263);
xnor U6430 (N_6430,N_6336,N_6272);
nand U6431 (N_6431,N_6298,N_6394);
and U6432 (N_6432,N_6300,N_6398);
or U6433 (N_6433,N_6375,N_6286);
and U6434 (N_6434,N_6357,N_6348);
nor U6435 (N_6435,N_6346,N_6275);
nand U6436 (N_6436,N_6260,N_6284);
or U6437 (N_6437,N_6301,N_6287);
or U6438 (N_6438,N_6363,N_6249);
nor U6439 (N_6439,N_6285,N_6309);
or U6440 (N_6440,N_6395,N_6270);
xor U6441 (N_6441,N_6323,N_6373);
nand U6442 (N_6442,N_6283,N_6267);
or U6443 (N_6443,N_6361,N_6386);
xnor U6444 (N_6444,N_6252,N_6277);
and U6445 (N_6445,N_6246,N_6389);
nor U6446 (N_6446,N_6364,N_6305);
xor U6447 (N_6447,N_6377,N_6383);
nand U6448 (N_6448,N_6330,N_6356);
xnor U6449 (N_6449,N_6385,N_6296);
or U6450 (N_6450,N_6353,N_6280);
nand U6451 (N_6451,N_6343,N_6380);
nand U6452 (N_6452,N_6316,N_6240);
or U6453 (N_6453,N_6319,N_6344);
xor U6454 (N_6454,N_6258,N_6331);
and U6455 (N_6455,N_6242,N_6247);
or U6456 (N_6456,N_6256,N_6369);
xnor U6457 (N_6457,N_6265,N_6392);
and U6458 (N_6458,N_6367,N_6376);
nand U6459 (N_6459,N_6355,N_6321);
and U6460 (N_6460,N_6350,N_6396);
or U6461 (N_6461,N_6352,N_6288);
and U6462 (N_6462,N_6312,N_6370);
xnor U6463 (N_6463,N_6366,N_6318);
and U6464 (N_6464,N_6241,N_6268);
or U6465 (N_6465,N_6304,N_6362);
and U6466 (N_6466,N_6329,N_6297);
and U6467 (N_6467,N_6337,N_6332);
nand U6468 (N_6468,N_6399,N_6262);
nand U6469 (N_6469,N_6244,N_6299);
xnor U6470 (N_6470,N_6306,N_6311);
and U6471 (N_6471,N_6281,N_6339);
nand U6472 (N_6472,N_6334,N_6291);
or U6473 (N_6473,N_6254,N_6261);
and U6474 (N_6474,N_6397,N_6245);
or U6475 (N_6475,N_6324,N_6379);
nor U6476 (N_6476,N_6341,N_6347);
or U6477 (N_6477,N_6292,N_6333);
nand U6478 (N_6478,N_6259,N_6271);
or U6479 (N_6479,N_6295,N_6384);
xnor U6480 (N_6480,N_6319,N_6360);
nor U6481 (N_6481,N_6323,N_6254);
and U6482 (N_6482,N_6269,N_6284);
nand U6483 (N_6483,N_6306,N_6249);
nand U6484 (N_6484,N_6337,N_6318);
xor U6485 (N_6485,N_6384,N_6385);
or U6486 (N_6486,N_6318,N_6298);
nor U6487 (N_6487,N_6305,N_6399);
or U6488 (N_6488,N_6256,N_6336);
nand U6489 (N_6489,N_6255,N_6293);
nor U6490 (N_6490,N_6348,N_6389);
nor U6491 (N_6491,N_6377,N_6352);
nor U6492 (N_6492,N_6382,N_6374);
xnor U6493 (N_6493,N_6260,N_6392);
and U6494 (N_6494,N_6393,N_6269);
nand U6495 (N_6495,N_6292,N_6341);
or U6496 (N_6496,N_6392,N_6247);
or U6497 (N_6497,N_6260,N_6305);
and U6498 (N_6498,N_6380,N_6317);
and U6499 (N_6499,N_6265,N_6290);
nor U6500 (N_6500,N_6284,N_6279);
and U6501 (N_6501,N_6272,N_6365);
and U6502 (N_6502,N_6250,N_6352);
and U6503 (N_6503,N_6245,N_6313);
and U6504 (N_6504,N_6254,N_6342);
nand U6505 (N_6505,N_6346,N_6298);
nand U6506 (N_6506,N_6373,N_6354);
nand U6507 (N_6507,N_6242,N_6262);
and U6508 (N_6508,N_6338,N_6365);
xor U6509 (N_6509,N_6294,N_6319);
or U6510 (N_6510,N_6263,N_6339);
nand U6511 (N_6511,N_6244,N_6329);
and U6512 (N_6512,N_6326,N_6241);
nand U6513 (N_6513,N_6379,N_6322);
and U6514 (N_6514,N_6298,N_6383);
xnor U6515 (N_6515,N_6345,N_6382);
xnor U6516 (N_6516,N_6313,N_6376);
nand U6517 (N_6517,N_6318,N_6273);
nor U6518 (N_6518,N_6305,N_6255);
and U6519 (N_6519,N_6360,N_6258);
or U6520 (N_6520,N_6286,N_6319);
nor U6521 (N_6521,N_6286,N_6267);
xnor U6522 (N_6522,N_6264,N_6294);
nand U6523 (N_6523,N_6358,N_6309);
xor U6524 (N_6524,N_6315,N_6246);
nor U6525 (N_6525,N_6364,N_6324);
xor U6526 (N_6526,N_6335,N_6241);
nand U6527 (N_6527,N_6334,N_6352);
nor U6528 (N_6528,N_6327,N_6328);
nand U6529 (N_6529,N_6377,N_6307);
and U6530 (N_6530,N_6337,N_6276);
or U6531 (N_6531,N_6253,N_6241);
nor U6532 (N_6532,N_6396,N_6392);
nor U6533 (N_6533,N_6287,N_6330);
and U6534 (N_6534,N_6284,N_6320);
or U6535 (N_6535,N_6326,N_6243);
xor U6536 (N_6536,N_6300,N_6342);
and U6537 (N_6537,N_6271,N_6322);
nand U6538 (N_6538,N_6399,N_6353);
and U6539 (N_6539,N_6387,N_6328);
and U6540 (N_6540,N_6306,N_6284);
and U6541 (N_6541,N_6321,N_6372);
or U6542 (N_6542,N_6366,N_6306);
nand U6543 (N_6543,N_6244,N_6258);
or U6544 (N_6544,N_6388,N_6289);
or U6545 (N_6545,N_6292,N_6346);
or U6546 (N_6546,N_6253,N_6245);
or U6547 (N_6547,N_6389,N_6378);
nor U6548 (N_6548,N_6288,N_6389);
or U6549 (N_6549,N_6380,N_6361);
or U6550 (N_6550,N_6279,N_6293);
nor U6551 (N_6551,N_6378,N_6339);
and U6552 (N_6552,N_6355,N_6250);
and U6553 (N_6553,N_6343,N_6327);
xnor U6554 (N_6554,N_6343,N_6260);
nand U6555 (N_6555,N_6397,N_6313);
and U6556 (N_6556,N_6316,N_6394);
and U6557 (N_6557,N_6296,N_6321);
nor U6558 (N_6558,N_6246,N_6337);
or U6559 (N_6559,N_6398,N_6297);
nand U6560 (N_6560,N_6424,N_6436);
nand U6561 (N_6561,N_6420,N_6421);
or U6562 (N_6562,N_6509,N_6423);
nor U6563 (N_6563,N_6512,N_6522);
nand U6564 (N_6564,N_6524,N_6534);
or U6565 (N_6565,N_6413,N_6495);
xnor U6566 (N_6566,N_6503,N_6549);
nand U6567 (N_6567,N_6441,N_6546);
nand U6568 (N_6568,N_6466,N_6543);
or U6569 (N_6569,N_6510,N_6540);
xnor U6570 (N_6570,N_6471,N_6453);
xnor U6571 (N_6571,N_6541,N_6462);
nand U6572 (N_6572,N_6508,N_6532);
and U6573 (N_6573,N_6446,N_6444);
xor U6574 (N_6574,N_6487,N_6435);
nand U6575 (N_6575,N_6499,N_6493);
or U6576 (N_6576,N_6430,N_6422);
nor U6577 (N_6577,N_6504,N_6431);
or U6578 (N_6578,N_6529,N_6555);
xnor U6579 (N_6579,N_6502,N_6456);
and U6580 (N_6580,N_6438,N_6498);
nor U6581 (N_6581,N_6440,N_6463);
nand U6582 (N_6582,N_6514,N_6511);
xnor U6583 (N_6583,N_6536,N_6559);
and U6584 (N_6584,N_6449,N_6507);
or U6585 (N_6585,N_6409,N_6486);
nand U6586 (N_6586,N_6458,N_6552);
nand U6587 (N_6587,N_6478,N_6537);
xor U6588 (N_6588,N_6544,N_6517);
nand U6589 (N_6589,N_6433,N_6400);
xnor U6590 (N_6590,N_6448,N_6489);
nand U6591 (N_6591,N_6501,N_6407);
nand U6592 (N_6592,N_6469,N_6452);
nor U6593 (N_6593,N_6538,N_6410);
nor U6594 (N_6594,N_6521,N_6465);
xor U6595 (N_6595,N_6557,N_6434);
nor U6596 (N_6596,N_6506,N_6548);
nor U6597 (N_6597,N_6530,N_6417);
nor U6598 (N_6598,N_6484,N_6526);
xor U6599 (N_6599,N_6445,N_6450);
or U6600 (N_6600,N_6490,N_6439);
nor U6601 (N_6601,N_6472,N_6419);
and U6602 (N_6602,N_6447,N_6513);
xor U6603 (N_6603,N_6406,N_6527);
and U6604 (N_6604,N_6418,N_6554);
and U6605 (N_6605,N_6467,N_6468);
xnor U6606 (N_6606,N_6459,N_6432);
or U6607 (N_6607,N_6525,N_6412);
nor U6608 (N_6608,N_6428,N_6500);
nand U6609 (N_6609,N_6482,N_6437);
xor U6610 (N_6610,N_6528,N_6483);
or U6611 (N_6611,N_6451,N_6551);
or U6612 (N_6612,N_6411,N_6556);
xor U6613 (N_6613,N_6455,N_6405);
nor U6614 (N_6614,N_6558,N_6416);
and U6615 (N_6615,N_6516,N_6518);
nand U6616 (N_6616,N_6425,N_6520);
nand U6617 (N_6617,N_6550,N_6539);
nand U6618 (N_6618,N_6408,N_6401);
nand U6619 (N_6619,N_6473,N_6429);
and U6620 (N_6620,N_6547,N_6491);
xnor U6621 (N_6621,N_6454,N_6404);
nand U6622 (N_6622,N_6496,N_6485);
nand U6623 (N_6623,N_6403,N_6531);
and U6624 (N_6624,N_6494,N_6480);
and U6625 (N_6625,N_6505,N_6460);
nand U6626 (N_6626,N_6545,N_6481);
xor U6627 (N_6627,N_6535,N_6492);
nor U6628 (N_6628,N_6479,N_6477);
and U6629 (N_6629,N_6553,N_6427);
xor U6630 (N_6630,N_6497,N_6523);
xnor U6631 (N_6631,N_6470,N_6402);
nand U6632 (N_6632,N_6542,N_6533);
xnor U6633 (N_6633,N_6415,N_6426);
and U6634 (N_6634,N_6475,N_6443);
or U6635 (N_6635,N_6414,N_6474);
nor U6636 (N_6636,N_6519,N_6488);
or U6637 (N_6637,N_6515,N_6442);
nor U6638 (N_6638,N_6457,N_6461);
xnor U6639 (N_6639,N_6464,N_6476);
and U6640 (N_6640,N_6527,N_6517);
nor U6641 (N_6641,N_6532,N_6446);
and U6642 (N_6642,N_6444,N_6519);
nor U6643 (N_6643,N_6554,N_6479);
nand U6644 (N_6644,N_6472,N_6525);
xor U6645 (N_6645,N_6484,N_6444);
xnor U6646 (N_6646,N_6416,N_6490);
nor U6647 (N_6647,N_6401,N_6426);
nor U6648 (N_6648,N_6401,N_6533);
or U6649 (N_6649,N_6477,N_6461);
nor U6650 (N_6650,N_6405,N_6555);
nor U6651 (N_6651,N_6542,N_6401);
or U6652 (N_6652,N_6447,N_6486);
nand U6653 (N_6653,N_6507,N_6527);
nor U6654 (N_6654,N_6553,N_6519);
nand U6655 (N_6655,N_6419,N_6412);
nand U6656 (N_6656,N_6476,N_6510);
or U6657 (N_6657,N_6441,N_6421);
nand U6658 (N_6658,N_6456,N_6513);
or U6659 (N_6659,N_6484,N_6476);
xnor U6660 (N_6660,N_6462,N_6488);
nor U6661 (N_6661,N_6475,N_6430);
nor U6662 (N_6662,N_6523,N_6457);
nand U6663 (N_6663,N_6553,N_6415);
and U6664 (N_6664,N_6420,N_6440);
or U6665 (N_6665,N_6431,N_6490);
nand U6666 (N_6666,N_6471,N_6493);
nor U6667 (N_6667,N_6473,N_6443);
or U6668 (N_6668,N_6413,N_6435);
and U6669 (N_6669,N_6469,N_6504);
or U6670 (N_6670,N_6535,N_6540);
xor U6671 (N_6671,N_6428,N_6457);
or U6672 (N_6672,N_6415,N_6465);
nor U6673 (N_6673,N_6526,N_6530);
and U6674 (N_6674,N_6401,N_6512);
or U6675 (N_6675,N_6456,N_6444);
nand U6676 (N_6676,N_6501,N_6465);
xor U6677 (N_6677,N_6413,N_6465);
nand U6678 (N_6678,N_6409,N_6437);
or U6679 (N_6679,N_6441,N_6519);
or U6680 (N_6680,N_6427,N_6483);
or U6681 (N_6681,N_6445,N_6409);
and U6682 (N_6682,N_6451,N_6549);
nor U6683 (N_6683,N_6546,N_6472);
xnor U6684 (N_6684,N_6442,N_6525);
and U6685 (N_6685,N_6422,N_6556);
or U6686 (N_6686,N_6452,N_6533);
and U6687 (N_6687,N_6549,N_6433);
nor U6688 (N_6688,N_6470,N_6550);
and U6689 (N_6689,N_6558,N_6443);
xnor U6690 (N_6690,N_6428,N_6481);
nor U6691 (N_6691,N_6424,N_6461);
nor U6692 (N_6692,N_6496,N_6526);
nor U6693 (N_6693,N_6471,N_6444);
nor U6694 (N_6694,N_6553,N_6490);
xor U6695 (N_6695,N_6487,N_6431);
and U6696 (N_6696,N_6538,N_6476);
and U6697 (N_6697,N_6419,N_6445);
nor U6698 (N_6698,N_6498,N_6474);
nand U6699 (N_6699,N_6499,N_6531);
nand U6700 (N_6700,N_6489,N_6422);
nand U6701 (N_6701,N_6441,N_6415);
and U6702 (N_6702,N_6532,N_6501);
and U6703 (N_6703,N_6470,N_6545);
xnor U6704 (N_6704,N_6487,N_6475);
and U6705 (N_6705,N_6515,N_6406);
nor U6706 (N_6706,N_6421,N_6424);
nand U6707 (N_6707,N_6454,N_6501);
or U6708 (N_6708,N_6440,N_6449);
nor U6709 (N_6709,N_6458,N_6467);
xor U6710 (N_6710,N_6417,N_6534);
nand U6711 (N_6711,N_6524,N_6432);
nor U6712 (N_6712,N_6547,N_6400);
or U6713 (N_6713,N_6460,N_6535);
xnor U6714 (N_6714,N_6515,N_6549);
or U6715 (N_6715,N_6516,N_6489);
or U6716 (N_6716,N_6462,N_6540);
nand U6717 (N_6717,N_6495,N_6453);
and U6718 (N_6718,N_6540,N_6474);
xor U6719 (N_6719,N_6406,N_6537);
xor U6720 (N_6720,N_6587,N_6605);
xor U6721 (N_6721,N_6654,N_6652);
and U6722 (N_6722,N_6707,N_6585);
and U6723 (N_6723,N_6598,N_6630);
xor U6724 (N_6724,N_6627,N_6581);
xor U6725 (N_6725,N_6676,N_6665);
nand U6726 (N_6726,N_6583,N_6604);
nor U6727 (N_6727,N_6616,N_6575);
nand U6728 (N_6728,N_6567,N_6675);
xnor U6729 (N_6729,N_6693,N_6618);
nor U6730 (N_6730,N_6625,N_6696);
nor U6731 (N_6731,N_6715,N_6572);
nor U6732 (N_6732,N_6642,N_6634);
and U6733 (N_6733,N_6574,N_6568);
or U6734 (N_6734,N_6713,N_6641);
nand U6735 (N_6735,N_6719,N_6580);
or U6736 (N_6736,N_6635,N_6599);
nor U6737 (N_6737,N_6695,N_6670);
or U6738 (N_6738,N_6661,N_6698);
nand U6739 (N_6739,N_6680,N_6623);
xnor U6740 (N_6740,N_6666,N_6699);
or U6741 (N_6741,N_6660,N_6667);
nor U6742 (N_6742,N_6613,N_6651);
xnor U6743 (N_6743,N_6702,N_6658);
xnor U6744 (N_6744,N_6579,N_6628);
or U6745 (N_6745,N_6638,N_6656);
nor U6746 (N_6746,N_6590,N_6571);
nand U6747 (N_6747,N_6570,N_6632);
nor U6748 (N_6748,N_6690,N_6601);
xnor U6749 (N_6749,N_6593,N_6566);
nand U6750 (N_6750,N_6683,N_6672);
nor U6751 (N_6751,N_6592,N_6608);
or U6752 (N_6752,N_6561,N_6615);
or U6753 (N_6753,N_6602,N_6711);
and U6754 (N_6754,N_6688,N_6614);
nor U6755 (N_6755,N_6603,N_6562);
nand U6756 (N_6756,N_6644,N_6584);
nor U6757 (N_6757,N_6563,N_6617);
nand U6758 (N_6758,N_6659,N_6708);
or U6759 (N_6759,N_6578,N_6620);
nand U6760 (N_6760,N_6685,N_6712);
xor U6761 (N_6761,N_6689,N_6637);
nand U6762 (N_6762,N_6704,N_6653);
xor U6763 (N_6763,N_6678,N_6714);
and U6764 (N_6764,N_6677,N_6569);
or U6765 (N_6765,N_6709,N_6646);
or U6766 (N_6766,N_6669,N_6629);
xnor U6767 (N_6767,N_6591,N_6684);
nand U6768 (N_6768,N_6560,N_6600);
nor U6769 (N_6769,N_6686,N_6662);
or U6770 (N_6770,N_6703,N_6694);
nand U6771 (N_6771,N_6682,N_6650);
nor U6772 (N_6772,N_6582,N_6612);
or U6773 (N_6773,N_6564,N_6664);
xnor U6774 (N_6774,N_6687,N_6588);
xnor U6775 (N_6775,N_6595,N_6586);
nor U6776 (N_6776,N_6668,N_6597);
xnor U6777 (N_6777,N_6643,N_6639);
nor U6778 (N_6778,N_6717,N_6631);
nor U6779 (N_6779,N_6671,N_6673);
xor U6780 (N_6780,N_6594,N_6710);
xnor U6781 (N_6781,N_6606,N_6622);
and U6782 (N_6782,N_6648,N_6640);
xor U6783 (N_6783,N_6691,N_6573);
nor U6784 (N_6784,N_6577,N_6645);
nand U6785 (N_6785,N_6636,N_6607);
xnor U6786 (N_6786,N_6609,N_6611);
and U6787 (N_6787,N_6576,N_6565);
nor U6788 (N_6788,N_6705,N_6663);
nor U6789 (N_6789,N_6706,N_6624);
nor U6790 (N_6790,N_6657,N_6692);
and U6791 (N_6791,N_6619,N_6610);
xor U6792 (N_6792,N_6681,N_6718);
xor U6793 (N_6793,N_6679,N_6647);
and U6794 (N_6794,N_6596,N_6633);
xnor U6795 (N_6795,N_6697,N_6621);
or U6796 (N_6796,N_6649,N_6716);
nor U6797 (N_6797,N_6589,N_6655);
nor U6798 (N_6798,N_6700,N_6701);
nor U6799 (N_6799,N_6626,N_6674);
and U6800 (N_6800,N_6564,N_6689);
nand U6801 (N_6801,N_6619,N_6631);
xnor U6802 (N_6802,N_6591,N_6614);
and U6803 (N_6803,N_6689,N_6571);
nor U6804 (N_6804,N_6632,N_6670);
xor U6805 (N_6805,N_6652,N_6653);
and U6806 (N_6806,N_6608,N_6625);
xor U6807 (N_6807,N_6584,N_6674);
nand U6808 (N_6808,N_6684,N_6564);
xor U6809 (N_6809,N_6568,N_6634);
and U6810 (N_6810,N_6704,N_6588);
nor U6811 (N_6811,N_6604,N_6582);
and U6812 (N_6812,N_6714,N_6595);
nor U6813 (N_6813,N_6617,N_6657);
nor U6814 (N_6814,N_6613,N_6621);
nand U6815 (N_6815,N_6674,N_6573);
xnor U6816 (N_6816,N_6625,N_6648);
or U6817 (N_6817,N_6648,N_6611);
nor U6818 (N_6818,N_6605,N_6630);
and U6819 (N_6819,N_6639,N_6700);
or U6820 (N_6820,N_6667,N_6614);
or U6821 (N_6821,N_6626,N_6630);
or U6822 (N_6822,N_6713,N_6665);
xnor U6823 (N_6823,N_6675,N_6615);
or U6824 (N_6824,N_6561,N_6592);
and U6825 (N_6825,N_6695,N_6621);
nor U6826 (N_6826,N_6708,N_6663);
nand U6827 (N_6827,N_6605,N_6676);
and U6828 (N_6828,N_6618,N_6591);
nor U6829 (N_6829,N_6573,N_6711);
or U6830 (N_6830,N_6571,N_6592);
or U6831 (N_6831,N_6699,N_6689);
and U6832 (N_6832,N_6619,N_6672);
or U6833 (N_6833,N_6684,N_6656);
or U6834 (N_6834,N_6659,N_6686);
nor U6835 (N_6835,N_6567,N_6658);
nor U6836 (N_6836,N_6596,N_6688);
and U6837 (N_6837,N_6578,N_6629);
or U6838 (N_6838,N_6703,N_6679);
and U6839 (N_6839,N_6613,N_6682);
nand U6840 (N_6840,N_6621,N_6704);
xnor U6841 (N_6841,N_6707,N_6567);
nand U6842 (N_6842,N_6619,N_6591);
nor U6843 (N_6843,N_6652,N_6590);
nand U6844 (N_6844,N_6665,N_6568);
nand U6845 (N_6845,N_6623,N_6638);
nand U6846 (N_6846,N_6649,N_6562);
nor U6847 (N_6847,N_6640,N_6639);
nor U6848 (N_6848,N_6631,N_6663);
or U6849 (N_6849,N_6588,N_6598);
nand U6850 (N_6850,N_6574,N_6702);
nand U6851 (N_6851,N_6642,N_6715);
nand U6852 (N_6852,N_6714,N_6591);
nor U6853 (N_6853,N_6709,N_6594);
and U6854 (N_6854,N_6703,N_6657);
nand U6855 (N_6855,N_6616,N_6612);
nor U6856 (N_6856,N_6579,N_6647);
or U6857 (N_6857,N_6649,N_6650);
nand U6858 (N_6858,N_6683,N_6688);
or U6859 (N_6859,N_6709,N_6624);
nand U6860 (N_6860,N_6704,N_6583);
nand U6861 (N_6861,N_6626,N_6663);
xor U6862 (N_6862,N_6702,N_6674);
and U6863 (N_6863,N_6655,N_6705);
xnor U6864 (N_6864,N_6632,N_6650);
xnor U6865 (N_6865,N_6605,N_6672);
nor U6866 (N_6866,N_6697,N_6691);
nand U6867 (N_6867,N_6561,N_6659);
nor U6868 (N_6868,N_6705,N_6648);
and U6869 (N_6869,N_6643,N_6624);
and U6870 (N_6870,N_6633,N_6614);
or U6871 (N_6871,N_6709,N_6569);
xor U6872 (N_6872,N_6621,N_6638);
nor U6873 (N_6873,N_6620,N_6599);
nor U6874 (N_6874,N_6702,N_6582);
nor U6875 (N_6875,N_6694,N_6587);
xor U6876 (N_6876,N_6667,N_6575);
or U6877 (N_6877,N_6589,N_6713);
and U6878 (N_6878,N_6635,N_6596);
xor U6879 (N_6879,N_6591,N_6710);
xor U6880 (N_6880,N_6812,N_6756);
xnor U6881 (N_6881,N_6854,N_6817);
and U6882 (N_6882,N_6748,N_6833);
and U6883 (N_6883,N_6722,N_6857);
or U6884 (N_6884,N_6770,N_6838);
xnor U6885 (N_6885,N_6777,N_6868);
or U6886 (N_6886,N_6768,N_6878);
nand U6887 (N_6887,N_6836,N_6736);
or U6888 (N_6888,N_6793,N_6775);
or U6889 (N_6889,N_6729,N_6753);
nor U6890 (N_6890,N_6747,N_6734);
xnor U6891 (N_6891,N_6835,N_6763);
nand U6892 (N_6892,N_6761,N_6843);
nor U6893 (N_6893,N_6735,N_6738);
nor U6894 (N_6894,N_6855,N_6828);
nor U6895 (N_6895,N_6787,N_6725);
xnor U6896 (N_6896,N_6877,N_6803);
nand U6897 (N_6897,N_6873,N_6824);
and U6898 (N_6898,N_6826,N_6851);
and U6899 (N_6899,N_6732,N_6808);
or U6900 (N_6900,N_6743,N_6823);
nor U6901 (N_6901,N_6807,N_6755);
or U6902 (N_6902,N_6754,N_6795);
or U6903 (N_6903,N_6765,N_6879);
nor U6904 (N_6904,N_6829,N_6850);
nand U6905 (N_6905,N_6794,N_6760);
nor U6906 (N_6906,N_6790,N_6841);
xor U6907 (N_6907,N_6783,N_6848);
xnor U6908 (N_6908,N_6757,N_6809);
nand U6909 (N_6909,N_6852,N_6774);
nand U6910 (N_6910,N_6860,N_6840);
and U6911 (N_6911,N_6786,N_6742);
xor U6912 (N_6912,N_6834,N_6832);
xnor U6913 (N_6913,N_6849,N_6781);
or U6914 (N_6914,N_6721,N_6731);
xnor U6915 (N_6915,N_6723,N_6737);
xnor U6916 (N_6916,N_6820,N_6875);
or U6917 (N_6917,N_6728,N_6865);
and U6918 (N_6918,N_6788,N_6845);
nand U6919 (N_6919,N_6806,N_6853);
or U6920 (N_6920,N_6750,N_6802);
or U6921 (N_6921,N_6741,N_6856);
nor U6922 (N_6922,N_6720,N_6846);
nand U6923 (N_6923,N_6815,N_6782);
and U6924 (N_6924,N_6827,N_6785);
nand U6925 (N_6925,N_6825,N_6800);
or U6926 (N_6926,N_6844,N_6767);
or U6927 (N_6927,N_6811,N_6810);
nand U6928 (N_6928,N_6780,N_6749);
or U6929 (N_6929,N_6822,N_6769);
nand U6930 (N_6930,N_6759,N_6789);
or U6931 (N_6931,N_6821,N_6746);
or U6932 (N_6932,N_6819,N_6816);
nor U6933 (N_6933,N_6814,N_6863);
or U6934 (N_6934,N_6799,N_6733);
and U6935 (N_6935,N_6758,N_6870);
or U6936 (N_6936,N_6764,N_6798);
xnor U6937 (N_6937,N_6779,N_6830);
xor U6938 (N_6938,N_6724,N_6797);
nand U6939 (N_6939,N_6778,N_6867);
or U6940 (N_6940,N_6858,N_6771);
or U6941 (N_6941,N_6871,N_6869);
nand U6942 (N_6942,N_6876,N_6859);
nand U6943 (N_6943,N_6813,N_6773);
nand U6944 (N_6944,N_6792,N_6791);
or U6945 (N_6945,N_6776,N_6762);
nand U6946 (N_6946,N_6784,N_6739);
nand U6947 (N_6947,N_6864,N_6751);
nor U6948 (N_6948,N_6740,N_6831);
and U6949 (N_6949,N_6842,N_6744);
nand U6950 (N_6950,N_6837,N_6874);
and U6951 (N_6951,N_6796,N_6766);
nand U6952 (N_6952,N_6839,N_6862);
xnor U6953 (N_6953,N_6861,N_6745);
and U6954 (N_6954,N_6818,N_6801);
xor U6955 (N_6955,N_6772,N_6805);
nor U6956 (N_6956,N_6752,N_6872);
nor U6957 (N_6957,N_6730,N_6804);
xnor U6958 (N_6958,N_6727,N_6847);
nand U6959 (N_6959,N_6866,N_6726);
and U6960 (N_6960,N_6832,N_6767);
xor U6961 (N_6961,N_6770,N_6763);
or U6962 (N_6962,N_6787,N_6752);
or U6963 (N_6963,N_6741,N_6770);
xnor U6964 (N_6964,N_6741,N_6758);
nand U6965 (N_6965,N_6758,N_6856);
nand U6966 (N_6966,N_6797,N_6740);
nor U6967 (N_6967,N_6804,N_6824);
and U6968 (N_6968,N_6823,N_6795);
and U6969 (N_6969,N_6770,N_6798);
or U6970 (N_6970,N_6829,N_6799);
nand U6971 (N_6971,N_6874,N_6722);
nor U6972 (N_6972,N_6726,N_6777);
xor U6973 (N_6973,N_6839,N_6845);
xnor U6974 (N_6974,N_6721,N_6733);
nand U6975 (N_6975,N_6767,N_6864);
xnor U6976 (N_6976,N_6724,N_6804);
and U6977 (N_6977,N_6867,N_6855);
nand U6978 (N_6978,N_6781,N_6744);
xor U6979 (N_6979,N_6752,N_6859);
nor U6980 (N_6980,N_6741,N_6752);
xnor U6981 (N_6981,N_6766,N_6849);
nor U6982 (N_6982,N_6824,N_6844);
or U6983 (N_6983,N_6856,N_6733);
nand U6984 (N_6984,N_6828,N_6772);
or U6985 (N_6985,N_6791,N_6813);
nand U6986 (N_6986,N_6771,N_6751);
nor U6987 (N_6987,N_6797,N_6766);
or U6988 (N_6988,N_6736,N_6870);
nor U6989 (N_6989,N_6758,N_6860);
nand U6990 (N_6990,N_6747,N_6735);
and U6991 (N_6991,N_6732,N_6816);
nor U6992 (N_6992,N_6735,N_6749);
nor U6993 (N_6993,N_6760,N_6736);
nand U6994 (N_6994,N_6854,N_6729);
or U6995 (N_6995,N_6745,N_6777);
and U6996 (N_6996,N_6764,N_6859);
and U6997 (N_6997,N_6847,N_6749);
and U6998 (N_6998,N_6794,N_6797);
xor U6999 (N_6999,N_6822,N_6786);
or U7000 (N_7000,N_6784,N_6793);
nor U7001 (N_7001,N_6858,N_6853);
xnor U7002 (N_7002,N_6838,N_6841);
and U7003 (N_7003,N_6803,N_6819);
nor U7004 (N_7004,N_6756,N_6833);
xor U7005 (N_7005,N_6808,N_6813);
and U7006 (N_7006,N_6865,N_6721);
and U7007 (N_7007,N_6765,N_6814);
nor U7008 (N_7008,N_6871,N_6737);
nand U7009 (N_7009,N_6747,N_6869);
xor U7010 (N_7010,N_6802,N_6843);
nor U7011 (N_7011,N_6727,N_6743);
xor U7012 (N_7012,N_6769,N_6780);
and U7013 (N_7013,N_6845,N_6841);
or U7014 (N_7014,N_6829,N_6746);
nand U7015 (N_7015,N_6876,N_6825);
nand U7016 (N_7016,N_6803,N_6757);
nor U7017 (N_7017,N_6826,N_6794);
nor U7018 (N_7018,N_6782,N_6740);
and U7019 (N_7019,N_6866,N_6827);
xor U7020 (N_7020,N_6847,N_6779);
nand U7021 (N_7021,N_6852,N_6810);
or U7022 (N_7022,N_6797,N_6755);
nand U7023 (N_7023,N_6832,N_6789);
nand U7024 (N_7024,N_6735,N_6755);
nor U7025 (N_7025,N_6804,N_6720);
xnor U7026 (N_7026,N_6818,N_6837);
xnor U7027 (N_7027,N_6871,N_6870);
or U7028 (N_7028,N_6822,N_6809);
and U7029 (N_7029,N_6732,N_6840);
xor U7030 (N_7030,N_6733,N_6845);
and U7031 (N_7031,N_6786,N_6813);
or U7032 (N_7032,N_6757,N_6832);
xnor U7033 (N_7033,N_6790,N_6741);
or U7034 (N_7034,N_6771,N_6865);
and U7035 (N_7035,N_6868,N_6736);
or U7036 (N_7036,N_6732,N_6772);
and U7037 (N_7037,N_6803,N_6728);
xor U7038 (N_7038,N_6859,N_6821);
xor U7039 (N_7039,N_6796,N_6801);
xor U7040 (N_7040,N_6984,N_6985);
xor U7041 (N_7041,N_6939,N_6941);
or U7042 (N_7042,N_6883,N_6956);
nand U7043 (N_7043,N_6909,N_7007);
and U7044 (N_7044,N_7006,N_6930);
nand U7045 (N_7045,N_6947,N_7009);
or U7046 (N_7046,N_7039,N_6949);
nand U7047 (N_7047,N_7038,N_6946);
or U7048 (N_7048,N_6994,N_6933);
nor U7049 (N_7049,N_6889,N_6921);
nand U7050 (N_7050,N_6961,N_6966);
or U7051 (N_7051,N_6928,N_6960);
nand U7052 (N_7052,N_6977,N_6901);
and U7053 (N_7053,N_6971,N_6979);
nand U7054 (N_7054,N_7024,N_6951);
xnor U7055 (N_7055,N_7031,N_6900);
nand U7056 (N_7056,N_6950,N_6888);
nor U7057 (N_7057,N_6915,N_7010);
xor U7058 (N_7058,N_6952,N_7028);
and U7059 (N_7059,N_6936,N_6998);
xnor U7060 (N_7060,N_6932,N_6982);
or U7061 (N_7061,N_7036,N_7027);
or U7062 (N_7062,N_6970,N_6990);
or U7063 (N_7063,N_6937,N_6974);
nand U7064 (N_7064,N_6934,N_7011);
xor U7065 (N_7065,N_6917,N_6954);
xnor U7066 (N_7066,N_6925,N_7015);
or U7067 (N_7067,N_6882,N_7021);
nor U7068 (N_7068,N_6938,N_6962);
or U7069 (N_7069,N_6926,N_6905);
and U7070 (N_7070,N_6992,N_6896);
and U7071 (N_7071,N_6927,N_6892);
nand U7072 (N_7072,N_7020,N_6986);
nor U7073 (N_7073,N_7029,N_6913);
or U7074 (N_7074,N_7004,N_6957);
and U7075 (N_7075,N_7016,N_6935);
or U7076 (N_7076,N_7005,N_6975);
or U7077 (N_7077,N_7035,N_6931);
nand U7078 (N_7078,N_6989,N_6923);
nor U7079 (N_7079,N_6967,N_7034);
or U7080 (N_7080,N_6953,N_6895);
or U7081 (N_7081,N_6916,N_6919);
nor U7082 (N_7082,N_7037,N_6884);
and U7083 (N_7083,N_6885,N_6991);
xnor U7084 (N_7084,N_7025,N_7003);
xor U7085 (N_7085,N_6891,N_6943);
nor U7086 (N_7086,N_6968,N_6983);
nand U7087 (N_7087,N_7014,N_6914);
xor U7088 (N_7088,N_6978,N_6940);
nand U7089 (N_7089,N_6886,N_6912);
nand U7090 (N_7090,N_6964,N_7000);
nor U7091 (N_7091,N_6997,N_7001);
and U7092 (N_7092,N_6944,N_7019);
nor U7093 (N_7093,N_6898,N_6887);
nor U7094 (N_7094,N_6881,N_6897);
nor U7095 (N_7095,N_6893,N_6920);
nor U7096 (N_7096,N_7018,N_6981);
xnor U7097 (N_7097,N_6948,N_6973);
xor U7098 (N_7098,N_6996,N_6894);
nand U7099 (N_7099,N_6999,N_7033);
nand U7100 (N_7100,N_6976,N_7012);
nand U7101 (N_7101,N_6910,N_6980);
xnor U7102 (N_7102,N_6958,N_6880);
and U7103 (N_7103,N_6906,N_7017);
or U7104 (N_7104,N_6945,N_6972);
and U7105 (N_7105,N_7022,N_6904);
and U7106 (N_7106,N_6929,N_6987);
xnor U7107 (N_7107,N_6903,N_7023);
and U7108 (N_7108,N_6995,N_7002);
or U7109 (N_7109,N_6988,N_6959);
or U7110 (N_7110,N_6907,N_7013);
nand U7111 (N_7111,N_6942,N_7008);
xor U7112 (N_7112,N_6963,N_6969);
xnor U7113 (N_7113,N_7032,N_6899);
xor U7114 (N_7114,N_6924,N_7030);
xnor U7115 (N_7115,N_6965,N_6911);
xor U7116 (N_7116,N_6918,N_6993);
nand U7117 (N_7117,N_7026,N_6922);
nand U7118 (N_7118,N_6902,N_6955);
nor U7119 (N_7119,N_6908,N_6890);
nor U7120 (N_7120,N_6922,N_7036);
xor U7121 (N_7121,N_6934,N_6968);
and U7122 (N_7122,N_7011,N_6939);
and U7123 (N_7123,N_6899,N_6895);
xor U7124 (N_7124,N_6942,N_6949);
nor U7125 (N_7125,N_6944,N_6913);
or U7126 (N_7126,N_6994,N_7013);
and U7127 (N_7127,N_6959,N_6949);
nor U7128 (N_7128,N_6906,N_7027);
nand U7129 (N_7129,N_6993,N_7002);
xnor U7130 (N_7130,N_6998,N_6890);
nor U7131 (N_7131,N_7007,N_6922);
or U7132 (N_7132,N_6913,N_6989);
and U7133 (N_7133,N_6893,N_6896);
and U7134 (N_7134,N_7004,N_6948);
or U7135 (N_7135,N_6898,N_7013);
or U7136 (N_7136,N_6970,N_6937);
or U7137 (N_7137,N_7028,N_6885);
nor U7138 (N_7138,N_6982,N_6909);
nand U7139 (N_7139,N_6949,N_7018);
and U7140 (N_7140,N_7011,N_6885);
nand U7141 (N_7141,N_6920,N_6912);
and U7142 (N_7142,N_6953,N_6946);
nor U7143 (N_7143,N_6985,N_6964);
nand U7144 (N_7144,N_7030,N_6918);
and U7145 (N_7145,N_6934,N_6953);
nand U7146 (N_7146,N_6909,N_7011);
xnor U7147 (N_7147,N_6957,N_7001);
nor U7148 (N_7148,N_7032,N_7018);
nor U7149 (N_7149,N_7033,N_6926);
or U7150 (N_7150,N_6938,N_6924);
nor U7151 (N_7151,N_7038,N_6893);
or U7152 (N_7152,N_7016,N_6938);
nor U7153 (N_7153,N_6897,N_6900);
and U7154 (N_7154,N_7001,N_6898);
or U7155 (N_7155,N_6962,N_6948);
or U7156 (N_7156,N_7001,N_6911);
or U7157 (N_7157,N_7002,N_6983);
and U7158 (N_7158,N_6976,N_6998);
nor U7159 (N_7159,N_6940,N_7028);
nor U7160 (N_7160,N_7018,N_7000);
or U7161 (N_7161,N_6947,N_6881);
or U7162 (N_7162,N_7009,N_6945);
or U7163 (N_7163,N_6916,N_6948);
xnor U7164 (N_7164,N_6979,N_6950);
xor U7165 (N_7165,N_7029,N_7009);
nor U7166 (N_7166,N_6902,N_7026);
nor U7167 (N_7167,N_6997,N_6966);
or U7168 (N_7168,N_6958,N_6969);
xnor U7169 (N_7169,N_6933,N_6912);
and U7170 (N_7170,N_6897,N_7026);
nor U7171 (N_7171,N_6917,N_7030);
nor U7172 (N_7172,N_6954,N_6956);
nor U7173 (N_7173,N_7023,N_6880);
and U7174 (N_7174,N_7039,N_6938);
nand U7175 (N_7175,N_7000,N_6952);
nand U7176 (N_7176,N_6939,N_7031);
xnor U7177 (N_7177,N_6963,N_6890);
xor U7178 (N_7178,N_6946,N_6925);
nor U7179 (N_7179,N_7037,N_6911);
nor U7180 (N_7180,N_6894,N_7026);
nand U7181 (N_7181,N_6919,N_7002);
or U7182 (N_7182,N_7019,N_6922);
and U7183 (N_7183,N_6989,N_6978);
xnor U7184 (N_7184,N_7028,N_6997);
and U7185 (N_7185,N_6987,N_6880);
or U7186 (N_7186,N_6908,N_7007);
xor U7187 (N_7187,N_7014,N_6979);
xnor U7188 (N_7188,N_6889,N_6975);
xnor U7189 (N_7189,N_6892,N_6999);
and U7190 (N_7190,N_6971,N_6900);
and U7191 (N_7191,N_6935,N_6901);
or U7192 (N_7192,N_7031,N_6882);
xor U7193 (N_7193,N_6893,N_6886);
nand U7194 (N_7194,N_7030,N_6989);
nand U7195 (N_7195,N_6993,N_6940);
xnor U7196 (N_7196,N_7018,N_6932);
nor U7197 (N_7197,N_6971,N_6973);
or U7198 (N_7198,N_6960,N_6954);
nand U7199 (N_7199,N_6927,N_6975);
and U7200 (N_7200,N_7051,N_7172);
or U7201 (N_7201,N_7116,N_7141);
or U7202 (N_7202,N_7056,N_7121);
nor U7203 (N_7203,N_7154,N_7081);
and U7204 (N_7204,N_7101,N_7112);
or U7205 (N_7205,N_7143,N_7097);
nand U7206 (N_7206,N_7067,N_7144);
nor U7207 (N_7207,N_7041,N_7174);
or U7208 (N_7208,N_7103,N_7178);
nand U7209 (N_7209,N_7155,N_7098);
xnor U7210 (N_7210,N_7196,N_7126);
xor U7211 (N_7211,N_7123,N_7107);
and U7212 (N_7212,N_7120,N_7104);
xnor U7213 (N_7213,N_7072,N_7160);
nor U7214 (N_7214,N_7170,N_7085);
xnor U7215 (N_7215,N_7193,N_7094);
and U7216 (N_7216,N_7158,N_7163);
xnor U7217 (N_7217,N_7054,N_7066);
or U7218 (N_7218,N_7052,N_7140);
nand U7219 (N_7219,N_7151,N_7093);
and U7220 (N_7220,N_7149,N_7086);
and U7221 (N_7221,N_7092,N_7148);
nand U7222 (N_7222,N_7164,N_7118);
xor U7223 (N_7223,N_7139,N_7059);
xor U7224 (N_7224,N_7062,N_7135);
nand U7225 (N_7225,N_7084,N_7064);
or U7226 (N_7226,N_7070,N_7156);
and U7227 (N_7227,N_7091,N_7082);
xnor U7228 (N_7228,N_7176,N_7069);
or U7229 (N_7229,N_7183,N_7113);
nor U7230 (N_7230,N_7175,N_7138);
and U7231 (N_7231,N_7169,N_7130);
nor U7232 (N_7232,N_7075,N_7105);
or U7233 (N_7233,N_7132,N_7087);
nand U7234 (N_7234,N_7061,N_7159);
xor U7235 (N_7235,N_7186,N_7142);
nor U7236 (N_7236,N_7182,N_7045);
xnor U7237 (N_7237,N_7194,N_7180);
xnor U7238 (N_7238,N_7044,N_7074);
nand U7239 (N_7239,N_7187,N_7189);
or U7240 (N_7240,N_7165,N_7137);
and U7241 (N_7241,N_7146,N_7134);
nor U7242 (N_7242,N_7109,N_7055);
and U7243 (N_7243,N_7049,N_7177);
and U7244 (N_7244,N_7150,N_7166);
or U7245 (N_7245,N_7131,N_7079);
xor U7246 (N_7246,N_7099,N_7171);
xnor U7247 (N_7247,N_7133,N_7157);
and U7248 (N_7248,N_7119,N_7089);
nor U7249 (N_7249,N_7073,N_7199);
or U7250 (N_7250,N_7108,N_7065);
nor U7251 (N_7251,N_7136,N_7167);
nor U7252 (N_7252,N_7161,N_7188);
and U7253 (N_7253,N_7198,N_7168);
and U7254 (N_7254,N_7185,N_7128);
nor U7255 (N_7255,N_7048,N_7096);
or U7256 (N_7256,N_7053,N_7173);
or U7257 (N_7257,N_7078,N_7114);
nor U7258 (N_7258,N_7077,N_7153);
xor U7259 (N_7259,N_7181,N_7063);
nor U7260 (N_7260,N_7076,N_7110);
and U7261 (N_7261,N_7095,N_7080);
xor U7262 (N_7262,N_7047,N_7058);
nor U7263 (N_7263,N_7179,N_7102);
nor U7264 (N_7264,N_7068,N_7083);
xnor U7265 (N_7265,N_7129,N_7115);
and U7266 (N_7266,N_7197,N_7050);
nor U7267 (N_7267,N_7192,N_7071);
nor U7268 (N_7268,N_7043,N_7127);
or U7269 (N_7269,N_7090,N_7125);
nand U7270 (N_7270,N_7088,N_7190);
and U7271 (N_7271,N_7191,N_7184);
xnor U7272 (N_7272,N_7124,N_7111);
and U7273 (N_7273,N_7057,N_7117);
or U7274 (N_7274,N_7122,N_7162);
nor U7275 (N_7275,N_7147,N_7046);
xnor U7276 (N_7276,N_7145,N_7060);
nor U7277 (N_7277,N_7040,N_7042);
and U7278 (N_7278,N_7195,N_7100);
and U7279 (N_7279,N_7152,N_7106);
or U7280 (N_7280,N_7183,N_7091);
nor U7281 (N_7281,N_7111,N_7057);
xor U7282 (N_7282,N_7188,N_7126);
or U7283 (N_7283,N_7070,N_7160);
or U7284 (N_7284,N_7145,N_7141);
or U7285 (N_7285,N_7197,N_7048);
and U7286 (N_7286,N_7158,N_7122);
nor U7287 (N_7287,N_7132,N_7121);
or U7288 (N_7288,N_7063,N_7080);
nand U7289 (N_7289,N_7087,N_7156);
nand U7290 (N_7290,N_7121,N_7192);
nand U7291 (N_7291,N_7048,N_7125);
xnor U7292 (N_7292,N_7144,N_7145);
and U7293 (N_7293,N_7072,N_7116);
and U7294 (N_7294,N_7045,N_7081);
nand U7295 (N_7295,N_7148,N_7091);
and U7296 (N_7296,N_7199,N_7101);
and U7297 (N_7297,N_7188,N_7140);
nand U7298 (N_7298,N_7040,N_7115);
or U7299 (N_7299,N_7064,N_7136);
nand U7300 (N_7300,N_7083,N_7074);
and U7301 (N_7301,N_7123,N_7053);
and U7302 (N_7302,N_7137,N_7132);
nand U7303 (N_7303,N_7147,N_7130);
and U7304 (N_7304,N_7042,N_7048);
xor U7305 (N_7305,N_7045,N_7084);
nand U7306 (N_7306,N_7165,N_7044);
xnor U7307 (N_7307,N_7118,N_7067);
xor U7308 (N_7308,N_7152,N_7071);
xor U7309 (N_7309,N_7181,N_7170);
nor U7310 (N_7310,N_7044,N_7066);
or U7311 (N_7311,N_7077,N_7104);
and U7312 (N_7312,N_7055,N_7063);
nor U7313 (N_7313,N_7175,N_7197);
or U7314 (N_7314,N_7188,N_7121);
or U7315 (N_7315,N_7041,N_7047);
and U7316 (N_7316,N_7198,N_7170);
nand U7317 (N_7317,N_7155,N_7152);
xor U7318 (N_7318,N_7187,N_7150);
nand U7319 (N_7319,N_7163,N_7091);
and U7320 (N_7320,N_7137,N_7140);
xnor U7321 (N_7321,N_7129,N_7164);
and U7322 (N_7322,N_7132,N_7129);
or U7323 (N_7323,N_7074,N_7050);
or U7324 (N_7324,N_7109,N_7087);
and U7325 (N_7325,N_7063,N_7145);
nand U7326 (N_7326,N_7052,N_7085);
nand U7327 (N_7327,N_7083,N_7098);
nor U7328 (N_7328,N_7053,N_7071);
nand U7329 (N_7329,N_7161,N_7186);
or U7330 (N_7330,N_7107,N_7166);
or U7331 (N_7331,N_7179,N_7074);
nor U7332 (N_7332,N_7085,N_7132);
and U7333 (N_7333,N_7156,N_7141);
nand U7334 (N_7334,N_7179,N_7059);
or U7335 (N_7335,N_7196,N_7150);
or U7336 (N_7336,N_7061,N_7173);
or U7337 (N_7337,N_7121,N_7041);
and U7338 (N_7338,N_7040,N_7089);
or U7339 (N_7339,N_7173,N_7051);
nor U7340 (N_7340,N_7064,N_7168);
nand U7341 (N_7341,N_7079,N_7139);
nor U7342 (N_7342,N_7144,N_7182);
xnor U7343 (N_7343,N_7163,N_7045);
and U7344 (N_7344,N_7180,N_7174);
and U7345 (N_7345,N_7120,N_7121);
and U7346 (N_7346,N_7130,N_7074);
nand U7347 (N_7347,N_7176,N_7159);
or U7348 (N_7348,N_7040,N_7155);
nand U7349 (N_7349,N_7094,N_7147);
or U7350 (N_7350,N_7079,N_7089);
xor U7351 (N_7351,N_7081,N_7098);
and U7352 (N_7352,N_7172,N_7090);
and U7353 (N_7353,N_7167,N_7079);
nand U7354 (N_7354,N_7103,N_7139);
nor U7355 (N_7355,N_7057,N_7137);
and U7356 (N_7356,N_7180,N_7098);
nand U7357 (N_7357,N_7105,N_7087);
nand U7358 (N_7358,N_7126,N_7045);
nor U7359 (N_7359,N_7087,N_7121);
nand U7360 (N_7360,N_7218,N_7352);
nand U7361 (N_7361,N_7293,N_7336);
nand U7362 (N_7362,N_7202,N_7251);
nor U7363 (N_7363,N_7328,N_7277);
nand U7364 (N_7364,N_7219,N_7340);
nand U7365 (N_7365,N_7294,N_7236);
nor U7366 (N_7366,N_7232,N_7215);
nand U7367 (N_7367,N_7306,N_7243);
nor U7368 (N_7368,N_7256,N_7272);
or U7369 (N_7369,N_7220,N_7229);
and U7370 (N_7370,N_7217,N_7212);
and U7371 (N_7371,N_7302,N_7273);
nor U7372 (N_7372,N_7319,N_7288);
or U7373 (N_7373,N_7206,N_7322);
and U7374 (N_7374,N_7201,N_7270);
nor U7375 (N_7375,N_7254,N_7292);
xnor U7376 (N_7376,N_7262,N_7300);
or U7377 (N_7377,N_7263,N_7305);
nand U7378 (N_7378,N_7303,N_7259);
nor U7379 (N_7379,N_7249,N_7241);
xnor U7380 (N_7380,N_7221,N_7320);
and U7381 (N_7381,N_7289,N_7280);
xor U7382 (N_7382,N_7250,N_7234);
nand U7383 (N_7383,N_7257,N_7346);
xnor U7384 (N_7384,N_7271,N_7237);
or U7385 (N_7385,N_7246,N_7313);
or U7386 (N_7386,N_7299,N_7327);
xor U7387 (N_7387,N_7356,N_7200);
or U7388 (N_7388,N_7248,N_7334);
nand U7389 (N_7389,N_7296,N_7285);
xor U7390 (N_7390,N_7351,N_7258);
nor U7391 (N_7391,N_7231,N_7337);
nor U7392 (N_7392,N_7211,N_7333);
or U7393 (N_7393,N_7216,N_7224);
and U7394 (N_7394,N_7233,N_7239);
or U7395 (N_7395,N_7307,N_7349);
xnor U7396 (N_7396,N_7255,N_7317);
or U7397 (N_7397,N_7311,N_7341);
or U7398 (N_7398,N_7261,N_7282);
or U7399 (N_7399,N_7310,N_7348);
or U7400 (N_7400,N_7284,N_7359);
xor U7401 (N_7401,N_7279,N_7324);
and U7402 (N_7402,N_7338,N_7358);
and U7403 (N_7403,N_7230,N_7223);
nor U7404 (N_7404,N_7286,N_7253);
and U7405 (N_7405,N_7344,N_7227);
xor U7406 (N_7406,N_7203,N_7308);
or U7407 (N_7407,N_7315,N_7268);
or U7408 (N_7408,N_7287,N_7316);
and U7409 (N_7409,N_7207,N_7332);
xor U7410 (N_7410,N_7321,N_7265);
nand U7411 (N_7411,N_7290,N_7213);
xnor U7412 (N_7412,N_7210,N_7335);
xnor U7413 (N_7413,N_7355,N_7252);
nand U7414 (N_7414,N_7240,N_7204);
nor U7415 (N_7415,N_7269,N_7222);
xnor U7416 (N_7416,N_7228,N_7330);
xnor U7417 (N_7417,N_7314,N_7347);
xor U7418 (N_7418,N_7242,N_7301);
nand U7419 (N_7419,N_7353,N_7331);
and U7420 (N_7420,N_7343,N_7245);
nand U7421 (N_7421,N_7298,N_7325);
xnor U7422 (N_7422,N_7297,N_7244);
nand U7423 (N_7423,N_7214,N_7208);
nor U7424 (N_7424,N_7238,N_7357);
nand U7425 (N_7425,N_7264,N_7309);
and U7426 (N_7426,N_7295,N_7304);
or U7427 (N_7427,N_7354,N_7281);
or U7428 (N_7428,N_7267,N_7283);
xor U7429 (N_7429,N_7275,N_7226);
and U7430 (N_7430,N_7339,N_7274);
and U7431 (N_7431,N_7350,N_7278);
nor U7432 (N_7432,N_7260,N_7225);
xnor U7433 (N_7433,N_7326,N_7291);
xnor U7434 (N_7434,N_7312,N_7342);
nor U7435 (N_7435,N_7329,N_7235);
and U7436 (N_7436,N_7318,N_7266);
and U7437 (N_7437,N_7205,N_7345);
or U7438 (N_7438,N_7323,N_7247);
nor U7439 (N_7439,N_7276,N_7209);
nand U7440 (N_7440,N_7251,N_7352);
nor U7441 (N_7441,N_7343,N_7351);
nor U7442 (N_7442,N_7333,N_7277);
nor U7443 (N_7443,N_7323,N_7296);
and U7444 (N_7444,N_7308,N_7311);
and U7445 (N_7445,N_7350,N_7344);
nand U7446 (N_7446,N_7212,N_7309);
nand U7447 (N_7447,N_7205,N_7323);
or U7448 (N_7448,N_7300,N_7276);
and U7449 (N_7449,N_7306,N_7251);
nand U7450 (N_7450,N_7201,N_7338);
nand U7451 (N_7451,N_7334,N_7291);
or U7452 (N_7452,N_7353,N_7279);
nor U7453 (N_7453,N_7293,N_7334);
nand U7454 (N_7454,N_7307,N_7319);
xor U7455 (N_7455,N_7349,N_7240);
nor U7456 (N_7456,N_7223,N_7290);
nand U7457 (N_7457,N_7285,N_7213);
xor U7458 (N_7458,N_7292,N_7259);
xor U7459 (N_7459,N_7225,N_7251);
xnor U7460 (N_7460,N_7331,N_7256);
xor U7461 (N_7461,N_7304,N_7359);
xor U7462 (N_7462,N_7240,N_7310);
or U7463 (N_7463,N_7311,N_7312);
and U7464 (N_7464,N_7242,N_7238);
nand U7465 (N_7465,N_7202,N_7314);
xor U7466 (N_7466,N_7297,N_7310);
nor U7467 (N_7467,N_7202,N_7280);
or U7468 (N_7468,N_7301,N_7253);
or U7469 (N_7469,N_7297,N_7335);
or U7470 (N_7470,N_7211,N_7297);
nor U7471 (N_7471,N_7314,N_7216);
xor U7472 (N_7472,N_7210,N_7263);
or U7473 (N_7473,N_7289,N_7300);
nand U7474 (N_7474,N_7352,N_7211);
and U7475 (N_7475,N_7254,N_7287);
xor U7476 (N_7476,N_7216,N_7345);
and U7477 (N_7477,N_7324,N_7269);
and U7478 (N_7478,N_7304,N_7246);
nand U7479 (N_7479,N_7314,N_7297);
nor U7480 (N_7480,N_7345,N_7291);
and U7481 (N_7481,N_7295,N_7213);
or U7482 (N_7482,N_7312,N_7203);
nand U7483 (N_7483,N_7322,N_7232);
and U7484 (N_7484,N_7314,N_7331);
or U7485 (N_7485,N_7336,N_7264);
or U7486 (N_7486,N_7333,N_7266);
nor U7487 (N_7487,N_7357,N_7335);
and U7488 (N_7488,N_7327,N_7319);
and U7489 (N_7489,N_7215,N_7206);
nand U7490 (N_7490,N_7252,N_7215);
or U7491 (N_7491,N_7338,N_7247);
xor U7492 (N_7492,N_7257,N_7291);
nand U7493 (N_7493,N_7280,N_7293);
and U7494 (N_7494,N_7205,N_7339);
or U7495 (N_7495,N_7203,N_7264);
nand U7496 (N_7496,N_7247,N_7260);
nand U7497 (N_7497,N_7322,N_7304);
nor U7498 (N_7498,N_7254,N_7319);
nor U7499 (N_7499,N_7310,N_7247);
xnor U7500 (N_7500,N_7352,N_7284);
or U7501 (N_7501,N_7305,N_7307);
and U7502 (N_7502,N_7300,N_7316);
nand U7503 (N_7503,N_7352,N_7238);
nand U7504 (N_7504,N_7255,N_7251);
nor U7505 (N_7505,N_7328,N_7278);
or U7506 (N_7506,N_7243,N_7218);
and U7507 (N_7507,N_7253,N_7256);
xnor U7508 (N_7508,N_7268,N_7238);
or U7509 (N_7509,N_7262,N_7349);
nand U7510 (N_7510,N_7331,N_7212);
and U7511 (N_7511,N_7220,N_7224);
or U7512 (N_7512,N_7270,N_7353);
or U7513 (N_7513,N_7205,N_7257);
or U7514 (N_7514,N_7221,N_7346);
nor U7515 (N_7515,N_7206,N_7253);
or U7516 (N_7516,N_7351,N_7210);
xor U7517 (N_7517,N_7295,N_7303);
nor U7518 (N_7518,N_7325,N_7251);
nor U7519 (N_7519,N_7258,N_7204);
xnor U7520 (N_7520,N_7485,N_7456);
nand U7521 (N_7521,N_7370,N_7504);
nor U7522 (N_7522,N_7373,N_7429);
xor U7523 (N_7523,N_7484,N_7483);
nand U7524 (N_7524,N_7479,N_7401);
and U7525 (N_7525,N_7469,N_7508);
or U7526 (N_7526,N_7482,N_7394);
nand U7527 (N_7527,N_7464,N_7408);
or U7528 (N_7528,N_7505,N_7512);
or U7529 (N_7529,N_7510,N_7441);
nand U7530 (N_7530,N_7473,N_7491);
and U7531 (N_7531,N_7434,N_7445);
or U7532 (N_7532,N_7371,N_7404);
nand U7533 (N_7533,N_7361,N_7486);
xnor U7534 (N_7534,N_7500,N_7514);
nor U7535 (N_7535,N_7474,N_7369);
nand U7536 (N_7536,N_7366,N_7495);
or U7537 (N_7537,N_7502,N_7431);
nand U7538 (N_7538,N_7470,N_7421);
or U7539 (N_7539,N_7409,N_7368);
or U7540 (N_7540,N_7415,N_7391);
or U7541 (N_7541,N_7390,N_7496);
or U7542 (N_7542,N_7438,N_7399);
nand U7543 (N_7543,N_7492,N_7403);
nor U7544 (N_7544,N_7416,N_7420);
or U7545 (N_7545,N_7396,N_7414);
nor U7546 (N_7546,N_7487,N_7515);
and U7547 (N_7547,N_7400,N_7519);
and U7548 (N_7548,N_7480,N_7364);
or U7549 (N_7549,N_7382,N_7406);
and U7550 (N_7550,N_7372,N_7516);
and U7551 (N_7551,N_7448,N_7365);
nand U7552 (N_7552,N_7446,N_7459);
and U7553 (N_7553,N_7466,N_7418);
or U7554 (N_7554,N_7439,N_7501);
nor U7555 (N_7555,N_7374,N_7509);
xor U7556 (N_7556,N_7385,N_7475);
nor U7557 (N_7557,N_7433,N_7503);
nor U7558 (N_7558,N_7497,N_7422);
nor U7559 (N_7559,N_7402,N_7413);
nand U7560 (N_7560,N_7379,N_7426);
nor U7561 (N_7561,N_7511,N_7481);
xnor U7562 (N_7562,N_7407,N_7463);
or U7563 (N_7563,N_7506,N_7455);
and U7564 (N_7564,N_7384,N_7452);
nor U7565 (N_7565,N_7398,N_7397);
xnor U7566 (N_7566,N_7363,N_7477);
nor U7567 (N_7567,N_7380,N_7378);
nand U7568 (N_7568,N_7412,N_7518);
and U7569 (N_7569,N_7517,N_7376);
nand U7570 (N_7570,N_7465,N_7388);
nor U7571 (N_7571,N_7423,N_7442);
or U7572 (N_7572,N_7471,N_7360);
nand U7573 (N_7573,N_7507,N_7461);
nand U7574 (N_7574,N_7478,N_7386);
nor U7575 (N_7575,N_7387,N_7488);
and U7576 (N_7576,N_7362,N_7460);
nor U7577 (N_7577,N_7513,N_7476);
and U7578 (N_7578,N_7417,N_7457);
or U7579 (N_7579,N_7432,N_7405);
or U7580 (N_7580,N_7427,N_7458);
nand U7581 (N_7581,N_7490,N_7410);
and U7582 (N_7582,N_7450,N_7411);
or U7583 (N_7583,N_7454,N_7462);
nor U7584 (N_7584,N_7444,N_7449);
nand U7585 (N_7585,N_7424,N_7472);
and U7586 (N_7586,N_7489,N_7428);
nor U7587 (N_7587,N_7493,N_7381);
xor U7588 (N_7588,N_7467,N_7430);
nor U7589 (N_7589,N_7498,N_7389);
nand U7590 (N_7590,N_7447,N_7395);
xor U7591 (N_7591,N_7468,N_7435);
or U7592 (N_7592,N_7499,N_7393);
and U7593 (N_7593,N_7425,N_7383);
or U7594 (N_7594,N_7377,N_7375);
or U7595 (N_7595,N_7437,N_7451);
nor U7596 (N_7596,N_7392,N_7419);
xor U7597 (N_7597,N_7494,N_7440);
nand U7598 (N_7598,N_7453,N_7436);
nor U7599 (N_7599,N_7443,N_7367);
and U7600 (N_7600,N_7370,N_7381);
nand U7601 (N_7601,N_7516,N_7417);
xnor U7602 (N_7602,N_7481,N_7513);
or U7603 (N_7603,N_7496,N_7479);
nor U7604 (N_7604,N_7409,N_7448);
nand U7605 (N_7605,N_7428,N_7455);
xor U7606 (N_7606,N_7405,N_7517);
nor U7607 (N_7607,N_7369,N_7506);
xor U7608 (N_7608,N_7510,N_7445);
nand U7609 (N_7609,N_7446,N_7447);
nand U7610 (N_7610,N_7404,N_7503);
nand U7611 (N_7611,N_7410,N_7456);
or U7612 (N_7612,N_7417,N_7393);
xor U7613 (N_7613,N_7473,N_7406);
and U7614 (N_7614,N_7444,N_7462);
and U7615 (N_7615,N_7411,N_7460);
nor U7616 (N_7616,N_7462,N_7486);
nor U7617 (N_7617,N_7515,N_7443);
or U7618 (N_7618,N_7432,N_7506);
nor U7619 (N_7619,N_7407,N_7424);
nor U7620 (N_7620,N_7517,N_7455);
nor U7621 (N_7621,N_7457,N_7391);
and U7622 (N_7622,N_7496,N_7378);
nor U7623 (N_7623,N_7405,N_7492);
xor U7624 (N_7624,N_7511,N_7415);
nor U7625 (N_7625,N_7494,N_7442);
nand U7626 (N_7626,N_7377,N_7379);
or U7627 (N_7627,N_7398,N_7459);
and U7628 (N_7628,N_7460,N_7468);
nor U7629 (N_7629,N_7429,N_7384);
nand U7630 (N_7630,N_7519,N_7406);
or U7631 (N_7631,N_7376,N_7430);
or U7632 (N_7632,N_7455,N_7480);
xor U7633 (N_7633,N_7486,N_7510);
nand U7634 (N_7634,N_7452,N_7450);
nand U7635 (N_7635,N_7399,N_7479);
or U7636 (N_7636,N_7387,N_7518);
xor U7637 (N_7637,N_7377,N_7495);
xor U7638 (N_7638,N_7422,N_7461);
xnor U7639 (N_7639,N_7453,N_7401);
or U7640 (N_7640,N_7498,N_7444);
nand U7641 (N_7641,N_7458,N_7447);
xor U7642 (N_7642,N_7391,N_7458);
xor U7643 (N_7643,N_7420,N_7474);
and U7644 (N_7644,N_7402,N_7393);
and U7645 (N_7645,N_7370,N_7492);
nor U7646 (N_7646,N_7458,N_7505);
or U7647 (N_7647,N_7407,N_7366);
xor U7648 (N_7648,N_7430,N_7478);
nand U7649 (N_7649,N_7384,N_7437);
xnor U7650 (N_7650,N_7421,N_7372);
nand U7651 (N_7651,N_7419,N_7493);
and U7652 (N_7652,N_7470,N_7418);
nor U7653 (N_7653,N_7504,N_7388);
or U7654 (N_7654,N_7427,N_7374);
and U7655 (N_7655,N_7491,N_7433);
xor U7656 (N_7656,N_7489,N_7444);
xor U7657 (N_7657,N_7370,N_7413);
nor U7658 (N_7658,N_7488,N_7482);
xor U7659 (N_7659,N_7488,N_7410);
and U7660 (N_7660,N_7422,N_7456);
or U7661 (N_7661,N_7407,N_7519);
nand U7662 (N_7662,N_7400,N_7508);
xnor U7663 (N_7663,N_7501,N_7502);
nand U7664 (N_7664,N_7439,N_7368);
or U7665 (N_7665,N_7515,N_7486);
xnor U7666 (N_7666,N_7516,N_7435);
xnor U7667 (N_7667,N_7402,N_7404);
nand U7668 (N_7668,N_7401,N_7466);
xor U7669 (N_7669,N_7402,N_7414);
xnor U7670 (N_7670,N_7512,N_7401);
nor U7671 (N_7671,N_7516,N_7453);
and U7672 (N_7672,N_7452,N_7512);
xor U7673 (N_7673,N_7463,N_7372);
nor U7674 (N_7674,N_7435,N_7433);
or U7675 (N_7675,N_7386,N_7374);
or U7676 (N_7676,N_7481,N_7382);
and U7677 (N_7677,N_7496,N_7425);
or U7678 (N_7678,N_7470,N_7378);
or U7679 (N_7679,N_7394,N_7516);
xnor U7680 (N_7680,N_7605,N_7607);
xnor U7681 (N_7681,N_7603,N_7630);
xor U7682 (N_7682,N_7601,N_7539);
or U7683 (N_7683,N_7676,N_7678);
xnor U7684 (N_7684,N_7589,N_7572);
and U7685 (N_7685,N_7663,N_7565);
nor U7686 (N_7686,N_7673,N_7664);
xor U7687 (N_7687,N_7626,N_7570);
and U7688 (N_7688,N_7583,N_7669);
nor U7689 (N_7689,N_7540,N_7606);
nor U7690 (N_7690,N_7580,N_7610);
and U7691 (N_7691,N_7616,N_7608);
xor U7692 (N_7692,N_7526,N_7615);
or U7693 (N_7693,N_7567,N_7552);
or U7694 (N_7694,N_7613,N_7535);
nor U7695 (N_7695,N_7592,N_7523);
nor U7696 (N_7696,N_7650,N_7633);
and U7697 (N_7697,N_7566,N_7550);
xnor U7698 (N_7698,N_7656,N_7623);
or U7699 (N_7699,N_7635,N_7679);
and U7700 (N_7700,N_7674,N_7600);
nand U7701 (N_7701,N_7581,N_7612);
and U7702 (N_7702,N_7555,N_7636);
or U7703 (N_7703,N_7662,N_7670);
nor U7704 (N_7704,N_7575,N_7548);
xor U7705 (N_7705,N_7668,N_7647);
nor U7706 (N_7706,N_7564,N_7631);
or U7707 (N_7707,N_7648,N_7598);
and U7708 (N_7708,N_7585,N_7624);
or U7709 (N_7709,N_7549,N_7594);
nor U7710 (N_7710,N_7595,N_7551);
or U7711 (N_7711,N_7641,N_7538);
xnor U7712 (N_7712,N_7541,N_7617);
nand U7713 (N_7713,N_7666,N_7671);
and U7714 (N_7714,N_7638,N_7659);
or U7715 (N_7715,N_7532,N_7536);
nor U7716 (N_7716,N_7556,N_7531);
nand U7717 (N_7717,N_7576,N_7542);
or U7718 (N_7718,N_7558,N_7563);
nand U7719 (N_7719,N_7599,N_7649);
xor U7720 (N_7720,N_7654,N_7597);
nand U7721 (N_7721,N_7578,N_7584);
xnor U7722 (N_7722,N_7561,N_7559);
nor U7723 (N_7723,N_7639,N_7562);
nand U7724 (N_7724,N_7568,N_7653);
nand U7725 (N_7725,N_7646,N_7618);
or U7726 (N_7726,N_7627,N_7620);
nand U7727 (N_7727,N_7672,N_7657);
xnor U7728 (N_7728,N_7590,N_7645);
or U7729 (N_7729,N_7553,N_7602);
nor U7730 (N_7730,N_7667,N_7521);
xor U7731 (N_7731,N_7614,N_7622);
nor U7732 (N_7732,N_7557,N_7644);
and U7733 (N_7733,N_7609,N_7632);
nand U7734 (N_7734,N_7529,N_7619);
nor U7735 (N_7735,N_7554,N_7591);
nor U7736 (N_7736,N_7588,N_7587);
and U7737 (N_7737,N_7628,N_7629);
nor U7738 (N_7738,N_7545,N_7577);
nand U7739 (N_7739,N_7582,N_7621);
and U7740 (N_7740,N_7528,N_7522);
and U7741 (N_7741,N_7544,N_7665);
nor U7742 (N_7742,N_7637,N_7651);
or U7743 (N_7743,N_7652,N_7569);
and U7744 (N_7744,N_7524,N_7675);
nor U7745 (N_7745,N_7579,N_7677);
nand U7746 (N_7746,N_7546,N_7625);
nand U7747 (N_7747,N_7574,N_7634);
or U7748 (N_7748,N_7593,N_7533);
xnor U7749 (N_7749,N_7527,N_7571);
nor U7750 (N_7750,N_7560,N_7658);
nand U7751 (N_7751,N_7547,N_7520);
and U7752 (N_7752,N_7661,N_7537);
or U7753 (N_7753,N_7660,N_7525);
or U7754 (N_7754,N_7530,N_7611);
nor U7755 (N_7755,N_7640,N_7643);
xnor U7756 (N_7756,N_7604,N_7586);
and U7757 (N_7757,N_7642,N_7596);
nand U7758 (N_7758,N_7655,N_7573);
nor U7759 (N_7759,N_7534,N_7543);
or U7760 (N_7760,N_7608,N_7585);
xnor U7761 (N_7761,N_7657,N_7624);
nand U7762 (N_7762,N_7662,N_7597);
nand U7763 (N_7763,N_7565,N_7668);
nand U7764 (N_7764,N_7664,N_7610);
nand U7765 (N_7765,N_7597,N_7542);
or U7766 (N_7766,N_7578,N_7619);
nor U7767 (N_7767,N_7643,N_7529);
or U7768 (N_7768,N_7632,N_7546);
nand U7769 (N_7769,N_7586,N_7602);
nand U7770 (N_7770,N_7660,N_7659);
nand U7771 (N_7771,N_7569,N_7635);
nor U7772 (N_7772,N_7597,N_7525);
and U7773 (N_7773,N_7621,N_7596);
nor U7774 (N_7774,N_7673,N_7654);
nor U7775 (N_7775,N_7646,N_7599);
and U7776 (N_7776,N_7618,N_7650);
and U7777 (N_7777,N_7611,N_7524);
and U7778 (N_7778,N_7679,N_7588);
and U7779 (N_7779,N_7572,N_7678);
xnor U7780 (N_7780,N_7585,N_7672);
or U7781 (N_7781,N_7636,N_7553);
or U7782 (N_7782,N_7562,N_7606);
or U7783 (N_7783,N_7604,N_7553);
xnor U7784 (N_7784,N_7626,N_7666);
xnor U7785 (N_7785,N_7569,N_7669);
and U7786 (N_7786,N_7631,N_7538);
or U7787 (N_7787,N_7570,N_7545);
nand U7788 (N_7788,N_7638,N_7584);
or U7789 (N_7789,N_7654,N_7664);
and U7790 (N_7790,N_7671,N_7607);
nand U7791 (N_7791,N_7602,N_7619);
nand U7792 (N_7792,N_7535,N_7653);
and U7793 (N_7793,N_7585,N_7588);
xor U7794 (N_7794,N_7619,N_7663);
and U7795 (N_7795,N_7673,N_7665);
or U7796 (N_7796,N_7539,N_7530);
nand U7797 (N_7797,N_7664,N_7589);
nand U7798 (N_7798,N_7668,N_7615);
and U7799 (N_7799,N_7613,N_7655);
xor U7800 (N_7800,N_7664,N_7646);
nand U7801 (N_7801,N_7658,N_7671);
or U7802 (N_7802,N_7622,N_7639);
xor U7803 (N_7803,N_7593,N_7558);
and U7804 (N_7804,N_7526,N_7668);
nor U7805 (N_7805,N_7651,N_7594);
nor U7806 (N_7806,N_7635,N_7644);
nor U7807 (N_7807,N_7595,N_7543);
nor U7808 (N_7808,N_7615,N_7555);
nor U7809 (N_7809,N_7583,N_7618);
nand U7810 (N_7810,N_7667,N_7548);
and U7811 (N_7811,N_7667,N_7658);
nand U7812 (N_7812,N_7530,N_7570);
or U7813 (N_7813,N_7673,N_7658);
nand U7814 (N_7814,N_7527,N_7638);
xnor U7815 (N_7815,N_7631,N_7654);
nand U7816 (N_7816,N_7618,N_7591);
or U7817 (N_7817,N_7660,N_7644);
or U7818 (N_7818,N_7615,N_7642);
or U7819 (N_7819,N_7528,N_7624);
nor U7820 (N_7820,N_7619,N_7645);
and U7821 (N_7821,N_7668,N_7530);
nand U7822 (N_7822,N_7653,N_7567);
or U7823 (N_7823,N_7635,N_7564);
and U7824 (N_7824,N_7663,N_7586);
xnor U7825 (N_7825,N_7632,N_7579);
nand U7826 (N_7826,N_7633,N_7587);
nand U7827 (N_7827,N_7548,N_7631);
or U7828 (N_7828,N_7549,N_7642);
or U7829 (N_7829,N_7565,N_7607);
and U7830 (N_7830,N_7659,N_7647);
or U7831 (N_7831,N_7630,N_7656);
nand U7832 (N_7832,N_7545,N_7603);
xnor U7833 (N_7833,N_7621,N_7614);
xnor U7834 (N_7834,N_7632,N_7635);
and U7835 (N_7835,N_7649,N_7626);
nand U7836 (N_7836,N_7538,N_7586);
xnor U7837 (N_7837,N_7654,N_7603);
or U7838 (N_7838,N_7562,N_7592);
nand U7839 (N_7839,N_7580,N_7617);
xor U7840 (N_7840,N_7680,N_7713);
or U7841 (N_7841,N_7793,N_7760);
nand U7842 (N_7842,N_7759,N_7748);
and U7843 (N_7843,N_7770,N_7826);
or U7844 (N_7844,N_7731,N_7730);
nand U7845 (N_7845,N_7720,N_7694);
nand U7846 (N_7846,N_7837,N_7792);
xnor U7847 (N_7847,N_7832,N_7754);
xnor U7848 (N_7848,N_7688,N_7802);
and U7849 (N_7849,N_7779,N_7810);
nand U7850 (N_7850,N_7708,N_7716);
xor U7851 (N_7851,N_7725,N_7796);
and U7852 (N_7852,N_7744,N_7797);
and U7853 (N_7853,N_7813,N_7738);
and U7854 (N_7854,N_7724,N_7767);
or U7855 (N_7855,N_7781,N_7714);
nor U7856 (N_7856,N_7681,N_7703);
nand U7857 (N_7857,N_7787,N_7717);
and U7858 (N_7858,N_7684,N_7762);
or U7859 (N_7859,N_7712,N_7686);
and U7860 (N_7860,N_7799,N_7822);
nand U7861 (N_7861,N_7682,N_7710);
nor U7862 (N_7862,N_7747,N_7752);
nor U7863 (N_7863,N_7758,N_7782);
nor U7864 (N_7864,N_7816,N_7778);
and U7865 (N_7865,N_7817,N_7791);
xnor U7866 (N_7866,N_7695,N_7701);
or U7867 (N_7867,N_7818,N_7709);
xor U7868 (N_7868,N_7711,N_7824);
nor U7869 (N_7869,N_7719,N_7765);
nor U7870 (N_7870,N_7803,N_7689);
or U7871 (N_7871,N_7735,N_7795);
xnor U7872 (N_7872,N_7789,N_7704);
or U7873 (N_7873,N_7788,N_7806);
and U7874 (N_7874,N_7728,N_7718);
or U7875 (N_7875,N_7838,N_7729);
and U7876 (N_7876,N_7707,N_7780);
nand U7877 (N_7877,N_7785,N_7819);
or U7878 (N_7878,N_7755,N_7739);
nor U7879 (N_7879,N_7798,N_7773);
nand U7880 (N_7880,N_7777,N_7732);
and U7881 (N_7881,N_7740,N_7727);
xnor U7882 (N_7882,N_7775,N_7699);
and U7883 (N_7883,N_7828,N_7702);
nand U7884 (N_7884,N_7763,N_7687);
and U7885 (N_7885,N_7746,N_7756);
and U7886 (N_7886,N_7742,N_7805);
and U7887 (N_7887,N_7726,N_7698);
nor U7888 (N_7888,N_7696,N_7804);
nand U7889 (N_7889,N_7691,N_7766);
nand U7890 (N_7890,N_7776,N_7723);
nor U7891 (N_7891,N_7825,N_7764);
and U7892 (N_7892,N_7750,N_7743);
and U7893 (N_7893,N_7812,N_7737);
xor U7894 (N_7894,N_7820,N_7706);
nand U7895 (N_7895,N_7734,N_7829);
xor U7896 (N_7896,N_7808,N_7839);
xnor U7897 (N_7897,N_7823,N_7692);
nand U7898 (N_7898,N_7700,N_7821);
and U7899 (N_7899,N_7790,N_7800);
nand U7900 (N_7900,N_7834,N_7807);
nor U7901 (N_7901,N_7809,N_7835);
nor U7902 (N_7902,N_7736,N_7715);
xnor U7903 (N_7903,N_7722,N_7794);
and U7904 (N_7904,N_7690,N_7786);
nor U7905 (N_7905,N_7811,N_7693);
xnor U7906 (N_7906,N_7830,N_7745);
nand U7907 (N_7907,N_7749,N_7705);
and U7908 (N_7908,N_7771,N_7827);
nor U7909 (N_7909,N_7761,N_7757);
and U7910 (N_7910,N_7721,N_7768);
xnor U7911 (N_7911,N_7836,N_7784);
xor U7912 (N_7912,N_7685,N_7774);
and U7913 (N_7913,N_7831,N_7814);
and U7914 (N_7914,N_7741,N_7769);
nor U7915 (N_7915,N_7683,N_7733);
nor U7916 (N_7916,N_7697,N_7833);
nand U7917 (N_7917,N_7753,N_7772);
or U7918 (N_7918,N_7815,N_7751);
nor U7919 (N_7919,N_7783,N_7801);
xnor U7920 (N_7920,N_7780,N_7786);
nor U7921 (N_7921,N_7829,N_7699);
xor U7922 (N_7922,N_7692,N_7811);
nor U7923 (N_7923,N_7759,N_7703);
or U7924 (N_7924,N_7829,N_7680);
nand U7925 (N_7925,N_7707,N_7824);
nand U7926 (N_7926,N_7770,N_7705);
xnor U7927 (N_7927,N_7689,N_7799);
and U7928 (N_7928,N_7681,N_7712);
nand U7929 (N_7929,N_7712,N_7825);
nor U7930 (N_7930,N_7693,N_7744);
and U7931 (N_7931,N_7685,N_7725);
and U7932 (N_7932,N_7693,N_7689);
nand U7933 (N_7933,N_7816,N_7709);
nand U7934 (N_7934,N_7754,N_7833);
nand U7935 (N_7935,N_7682,N_7815);
or U7936 (N_7936,N_7806,N_7803);
or U7937 (N_7937,N_7737,N_7690);
nor U7938 (N_7938,N_7788,N_7763);
or U7939 (N_7939,N_7782,N_7750);
nand U7940 (N_7940,N_7834,N_7823);
nand U7941 (N_7941,N_7832,N_7682);
and U7942 (N_7942,N_7742,N_7726);
nand U7943 (N_7943,N_7808,N_7795);
nand U7944 (N_7944,N_7804,N_7719);
xnor U7945 (N_7945,N_7818,N_7696);
and U7946 (N_7946,N_7687,N_7760);
and U7947 (N_7947,N_7734,N_7816);
or U7948 (N_7948,N_7689,N_7762);
or U7949 (N_7949,N_7719,N_7724);
xnor U7950 (N_7950,N_7691,N_7835);
nor U7951 (N_7951,N_7746,N_7686);
nor U7952 (N_7952,N_7821,N_7812);
xor U7953 (N_7953,N_7711,N_7804);
and U7954 (N_7954,N_7800,N_7681);
nor U7955 (N_7955,N_7799,N_7716);
xnor U7956 (N_7956,N_7728,N_7801);
xnor U7957 (N_7957,N_7737,N_7795);
xnor U7958 (N_7958,N_7796,N_7759);
xnor U7959 (N_7959,N_7806,N_7694);
nand U7960 (N_7960,N_7763,N_7685);
nor U7961 (N_7961,N_7824,N_7832);
nand U7962 (N_7962,N_7777,N_7764);
xnor U7963 (N_7963,N_7771,N_7807);
and U7964 (N_7964,N_7762,N_7729);
xor U7965 (N_7965,N_7815,N_7746);
and U7966 (N_7966,N_7742,N_7715);
nor U7967 (N_7967,N_7735,N_7765);
xor U7968 (N_7968,N_7702,N_7711);
nand U7969 (N_7969,N_7825,N_7778);
or U7970 (N_7970,N_7733,N_7794);
nor U7971 (N_7971,N_7742,N_7826);
and U7972 (N_7972,N_7691,N_7792);
nor U7973 (N_7973,N_7745,N_7770);
or U7974 (N_7974,N_7827,N_7705);
or U7975 (N_7975,N_7791,N_7746);
xor U7976 (N_7976,N_7725,N_7789);
or U7977 (N_7977,N_7777,N_7731);
nor U7978 (N_7978,N_7749,N_7683);
nand U7979 (N_7979,N_7707,N_7719);
and U7980 (N_7980,N_7708,N_7688);
or U7981 (N_7981,N_7745,N_7720);
nand U7982 (N_7982,N_7687,N_7776);
nand U7983 (N_7983,N_7686,N_7818);
nor U7984 (N_7984,N_7683,N_7709);
and U7985 (N_7985,N_7688,N_7698);
or U7986 (N_7986,N_7753,N_7686);
xor U7987 (N_7987,N_7720,N_7741);
and U7988 (N_7988,N_7702,N_7713);
or U7989 (N_7989,N_7828,N_7754);
nor U7990 (N_7990,N_7789,N_7680);
xnor U7991 (N_7991,N_7798,N_7815);
and U7992 (N_7992,N_7823,N_7802);
xor U7993 (N_7993,N_7685,N_7824);
nand U7994 (N_7994,N_7826,N_7792);
xnor U7995 (N_7995,N_7728,N_7733);
or U7996 (N_7996,N_7789,N_7833);
nor U7997 (N_7997,N_7771,N_7838);
nor U7998 (N_7998,N_7785,N_7709);
and U7999 (N_7999,N_7838,N_7832);
xor U8000 (N_8000,N_7937,N_7852);
xnor U8001 (N_8001,N_7878,N_7995);
xnor U8002 (N_8002,N_7926,N_7901);
nor U8003 (N_8003,N_7868,N_7961);
and U8004 (N_8004,N_7934,N_7996);
and U8005 (N_8005,N_7844,N_7975);
or U8006 (N_8006,N_7988,N_7883);
xnor U8007 (N_8007,N_7921,N_7923);
nand U8008 (N_8008,N_7889,N_7971);
and U8009 (N_8009,N_7997,N_7873);
nor U8010 (N_8010,N_7925,N_7879);
nand U8011 (N_8011,N_7893,N_7900);
xnor U8012 (N_8012,N_7843,N_7966);
nand U8013 (N_8013,N_7933,N_7951);
or U8014 (N_8014,N_7936,N_7977);
xnor U8015 (N_8015,N_7871,N_7916);
nand U8016 (N_8016,N_7944,N_7919);
and U8017 (N_8017,N_7981,N_7987);
or U8018 (N_8018,N_7902,N_7954);
nor U8019 (N_8019,N_7858,N_7970);
nor U8020 (N_8020,N_7999,N_7924);
nand U8021 (N_8021,N_7845,N_7976);
or U8022 (N_8022,N_7892,N_7956);
xnor U8023 (N_8023,N_7910,N_7959);
and U8024 (N_8024,N_7982,N_7905);
and U8025 (N_8025,N_7854,N_7891);
nand U8026 (N_8026,N_7938,N_7840);
xor U8027 (N_8027,N_7855,N_7940);
xor U8028 (N_8028,N_7967,N_7918);
and U8029 (N_8029,N_7880,N_7946);
nand U8030 (N_8030,N_7897,N_7890);
xnor U8031 (N_8031,N_7895,N_7853);
nand U8032 (N_8032,N_7964,N_7952);
nor U8033 (N_8033,N_7841,N_7915);
xor U8034 (N_8034,N_7958,N_7948);
xnor U8035 (N_8035,N_7993,N_7887);
or U8036 (N_8036,N_7888,N_7908);
nor U8037 (N_8037,N_7932,N_7943);
nand U8038 (N_8038,N_7973,N_7986);
xnor U8039 (N_8039,N_7864,N_7985);
nand U8040 (N_8040,N_7896,N_7857);
nand U8041 (N_8041,N_7990,N_7885);
xnor U8042 (N_8042,N_7904,N_7945);
nand U8043 (N_8043,N_7979,N_7863);
nor U8044 (N_8044,N_7906,N_7877);
xnor U8045 (N_8045,N_7927,N_7969);
and U8046 (N_8046,N_7984,N_7968);
and U8047 (N_8047,N_7869,N_7872);
nor U8048 (N_8048,N_7917,N_7862);
and U8049 (N_8049,N_7929,N_7874);
nor U8050 (N_8050,N_7875,N_7939);
nor U8051 (N_8051,N_7953,N_7886);
and U8052 (N_8052,N_7920,N_7931);
nand U8053 (N_8053,N_7860,N_7859);
nor U8054 (N_8054,N_7898,N_7846);
nor U8055 (N_8055,N_7955,N_7903);
nor U8056 (N_8056,N_7870,N_7957);
or U8057 (N_8057,N_7941,N_7928);
nand U8058 (N_8058,N_7912,N_7978);
nand U8059 (N_8059,N_7851,N_7861);
and U8060 (N_8060,N_7949,N_7849);
nand U8061 (N_8061,N_7842,N_7980);
xnor U8062 (N_8062,N_7962,N_7991);
and U8063 (N_8063,N_7907,N_7876);
xor U8064 (N_8064,N_7913,N_7856);
xor U8065 (N_8065,N_7881,N_7847);
nand U8066 (N_8066,N_7899,N_7884);
nand U8067 (N_8067,N_7909,N_7983);
and U8068 (N_8068,N_7992,N_7935);
nor U8069 (N_8069,N_7911,N_7998);
xnor U8070 (N_8070,N_7914,N_7850);
xnor U8071 (N_8071,N_7930,N_7848);
nor U8072 (N_8072,N_7965,N_7972);
xnor U8073 (N_8073,N_7947,N_7942);
or U8074 (N_8074,N_7989,N_7963);
or U8075 (N_8075,N_7922,N_7894);
or U8076 (N_8076,N_7865,N_7950);
nor U8077 (N_8077,N_7867,N_7866);
or U8078 (N_8078,N_7974,N_7994);
and U8079 (N_8079,N_7882,N_7960);
nand U8080 (N_8080,N_7917,N_7972);
or U8081 (N_8081,N_7940,N_7938);
nand U8082 (N_8082,N_7892,N_7916);
or U8083 (N_8083,N_7897,N_7941);
nand U8084 (N_8084,N_7878,N_7947);
or U8085 (N_8085,N_7871,N_7908);
nand U8086 (N_8086,N_7958,N_7935);
nand U8087 (N_8087,N_7866,N_7851);
nand U8088 (N_8088,N_7844,N_7958);
nor U8089 (N_8089,N_7963,N_7861);
and U8090 (N_8090,N_7975,N_7989);
or U8091 (N_8091,N_7906,N_7853);
and U8092 (N_8092,N_7944,N_7975);
or U8093 (N_8093,N_7903,N_7846);
or U8094 (N_8094,N_7924,N_7970);
nand U8095 (N_8095,N_7855,N_7942);
xnor U8096 (N_8096,N_7876,N_7914);
nor U8097 (N_8097,N_7871,N_7975);
nand U8098 (N_8098,N_7899,N_7922);
nand U8099 (N_8099,N_7870,N_7932);
xor U8100 (N_8100,N_7966,N_7948);
nor U8101 (N_8101,N_7926,N_7915);
or U8102 (N_8102,N_7861,N_7962);
nor U8103 (N_8103,N_7952,N_7936);
xnor U8104 (N_8104,N_7963,N_7848);
nand U8105 (N_8105,N_7955,N_7998);
nand U8106 (N_8106,N_7925,N_7874);
nor U8107 (N_8107,N_7876,N_7922);
xor U8108 (N_8108,N_7976,N_7989);
nor U8109 (N_8109,N_7906,N_7845);
nand U8110 (N_8110,N_7985,N_7854);
and U8111 (N_8111,N_7859,N_7956);
nor U8112 (N_8112,N_7866,N_7901);
nand U8113 (N_8113,N_7895,N_7997);
xnor U8114 (N_8114,N_7910,N_7985);
xor U8115 (N_8115,N_7873,N_7864);
or U8116 (N_8116,N_7959,N_7855);
or U8117 (N_8117,N_7842,N_7964);
and U8118 (N_8118,N_7907,N_7911);
xor U8119 (N_8119,N_7880,N_7873);
nor U8120 (N_8120,N_7969,N_7894);
nor U8121 (N_8121,N_7996,N_7903);
nor U8122 (N_8122,N_7985,N_7942);
or U8123 (N_8123,N_7870,N_7986);
xnor U8124 (N_8124,N_7879,N_7976);
and U8125 (N_8125,N_7956,N_7870);
nor U8126 (N_8126,N_7870,N_7893);
xor U8127 (N_8127,N_7854,N_7863);
nand U8128 (N_8128,N_7970,N_7908);
and U8129 (N_8129,N_7864,N_7861);
nand U8130 (N_8130,N_7925,N_7918);
and U8131 (N_8131,N_7923,N_7925);
and U8132 (N_8132,N_7905,N_7993);
xnor U8133 (N_8133,N_7989,N_7992);
and U8134 (N_8134,N_7927,N_7975);
and U8135 (N_8135,N_7989,N_7919);
and U8136 (N_8136,N_7920,N_7887);
and U8137 (N_8137,N_7903,N_7945);
nand U8138 (N_8138,N_7840,N_7983);
xor U8139 (N_8139,N_7994,N_7942);
and U8140 (N_8140,N_7898,N_7859);
nor U8141 (N_8141,N_7892,N_7860);
nand U8142 (N_8142,N_7847,N_7912);
and U8143 (N_8143,N_7860,N_7939);
xnor U8144 (N_8144,N_7958,N_7954);
or U8145 (N_8145,N_7913,N_7961);
xnor U8146 (N_8146,N_7925,N_7969);
nor U8147 (N_8147,N_7922,N_7907);
nand U8148 (N_8148,N_7933,N_7961);
xor U8149 (N_8149,N_7987,N_7854);
xor U8150 (N_8150,N_7887,N_7845);
and U8151 (N_8151,N_7936,N_7883);
nor U8152 (N_8152,N_7993,N_7931);
xor U8153 (N_8153,N_7905,N_7850);
nor U8154 (N_8154,N_7951,N_7963);
xor U8155 (N_8155,N_7863,N_7906);
or U8156 (N_8156,N_7868,N_7894);
and U8157 (N_8157,N_7900,N_7876);
or U8158 (N_8158,N_7871,N_7968);
or U8159 (N_8159,N_7884,N_7932);
xnor U8160 (N_8160,N_8029,N_8036);
and U8161 (N_8161,N_8144,N_8138);
and U8162 (N_8162,N_8047,N_8002);
nand U8163 (N_8163,N_8026,N_8063);
or U8164 (N_8164,N_8058,N_8121);
or U8165 (N_8165,N_8122,N_8021);
and U8166 (N_8166,N_8103,N_8046);
and U8167 (N_8167,N_8133,N_8069);
or U8168 (N_8168,N_8023,N_8132);
and U8169 (N_8169,N_8085,N_8042);
or U8170 (N_8170,N_8120,N_8020);
nand U8171 (N_8171,N_8080,N_8147);
nand U8172 (N_8172,N_8106,N_8072);
xnor U8173 (N_8173,N_8115,N_8093);
nor U8174 (N_8174,N_8001,N_8139);
nand U8175 (N_8175,N_8135,N_8044);
or U8176 (N_8176,N_8056,N_8073);
nand U8177 (N_8177,N_8079,N_8130);
xnor U8178 (N_8178,N_8030,N_8095);
nand U8179 (N_8179,N_8015,N_8022);
nand U8180 (N_8180,N_8101,N_8082);
and U8181 (N_8181,N_8158,N_8051);
and U8182 (N_8182,N_8146,N_8075);
or U8183 (N_8183,N_8127,N_8066);
nor U8184 (N_8184,N_8154,N_8092);
nand U8185 (N_8185,N_8113,N_8025);
and U8186 (N_8186,N_8007,N_8110);
xor U8187 (N_8187,N_8083,N_8009);
nand U8188 (N_8188,N_8142,N_8054);
xor U8189 (N_8189,N_8091,N_8011);
or U8190 (N_8190,N_8149,N_8043);
and U8191 (N_8191,N_8151,N_8145);
nand U8192 (N_8192,N_8057,N_8157);
nand U8193 (N_8193,N_8018,N_8140);
and U8194 (N_8194,N_8109,N_8003);
and U8195 (N_8195,N_8153,N_8148);
nand U8196 (N_8196,N_8039,N_8125);
or U8197 (N_8197,N_8071,N_8077);
or U8198 (N_8198,N_8027,N_8064);
and U8199 (N_8199,N_8116,N_8137);
nand U8200 (N_8200,N_8035,N_8098);
nand U8201 (N_8201,N_8010,N_8108);
and U8202 (N_8202,N_8076,N_8034);
nor U8203 (N_8203,N_8104,N_8031);
nand U8204 (N_8204,N_8152,N_8081);
xnor U8205 (N_8205,N_8059,N_8037);
or U8206 (N_8206,N_8105,N_8065);
nand U8207 (N_8207,N_8117,N_8004);
xor U8208 (N_8208,N_8124,N_8061);
nand U8209 (N_8209,N_8159,N_8074);
nor U8210 (N_8210,N_8041,N_8045);
or U8211 (N_8211,N_8123,N_8016);
or U8212 (N_8212,N_8099,N_8012);
nand U8213 (N_8213,N_8067,N_8032);
nor U8214 (N_8214,N_8006,N_8107);
xor U8215 (N_8215,N_8052,N_8048);
nor U8216 (N_8216,N_8134,N_8000);
and U8217 (N_8217,N_8033,N_8097);
nor U8218 (N_8218,N_8129,N_8090);
nand U8219 (N_8219,N_8053,N_8143);
and U8220 (N_8220,N_8155,N_8049);
nor U8221 (N_8221,N_8084,N_8005);
xor U8222 (N_8222,N_8094,N_8096);
xnor U8223 (N_8223,N_8119,N_8014);
xor U8224 (N_8224,N_8060,N_8038);
nor U8225 (N_8225,N_8111,N_8017);
nand U8226 (N_8226,N_8086,N_8114);
nor U8227 (N_8227,N_8126,N_8070);
nand U8228 (N_8228,N_8055,N_8062);
xor U8229 (N_8229,N_8128,N_8102);
xor U8230 (N_8230,N_8141,N_8008);
or U8231 (N_8231,N_8089,N_8100);
nor U8232 (N_8232,N_8028,N_8013);
and U8233 (N_8233,N_8040,N_8087);
nor U8234 (N_8234,N_8088,N_8078);
xor U8235 (N_8235,N_8150,N_8019);
nand U8236 (N_8236,N_8136,N_8156);
nor U8237 (N_8237,N_8050,N_8112);
nor U8238 (N_8238,N_8131,N_8118);
and U8239 (N_8239,N_8068,N_8024);
xor U8240 (N_8240,N_8018,N_8151);
xor U8241 (N_8241,N_8150,N_8028);
nor U8242 (N_8242,N_8130,N_8145);
nor U8243 (N_8243,N_8086,N_8102);
or U8244 (N_8244,N_8136,N_8103);
nor U8245 (N_8245,N_8009,N_8059);
nor U8246 (N_8246,N_8087,N_8060);
nand U8247 (N_8247,N_8140,N_8086);
nand U8248 (N_8248,N_8061,N_8014);
and U8249 (N_8249,N_8051,N_8052);
nor U8250 (N_8250,N_8150,N_8095);
nand U8251 (N_8251,N_8076,N_8147);
and U8252 (N_8252,N_8144,N_8014);
or U8253 (N_8253,N_8069,N_8027);
or U8254 (N_8254,N_8094,N_8105);
and U8255 (N_8255,N_8140,N_8007);
nor U8256 (N_8256,N_8104,N_8149);
nor U8257 (N_8257,N_8021,N_8057);
nor U8258 (N_8258,N_8056,N_8133);
nor U8259 (N_8259,N_8082,N_8154);
nor U8260 (N_8260,N_8101,N_8105);
xnor U8261 (N_8261,N_8050,N_8089);
nor U8262 (N_8262,N_8085,N_8150);
nor U8263 (N_8263,N_8118,N_8016);
or U8264 (N_8264,N_8004,N_8079);
nand U8265 (N_8265,N_8002,N_8121);
and U8266 (N_8266,N_8069,N_8094);
nor U8267 (N_8267,N_8121,N_8008);
nand U8268 (N_8268,N_8035,N_8112);
xor U8269 (N_8269,N_8021,N_8114);
xor U8270 (N_8270,N_8005,N_8109);
or U8271 (N_8271,N_8145,N_8023);
and U8272 (N_8272,N_8102,N_8117);
nor U8273 (N_8273,N_8061,N_8096);
nor U8274 (N_8274,N_8078,N_8144);
nand U8275 (N_8275,N_8095,N_8107);
nand U8276 (N_8276,N_8118,N_8142);
xor U8277 (N_8277,N_8088,N_8049);
nand U8278 (N_8278,N_8078,N_8082);
nand U8279 (N_8279,N_8113,N_8157);
nor U8280 (N_8280,N_8017,N_8009);
nand U8281 (N_8281,N_8051,N_8084);
or U8282 (N_8282,N_8045,N_8053);
xor U8283 (N_8283,N_8008,N_8084);
and U8284 (N_8284,N_8135,N_8040);
nor U8285 (N_8285,N_8024,N_8048);
nor U8286 (N_8286,N_8015,N_8103);
and U8287 (N_8287,N_8033,N_8158);
nor U8288 (N_8288,N_8000,N_8118);
or U8289 (N_8289,N_8053,N_8123);
and U8290 (N_8290,N_8131,N_8084);
nor U8291 (N_8291,N_8144,N_8147);
nor U8292 (N_8292,N_8057,N_8039);
or U8293 (N_8293,N_8029,N_8152);
and U8294 (N_8294,N_8101,N_8063);
nor U8295 (N_8295,N_8159,N_8147);
nor U8296 (N_8296,N_8086,N_8093);
nor U8297 (N_8297,N_8040,N_8061);
nand U8298 (N_8298,N_8155,N_8129);
nor U8299 (N_8299,N_8024,N_8112);
and U8300 (N_8300,N_8139,N_8130);
and U8301 (N_8301,N_8083,N_8019);
nand U8302 (N_8302,N_8105,N_8111);
or U8303 (N_8303,N_8062,N_8121);
nand U8304 (N_8304,N_8053,N_8075);
nor U8305 (N_8305,N_8010,N_8079);
or U8306 (N_8306,N_8123,N_8055);
or U8307 (N_8307,N_8089,N_8144);
or U8308 (N_8308,N_8134,N_8086);
xor U8309 (N_8309,N_8020,N_8076);
xor U8310 (N_8310,N_8088,N_8091);
nor U8311 (N_8311,N_8086,N_8158);
or U8312 (N_8312,N_8137,N_8072);
nand U8313 (N_8313,N_8100,N_8029);
nor U8314 (N_8314,N_8158,N_8127);
and U8315 (N_8315,N_8140,N_8029);
nor U8316 (N_8316,N_8037,N_8133);
nand U8317 (N_8317,N_8073,N_8130);
xnor U8318 (N_8318,N_8153,N_8030);
nand U8319 (N_8319,N_8002,N_8061);
nor U8320 (N_8320,N_8222,N_8190);
nand U8321 (N_8321,N_8292,N_8239);
nand U8322 (N_8322,N_8195,N_8275);
nand U8323 (N_8323,N_8290,N_8219);
and U8324 (N_8324,N_8167,N_8287);
and U8325 (N_8325,N_8231,N_8170);
and U8326 (N_8326,N_8210,N_8197);
or U8327 (N_8327,N_8270,N_8297);
nor U8328 (N_8328,N_8161,N_8244);
xnor U8329 (N_8329,N_8178,N_8160);
xor U8330 (N_8330,N_8173,N_8237);
nand U8331 (N_8331,N_8256,N_8242);
nand U8332 (N_8332,N_8207,N_8313);
nor U8333 (N_8333,N_8229,N_8276);
xor U8334 (N_8334,N_8204,N_8296);
nor U8335 (N_8335,N_8246,N_8234);
and U8336 (N_8336,N_8241,N_8230);
xor U8337 (N_8337,N_8303,N_8250);
nor U8338 (N_8338,N_8315,N_8221);
xnor U8339 (N_8339,N_8310,N_8214);
nand U8340 (N_8340,N_8181,N_8232);
nor U8341 (N_8341,N_8235,N_8259);
nor U8342 (N_8342,N_8304,N_8286);
or U8343 (N_8343,N_8257,N_8299);
nand U8344 (N_8344,N_8164,N_8288);
or U8345 (N_8345,N_8266,N_8278);
nor U8346 (N_8346,N_8179,N_8215);
nand U8347 (N_8347,N_8206,N_8284);
or U8348 (N_8348,N_8177,N_8260);
xor U8349 (N_8349,N_8302,N_8208);
nor U8350 (N_8350,N_8265,N_8247);
xnor U8351 (N_8351,N_8258,N_8238);
and U8352 (N_8352,N_8166,N_8171);
or U8353 (N_8353,N_8316,N_8306);
nor U8354 (N_8354,N_8199,N_8193);
and U8355 (N_8355,N_8174,N_8245);
or U8356 (N_8356,N_8311,N_8205);
nand U8357 (N_8357,N_8298,N_8200);
or U8358 (N_8358,N_8217,N_8180);
or U8359 (N_8359,N_8243,N_8182);
nor U8360 (N_8360,N_8312,N_8279);
nor U8361 (N_8361,N_8262,N_8189);
xor U8362 (N_8362,N_8273,N_8175);
nand U8363 (N_8363,N_8224,N_8196);
or U8364 (N_8364,N_8263,N_8213);
or U8365 (N_8365,N_8192,N_8209);
and U8366 (N_8366,N_8252,N_8248);
nand U8367 (N_8367,N_8283,N_8240);
and U8368 (N_8368,N_8317,N_8253);
nor U8369 (N_8369,N_8285,N_8227);
nor U8370 (N_8370,N_8194,N_8289);
xnor U8371 (N_8371,N_8255,N_8233);
or U8372 (N_8372,N_8163,N_8269);
xnor U8373 (N_8373,N_8307,N_8271);
or U8374 (N_8374,N_8293,N_8198);
nand U8375 (N_8375,N_8291,N_8191);
nor U8376 (N_8376,N_8264,N_8282);
and U8377 (N_8377,N_8186,N_8162);
or U8378 (N_8378,N_8201,N_8280);
nand U8379 (N_8379,N_8176,N_8185);
or U8380 (N_8380,N_8172,N_8277);
nor U8381 (N_8381,N_8274,N_8261);
or U8382 (N_8382,N_8268,N_8295);
and U8383 (N_8383,N_8294,N_8203);
nor U8384 (N_8384,N_8249,N_8308);
and U8385 (N_8385,N_8165,N_8305);
xnor U8386 (N_8386,N_8168,N_8187);
xor U8387 (N_8387,N_8301,N_8236);
nand U8388 (N_8388,N_8202,N_8220);
and U8389 (N_8389,N_8254,N_8216);
nand U8390 (N_8390,N_8281,N_8272);
nand U8391 (N_8391,N_8319,N_8184);
xor U8392 (N_8392,N_8169,N_8218);
and U8393 (N_8393,N_8228,N_8183);
xnor U8394 (N_8394,N_8267,N_8225);
nand U8395 (N_8395,N_8223,N_8309);
or U8396 (N_8396,N_8226,N_8318);
nor U8397 (N_8397,N_8212,N_8211);
or U8398 (N_8398,N_8251,N_8300);
xnor U8399 (N_8399,N_8188,N_8314);
xnor U8400 (N_8400,N_8235,N_8223);
nor U8401 (N_8401,N_8278,N_8175);
nand U8402 (N_8402,N_8246,N_8268);
nor U8403 (N_8403,N_8257,N_8307);
nor U8404 (N_8404,N_8208,N_8233);
xnor U8405 (N_8405,N_8300,N_8216);
nor U8406 (N_8406,N_8177,N_8165);
xor U8407 (N_8407,N_8199,N_8276);
xnor U8408 (N_8408,N_8242,N_8188);
and U8409 (N_8409,N_8253,N_8173);
nand U8410 (N_8410,N_8161,N_8273);
and U8411 (N_8411,N_8258,N_8187);
xor U8412 (N_8412,N_8193,N_8175);
xnor U8413 (N_8413,N_8183,N_8255);
nor U8414 (N_8414,N_8301,N_8262);
and U8415 (N_8415,N_8311,N_8177);
nand U8416 (N_8416,N_8168,N_8196);
nand U8417 (N_8417,N_8290,N_8235);
or U8418 (N_8418,N_8182,N_8178);
xnor U8419 (N_8419,N_8251,N_8267);
xnor U8420 (N_8420,N_8318,N_8311);
nand U8421 (N_8421,N_8201,N_8213);
or U8422 (N_8422,N_8243,N_8224);
and U8423 (N_8423,N_8181,N_8290);
xnor U8424 (N_8424,N_8194,N_8278);
and U8425 (N_8425,N_8248,N_8167);
or U8426 (N_8426,N_8186,N_8274);
xnor U8427 (N_8427,N_8314,N_8236);
nand U8428 (N_8428,N_8265,N_8171);
or U8429 (N_8429,N_8268,N_8236);
xor U8430 (N_8430,N_8224,N_8296);
nor U8431 (N_8431,N_8267,N_8190);
nand U8432 (N_8432,N_8233,N_8224);
and U8433 (N_8433,N_8165,N_8193);
nand U8434 (N_8434,N_8245,N_8242);
nor U8435 (N_8435,N_8182,N_8293);
nand U8436 (N_8436,N_8252,N_8194);
or U8437 (N_8437,N_8211,N_8215);
and U8438 (N_8438,N_8224,N_8249);
and U8439 (N_8439,N_8241,N_8168);
xor U8440 (N_8440,N_8172,N_8211);
xnor U8441 (N_8441,N_8237,N_8287);
and U8442 (N_8442,N_8219,N_8171);
and U8443 (N_8443,N_8248,N_8270);
xor U8444 (N_8444,N_8297,N_8163);
and U8445 (N_8445,N_8183,N_8180);
xnor U8446 (N_8446,N_8251,N_8208);
nand U8447 (N_8447,N_8239,N_8169);
nor U8448 (N_8448,N_8260,N_8305);
or U8449 (N_8449,N_8265,N_8236);
and U8450 (N_8450,N_8254,N_8308);
nand U8451 (N_8451,N_8299,N_8217);
nand U8452 (N_8452,N_8184,N_8253);
or U8453 (N_8453,N_8206,N_8264);
or U8454 (N_8454,N_8177,N_8251);
nand U8455 (N_8455,N_8183,N_8286);
xor U8456 (N_8456,N_8308,N_8267);
nand U8457 (N_8457,N_8315,N_8163);
nand U8458 (N_8458,N_8221,N_8219);
nor U8459 (N_8459,N_8213,N_8316);
and U8460 (N_8460,N_8233,N_8209);
nor U8461 (N_8461,N_8272,N_8316);
and U8462 (N_8462,N_8318,N_8298);
xor U8463 (N_8463,N_8310,N_8217);
and U8464 (N_8464,N_8240,N_8299);
and U8465 (N_8465,N_8223,N_8251);
nor U8466 (N_8466,N_8166,N_8226);
nor U8467 (N_8467,N_8316,N_8192);
nand U8468 (N_8468,N_8300,N_8298);
and U8469 (N_8469,N_8285,N_8188);
nor U8470 (N_8470,N_8163,N_8314);
and U8471 (N_8471,N_8275,N_8249);
xnor U8472 (N_8472,N_8190,N_8162);
or U8473 (N_8473,N_8180,N_8282);
xnor U8474 (N_8474,N_8214,N_8195);
or U8475 (N_8475,N_8220,N_8227);
nand U8476 (N_8476,N_8280,N_8240);
nand U8477 (N_8477,N_8172,N_8199);
and U8478 (N_8478,N_8312,N_8168);
nand U8479 (N_8479,N_8239,N_8258);
nand U8480 (N_8480,N_8438,N_8341);
nor U8481 (N_8481,N_8434,N_8420);
and U8482 (N_8482,N_8346,N_8334);
xor U8483 (N_8483,N_8469,N_8391);
nor U8484 (N_8484,N_8363,N_8451);
and U8485 (N_8485,N_8471,N_8418);
or U8486 (N_8486,N_8407,N_8394);
xor U8487 (N_8487,N_8321,N_8376);
nand U8488 (N_8488,N_8326,N_8406);
nand U8489 (N_8489,N_8371,N_8340);
or U8490 (N_8490,N_8343,N_8364);
or U8491 (N_8491,N_8479,N_8408);
nand U8492 (N_8492,N_8467,N_8424);
or U8493 (N_8493,N_8421,N_8413);
xnor U8494 (N_8494,N_8444,N_8445);
and U8495 (N_8495,N_8373,N_8442);
nor U8496 (N_8496,N_8349,N_8372);
nand U8497 (N_8497,N_8475,N_8459);
nor U8498 (N_8498,N_8377,N_8403);
nand U8499 (N_8499,N_8392,N_8390);
or U8500 (N_8500,N_8379,N_8337);
or U8501 (N_8501,N_8472,N_8374);
nor U8502 (N_8502,N_8370,N_8468);
or U8503 (N_8503,N_8386,N_8339);
or U8504 (N_8504,N_8345,N_8449);
or U8505 (N_8505,N_8415,N_8430);
or U8506 (N_8506,N_8362,N_8432);
nor U8507 (N_8507,N_8455,N_8387);
and U8508 (N_8508,N_8431,N_8401);
nand U8509 (N_8509,N_8375,N_8457);
xnor U8510 (N_8510,N_8325,N_8476);
or U8511 (N_8511,N_8478,N_8350);
and U8512 (N_8512,N_8440,N_8448);
or U8513 (N_8513,N_8351,N_8410);
and U8514 (N_8514,N_8389,N_8331);
nand U8515 (N_8515,N_8395,N_8416);
nand U8516 (N_8516,N_8384,N_8393);
nand U8517 (N_8517,N_8453,N_8464);
xor U8518 (N_8518,N_8433,N_8366);
or U8519 (N_8519,N_8458,N_8354);
or U8520 (N_8520,N_8419,N_8355);
and U8521 (N_8521,N_8404,N_8474);
or U8522 (N_8522,N_8398,N_8439);
nor U8523 (N_8523,N_8436,N_8347);
nor U8524 (N_8524,N_8443,N_8369);
xor U8525 (N_8525,N_8462,N_8332);
xnor U8526 (N_8526,N_8428,N_8423);
and U8527 (N_8527,N_8417,N_8473);
nand U8528 (N_8528,N_8409,N_8367);
nor U8529 (N_8529,N_8353,N_8335);
or U8530 (N_8530,N_8466,N_8338);
or U8531 (N_8531,N_8356,N_8402);
xnor U8532 (N_8532,N_8470,N_8437);
nand U8533 (N_8533,N_8422,N_8460);
or U8534 (N_8534,N_8429,N_8465);
or U8535 (N_8535,N_8359,N_8322);
nand U8536 (N_8536,N_8324,N_8441);
nor U8537 (N_8537,N_8358,N_8382);
or U8538 (N_8538,N_8452,N_8385);
or U8539 (N_8539,N_8396,N_8344);
xnor U8540 (N_8540,N_8477,N_8463);
or U8541 (N_8541,N_8365,N_8388);
nor U8542 (N_8542,N_8414,N_8336);
and U8543 (N_8543,N_8342,N_8397);
or U8544 (N_8544,N_8405,N_8411);
nor U8545 (N_8545,N_8461,N_8400);
nand U8546 (N_8546,N_8454,N_8412);
nor U8547 (N_8547,N_8435,N_8427);
nand U8548 (N_8548,N_8446,N_8383);
nand U8549 (N_8549,N_8323,N_8450);
nor U8550 (N_8550,N_8327,N_8330);
nor U8551 (N_8551,N_8399,N_8426);
and U8552 (N_8552,N_8357,N_8328);
xor U8553 (N_8553,N_8381,N_8447);
and U8554 (N_8554,N_8333,N_8361);
or U8555 (N_8555,N_8329,N_8425);
nor U8556 (N_8556,N_8352,N_8360);
xnor U8557 (N_8557,N_8378,N_8380);
xor U8558 (N_8558,N_8320,N_8456);
nor U8559 (N_8559,N_8368,N_8348);
and U8560 (N_8560,N_8418,N_8326);
xnor U8561 (N_8561,N_8418,N_8394);
or U8562 (N_8562,N_8377,N_8458);
or U8563 (N_8563,N_8323,N_8327);
and U8564 (N_8564,N_8323,N_8424);
and U8565 (N_8565,N_8349,N_8474);
xnor U8566 (N_8566,N_8321,N_8368);
nor U8567 (N_8567,N_8451,N_8456);
or U8568 (N_8568,N_8375,N_8430);
or U8569 (N_8569,N_8360,N_8335);
xnor U8570 (N_8570,N_8425,N_8400);
nor U8571 (N_8571,N_8425,N_8452);
nor U8572 (N_8572,N_8363,N_8388);
nand U8573 (N_8573,N_8331,N_8434);
xor U8574 (N_8574,N_8373,N_8431);
nand U8575 (N_8575,N_8391,N_8385);
nor U8576 (N_8576,N_8404,N_8339);
or U8577 (N_8577,N_8371,N_8401);
and U8578 (N_8578,N_8466,N_8321);
nand U8579 (N_8579,N_8463,N_8478);
xor U8580 (N_8580,N_8417,N_8465);
nor U8581 (N_8581,N_8456,N_8333);
or U8582 (N_8582,N_8390,N_8462);
and U8583 (N_8583,N_8370,N_8419);
nor U8584 (N_8584,N_8395,N_8347);
nand U8585 (N_8585,N_8362,N_8360);
xnor U8586 (N_8586,N_8466,N_8340);
and U8587 (N_8587,N_8373,N_8439);
nor U8588 (N_8588,N_8475,N_8346);
and U8589 (N_8589,N_8344,N_8457);
nand U8590 (N_8590,N_8355,N_8399);
and U8591 (N_8591,N_8478,N_8330);
nand U8592 (N_8592,N_8369,N_8426);
nor U8593 (N_8593,N_8332,N_8476);
nand U8594 (N_8594,N_8429,N_8385);
or U8595 (N_8595,N_8430,N_8341);
nor U8596 (N_8596,N_8461,N_8471);
nand U8597 (N_8597,N_8445,N_8350);
nor U8598 (N_8598,N_8337,N_8342);
or U8599 (N_8599,N_8479,N_8388);
xor U8600 (N_8600,N_8382,N_8347);
and U8601 (N_8601,N_8427,N_8347);
and U8602 (N_8602,N_8327,N_8440);
or U8603 (N_8603,N_8463,N_8379);
xnor U8604 (N_8604,N_8383,N_8342);
or U8605 (N_8605,N_8332,N_8380);
xor U8606 (N_8606,N_8328,N_8361);
nand U8607 (N_8607,N_8332,N_8460);
nor U8608 (N_8608,N_8394,N_8475);
xor U8609 (N_8609,N_8453,N_8445);
or U8610 (N_8610,N_8420,N_8350);
xnor U8611 (N_8611,N_8375,N_8345);
or U8612 (N_8612,N_8460,N_8414);
nor U8613 (N_8613,N_8327,N_8345);
and U8614 (N_8614,N_8382,N_8342);
nor U8615 (N_8615,N_8477,N_8428);
or U8616 (N_8616,N_8476,N_8364);
nand U8617 (N_8617,N_8453,N_8354);
nor U8618 (N_8618,N_8373,N_8428);
nand U8619 (N_8619,N_8417,N_8371);
nor U8620 (N_8620,N_8447,N_8408);
and U8621 (N_8621,N_8453,N_8350);
nand U8622 (N_8622,N_8328,N_8373);
or U8623 (N_8623,N_8376,N_8373);
xor U8624 (N_8624,N_8341,N_8452);
xor U8625 (N_8625,N_8401,N_8414);
and U8626 (N_8626,N_8331,N_8413);
nor U8627 (N_8627,N_8403,N_8476);
nand U8628 (N_8628,N_8382,N_8391);
or U8629 (N_8629,N_8366,N_8324);
xor U8630 (N_8630,N_8476,N_8409);
or U8631 (N_8631,N_8373,N_8478);
nor U8632 (N_8632,N_8324,N_8364);
nor U8633 (N_8633,N_8405,N_8367);
nor U8634 (N_8634,N_8348,N_8414);
or U8635 (N_8635,N_8398,N_8422);
or U8636 (N_8636,N_8337,N_8384);
or U8637 (N_8637,N_8356,N_8424);
nor U8638 (N_8638,N_8361,N_8404);
nor U8639 (N_8639,N_8421,N_8432);
and U8640 (N_8640,N_8557,N_8535);
and U8641 (N_8641,N_8517,N_8508);
and U8642 (N_8642,N_8540,N_8481);
and U8643 (N_8643,N_8631,N_8581);
nor U8644 (N_8644,N_8534,N_8525);
nand U8645 (N_8645,N_8612,N_8602);
or U8646 (N_8646,N_8635,N_8552);
and U8647 (N_8647,N_8561,N_8521);
nor U8648 (N_8648,N_8571,N_8502);
nor U8649 (N_8649,N_8568,N_8487);
nand U8650 (N_8650,N_8596,N_8504);
nor U8651 (N_8651,N_8514,N_8501);
or U8652 (N_8652,N_8606,N_8522);
nand U8653 (N_8653,N_8579,N_8482);
nand U8654 (N_8654,N_8513,N_8529);
or U8655 (N_8655,N_8630,N_8632);
or U8656 (N_8656,N_8576,N_8597);
xor U8657 (N_8657,N_8621,N_8609);
and U8658 (N_8658,N_8503,N_8492);
or U8659 (N_8659,N_8589,N_8528);
or U8660 (N_8660,N_8623,N_8572);
and U8661 (N_8661,N_8603,N_8499);
and U8662 (N_8662,N_8559,N_8539);
xor U8663 (N_8663,N_8553,N_8637);
or U8664 (N_8664,N_8538,N_8560);
nand U8665 (N_8665,N_8626,N_8537);
and U8666 (N_8666,N_8544,N_8498);
nand U8667 (N_8667,N_8566,N_8532);
xnor U8668 (N_8668,N_8491,N_8512);
or U8669 (N_8669,N_8614,N_8564);
and U8670 (N_8670,N_8556,N_8554);
nor U8671 (N_8671,N_8613,N_8531);
nor U8672 (N_8672,N_8628,N_8583);
xor U8673 (N_8673,N_8541,N_8578);
nand U8674 (N_8674,N_8598,N_8573);
or U8675 (N_8675,N_8618,N_8524);
or U8676 (N_8676,N_8625,N_8616);
nand U8677 (N_8677,N_8507,N_8530);
and U8678 (N_8678,N_8611,N_8627);
nor U8679 (N_8679,N_8518,N_8629);
nand U8680 (N_8680,N_8577,N_8563);
nor U8681 (N_8681,N_8523,N_8569);
and U8682 (N_8682,N_8550,N_8496);
and U8683 (N_8683,N_8584,N_8548);
or U8684 (N_8684,N_8497,N_8588);
nor U8685 (N_8685,N_8526,N_8565);
and U8686 (N_8686,N_8536,N_8510);
or U8687 (N_8687,N_8505,N_8533);
xnor U8688 (N_8688,N_8546,N_8634);
nor U8689 (N_8689,N_8620,N_8586);
nand U8690 (N_8690,N_8490,N_8567);
xnor U8691 (N_8691,N_8615,N_8604);
and U8692 (N_8692,N_8527,N_8608);
nor U8693 (N_8693,N_8639,N_8519);
xor U8694 (N_8694,N_8617,N_8574);
or U8695 (N_8695,N_8551,N_8595);
or U8696 (N_8696,N_8506,N_8580);
nand U8697 (N_8697,N_8545,N_8494);
nor U8698 (N_8698,N_8516,N_8622);
nor U8699 (N_8699,N_8558,N_8562);
xnor U8700 (N_8700,N_8601,N_8591);
nor U8701 (N_8701,N_8570,N_8509);
nor U8702 (N_8702,N_8484,N_8593);
or U8703 (N_8703,N_8493,N_8511);
nor U8704 (N_8704,N_8619,N_8587);
or U8705 (N_8705,N_8485,N_8599);
and U8706 (N_8706,N_8488,N_8500);
xor U8707 (N_8707,N_8575,N_8624);
xnor U8708 (N_8708,N_8495,N_8590);
nand U8709 (N_8709,N_8549,N_8520);
and U8710 (N_8710,N_8542,N_8555);
xor U8711 (N_8711,N_8486,N_8515);
and U8712 (N_8712,N_8610,N_8592);
xor U8713 (N_8713,N_8605,N_8489);
nand U8714 (N_8714,N_8633,N_8480);
nand U8715 (N_8715,N_8585,N_8636);
and U8716 (N_8716,N_8582,N_8543);
or U8717 (N_8717,N_8638,N_8594);
or U8718 (N_8718,N_8547,N_8483);
nor U8719 (N_8719,N_8600,N_8607);
xnor U8720 (N_8720,N_8539,N_8601);
nand U8721 (N_8721,N_8520,N_8621);
nand U8722 (N_8722,N_8484,N_8507);
or U8723 (N_8723,N_8529,N_8549);
xnor U8724 (N_8724,N_8526,N_8564);
nor U8725 (N_8725,N_8541,N_8538);
and U8726 (N_8726,N_8534,N_8579);
or U8727 (N_8727,N_8486,N_8605);
nor U8728 (N_8728,N_8587,N_8638);
or U8729 (N_8729,N_8523,N_8632);
nand U8730 (N_8730,N_8506,N_8512);
or U8731 (N_8731,N_8517,N_8527);
nor U8732 (N_8732,N_8630,N_8586);
nand U8733 (N_8733,N_8513,N_8635);
xor U8734 (N_8734,N_8511,N_8537);
or U8735 (N_8735,N_8507,N_8556);
xnor U8736 (N_8736,N_8568,N_8544);
xnor U8737 (N_8737,N_8556,N_8593);
and U8738 (N_8738,N_8519,N_8624);
nor U8739 (N_8739,N_8552,N_8483);
xor U8740 (N_8740,N_8537,N_8502);
or U8741 (N_8741,N_8546,N_8562);
or U8742 (N_8742,N_8559,N_8482);
nor U8743 (N_8743,N_8617,N_8538);
nor U8744 (N_8744,N_8617,N_8575);
nor U8745 (N_8745,N_8633,N_8513);
xor U8746 (N_8746,N_8517,N_8501);
xor U8747 (N_8747,N_8523,N_8564);
or U8748 (N_8748,N_8568,N_8541);
nor U8749 (N_8749,N_8613,N_8632);
xnor U8750 (N_8750,N_8609,N_8632);
nand U8751 (N_8751,N_8531,N_8483);
nand U8752 (N_8752,N_8518,N_8617);
or U8753 (N_8753,N_8508,N_8584);
xor U8754 (N_8754,N_8612,N_8569);
or U8755 (N_8755,N_8547,N_8600);
and U8756 (N_8756,N_8497,N_8557);
or U8757 (N_8757,N_8539,N_8556);
xnor U8758 (N_8758,N_8555,N_8500);
xnor U8759 (N_8759,N_8586,N_8526);
nor U8760 (N_8760,N_8487,N_8611);
and U8761 (N_8761,N_8614,N_8552);
xnor U8762 (N_8762,N_8637,N_8591);
and U8763 (N_8763,N_8559,N_8626);
nand U8764 (N_8764,N_8615,N_8492);
and U8765 (N_8765,N_8555,N_8584);
xnor U8766 (N_8766,N_8561,N_8596);
and U8767 (N_8767,N_8562,N_8519);
or U8768 (N_8768,N_8604,N_8595);
xor U8769 (N_8769,N_8515,N_8549);
and U8770 (N_8770,N_8500,N_8537);
xor U8771 (N_8771,N_8550,N_8518);
xnor U8772 (N_8772,N_8602,N_8527);
or U8773 (N_8773,N_8493,N_8603);
xnor U8774 (N_8774,N_8527,N_8585);
nand U8775 (N_8775,N_8484,N_8519);
xnor U8776 (N_8776,N_8595,N_8504);
nor U8777 (N_8777,N_8495,N_8547);
nor U8778 (N_8778,N_8603,N_8583);
nand U8779 (N_8779,N_8551,N_8634);
nand U8780 (N_8780,N_8636,N_8616);
nand U8781 (N_8781,N_8586,N_8614);
xor U8782 (N_8782,N_8495,N_8494);
and U8783 (N_8783,N_8579,N_8624);
or U8784 (N_8784,N_8504,N_8556);
and U8785 (N_8785,N_8543,N_8498);
nor U8786 (N_8786,N_8615,N_8536);
and U8787 (N_8787,N_8559,N_8533);
nand U8788 (N_8788,N_8538,N_8629);
or U8789 (N_8789,N_8539,N_8513);
xnor U8790 (N_8790,N_8557,N_8570);
xnor U8791 (N_8791,N_8548,N_8492);
nand U8792 (N_8792,N_8521,N_8554);
nor U8793 (N_8793,N_8589,N_8549);
xor U8794 (N_8794,N_8559,N_8639);
or U8795 (N_8795,N_8629,N_8564);
or U8796 (N_8796,N_8585,N_8635);
nand U8797 (N_8797,N_8568,N_8495);
or U8798 (N_8798,N_8605,N_8603);
and U8799 (N_8799,N_8630,N_8615);
or U8800 (N_8800,N_8714,N_8753);
xnor U8801 (N_8801,N_8759,N_8787);
xnor U8802 (N_8802,N_8725,N_8688);
nor U8803 (N_8803,N_8703,N_8773);
nor U8804 (N_8804,N_8648,N_8670);
or U8805 (N_8805,N_8765,N_8678);
nand U8806 (N_8806,N_8763,N_8727);
nor U8807 (N_8807,N_8656,N_8646);
xor U8808 (N_8808,N_8724,N_8658);
and U8809 (N_8809,N_8689,N_8743);
nor U8810 (N_8810,N_8739,N_8662);
xnor U8811 (N_8811,N_8708,N_8695);
nand U8812 (N_8812,N_8780,N_8660);
or U8813 (N_8813,N_8666,N_8653);
and U8814 (N_8814,N_8683,N_8735);
or U8815 (N_8815,N_8737,N_8652);
nor U8816 (N_8816,N_8779,N_8760);
and U8817 (N_8817,N_8702,N_8681);
nor U8818 (N_8818,N_8676,N_8645);
nand U8819 (N_8819,N_8642,N_8734);
nor U8820 (N_8820,N_8778,N_8793);
nor U8821 (N_8821,N_8748,N_8783);
or U8822 (N_8822,N_8694,N_8716);
nand U8823 (N_8823,N_8752,N_8758);
or U8824 (N_8824,N_8788,N_8697);
and U8825 (N_8825,N_8671,N_8796);
nand U8826 (N_8826,N_8731,N_8757);
or U8827 (N_8827,N_8649,N_8647);
nand U8828 (N_8828,N_8691,N_8718);
xor U8829 (N_8829,N_8685,N_8746);
and U8830 (N_8830,N_8749,N_8712);
or U8831 (N_8831,N_8770,N_8742);
nor U8832 (N_8832,N_8700,N_8730);
nor U8833 (N_8833,N_8684,N_8669);
and U8834 (N_8834,N_8672,N_8687);
xnor U8835 (N_8835,N_8772,N_8792);
xor U8836 (N_8836,N_8761,N_8767);
nor U8837 (N_8837,N_8696,N_8799);
xor U8838 (N_8838,N_8795,N_8728);
or U8839 (N_8839,N_8677,N_8690);
nand U8840 (N_8840,N_8794,N_8747);
nand U8841 (N_8841,N_8679,N_8674);
xor U8842 (N_8842,N_8673,N_8651);
nand U8843 (N_8843,N_8709,N_8657);
nand U8844 (N_8844,N_8692,N_8711);
and U8845 (N_8845,N_8717,N_8754);
xnor U8846 (N_8846,N_8650,N_8776);
or U8847 (N_8847,N_8721,N_8644);
and U8848 (N_8848,N_8664,N_8750);
nand U8849 (N_8849,N_8667,N_8741);
xnor U8850 (N_8850,N_8661,N_8707);
nor U8851 (N_8851,N_8715,N_8798);
xor U8852 (N_8852,N_8781,N_8693);
nand U8853 (N_8853,N_8641,N_8797);
and U8854 (N_8854,N_8789,N_8755);
nand U8855 (N_8855,N_8777,N_8768);
nor U8856 (N_8856,N_8726,N_8675);
and U8857 (N_8857,N_8665,N_8720);
nand U8858 (N_8858,N_8732,N_8699);
nor U8859 (N_8859,N_8784,N_8706);
nor U8860 (N_8860,N_8668,N_8719);
or U8861 (N_8861,N_8713,N_8771);
xor U8862 (N_8862,N_8698,N_8722);
and U8863 (N_8863,N_8791,N_8786);
or U8864 (N_8864,N_8762,N_8782);
or U8865 (N_8865,N_8751,N_8736);
nor U8866 (N_8866,N_8733,N_8744);
and U8867 (N_8867,N_8729,N_8769);
or U8868 (N_8868,N_8686,N_8659);
xor U8869 (N_8869,N_8723,N_8790);
or U8870 (N_8870,N_8745,N_8775);
nand U8871 (N_8871,N_8704,N_8682);
xor U8872 (N_8872,N_8680,N_8710);
xor U8873 (N_8873,N_8738,N_8701);
xor U8874 (N_8874,N_8764,N_8654);
nand U8875 (N_8875,N_8640,N_8655);
nand U8876 (N_8876,N_8705,N_8774);
nor U8877 (N_8877,N_8785,N_8740);
nor U8878 (N_8878,N_8766,N_8663);
nand U8879 (N_8879,N_8756,N_8643);
or U8880 (N_8880,N_8652,N_8672);
nor U8881 (N_8881,N_8793,N_8798);
nand U8882 (N_8882,N_8645,N_8714);
nand U8883 (N_8883,N_8750,N_8715);
and U8884 (N_8884,N_8657,N_8688);
nand U8885 (N_8885,N_8704,N_8788);
or U8886 (N_8886,N_8799,N_8681);
or U8887 (N_8887,N_8688,N_8649);
xor U8888 (N_8888,N_8691,N_8785);
nand U8889 (N_8889,N_8724,N_8738);
nand U8890 (N_8890,N_8715,N_8703);
or U8891 (N_8891,N_8666,N_8702);
xor U8892 (N_8892,N_8692,N_8729);
nand U8893 (N_8893,N_8732,N_8772);
or U8894 (N_8894,N_8707,N_8771);
nor U8895 (N_8895,N_8790,N_8681);
and U8896 (N_8896,N_8733,N_8721);
nand U8897 (N_8897,N_8670,N_8793);
or U8898 (N_8898,N_8730,N_8767);
nor U8899 (N_8899,N_8741,N_8725);
and U8900 (N_8900,N_8775,N_8682);
xor U8901 (N_8901,N_8708,N_8789);
or U8902 (N_8902,N_8658,N_8746);
or U8903 (N_8903,N_8663,N_8770);
xor U8904 (N_8904,N_8669,N_8782);
nor U8905 (N_8905,N_8793,N_8731);
nand U8906 (N_8906,N_8799,N_8777);
or U8907 (N_8907,N_8649,N_8732);
and U8908 (N_8908,N_8728,N_8675);
nor U8909 (N_8909,N_8731,N_8713);
nand U8910 (N_8910,N_8706,N_8672);
nor U8911 (N_8911,N_8660,N_8693);
nor U8912 (N_8912,N_8648,N_8747);
xnor U8913 (N_8913,N_8659,N_8718);
nor U8914 (N_8914,N_8723,N_8654);
or U8915 (N_8915,N_8670,N_8688);
or U8916 (N_8916,N_8798,N_8685);
and U8917 (N_8917,N_8780,N_8761);
and U8918 (N_8918,N_8731,N_8677);
or U8919 (N_8919,N_8660,N_8773);
nand U8920 (N_8920,N_8718,N_8797);
and U8921 (N_8921,N_8719,N_8643);
xnor U8922 (N_8922,N_8700,N_8758);
or U8923 (N_8923,N_8709,N_8645);
or U8924 (N_8924,N_8772,N_8686);
nor U8925 (N_8925,N_8733,N_8656);
xor U8926 (N_8926,N_8740,N_8713);
nor U8927 (N_8927,N_8686,N_8700);
xnor U8928 (N_8928,N_8655,N_8754);
nand U8929 (N_8929,N_8794,N_8670);
xor U8930 (N_8930,N_8754,N_8669);
and U8931 (N_8931,N_8758,N_8648);
xor U8932 (N_8932,N_8642,N_8784);
nor U8933 (N_8933,N_8789,N_8748);
xnor U8934 (N_8934,N_8674,N_8686);
xor U8935 (N_8935,N_8784,N_8645);
nor U8936 (N_8936,N_8792,N_8718);
nor U8937 (N_8937,N_8656,N_8759);
or U8938 (N_8938,N_8641,N_8758);
or U8939 (N_8939,N_8678,N_8641);
nor U8940 (N_8940,N_8727,N_8674);
xnor U8941 (N_8941,N_8647,N_8780);
nor U8942 (N_8942,N_8761,N_8748);
nor U8943 (N_8943,N_8731,N_8740);
nor U8944 (N_8944,N_8668,N_8720);
nor U8945 (N_8945,N_8649,N_8752);
and U8946 (N_8946,N_8664,N_8751);
or U8947 (N_8947,N_8695,N_8666);
xor U8948 (N_8948,N_8699,N_8798);
and U8949 (N_8949,N_8772,N_8724);
nand U8950 (N_8950,N_8686,N_8684);
or U8951 (N_8951,N_8783,N_8674);
xor U8952 (N_8952,N_8791,N_8782);
nor U8953 (N_8953,N_8664,N_8690);
or U8954 (N_8954,N_8794,N_8684);
nand U8955 (N_8955,N_8709,N_8758);
xor U8956 (N_8956,N_8770,N_8679);
and U8957 (N_8957,N_8646,N_8694);
nor U8958 (N_8958,N_8732,N_8709);
xnor U8959 (N_8959,N_8650,N_8662);
nand U8960 (N_8960,N_8810,N_8911);
or U8961 (N_8961,N_8862,N_8924);
and U8962 (N_8962,N_8825,N_8883);
xor U8963 (N_8963,N_8942,N_8820);
nor U8964 (N_8964,N_8807,N_8811);
and U8965 (N_8965,N_8945,N_8834);
xor U8966 (N_8966,N_8958,N_8946);
and U8967 (N_8967,N_8907,N_8879);
nor U8968 (N_8968,N_8864,N_8860);
nor U8969 (N_8969,N_8804,N_8902);
xnor U8970 (N_8970,N_8900,N_8812);
and U8971 (N_8971,N_8857,N_8826);
nand U8972 (N_8972,N_8899,N_8832);
nand U8973 (N_8973,N_8872,N_8819);
or U8974 (N_8974,N_8829,N_8806);
nand U8975 (N_8975,N_8897,N_8903);
or U8976 (N_8976,N_8861,N_8957);
nand U8977 (N_8977,N_8931,N_8888);
and U8978 (N_8978,N_8821,N_8892);
nand U8979 (N_8979,N_8882,N_8837);
nor U8980 (N_8980,N_8893,N_8853);
nand U8981 (N_8981,N_8841,N_8851);
or U8982 (N_8982,N_8865,N_8896);
nand U8983 (N_8983,N_8874,N_8824);
and U8984 (N_8984,N_8828,N_8930);
and U8985 (N_8985,N_8953,N_8939);
and U8986 (N_8986,N_8870,N_8955);
or U8987 (N_8987,N_8923,N_8836);
nor U8988 (N_8988,N_8854,N_8915);
nand U8989 (N_8989,N_8875,N_8920);
nand U8990 (N_8990,N_8885,N_8910);
or U8991 (N_8991,N_8863,N_8928);
nand U8992 (N_8992,N_8952,N_8889);
nand U8993 (N_8993,N_8926,N_8941);
and U8994 (N_8994,N_8919,N_8936);
nand U8995 (N_8995,N_8849,N_8816);
or U8996 (N_8996,N_8918,N_8839);
xor U8997 (N_8997,N_8814,N_8881);
or U8998 (N_8998,N_8867,N_8947);
and U8999 (N_8999,N_8925,N_8845);
xor U9000 (N_9000,N_8948,N_8800);
or U9001 (N_9001,N_8950,N_8934);
xnor U9002 (N_9002,N_8871,N_8884);
or U9003 (N_9003,N_8833,N_8949);
or U9004 (N_9004,N_8908,N_8886);
nor U9005 (N_9005,N_8842,N_8940);
xnor U9006 (N_9006,N_8831,N_8951);
and U9007 (N_9007,N_8823,N_8916);
or U9008 (N_9008,N_8901,N_8921);
nand U9009 (N_9009,N_8847,N_8817);
xor U9010 (N_9010,N_8898,N_8848);
nor U9011 (N_9011,N_8944,N_8933);
xor U9012 (N_9012,N_8868,N_8873);
and U9013 (N_9013,N_8912,N_8943);
xor U9014 (N_9014,N_8869,N_8809);
or U9015 (N_9015,N_8866,N_8852);
nor U9016 (N_9016,N_8935,N_8805);
nand U9017 (N_9017,N_8878,N_8813);
or U9018 (N_9018,N_8876,N_8818);
and U9019 (N_9019,N_8906,N_8956);
nor U9020 (N_9020,N_8856,N_8927);
xnor U9021 (N_9021,N_8855,N_8929);
xor U9022 (N_9022,N_8880,N_8914);
xor U9023 (N_9023,N_8815,N_8844);
and U9024 (N_9024,N_8938,N_8905);
xnor U9025 (N_9025,N_8803,N_8877);
and U9026 (N_9026,N_8827,N_8894);
or U9027 (N_9027,N_8890,N_8840);
nand U9028 (N_9028,N_8909,N_8895);
nand U9029 (N_9029,N_8959,N_8808);
xor U9030 (N_9030,N_8887,N_8922);
xor U9031 (N_9031,N_8932,N_8859);
and U9032 (N_9032,N_8846,N_8822);
or U9033 (N_9033,N_8801,N_8830);
or U9034 (N_9034,N_8858,N_8838);
and U9035 (N_9035,N_8913,N_8850);
xor U9036 (N_9036,N_8835,N_8843);
nand U9037 (N_9037,N_8917,N_8937);
nor U9038 (N_9038,N_8954,N_8802);
or U9039 (N_9039,N_8904,N_8891);
xor U9040 (N_9040,N_8837,N_8920);
nand U9041 (N_9041,N_8953,N_8936);
xor U9042 (N_9042,N_8821,N_8840);
and U9043 (N_9043,N_8822,N_8957);
nor U9044 (N_9044,N_8959,N_8847);
and U9045 (N_9045,N_8847,N_8844);
nand U9046 (N_9046,N_8873,N_8836);
xor U9047 (N_9047,N_8957,N_8890);
nand U9048 (N_9048,N_8930,N_8808);
nand U9049 (N_9049,N_8861,N_8842);
xnor U9050 (N_9050,N_8829,N_8860);
nand U9051 (N_9051,N_8932,N_8807);
nor U9052 (N_9052,N_8820,N_8925);
nor U9053 (N_9053,N_8897,N_8840);
or U9054 (N_9054,N_8904,N_8876);
and U9055 (N_9055,N_8883,N_8899);
xor U9056 (N_9056,N_8925,N_8935);
and U9057 (N_9057,N_8916,N_8929);
nor U9058 (N_9058,N_8942,N_8892);
xnor U9059 (N_9059,N_8909,N_8924);
nor U9060 (N_9060,N_8801,N_8931);
and U9061 (N_9061,N_8887,N_8808);
nor U9062 (N_9062,N_8868,N_8882);
xor U9063 (N_9063,N_8823,N_8878);
xor U9064 (N_9064,N_8930,N_8883);
nor U9065 (N_9065,N_8820,N_8959);
and U9066 (N_9066,N_8840,N_8921);
and U9067 (N_9067,N_8875,N_8945);
nor U9068 (N_9068,N_8899,N_8958);
nand U9069 (N_9069,N_8858,N_8924);
xor U9070 (N_9070,N_8896,N_8846);
xor U9071 (N_9071,N_8936,N_8869);
nor U9072 (N_9072,N_8854,N_8958);
nor U9073 (N_9073,N_8911,N_8929);
and U9074 (N_9074,N_8882,N_8881);
nand U9075 (N_9075,N_8947,N_8809);
xnor U9076 (N_9076,N_8870,N_8929);
nand U9077 (N_9077,N_8821,N_8857);
or U9078 (N_9078,N_8946,N_8841);
and U9079 (N_9079,N_8932,N_8940);
or U9080 (N_9080,N_8945,N_8826);
and U9081 (N_9081,N_8944,N_8840);
nand U9082 (N_9082,N_8853,N_8868);
or U9083 (N_9083,N_8869,N_8921);
xnor U9084 (N_9084,N_8883,N_8874);
nand U9085 (N_9085,N_8916,N_8909);
and U9086 (N_9086,N_8909,N_8854);
or U9087 (N_9087,N_8884,N_8877);
and U9088 (N_9088,N_8818,N_8822);
and U9089 (N_9089,N_8843,N_8921);
and U9090 (N_9090,N_8921,N_8821);
xnor U9091 (N_9091,N_8870,N_8947);
or U9092 (N_9092,N_8889,N_8931);
nand U9093 (N_9093,N_8803,N_8849);
nor U9094 (N_9094,N_8843,N_8874);
nor U9095 (N_9095,N_8885,N_8954);
xor U9096 (N_9096,N_8802,N_8929);
nand U9097 (N_9097,N_8824,N_8919);
or U9098 (N_9098,N_8911,N_8913);
nor U9099 (N_9099,N_8845,N_8888);
or U9100 (N_9100,N_8854,N_8850);
and U9101 (N_9101,N_8868,N_8885);
nor U9102 (N_9102,N_8951,N_8880);
nor U9103 (N_9103,N_8865,N_8815);
nand U9104 (N_9104,N_8945,N_8848);
and U9105 (N_9105,N_8855,N_8811);
xnor U9106 (N_9106,N_8899,N_8864);
xor U9107 (N_9107,N_8883,N_8819);
and U9108 (N_9108,N_8826,N_8919);
nor U9109 (N_9109,N_8833,N_8933);
or U9110 (N_9110,N_8872,N_8918);
nand U9111 (N_9111,N_8946,N_8833);
or U9112 (N_9112,N_8895,N_8859);
or U9113 (N_9113,N_8884,N_8860);
nor U9114 (N_9114,N_8901,N_8822);
nand U9115 (N_9115,N_8808,N_8928);
nor U9116 (N_9116,N_8807,N_8837);
nor U9117 (N_9117,N_8906,N_8939);
or U9118 (N_9118,N_8949,N_8928);
or U9119 (N_9119,N_8954,N_8929);
xnor U9120 (N_9120,N_8994,N_9082);
xor U9121 (N_9121,N_8978,N_9009);
xnor U9122 (N_9122,N_9045,N_8975);
and U9123 (N_9123,N_9097,N_9098);
or U9124 (N_9124,N_9085,N_8972);
nand U9125 (N_9125,N_8968,N_9003);
xnor U9126 (N_9126,N_9100,N_9105);
xnor U9127 (N_9127,N_9078,N_9093);
and U9128 (N_9128,N_9095,N_8961);
nand U9129 (N_9129,N_9090,N_9013);
xor U9130 (N_9130,N_8982,N_9116);
or U9131 (N_9131,N_9002,N_9083);
and U9132 (N_9132,N_8990,N_9033);
xor U9133 (N_9133,N_9055,N_8979);
or U9134 (N_9134,N_9005,N_9057);
nand U9135 (N_9135,N_9014,N_9106);
nand U9136 (N_9136,N_8998,N_9065);
nor U9137 (N_9137,N_9008,N_9081);
nor U9138 (N_9138,N_9023,N_9018);
xor U9139 (N_9139,N_9086,N_9034);
nand U9140 (N_9140,N_9104,N_9041);
nand U9141 (N_9141,N_9077,N_8993);
nand U9142 (N_9142,N_9056,N_9007);
nor U9143 (N_9143,N_8962,N_9028);
nand U9144 (N_9144,N_9042,N_8988);
nand U9145 (N_9145,N_9012,N_9068);
xnor U9146 (N_9146,N_8970,N_8984);
and U9147 (N_9147,N_9052,N_9109);
or U9148 (N_9148,N_8997,N_8985);
nand U9149 (N_9149,N_9072,N_9108);
xnor U9150 (N_9150,N_8986,N_9073);
nand U9151 (N_9151,N_9029,N_9017);
nor U9152 (N_9152,N_9020,N_9076);
xnor U9153 (N_9153,N_9080,N_9015);
nor U9154 (N_9154,N_9043,N_9091);
nor U9155 (N_9155,N_9038,N_9069);
nand U9156 (N_9156,N_9026,N_9046);
nand U9157 (N_9157,N_8992,N_8971);
xnor U9158 (N_9158,N_8963,N_9062);
xnor U9159 (N_9159,N_8977,N_9054);
or U9160 (N_9160,N_9044,N_8987);
nor U9161 (N_9161,N_9075,N_8983);
or U9162 (N_9162,N_9032,N_8995);
xnor U9163 (N_9163,N_9113,N_9067);
and U9164 (N_9164,N_9049,N_8981);
nor U9165 (N_9165,N_9074,N_8960);
nor U9166 (N_9166,N_9051,N_8966);
or U9167 (N_9167,N_9115,N_9117);
nand U9168 (N_9168,N_9101,N_9011);
and U9169 (N_9169,N_9006,N_9016);
and U9170 (N_9170,N_8973,N_9110);
or U9171 (N_9171,N_9022,N_9070);
and U9172 (N_9172,N_9060,N_9099);
nand U9173 (N_9173,N_9066,N_9050);
or U9174 (N_9174,N_9089,N_9084);
xnor U9175 (N_9175,N_9030,N_9061);
nor U9176 (N_9176,N_9001,N_8967);
nand U9177 (N_9177,N_9059,N_8991);
and U9178 (N_9178,N_8980,N_9000);
nor U9179 (N_9179,N_9021,N_8969);
nand U9180 (N_9180,N_9058,N_8976);
nor U9181 (N_9181,N_9071,N_8989);
nand U9182 (N_9182,N_9031,N_9027);
xor U9183 (N_9183,N_9092,N_9112);
or U9184 (N_9184,N_9039,N_9088);
and U9185 (N_9185,N_9111,N_9118);
nor U9186 (N_9186,N_9040,N_9096);
nand U9187 (N_9187,N_9036,N_9048);
nand U9188 (N_9188,N_9094,N_9035);
xnor U9189 (N_9189,N_9102,N_9063);
or U9190 (N_9190,N_8965,N_9053);
xor U9191 (N_9191,N_9010,N_8996);
nor U9192 (N_9192,N_9019,N_9079);
nand U9193 (N_9193,N_8974,N_9024);
xnor U9194 (N_9194,N_9103,N_9107);
nor U9195 (N_9195,N_9064,N_9047);
xor U9196 (N_9196,N_9087,N_9114);
nor U9197 (N_9197,N_9004,N_8964);
xor U9198 (N_9198,N_9037,N_9119);
or U9199 (N_9199,N_9025,N_8999);
or U9200 (N_9200,N_8960,N_9019);
xor U9201 (N_9201,N_9011,N_9092);
or U9202 (N_9202,N_9055,N_9099);
nor U9203 (N_9203,N_8965,N_9008);
and U9204 (N_9204,N_9050,N_9021);
and U9205 (N_9205,N_9053,N_9103);
nor U9206 (N_9206,N_9106,N_9094);
nand U9207 (N_9207,N_9089,N_9001);
and U9208 (N_9208,N_8964,N_9114);
xnor U9209 (N_9209,N_9037,N_9028);
xnor U9210 (N_9210,N_9058,N_8997);
and U9211 (N_9211,N_9067,N_9087);
or U9212 (N_9212,N_8997,N_8964);
nor U9213 (N_9213,N_9000,N_9078);
and U9214 (N_9214,N_9030,N_9074);
nor U9215 (N_9215,N_8977,N_9107);
or U9216 (N_9216,N_9028,N_9015);
nand U9217 (N_9217,N_9010,N_9070);
and U9218 (N_9218,N_9056,N_9082);
xnor U9219 (N_9219,N_8999,N_9009);
nor U9220 (N_9220,N_9038,N_9048);
or U9221 (N_9221,N_9086,N_9083);
xnor U9222 (N_9222,N_8960,N_9023);
or U9223 (N_9223,N_9040,N_9012);
nor U9224 (N_9224,N_9117,N_8996);
or U9225 (N_9225,N_9035,N_9026);
or U9226 (N_9226,N_8985,N_9059);
and U9227 (N_9227,N_9070,N_9068);
and U9228 (N_9228,N_9031,N_9000);
and U9229 (N_9229,N_9006,N_9068);
nand U9230 (N_9230,N_9108,N_9029);
xnor U9231 (N_9231,N_9078,N_9062);
nand U9232 (N_9232,N_9080,N_9044);
or U9233 (N_9233,N_9051,N_9013);
xnor U9234 (N_9234,N_8989,N_9056);
nand U9235 (N_9235,N_9076,N_9034);
or U9236 (N_9236,N_8999,N_9004);
xnor U9237 (N_9237,N_9069,N_9048);
nand U9238 (N_9238,N_8978,N_9019);
or U9239 (N_9239,N_8988,N_9057);
and U9240 (N_9240,N_9064,N_8962);
nand U9241 (N_9241,N_9097,N_8992);
nand U9242 (N_9242,N_8997,N_9095);
or U9243 (N_9243,N_9039,N_9083);
and U9244 (N_9244,N_9013,N_8977);
nor U9245 (N_9245,N_9081,N_9005);
xor U9246 (N_9246,N_9070,N_9013);
xnor U9247 (N_9247,N_8989,N_9086);
xnor U9248 (N_9248,N_9094,N_9075);
nor U9249 (N_9249,N_9113,N_9048);
nor U9250 (N_9250,N_9037,N_9014);
nor U9251 (N_9251,N_9027,N_9020);
nor U9252 (N_9252,N_9104,N_9076);
nand U9253 (N_9253,N_9084,N_9088);
or U9254 (N_9254,N_9002,N_9044);
nand U9255 (N_9255,N_9081,N_8985);
and U9256 (N_9256,N_9040,N_8980);
or U9257 (N_9257,N_9105,N_9073);
xor U9258 (N_9258,N_8994,N_8981);
and U9259 (N_9259,N_9087,N_9077);
or U9260 (N_9260,N_8994,N_9053);
nor U9261 (N_9261,N_9068,N_9058);
and U9262 (N_9262,N_9072,N_9110);
or U9263 (N_9263,N_8969,N_9053);
nand U9264 (N_9264,N_9082,N_9079);
nor U9265 (N_9265,N_9111,N_9025);
xnor U9266 (N_9266,N_9008,N_9023);
and U9267 (N_9267,N_8972,N_9011);
and U9268 (N_9268,N_9055,N_9024);
and U9269 (N_9269,N_9049,N_9078);
nand U9270 (N_9270,N_9008,N_9118);
and U9271 (N_9271,N_9051,N_9005);
and U9272 (N_9272,N_9071,N_8968);
and U9273 (N_9273,N_9110,N_9019);
nand U9274 (N_9274,N_8976,N_9012);
xnor U9275 (N_9275,N_9110,N_9117);
or U9276 (N_9276,N_9087,N_8982);
or U9277 (N_9277,N_8965,N_9101);
nand U9278 (N_9278,N_9113,N_9105);
nand U9279 (N_9279,N_9044,N_8968);
and U9280 (N_9280,N_9138,N_9206);
nor U9281 (N_9281,N_9229,N_9220);
nor U9282 (N_9282,N_9277,N_9241);
or U9283 (N_9283,N_9125,N_9208);
nor U9284 (N_9284,N_9195,N_9260);
and U9285 (N_9285,N_9197,N_9278);
nand U9286 (N_9286,N_9211,N_9154);
nor U9287 (N_9287,N_9198,N_9132);
xnor U9288 (N_9288,N_9262,N_9143);
xor U9289 (N_9289,N_9164,N_9237);
and U9290 (N_9290,N_9120,N_9231);
xnor U9291 (N_9291,N_9163,N_9140);
xor U9292 (N_9292,N_9236,N_9274);
and U9293 (N_9293,N_9235,N_9176);
nand U9294 (N_9294,N_9279,N_9142);
nor U9295 (N_9295,N_9127,N_9152);
and U9296 (N_9296,N_9203,N_9123);
nand U9297 (N_9297,N_9188,N_9253);
nor U9298 (N_9298,N_9190,N_9248);
xor U9299 (N_9299,N_9269,N_9160);
or U9300 (N_9300,N_9135,N_9240);
or U9301 (N_9301,N_9234,N_9146);
nor U9302 (N_9302,N_9230,N_9252);
xor U9303 (N_9303,N_9182,N_9162);
nand U9304 (N_9304,N_9180,N_9124);
or U9305 (N_9305,N_9187,N_9128);
or U9306 (N_9306,N_9157,N_9136);
nor U9307 (N_9307,N_9247,N_9225);
nor U9308 (N_9308,N_9226,N_9172);
xnor U9309 (N_9309,N_9168,N_9242);
or U9310 (N_9310,N_9199,N_9178);
xor U9311 (N_9311,N_9192,N_9181);
and U9312 (N_9312,N_9244,N_9175);
nor U9313 (N_9313,N_9141,N_9239);
nor U9314 (N_9314,N_9232,N_9272);
and U9315 (N_9315,N_9167,N_9243);
xor U9316 (N_9316,N_9270,N_9144);
nand U9317 (N_9317,N_9215,N_9165);
and U9318 (N_9318,N_9191,N_9149);
nand U9319 (N_9319,N_9122,N_9189);
nand U9320 (N_9320,N_9169,N_9256);
nor U9321 (N_9321,N_9201,N_9219);
nand U9322 (N_9322,N_9156,N_9202);
xnor U9323 (N_9323,N_9193,N_9261);
nand U9324 (N_9324,N_9158,N_9209);
nand U9325 (N_9325,N_9233,N_9151);
nand U9326 (N_9326,N_9216,N_9224);
and U9327 (N_9327,N_9258,N_9200);
and U9328 (N_9328,N_9223,N_9271);
xor U9329 (N_9329,N_9179,N_9121);
or U9330 (N_9330,N_9196,N_9266);
nor U9331 (N_9331,N_9155,N_9228);
and U9332 (N_9332,N_9177,N_9249);
nor U9333 (N_9333,N_9159,N_9254);
xnor U9334 (N_9334,N_9245,N_9130);
or U9335 (N_9335,N_9148,N_9227);
nor U9336 (N_9336,N_9133,N_9161);
nand U9337 (N_9337,N_9210,N_9218);
nand U9338 (N_9338,N_9250,N_9194);
or U9339 (N_9339,N_9263,N_9217);
xnor U9340 (N_9340,N_9273,N_9145);
nor U9341 (N_9341,N_9126,N_9212);
nand U9342 (N_9342,N_9222,N_9137);
or U9343 (N_9343,N_9153,N_9204);
xnor U9344 (N_9344,N_9257,N_9259);
and U9345 (N_9345,N_9183,N_9170);
xnor U9346 (N_9346,N_9166,N_9131);
xnor U9347 (N_9347,N_9276,N_9171);
and U9348 (N_9348,N_9214,N_9186);
nor U9349 (N_9349,N_9205,N_9174);
nor U9350 (N_9350,N_9251,N_9221);
xor U9351 (N_9351,N_9207,N_9147);
nor U9352 (N_9352,N_9134,N_9150);
nand U9353 (N_9353,N_9246,N_9255);
xor U9354 (N_9354,N_9264,N_9185);
and U9355 (N_9355,N_9265,N_9184);
xnor U9356 (N_9356,N_9129,N_9238);
nand U9357 (N_9357,N_9267,N_9139);
nor U9358 (N_9358,N_9268,N_9213);
nand U9359 (N_9359,N_9275,N_9173);
nand U9360 (N_9360,N_9182,N_9127);
xnor U9361 (N_9361,N_9226,N_9233);
nand U9362 (N_9362,N_9123,N_9183);
and U9363 (N_9363,N_9239,N_9165);
nor U9364 (N_9364,N_9255,N_9268);
or U9365 (N_9365,N_9174,N_9206);
xor U9366 (N_9366,N_9157,N_9279);
or U9367 (N_9367,N_9253,N_9270);
xnor U9368 (N_9368,N_9270,N_9250);
nand U9369 (N_9369,N_9251,N_9266);
and U9370 (N_9370,N_9199,N_9177);
xnor U9371 (N_9371,N_9234,N_9236);
or U9372 (N_9372,N_9151,N_9244);
and U9373 (N_9373,N_9259,N_9168);
xnor U9374 (N_9374,N_9244,N_9216);
or U9375 (N_9375,N_9220,N_9234);
nor U9376 (N_9376,N_9152,N_9190);
and U9377 (N_9377,N_9224,N_9264);
nand U9378 (N_9378,N_9136,N_9134);
or U9379 (N_9379,N_9148,N_9237);
xor U9380 (N_9380,N_9226,N_9237);
xor U9381 (N_9381,N_9195,N_9170);
nor U9382 (N_9382,N_9173,N_9124);
or U9383 (N_9383,N_9143,N_9243);
nor U9384 (N_9384,N_9250,N_9125);
or U9385 (N_9385,N_9144,N_9150);
and U9386 (N_9386,N_9266,N_9180);
nor U9387 (N_9387,N_9146,N_9141);
or U9388 (N_9388,N_9240,N_9151);
xnor U9389 (N_9389,N_9230,N_9183);
or U9390 (N_9390,N_9212,N_9173);
nor U9391 (N_9391,N_9182,N_9169);
nor U9392 (N_9392,N_9131,N_9188);
nand U9393 (N_9393,N_9231,N_9161);
xnor U9394 (N_9394,N_9162,N_9214);
or U9395 (N_9395,N_9187,N_9150);
nor U9396 (N_9396,N_9194,N_9197);
xnor U9397 (N_9397,N_9277,N_9207);
nor U9398 (N_9398,N_9160,N_9178);
xnor U9399 (N_9399,N_9238,N_9214);
nor U9400 (N_9400,N_9223,N_9181);
xor U9401 (N_9401,N_9249,N_9159);
nand U9402 (N_9402,N_9274,N_9211);
and U9403 (N_9403,N_9152,N_9177);
nor U9404 (N_9404,N_9221,N_9228);
and U9405 (N_9405,N_9155,N_9186);
nand U9406 (N_9406,N_9125,N_9145);
nor U9407 (N_9407,N_9205,N_9259);
nand U9408 (N_9408,N_9184,N_9192);
nand U9409 (N_9409,N_9251,N_9172);
xor U9410 (N_9410,N_9221,N_9197);
and U9411 (N_9411,N_9144,N_9131);
nand U9412 (N_9412,N_9180,N_9232);
or U9413 (N_9413,N_9159,N_9192);
and U9414 (N_9414,N_9178,N_9187);
or U9415 (N_9415,N_9248,N_9125);
nor U9416 (N_9416,N_9204,N_9159);
or U9417 (N_9417,N_9216,N_9152);
and U9418 (N_9418,N_9212,N_9236);
xnor U9419 (N_9419,N_9255,N_9216);
or U9420 (N_9420,N_9174,N_9197);
and U9421 (N_9421,N_9258,N_9202);
nor U9422 (N_9422,N_9274,N_9209);
nor U9423 (N_9423,N_9242,N_9136);
nand U9424 (N_9424,N_9254,N_9123);
nand U9425 (N_9425,N_9232,N_9255);
and U9426 (N_9426,N_9277,N_9124);
nor U9427 (N_9427,N_9275,N_9154);
nor U9428 (N_9428,N_9161,N_9175);
and U9429 (N_9429,N_9204,N_9165);
xor U9430 (N_9430,N_9208,N_9209);
xor U9431 (N_9431,N_9209,N_9178);
nand U9432 (N_9432,N_9169,N_9167);
and U9433 (N_9433,N_9131,N_9253);
nand U9434 (N_9434,N_9186,N_9128);
and U9435 (N_9435,N_9131,N_9150);
or U9436 (N_9436,N_9212,N_9195);
or U9437 (N_9437,N_9262,N_9157);
nor U9438 (N_9438,N_9122,N_9180);
nand U9439 (N_9439,N_9225,N_9193);
nor U9440 (N_9440,N_9315,N_9360);
and U9441 (N_9441,N_9397,N_9425);
nand U9442 (N_9442,N_9293,N_9319);
and U9443 (N_9443,N_9332,N_9282);
xor U9444 (N_9444,N_9409,N_9426);
nor U9445 (N_9445,N_9393,N_9390);
nand U9446 (N_9446,N_9311,N_9297);
and U9447 (N_9447,N_9404,N_9334);
or U9448 (N_9448,N_9417,N_9364);
and U9449 (N_9449,N_9400,N_9370);
nor U9450 (N_9450,N_9424,N_9321);
xor U9451 (N_9451,N_9378,N_9421);
xor U9452 (N_9452,N_9356,N_9423);
nor U9453 (N_9453,N_9304,N_9434);
xor U9454 (N_9454,N_9373,N_9392);
xnor U9455 (N_9455,N_9386,N_9317);
or U9456 (N_9456,N_9388,N_9380);
xnor U9457 (N_9457,N_9318,N_9344);
or U9458 (N_9458,N_9357,N_9303);
xor U9459 (N_9459,N_9292,N_9310);
nand U9460 (N_9460,N_9377,N_9411);
or U9461 (N_9461,N_9387,N_9384);
and U9462 (N_9462,N_9432,N_9312);
nor U9463 (N_9463,N_9306,N_9322);
or U9464 (N_9464,N_9340,N_9412);
nor U9465 (N_9465,N_9283,N_9428);
xor U9466 (N_9466,N_9301,N_9307);
xor U9467 (N_9467,N_9420,N_9399);
and U9468 (N_9468,N_9398,N_9294);
or U9469 (N_9469,N_9338,N_9427);
or U9470 (N_9470,N_9381,N_9407);
nor U9471 (N_9471,N_9406,N_9359);
and U9472 (N_9472,N_9413,N_9436);
nor U9473 (N_9473,N_9401,N_9410);
and U9474 (N_9474,N_9365,N_9350);
or U9475 (N_9475,N_9419,N_9366);
nor U9476 (N_9476,N_9362,N_9439);
and U9477 (N_9477,N_9438,N_9351);
nand U9478 (N_9478,N_9313,N_9382);
nand U9479 (N_9479,N_9352,N_9355);
nand U9480 (N_9480,N_9309,N_9349);
nor U9481 (N_9481,N_9302,N_9323);
xnor U9482 (N_9482,N_9363,N_9286);
or U9483 (N_9483,N_9358,N_9375);
xnor U9484 (N_9484,N_9314,N_9422);
nand U9485 (N_9485,N_9374,N_9430);
xor U9486 (N_9486,N_9339,N_9371);
and U9487 (N_9487,N_9433,N_9284);
xor U9488 (N_9488,N_9348,N_9431);
nand U9489 (N_9489,N_9330,N_9394);
and U9490 (N_9490,N_9345,N_9300);
nor U9491 (N_9491,N_9368,N_9408);
and U9492 (N_9492,N_9435,N_9395);
and U9493 (N_9493,N_9403,N_9379);
and U9494 (N_9494,N_9429,N_9324);
xnor U9495 (N_9495,N_9287,N_9316);
or U9496 (N_9496,N_9320,N_9329);
nor U9497 (N_9497,N_9291,N_9347);
and U9498 (N_9498,N_9369,N_9396);
xor U9499 (N_9499,N_9353,N_9372);
or U9500 (N_9500,N_9326,N_9325);
xor U9501 (N_9501,N_9346,N_9289);
xnor U9502 (N_9502,N_9361,N_9288);
and U9503 (N_9503,N_9333,N_9336);
and U9504 (N_9504,N_9437,N_9299);
or U9505 (N_9505,N_9414,N_9389);
or U9506 (N_9506,N_9415,N_9327);
xnor U9507 (N_9507,N_9298,N_9376);
or U9508 (N_9508,N_9418,N_9337);
nand U9509 (N_9509,N_9308,N_9296);
xnor U9510 (N_9510,N_9343,N_9285);
or U9511 (N_9511,N_9335,N_9354);
xor U9512 (N_9512,N_9341,N_9290);
or U9513 (N_9513,N_9328,N_9367);
nand U9514 (N_9514,N_9295,N_9402);
and U9515 (N_9515,N_9405,N_9416);
and U9516 (N_9516,N_9342,N_9305);
or U9517 (N_9517,N_9391,N_9383);
nor U9518 (N_9518,N_9280,N_9331);
nor U9519 (N_9519,N_9281,N_9385);
and U9520 (N_9520,N_9368,N_9358);
nor U9521 (N_9521,N_9307,N_9382);
xnor U9522 (N_9522,N_9343,N_9342);
or U9523 (N_9523,N_9395,N_9437);
nor U9524 (N_9524,N_9283,N_9390);
xnor U9525 (N_9525,N_9362,N_9416);
xor U9526 (N_9526,N_9435,N_9342);
and U9527 (N_9527,N_9318,N_9365);
nor U9528 (N_9528,N_9366,N_9360);
nor U9529 (N_9529,N_9305,N_9391);
and U9530 (N_9530,N_9303,N_9300);
or U9531 (N_9531,N_9399,N_9346);
or U9532 (N_9532,N_9362,N_9389);
and U9533 (N_9533,N_9427,N_9327);
and U9534 (N_9534,N_9421,N_9361);
nor U9535 (N_9535,N_9357,N_9405);
xor U9536 (N_9536,N_9387,N_9430);
nor U9537 (N_9537,N_9320,N_9369);
nor U9538 (N_9538,N_9395,N_9411);
xor U9539 (N_9539,N_9421,N_9381);
or U9540 (N_9540,N_9298,N_9396);
xor U9541 (N_9541,N_9311,N_9350);
nand U9542 (N_9542,N_9374,N_9313);
nand U9543 (N_9543,N_9388,N_9327);
nor U9544 (N_9544,N_9430,N_9366);
nor U9545 (N_9545,N_9417,N_9360);
xnor U9546 (N_9546,N_9308,N_9303);
or U9547 (N_9547,N_9300,N_9396);
and U9548 (N_9548,N_9414,N_9439);
nand U9549 (N_9549,N_9339,N_9439);
or U9550 (N_9550,N_9371,N_9394);
nand U9551 (N_9551,N_9391,N_9318);
nor U9552 (N_9552,N_9288,N_9387);
or U9553 (N_9553,N_9393,N_9435);
and U9554 (N_9554,N_9403,N_9336);
and U9555 (N_9555,N_9286,N_9288);
nor U9556 (N_9556,N_9357,N_9412);
xor U9557 (N_9557,N_9338,N_9390);
nor U9558 (N_9558,N_9307,N_9385);
xnor U9559 (N_9559,N_9426,N_9388);
and U9560 (N_9560,N_9383,N_9335);
and U9561 (N_9561,N_9282,N_9384);
and U9562 (N_9562,N_9345,N_9285);
and U9563 (N_9563,N_9412,N_9333);
and U9564 (N_9564,N_9315,N_9409);
nand U9565 (N_9565,N_9353,N_9405);
and U9566 (N_9566,N_9349,N_9358);
xor U9567 (N_9567,N_9308,N_9426);
nor U9568 (N_9568,N_9380,N_9300);
xnor U9569 (N_9569,N_9372,N_9306);
xnor U9570 (N_9570,N_9390,N_9408);
xnor U9571 (N_9571,N_9394,N_9396);
xnor U9572 (N_9572,N_9380,N_9308);
nand U9573 (N_9573,N_9346,N_9324);
nor U9574 (N_9574,N_9416,N_9352);
xor U9575 (N_9575,N_9282,N_9292);
nand U9576 (N_9576,N_9350,N_9308);
nor U9577 (N_9577,N_9345,N_9342);
nor U9578 (N_9578,N_9395,N_9335);
nor U9579 (N_9579,N_9325,N_9294);
nor U9580 (N_9580,N_9365,N_9302);
nor U9581 (N_9581,N_9379,N_9391);
nor U9582 (N_9582,N_9361,N_9357);
or U9583 (N_9583,N_9333,N_9433);
xor U9584 (N_9584,N_9384,N_9330);
nor U9585 (N_9585,N_9399,N_9324);
nand U9586 (N_9586,N_9321,N_9397);
nor U9587 (N_9587,N_9394,N_9339);
and U9588 (N_9588,N_9353,N_9282);
nor U9589 (N_9589,N_9311,N_9285);
and U9590 (N_9590,N_9434,N_9343);
or U9591 (N_9591,N_9347,N_9327);
xor U9592 (N_9592,N_9294,N_9317);
nand U9593 (N_9593,N_9282,N_9336);
or U9594 (N_9594,N_9364,N_9322);
nand U9595 (N_9595,N_9290,N_9319);
nand U9596 (N_9596,N_9329,N_9348);
nor U9597 (N_9597,N_9390,N_9422);
nor U9598 (N_9598,N_9376,N_9354);
nand U9599 (N_9599,N_9425,N_9378);
and U9600 (N_9600,N_9538,N_9467);
xnor U9601 (N_9601,N_9461,N_9471);
and U9602 (N_9602,N_9591,N_9553);
and U9603 (N_9603,N_9491,N_9457);
nand U9604 (N_9604,N_9589,N_9545);
nand U9605 (N_9605,N_9513,N_9597);
xor U9606 (N_9606,N_9547,N_9444);
xnor U9607 (N_9607,N_9478,N_9494);
and U9608 (N_9608,N_9532,N_9537);
or U9609 (N_9609,N_9512,N_9511);
xnor U9610 (N_9610,N_9558,N_9463);
nand U9611 (N_9611,N_9448,N_9507);
xnor U9612 (N_9612,N_9549,N_9498);
xor U9613 (N_9613,N_9514,N_9524);
nor U9614 (N_9614,N_9470,N_9529);
and U9615 (N_9615,N_9520,N_9517);
nor U9616 (N_9616,N_9590,N_9446);
xnor U9617 (N_9617,N_9577,N_9581);
or U9618 (N_9618,N_9540,N_9550);
nand U9619 (N_9619,N_9502,N_9447);
nand U9620 (N_9620,N_9489,N_9536);
nor U9621 (N_9621,N_9587,N_9556);
or U9622 (N_9622,N_9569,N_9533);
and U9623 (N_9623,N_9560,N_9506);
and U9624 (N_9624,N_9563,N_9504);
or U9625 (N_9625,N_9598,N_9440);
xor U9626 (N_9626,N_9528,N_9466);
xnor U9627 (N_9627,N_9501,N_9499);
nand U9628 (N_9628,N_9573,N_9548);
and U9629 (N_9629,N_9594,N_9472);
nor U9630 (N_9630,N_9441,N_9580);
or U9631 (N_9631,N_9542,N_9454);
xnor U9632 (N_9632,N_9488,N_9572);
xnor U9633 (N_9633,N_9571,N_9453);
nand U9634 (N_9634,N_9493,N_9552);
nor U9635 (N_9635,N_9445,N_9481);
nor U9636 (N_9636,N_9592,N_9442);
nor U9637 (N_9637,N_9518,N_9588);
and U9638 (N_9638,N_9450,N_9586);
or U9639 (N_9639,N_9460,N_9585);
xnor U9640 (N_9640,N_9599,N_9530);
nand U9641 (N_9641,N_9557,N_9566);
and U9642 (N_9642,N_9579,N_9508);
nor U9643 (N_9643,N_9469,N_9593);
and U9644 (N_9644,N_9495,N_9525);
or U9645 (N_9645,N_9531,N_9468);
xnor U9646 (N_9646,N_9459,N_9496);
and U9647 (N_9647,N_9465,N_9564);
or U9648 (N_9648,N_9596,N_9497);
xor U9649 (N_9649,N_9568,N_9526);
or U9650 (N_9650,N_9551,N_9474);
xor U9651 (N_9651,N_9559,N_9522);
nand U9652 (N_9652,N_9455,N_9595);
nor U9653 (N_9653,N_9503,N_9574);
and U9654 (N_9654,N_9487,N_9578);
or U9655 (N_9655,N_9484,N_9541);
nand U9656 (N_9656,N_9544,N_9443);
nor U9657 (N_9657,N_9485,N_9554);
or U9658 (N_9658,N_9575,N_9539);
and U9659 (N_9659,N_9546,N_9482);
nand U9660 (N_9660,N_9500,N_9521);
nand U9661 (N_9661,N_9583,N_9458);
nand U9662 (N_9662,N_9505,N_9555);
and U9663 (N_9663,N_9476,N_9567);
xnor U9664 (N_9664,N_9473,N_9543);
nand U9665 (N_9665,N_9535,N_9519);
or U9666 (N_9666,N_9534,N_9490);
nor U9667 (N_9667,N_9527,N_9449);
and U9668 (N_9668,N_9582,N_9584);
xnor U9669 (N_9669,N_9486,N_9576);
xnor U9670 (N_9670,N_9452,N_9456);
nor U9671 (N_9671,N_9570,N_9462);
nor U9672 (N_9672,N_9516,N_9483);
nor U9673 (N_9673,N_9510,N_9523);
or U9674 (N_9674,N_9451,N_9477);
or U9675 (N_9675,N_9480,N_9509);
xor U9676 (N_9676,N_9479,N_9464);
xor U9677 (N_9677,N_9562,N_9475);
or U9678 (N_9678,N_9561,N_9515);
nor U9679 (N_9679,N_9492,N_9565);
nor U9680 (N_9680,N_9518,N_9536);
nor U9681 (N_9681,N_9574,N_9544);
xor U9682 (N_9682,N_9522,N_9593);
nor U9683 (N_9683,N_9463,N_9440);
and U9684 (N_9684,N_9476,N_9504);
nand U9685 (N_9685,N_9464,N_9457);
and U9686 (N_9686,N_9508,N_9460);
or U9687 (N_9687,N_9555,N_9474);
nor U9688 (N_9688,N_9591,N_9530);
xnor U9689 (N_9689,N_9596,N_9460);
or U9690 (N_9690,N_9590,N_9523);
xnor U9691 (N_9691,N_9595,N_9486);
nor U9692 (N_9692,N_9547,N_9584);
xnor U9693 (N_9693,N_9583,N_9562);
or U9694 (N_9694,N_9544,N_9474);
xnor U9695 (N_9695,N_9480,N_9470);
nand U9696 (N_9696,N_9522,N_9471);
or U9697 (N_9697,N_9557,N_9501);
nor U9698 (N_9698,N_9561,N_9548);
nand U9699 (N_9699,N_9545,N_9541);
nor U9700 (N_9700,N_9547,N_9450);
and U9701 (N_9701,N_9498,N_9585);
xor U9702 (N_9702,N_9510,N_9558);
xor U9703 (N_9703,N_9520,N_9440);
nor U9704 (N_9704,N_9530,N_9587);
or U9705 (N_9705,N_9483,N_9459);
nor U9706 (N_9706,N_9562,N_9510);
or U9707 (N_9707,N_9514,N_9444);
nor U9708 (N_9708,N_9513,N_9444);
nand U9709 (N_9709,N_9476,N_9453);
nor U9710 (N_9710,N_9575,N_9489);
or U9711 (N_9711,N_9484,N_9576);
nor U9712 (N_9712,N_9506,N_9477);
nor U9713 (N_9713,N_9505,N_9519);
nand U9714 (N_9714,N_9517,N_9538);
or U9715 (N_9715,N_9483,N_9449);
xor U9716 (N_9716,N_9478,N_9450);
or U9717 (N_9717,N_9546,N_9458);
and U9718 (N_9718,N_9461,N_9587);
xor U9719 (N_9719,N_9595,N_9556);
nand U9720 (N_9720,N_9560,N_9566);
nand U9721 (N_9721,N_9523,N_9448);
nand U9722 (N_9722,N_9511,N_9581);
and U9723 (N_9723,N_9449,N_9532);
or U9724 (N_9724,N_9537,N_9445);
nor U9725 (N_9725,N_9534,N_9515);
xnor U9726 (N_9726,N_9440,N_9590);
and U9727 (N_9727,N_9534,N_9460);
nor U9728 (N_9728,N_9522,N_9577);
nand U9729 (N_9729,N_9593,N_9470);
nand U9730 (N_9730,N_9457,N_9463);
xnor U9731 (N_9731,N_9597,N_9487);
and U9732 (N_9732,N_9568,N_9469);
nor U9733 (N_9733,N_9518,N_9599);
nor U9734 (N_9734,N_9579,N_9454);
nand U9735 (N_9735,N_9448,N_9566);
nand U9736 (N_9736,N_9502,N_9570);
or U9737 (N_9737,N_9455,N_9545);
or U9738 (N_9738,N_9521,N_9587);
nand U9739 (N_9739,N_9483,N_9524);
or U9740 (N_9740,N_9504,N_9522);
nor U9741 (N_9741,N_9455,N_9567);
or U9742 (N_9742,N_9465,N_9575);
nor U9743 (N_9743,N_9571,N_9474);
and U9744 (N_9744,N_9558,N_9585);
or U9745 (N_9745,N_9548,N_9522);
nand U9746 (N_9746,N_9597,N_9464);
xnor U9747 (N_9747,N_9583,N_9545);
and U9748 (N_9748,N_9584,N_9451);
nand U9749 (N_9749,N_9484,N_9477);
nor U9750 (N_9750,N_9594,N_9557);
and U9751 (N_9751,N_9462,N_9457);
or U9752 (N_9752,N_9475,N_9478);
xor U9753 (N_9753,N_9482,N_9477);
and U9754 (N_9754,N_9513,N_9512);
and U9755 (N_9755,N_9523,N_9466);
and U9756 (N_9756,N_9467,N_9570);
and U9757 (N_9757,N_9517,N_9586);
nor U9758 (N_9758,N_9585,N_9522);
xnor U9759 (N_9759,N_9577,N_9540);
or U9760 (N_9760,N_9631,N_9742);
and U9761 (N_9761,N_9601,N_9643);
or U9762 (N_9762,N_9620,N_9730);
xnor U9763 (N_9763,N_9659,N_9625);
nor U9764 (N_9764,N_9663,N_9606);
nand U9765 (N_9765,N_9657,N_9682);
or U9766 (N_9766,N_9607,N_9621);
nor U9767 (N_9767,N_9691,N_9604);
nor U9768 (N_9768,N_9751,N_9628);
or U9769 (N_9769,N_9603,N_9616);
nand U9770 (N_9770,N_9677,N_9695);
xor U9771 (N_9771,N_9684,N_9726);
xnor U9772 (N_9772,N_9735,N_9623);
nor U9773 (N_9773,N_9741,N_9750);
or U9774 (N_9774,N_9727,N_9674);
or U9775 (N_9775,N_9755,N_9634);
or U9776 (N_9776,N_9715,N_9708);
and U9777 (N_9777,N_9645,N_9641);
and U9778 (N_9778,N_9738,N_9692);
and U9779 (N_9779,N_9748,N_9629);
xor U9780 (N_9780,N_9752,N_9700);
nand U9781 (N_9781,N_9729,N_9679);
or U9782 (N_9782,N_9626,N_9611);
nor U9783 (N_9783,N_9705,N_9711);
nor U9784 (N_9784,N_9732,N_9608);
xnor U9785 (N_9785,N_9714,N_9671);
nor U9786 (N_9786,N_9661,N_9668);
xnor U9787 (N_9787,N_9736,N_9644);
or U9788 (N_9788,N_9722,N_9652);
nand U9789 (N_9789,N_9747,N_9651);
or U9790 (N_9790,N_9706,N_9737);
nor U9791 (N_9791,N_9709,N_9694);
and U9792 (N_9792,N_9753,N_9724);
and U9793 (N_9793,N_9609,N_9749);
nand U9794 (N_9794,N_9710,N_9685);
or U9795 (N_9795,N_9669,N_9618);
or U9796 (N_9796,N_9642,N_9624);
nor U9797 (N_9797,N_9719,N_9615);
xor U9798 (N_9798,N_9600,N_9648);
or U9799 (N_9799,N_9758,N_9650);
nor U9800 (N_9800,N_9656,N_9658);
and U9801 (N_9801,N_9731,N_9639);
nand U9802 (N_9802,N_9687,N_9667);
and U9803 (N_9803,N_9712,N_9720);
or U9804 (N_9804,N_9632,N_9713);
xnor U9805 (N_9805,N_9745,N_9670);
nand U9806 (N_9806,N_9665,N_9686);
nor U9807 (N_9807,N_9740,N_9699);
and U9808 (N_9808,N_9718,N_9683);
nand U9809 (N_9809,N_9637,N_9614);
xor U9810 (N_9810,N_9676,N_9734);
nand U9811 (N_9811,N_9690,N_9653);
or U9812 (N_9812,N_9757,N_9759);
or U9813 (N_9813,N_9696,N_9630);
xnor U9814 (N_9814,N_9617,N_9725);
nor U9815 (N_9815,N_9647,N_9743);
or U9816 (N_9816,N_9664,N_9716);
or U9817 (N_9817,N_9633,N_9612);
or U9818 (N_9818,N_9649,N_9754);
nand U9819 (N_9819,N_9689,N_9646);
and U9820 (N_9820,N_9602,N_9635);
nor U9821 (N_9821,N_9680,N_9638);
nor U9822 (N_9822,N_9640,N_9688);
nor U9823 (N_9823,N_9655,N_9654);
nor U9824 (N_9824,N_9666,N_9707);
and U9825 (N_9825,N_9756,N_9627);
and U9826 (N_9826,N_9610,N_9673);
nor U9827 (N_9827,N_9739,N_9703);
and U9828 (N_9828,N_9701,N_9723);
xor U9829 (N_9829,N_9721,N_9681);
nor U9830 (N_9830,N_9717,N_9613);
nor U9831 (N_9831,N_9744,N_9702);
or U9832 (N_9832,N_9698,N_9697);
and U9833 (N_9833,N_9678,N_9672);
nor U9834 (N_9834,N_9622,N_9704);
xnor U9835 (N_9835,N_9660,N_9733);
nor U9836 (N_9836,N_9693,N_9636);
or U9837 (N_9837,N_9675,N_9728);
and U9838 (N_9838,N_9605,N_9619);
xor U9839 (N_9839,N_9746,N_9662);
or U9840 (N_9840,N_9741,N_9755);
nand U9841 (N_9841,N_9626,N_9714);
or U9842 (N_9842,N_9607,N_9616);
nor U9843 (N_9843,N_9721,N_9658);
xor U9844 (N_9844,N_9738,N_9601);
and U9845 (N_9845,N_9698,N_9691);
nor U9846 (N_9846,N_9754,N_9733);
and U9847 (N_9847,N_9738,N_9743);
xnor U9848 (N_9848,N_9695,N_9748);
or U9849 (N_9849,N_9652,N_9744);
xor U9850 (N_9850,N_9639,N_9626);
xnor U9851 (N_9851,N_9614,N_9733);
nor U9852 (N_9852,N_9653,N_9737);
nor U9853 (N_9853,N_9745,N_9759);
nor U9854 (N_9854,N_9741,N_9600);
nand U9855 (N_9855,N_9678,N_9606);
xor U9856 (N_9856,N_9686,N_9618);
nand U9857 (N_9857,N_9691,N_9608);
and U9858 (N_9858,N_9606,N_9699);
or U9859 (N_9859,N_9699,N_9621);
nor U9860 (N_9860,N_9678,N_9630);
xor U9861 (N_9861,N_9609,N_9666);
xnor U9862 (N_9862,N_9602,N_9688);
or U9863 (N_9863,N_9736,N_9757);
nor U9864 (N_9864,N_9719,N_9728);
nand U9865 (N_9865,N_9602,N_9756);
or U9866 (N_9866,N_9632,N_9625);
nand U9867 (N_9867,N_9673,N_9682);
nor U9868 (N_9868,N_9619,N_9685);
or U9869 (N_9869,N_9662,N_9702);
nor U9870 (N_9870,N_9724,N_9676);
or U9871 (N_9871,N_9620,N_9722);
or U9872 (N_9872,N_9677,N_9647);
and U9873 (N_9873,N_9655,N_9662);
nand U9874 (N_9874,N_9722,N_9732);
or U9875 (N_9875,N_9660,N_9730);
xor U9876 (N_9876,N_9658,N_9672);
and U9877 (N_9877,N_9709,N_9748);
and U9878 (N_9878,N_9646,N_9626);
nand U9879 (N_9879,N_9727,N_9755);
nor U9880 (N_9880,N_9744,N_9669);
xor U9881 (N_9881,N_9615,N_9685);
and U9882 (N_9882,N_9661,N_9739);
and U9883 (N_9883,N_9673,N_9660);
or U9884 (N_9884,N_9747,N_9606);
xor U9885 (N_9885,N_9683,N_9679);
or U9886 (N_9886,N_9755,N_9664);
nor U9887 (N_9887,N_9610,N_9637);
nand U9888 (N_9888,N_9628,N_9724);
and U9889 (N_9889,N_9661,N_9730);
or U9890 (N_9890,N_9643,N_9714);
and U9891 (N_9891,N_9710,N_9688);
or U9892 (N_9892,N_9686,N_9663);
nor U9893 (N_9893,N_9699,N_9716);
nor U9894 (N_9894,N_9750,N_9632);
nand U9895 (N_9895,N_9628,N_9758);
nand U9896 (N_9896,N_9648,N_9660);
nand U9897 (N_9897,N_9635,N_9679);
nand U9898 (N_9898,N_9671,N_9651);
xor U9899 (N_9899,N_9667,N_9712);
nor U9900 (N_9900,N_9670,N_9625);
xor U9901 (N_9901,N_9696,N_9636);
or U9902 (N_9902,N_9617,N_9758);
or U9903 (N_9903,N_9757,N_9604);
or U9904 (N_9904,N_9743,N_9650);
and U9905 (N_9905,N_9648,N_9646);
nor U9906 (N_9906,N_9611,N_9699);
nand U9907 (N_9907,N_9628,N_9612);
or U9908 (N_9908,N_9740,N_9621);
xnor U9909 (N_9909,N_9666,N_9675);
nor U9910 (N_9910,N_9671,N_9748);
xor U9911 (N_9911,N_9701,N_9647);
xnor U9912 (N_9912,N_9703,N_9728);
and U9913 (N_9913,N_9605,N_9675);
and U9914 (N_9914,N_9641,N_9665);
xnor U9915 (N_9915,N_9754,N_9751);
nand U9916 (N_9916,N_9674,N_9621);
or U9917 (N_9917,N_9696,N_9715);
xor U9918 (N_9918,N_9659,N_9613);
or U9919 (N_9919,N_9755,N_9747);
and U9920 (N_9920,N_9812,N_9770);
or U9921 (N_9921,N_9918,N_9876);
nor U9922 (N_9922,N_9909,N_9878);
or U9923 (N_9923,N_9892,N_9877);
nand U9924 (N_9924,N_9888,N_9788);
or U9925 (N_9925,N_9791,N_9882);
and U9926 (N_9926,N_9919,N_9911);
nand U9927 (N_9927,N_9836,N_9815);
nand U9928 (N_9928,N_9852,N_9845);
xor U9929 (N_9929,N_9792,N_9841);
and U9930 (N_9930,N_9829,N_9903);
and U9931 (N_9931,N_9899,N_9783);
xnor U9932 (N_9932,N_9779,N_9814);
xnor U9933 (N_9933,N_9912,N_9823);
or U9934 (N_9934,N_9794,N_9879);
nor U9935 (N_9935,N_9799,N_9910);
nor U9936 (N_9936,N_9835,N_9828);
or U9937 (N_9937,N_9802,N_9913);
and U9938 (N_9938,N_9781,N_9874);
xor U9939 (N_9939,N_9858,N_9824);
xor U9940 (N_9940,N_9797,N_9895);
xnor U9941 (N_9941,N_9864,N_9855);
and U9942 (N_9942,N_9856,N_9796);
or U9943 (N_9943,N_9851,N_9771);
and U9944 (N_9944,N_9847,N_9793);
and U9945 (N_9945,N_9893,N_9857);
nand U9946 (N_9946,N_9904,N_9880);
xor U9947 (N_9947,N_9822,N_9811);
nor U9948 (N_9948,N_9780,N_9839);
xor U9949 (N_9949,N_9821,N_9804);
or U9950 (N_9950,N_9827,N_9833);
xnor U9951 (N_9951,N_9881,N_9891);
nor U9952 (N_9952,N_9782,N_9831);
xor U9953 (N_9953,N_9901,N_9898);
nand U9954 (N_9954,N_9889,N_9907);
xor U9955 (N_9955,N_9848,N_9817);
xor U9956 (N_9956,N_9885,N_9853);
and U9957 (N_9957,N_9768,N_9832);
nand U9958 (N_9958,N_9860,N_9830);
nand U9959 (N_9959,N_9764,N_9834);
nor U9960 (N_9960,N_9837,N_9862);
and U9961 (N_9961,N_9813,N_9766);
and U9962 (N_9962,N_9820,N_9914);
or U9963 (N_9963,N_9865,N_9850);
and U9964 (N_9964,N_9777,N_9803);
and U9965 (N_9965,N_9840,N_9810);
or U9966 (N_9966,N_9897,N_9890);
nand U9967 (N_9967,N_9775,N_9884);
nor U9968 (N_9968,N_9762,N_9805);
xor U9969 (N_9969,N_9763,N_9808);
and U9970 (N_9970,N_9786,N_9867);
or U9971 (N_9971,N_9859,N_9844);
nand U9972 (N_9972,N_9789,N_9769);
or U9973 (N_9973,N_9846,N_9870);
xor U9974 (N_9974,N_9798,N_9790);
nor U9975 (N_9975,N_9787,N_9871);
or U9976 (N_9976,N_9869,N_9816);
and U9977 (N_9977,N_9806,N_9905);
nand U9978 (N_9978,N_9887,N_9801);
or U9979 (N_9979,N_9906,N_9886);
and U9980 (N_9980,N_9826,N_9875);
xor U9981 (N_9981,N_9917,N_9785);
nor U9982 (N_9982,N_9773,N_9854);
and U9983 (N_9983,N_9795,N_9776);
nor U9984 (N_9984,N_9778,N_9761);
xor U9985 (N_9985,N_9863,N_9873);
or U9986 (N_9986,N_9915,N_9843);
or U9987 (N_9987,N_9772,N_9916);
and U9988 (N_9988,N_9894,N_9861);
xor U9989 (N_9989,N_9849,N_9809);
xnor U9990 (N_9990,N_9765,N_9818);
nand U9991 (N_9991,N_9838,N_9868);
nor U9992 (N_9992,N_9842,N_9784);
xor U9993 (N_9993,N_9883,N_9902);
xnor U9994 (N_9994,N_9900,N_9866);
and U9995 (N_9995,N_9825,N_9774);
and U9996 (N_9996,N_9760,N_9908);
or U9997 (N_9997,N_9767,N_9819);
nand U9998 (N_9998,N_9896,N_9800);
xnor U9999 (N_9999,N_9807,N_9872);
or U10000 (N_10000,N_9839,N_9861);
or U10001 (N_10001,N_9883,N_9800);
xor U10002 (N_10002,N_9878,N_9888);
nor U10003 (N_10003,N_9831,N_9879);
and U10004 (N_10004,N_9873,N_9796);
xnor U10005 (N_10005,N_9917,N_9795);
xor U10006 (N_10006,N_9762,N_9883);
and U10007 (N_10007,N_9775,N_9877);
and U10008 (N_10008,N_9876,N_9799);
nand U10009 (N_10009,N_9763,N_9820);
and U10010 (N_10010,N_9839,N_9870);
xor U10011 (N_10011,N_9760,N_9779);
or U10012 (N_10012,N_9880,N_9839);
nor U10013 (N_10013,N_9899,N_9792);
or U10014 (N_10014,N_9916,N_9895);
and U10015 (N_10015,N_9877,N_9867);
xnor U10016 (N_10016,N_9794,N_9914);
nand U10017 (N_10017,N_9859,N_9826);
nor U10018 (N_10018,N_9794,N_9906);
and U10019 (N_10019,N_9859,N_9916);
or U10020 (N_10020,N_9770,N_9912);
or U10021 (N_10021,N_9905,N_9836);
nor U10022 (N_10022,N_9833,N_9811);
nor U10023 (N_10023,N_9871,N_9840);
nor U10024 (N_10024,N_9844,N_9898);
xnor U10025 (N_10025,N_9848,N_9768);
or U10026 (N_10026,N_9904,N_9898);
nand U10027 (N_10027,N_9918,N_9837);
xnor U10028 (N_10028,N_9766,N_9872);
and U10029 (N_10029,N_9809,N_9817);
and U10030 (N_10030,N_9822,N_9825);
or U10031 (N_10031,N_9861,N_9911);
xor U10032 (N_10032,N_9809,N_9816);
xor U10033 (N_10033,N_9793,N_9892);
xor U10034 (N_10034,N_9901,N_9845);
xor U10035 (N_10035,N_9900,N_9811);
or U10036 (N_10036,N_9821,N_9780);
xor U10037 (N_10037,N_9821,N_9850);
and U10038 (N_10038,N_9832,N_9780);
nor U10039 (N_10039,N_9812,N_9791);
nand U10040 (N_10040,N_9792,N_9867);
nor U10041 (N_10041,N_9766,N_9769);
nor U10042 (N_10042,N_9802,N_9839);
or U10043 (N_10043,N_9870,N_9783);
or U10044 (N_10044,N_9907,N_9819);
or U10045 (N_10045,N_9818,N_9899);
xnor U10046 (N_10046,N_9822,N_9799);
xor U10047 (N_10047,N_9871,N_9875);
or U10048 (N_10048,N_9785,N_9901);
nand U10049 (N_10049,N_9770,N_9809);
or U10050 (N_10050,N_9912,N_9907);
nor U10051 (N_10051,N_9780,N_9797);
and U10052 (N_10052,N_9813,N_9839);
and U10053 (N_10053,N_9882,N_9800);
and U10054 (N_10054,N_9828,N_9858);
nor U10055 (N_10055,N_9814,N_9872);
nor U10056 (N_10056,N_9800,N_9838);
nand U10057 (N_10057,N_9785,N_9845);
or U10058 (N_10058,N_9840,N_9830);
or U10059 (N_10059,N_9829,N_9880);
or U10060 (N_10060,N_9762,N_9873);
nand U10061 (N_10061,N_9827,N_9785);
xnor U10062 (N_10062,N_9889,N_9905);
and U10063 (N_10063,N_9764,N_9785);
and U10064 (N_10064,N_9869,N_9814);
or U10065 (N_10065,N_9793,N_9762);
xor U10066 (N_10066,N_9891,N_9872);
and U10067 (N_10067,N_9844,N_9852);
xor U10068 (N_10068,N_9803,N_9901);
nor U10069 (N_10069,N_9911,N_9812);
nand U10070 (N_10070,N_9865,N_9868);
nor U10071 (N_10071,N_9882,N_9905);
xor U10072 (N_10072,N_9853,N_9823);
or U10073 (N_10073,N_9780,N_9849);
nor U10074 (N_10074,N_9767,N_9860);
xnor U10075 (N_10075,N_9886,N_9904);
and U10076 (N_10076,N_9767,N_9873);
and U10077 (N_10077,N_9780,N_9880);
or U10078 (N_10078,N_9835,N_9813);
nor U10079 (N_10079,N_9825,N_9882);
or U10080 (N_10080,N_9988,N_10045);
xnor U10081 (N_10081,N_10054,N_10007);
xnor U10082 (N_10082,N_10035,N_10021);
nand U10083 (N_10083,N_10051,N_10027);
xor U10084 (N_10084,N_10002,N_10019);
or U10085 (N_10085,N_10033,N_10005);
nor U10086 (N_10086,N_9947,N_10048);
xor U10087 (N_10087,N_9984,N_10065);
nor U10088 (N_10088,N_10077,N_10026);
nor U10089 (N_10089,N_10046,N_10052);
nor U10090 (N_10090,N_10024,N_9926);
and U10091 (N_10091,N_9945,N_9959);
xnor U10092 (N_10092,N_10059,N_9982);
nand U10093 (N_10093,N_10008,N_10075);
or U10094 (N_10094,N_10057,N_9925);
and U10095 (N_10095,N_10062,N_9936);
and U10096 (N_10096,N_9941,N_9973);
nor U10097 (N_10097,N_10061,N_9946);
or U10098 (N_10098,N_10001,N_9944);
or U10099 (N_10099,N_10072,N_10055);
nand U10100 (N_10100,N_9922,N_9920);
and U10101 (N_10101,N_9989,N_9937);
or U10102 (N_10102,N_9995,N_10017);
or U10103 (N_10103,N_9971,N_9994);
or U10104 (N_10104,N_9928,N_10011);
nand U10105 (N_10105,N_10040,N_9921);
nor U10106 (N_10106,N_10047,N_9997);
nand U10107 (N_10107,N_9951,N_9975);
and U10108 (N_10108,N_9991,N_9955);
and U10109 (N_10109,N_10004,N_9929);
nor U10110 (N_10110,N_9977,N_10043);
and U10111 (N_10111,N_10073,N_9967);
xor U10112 (N_10112,N_10003,N_9957);
and U10113 (N_10113,N_10066,N_10069);
nand U10114 (N_10114,N_10018,N_9999);
xnor U10115 (N_10115,N_10034,N_10060);
nor U10116 (N_10116,N_9996,N_9968);
nand U10117 (N_10117,N_10042,N_10041);
or U10118 (N_10118,N_9962,N_9979);
nor U10119 (N_10119,N_10078,N_9940);
and U10120 (N_10120,N_10070,N_9958);
xor U10121 (N_10121,N_10063,N_9956);
or U10122 (N_10122,N_9950,N_9980);
nand U10123 (N_10123,N_9938,N_9933);
and U10124 (N_10124,N_10076,N_9990);
xor U10125 (N_10125,N_10022,N_10074);
xor U10126 (N_10126,N_9983,N_10030);
xor U10127 (N_10127,N_10079,N_10009);
or U10128 (N_10128,N_10064,N_10038);
nand U10129 (N_10129,N_9992,N_10037);
or U10130 (N_10130,N_9998,N_9939);
nor U10131 (N_10131,N_9960,N_10012);
or U10132 (N_10132,N_10031,N_10049);
xor U10133 (N_10133,N_9961,N_9942);
and U10134 (N_10134,N_9981,N_9954);
nand U10135 (N_10135,N_10067,N_9924);
and U10136 (N_10136,N_9985,N_9966);
or U10137 (N_10137,N_9948,N_10015);
nand U10138 (N_10138,N_10016,N_9932);
nor U10139 (N_10139,N_10025,N_10056);
nand U10140 (N_10140,N_9935,N_10028);
nor U10141 (N_10141,N_9976,N_10013);
nand U10142 (N_10142,N_9952,N_9965);
nor U10143 (N_10143,N_10036,N_9943);
nand U10144 (N_10144,N_10039,N_9986);
nor U10145 (N_10145,N_9987,N_10000);
nand U10146 (N_10146,N_9970,N_9978);
and U10147 (N_10147,N_10032,N_10006);
nand U10148 (N_10148,N_9949,N_9927);
nor U10149 (N_10149,N_10071,N_10068);
xor U10150 (N_10150,N_10044,N_9969);
and U10151 (N_10151,N_9974,N_9963);
or U10152 (N_10152,N_10020,N_10010);
and U10153 (N_10153,N_10014,N_9931);
or U10154 (N_10154,N_10029,N_10050);
and U10155 (N_10155,N_9993,N_9972);
or U10156 (N_10156,N_10023,N_9930);
xnor U10157 (N_10157,N_9934,N_10053);
nor U10158 (N_10158,N_10058,N_9964);
and U10159 (N_10159,N_9953,N_9923);
or U10160 (N_10160,N_10072,N_9926);
nor U10161 (N_10161,N_9941,N_9975);
and U10162 (N_10162,N_9962,N_10027);
xor U10163 (N_10163,N_9960,N_9980);
and U10164 (N_10164,N_9930,N_9956);
nand U10165 (N_10165,N_10017,N_9965);
nand U10166 (N_10166,N_10045,N_9934);
or U10167 (N_10167,N_9996,N_9936);
and U10168 (N_10168,N_9966,N_9938);
and U10169 (N_10169,N_9955,N_9990);
nor U10170 (N_10170,N_9987,N_9947);
nand U10171 (N_10171,N_9957,N_10014);
and U10172 (N_10172,N_9962,N_9954);
xor U10173 (N_10173,N_9997,N_9921);
nor U10174 (N_10174,N_10019,N_9936);
or U10175 (N_10175,N_10027,N_9958);
and U10176 (N_10176,N_9993,N_9995);
nor U10177 (N_10177,N_10012,N_9936);
and U10178 (N_10178,N_10030,N_10011);
and U10179 (N_10179,N_9973,N_9934);
nor U10180 (N_10180,N_10069,N_9997);
nand U10181 (N_10181,N_10054,N_9926);
xnor U10182 (N_10182,N_10034,N_9926);
and U10183 (N_10183,N_9969,N_9962);
and U10184 (N_10184,N_10077,N_9961);
nor U10185 (N_10185,N_10071,N_9935);
or U10186 (N_10186,N_10015,N_9929);
and U10187 (N_10187,N_10062,N_9925);
xnor U10188 (N_10188,N_9999,N_9988);
and U10189 (N_10189,N_9937,N_10000);
and U10190 (N_10190,N_9935,N_9975);
nor U10191 (N_10191,N_10073,N_10007);
xor U10192 (N_10192,N_9943,N_9937);
or U10193 (N_10193,N_10038,N_10079);
and U10194 (N_10194,N_9990,N_10050);
nand U10195 (N_10195,N_10071,N_10054);
nor U10196 (N_10196,N_10013,N_10068);
or U10197 (N_10197,N_9972,N_10054);
and U10198 (N_10198,N_9997,N_10065);
nand U10199 (N_10199,N_10077,N_9937);
nor U10200 (N_10200,N_10062,N_9998);
nand U10201 (N_10201,N_10019,N_10043);
nor U10202 (N_10202,N_9991,N_10047);
xor U10203 (N_10203,N_10044,N_10006);
nor U10204 (N_10204,N_9966,N_9939);
xnor U10205 (N_10205,N_9998,N_10010);
or U10206 (N_10206,N_9965,N_9935);
xor U10207 (N_10207,N_9975,N_10024);
nand U10208 (N_10208,N_10034,N_10054);
and U10209 (N_10209,N_9920,N_9993);
nand U10210 (N_10210,N_10019,N_9987);
or U10211 (N_10211,N_10048,N_10046);
nand U10212 (N_10212,N_9964,N_10025);
nand U10213 (N_10213,N_10011,N_10068);
nand U10214 (N_10214,N_9959,N_9936);
or U10215 (N_10215,N_9930,N_10004);
xnor U10216 (N_10216,N_10033,N_10051);
xor U10217 (N_10217,N_9977,N_10014);
and U10218 (N_10218,N_9964,N_10077);
or U10219 (N_10219,N_9923,N_10066);
nand U10220 (N_10220,N_10075,N_10065);
xnor U10221 (N_10221,N_10062,N_10006);
and U10222 (N_10222,N_10036,N_9945);
or U10223 (N_10223,N_9972,N_10008);
nand U10224 (N_10224,N_9934,N_9969);
and U10225 (N_10225,N_10000,N_10064);
or U10226 (N_10226,N_10007,N_9997);
or U10227 (N_10227,N_9990,N_10009);
nand U10228 (N_10228,N_9998,N_9929);
xor U10229 (N_10229,N_10068,N_9924);
or U10230 (N_10230,N_9921,N_9943);
nand U10231 (N_10231,N_10060,N_10035);
nor U10232 (N_10232,N_9958,N_10011);
nand U10233 (N_10233,N_9927,N_9945);
or U10234 (N_10234,N_10045,N_10077);
and U10235 (N_10235,N_9968,N_10005);
nand U10236 (N_10236,N_10023,N_9956);
xor U10237 (N_10237,N_10071,N_9996);
nor U10238 (N_10238,N_9945,N_10074);
nor U10239 (N_10239,N_9978,N_9920);
and U10240 (N_10240,N_10157,N_10171);
nand U10241 (N_10241,N_10095,N_10212);
or U10242 (N_10242,N_10085,N_10197);
nand U10243 (N_10243,N_10227,N_10082);
nor U10244 (N_10244,N_10107,N_10218);
or U10245 (N_10245,N_10204,N_10092);
nand U10246 (N_10246,N_10113,N_10229);
and U10247 (N_10247,N_10205,N_10210);
and U10248 (N_10248,N_10146,N_10083);
and U10249 (N_10249,N_10108,N_10187);
nand U10250 (N_10250,N_10109,N_10087);
and U10251 (N_10251,N_10167,N_10144);
nor U10252 (N_10252,N_10216,N_10202);
nand U10253 (N_10253,N_10156,N_10117);
nor U10254 (N_10254,N_10114,N_10172);
and U10255 (N_10255,N_10173,N_10236);
nor U10256 (N_10256,N_10192,N_10217);
nor U10257 (N_10257,N_10220,N_10132);
or U10258 (N_10258,N_10176,N_10221);
nand U10259 (N_10259,N_10089,N_10198);
nor U10260 (N_10260,N_10189,N_10104);
xor U10261 (N_10261,N_10159,N_10102);
or U10262 (N_10262,N_10147,N_10224);
xnor U10263 (N_10263,N_10097,N_10143);
nor U10264 (N_10264,N_10105,N_10090);
xnor U10265 (N_10265,N_10134,N_10124);
nor U10266 (N_10266,N_10211,N_10100);
nand U10267 (N_10267,N_10174,N_10206);
nand U10268 (N_10268,N_10088,N_10162);
nor U10269 (N_10269,N_10209,N_10094);
and U10270 (N_10270,N_10178,N_10101);
xnor U10271 (N_10271,N_10148,N_10128);
nor U10272 (N_10272,N_10131,N_10184);
and U10273 (N_10273,N_10234,N_10133);
xnor U10274 (N_10274,N_10141,N_10233);
nor U10275 (N_10275,N_10235,N_10179);
and U10276 (N_10276,N_10231,N_10135);
nand U10277 (N_10277,N_10194,N_10130);
and U10278 (N_10278,N_10190,N_10228);
or U10279 (N_10279,N_10181,N_10145);
and U10280 (N_10280,N_10196,N_10180);
and U10281 (N_10281,N_10098,N_10084);
xnor U10282 (N_10282,N_10142,N_10219);
nand U10283 (N_10283,N_10086,N_10199);
xnor U10284 (N_10284,N_10140,N_10093);
xor U10285 (N_10285,N_10116,N_10164);
or U10286 (N_10286,N_10081,N_10155);
and U10287 (N_10287,N_10185,N_10232);
xor U10288 (N_10288,N_10123,N_10126);
or U10289 (N_10289,N_10207,N_10165);
and U10290 (N_10290,N_10106,N_10151);
or U10291 (N_10291,N_10200,N_10203);
or U10292 (N_10292,N_10139,N_10183);
or U10293 (N_10293,N_10137,N_10091);
nand U10294 (N_10294,N_10175,N_10127);
nand U10295 (N_10295,N_10166,N_10096);
xnor U10296 (N_10296,N_10080,N_10153);
nand U10297 (N_10297,N_10103,N_10169);
or U10298 (N_10298,N_10188,N_10099);
and U10299 (N_10299,N_10230,N_10239);
and U10300 (N_10300,N_10115,N_10223);
nor U10301 (N_10301,N_10193,N_10119);
and U10302 (N_10302,N_10111,N_10160);
and U10303 (N_10303,N_10215,N_10186);
nor U10304 (N_10304,N_10136,N_10138);
and U10305 (N_10305,N_10154,N_10129);
nor U10306 (N_10306,N_10149,N_10222);
or U10307 (N_10307,N_10150,N_10177);
nor U10308 (N_10308,N_10182,N_10110);
nand U10309 (N_10309,N_10237,N_10225);
nand U10310 (N_10310,N_10122,N_10112);
nor U10311 (N_10311,N_10152,N_10170);
or U10312 (N_10312,N_10208,N_10191);
xor U10313 (N_10313,N_10214,N_10195);
xnor U10314 (N_10314,N_10161,N_10158);
xor U10315 (N_10315,N_10118,N_10238);
or U10316 (N_10316,N_10125,N_10226);
nand U10317 (N_10317,N_10168,N_10213);
nand U10318 (N_10318,N_10201,N_10120);
nor U10319 (N_10319,N_10121,N_10163);
xnor U10320 (N_10320,N_10084,N_10178);
xor U10321 (N_10321,N_10226,N_10196);
and U10322 (N_10322,N_10238,N_10201);
nand U10323 (N_10323,N_10102,N_10129);
or U10324 (N_10324,N_10084,N_10182);
xor U10325 (N_10325,N_10134,N_10232);
xor U10326 (N_10326,N_10213,N_10228);
or U10327 (N_10327,N_10234,N_10127);
nor U10328 (N_10328,N_10222,N_10230);
xnor U10329 (N_10329,N_10095,N_10137);
nand U10330 (N_10330,N_10105,N_10176);
nand U10331 (N_10331,N_10176,N_10112);
nor U10332 (N_10332,N_10103,N_10127);
or U10333 (N_10333,N_10102,N_10190);
xor U10334 (N_10334,N_10178,N_10080);
nor U10335 (N_10335,N_10142,N_10090);
xor U10336 (N_10336,N_10108,N_10223);
or U10337 (N_10337,N_10131,N_10130);
xor U10338 (N_10338,N_10099,N_10135);
xnor U10339 (N_10339,N_10096,N_10181);
and U10340 (N_10340,N_10212,N_10122);
xnor U10341 (N_10341,N_10178,N_10203);
or U10342 (N_10342,N_10190,N_10231);
and U10343 (N_10343,N_10111,N_10129);
and U10344 (N_10344,N_10084,N_10158);
nor U10345 (N_10345,N_10107,N_10091);
or U10346 (N_10346,N_10223,N_10183);
or U10347 (N_10347,N_10131,N_10190);
or U10348 (N_10348,N_10119,N_10141);
nor U10349 (N_10349,N_10158,N_10237);
and U10350 (N_10350,N_10092,N_10219);
xor U10351 (N_10351,N_10188,N_10189);
nand U10352 (N_10352,N_10215,N_10188);
nand U10353 (N_10353,N_10087,N_10192);
nor U10354 (N_10354,N_10188,N_10194);
nor U10355 (N_10355,N_10173,N_10223);
and U10356 (N_10356,N_10156,N_10179);
and U10357 (N_10357,N_10138,N_10195);
xnor U10358 (N_10358,N_10237,N_10202);
xnor U10359 (N_10359,N_10191,N_10143);
or U10360 (N_10360,N_10162,N_10169);
xnor U10361 (N_10361,N_10226,N_10158);
and U10362 (N_10362,N_10102,N_10153);
nor U10363 (N_10363,N_10104,N_10106);
xnor U10364 (N_10364,N_10227,N_10165);
xnor U10365 (N_10365,N_10160,N_10098);
nor U10366 (N_10366,N_10128,N_10228);
nor U10367 (N_10367,N_10176,N_10203);
and U10368 (N_10368,N_10091,N_10090);
and U10369 (N_10369,N_10172,N_10103);
and U10370 (N_10370,N_10239,N_10222);
or U10371 (N_10371,N_10125,N_10143);
and U10372 (N_10372,N_10104,N_10098);
or U10373 (N_10373,N_10205,N_10172);
or U10374 (N_10374,N_10218,N_10224);
nor U10375 (N_10375,N_10193,N_10126);
nand U10376 (N_10376,N_10166,N_10157);
and U10377 (N_10377,N_10103,N_10131);
xor U10378 (N_10378,N_10188,N_10166);
nor U10379 (N_10379,N_10170,N_10145);
nand U10380 (N_10380,N_10224,N_10158);
nor U10381 (N_10381,N_10230,N_10197);
xnor U10382 (N_10382,N_10111,N_10176);
xor U10383 (N_10383,N_10179,N_10097);
and U10384 (N_10384,N_10220,N_10224);
and U10385 (N_10385,N_10168,N_10113);
nor U10386 (N_10386,N_10206,N_10193);
nor U10387 (N_10387,N_10121,N_10215);
xnor U10388 (N_10388,N_10170,N_10106);
or U10389 (N_10389,N_10144,N_10115);
xor U10390 (N_10390,N_10211,N_10192);
xnor U10391 (N_10391,N_10184,N_10155);
nor U10392 (N_10392,N_10147,N_10135);
and U10393 (N_10393,N_10199,N_10084);
or U10394 (N_10394,N_10234,N_10167);
nand U10395 (N_10395,N_10095,N_10229);
nand U10396 (N_10396,N_10141,N_10142);
and U10397 (N_10397,N_10181,N_10198);
nand U10398 (N_10398,N_10213,N_10214);
nand U10399 (N_10399,N_10187,N_10170);
or U10400 (N_10400,N_10303,N_10318);
or U10401 (N_10401,N_10242,N_10324);
nor U10402 (N_10402,N_10397,N_10337);
or U10403 (N_10403,N_10368,N_10361);
nor U10404 (N_10404,N_10256,N_10321);
or U10405 (N_10405,N_10312,N_10369);
and U10406 (N_10406,N_10243,N_10354);
and U10407 (N_10407,N_10394,N_10391);
xnor U10408 (N_10408,N_10356,N_10349);
nand U10409 (N_10409,N_10373,N_10363);
and U10410 (N_10410,N_10320,N_10286);
or U10411 (N_10411,N_10390,N_10270);
nand U10412 (N_10412,N_10298,N_10342);
nor U10413 (N_10413,N_10291,N_10310);
nor U10414 (N_10414,N_10307,N_10241);
xor U10415 (N_10415,N_10305,N_10374);
xor U10416 (N_10416,N_10336,N_10268);
xnor U10417 (N_10417,N_10319,N_10365);
nand U10418 (N_10418,N_10383,N_10387);
and U10419 (N_10419,N_10289,N_10309);
nor U10420 (N_10420,N_10250,N_10316);
xor U10421 (N_10421,N_10251,N_10345);
nand U10422 (N_10422,N_10267,N_10258);
nor U10423 (N_10423,N_10366,N_10295);
nor U10424 (N_10424,N_10264,N_10327);
xnor U10425 (N_10425,N_10274,N_10347);
nand U10426 (N_10426,N_10352,N_10380);
or U10427 (N_10427,N_10334,N_10381);
nor U10428 (N_10428,N_10371,N_10364);
xor U10429 (N_10429,N_10370,N_10377);
or U10430 (N_10430,N_10362,N_10263);
nand U10431 (N_10431,N_10276,N_10300);
or U10432 (N_10432,N_10357,N_10341);
and U10433 (N_10433,N_10389,N_10294);
nand U10434 (N_10434,N_10340,N_10375);
or U10435 (N_10435,N_10313,N_10292);
xnor U10436 (N_10436,N_10285,N_10245);
nand U10437 (N_10437,N_10244,N_10266);
nor U10438 (N_10438,N_10360,N_10265);
nor U10439 (N_10439,N_10252,N_10398);
or U10440 (N_10440,N_10314,N_10288);
or U10441 (N_10441,N_10344,N_10297);
xnor U10442 (N_10442,N_10322,N_10240);
xnor U10443 (N_10443,N_10283,N_10399);
xnor U10444 (N_10444,N_10287,N_10351);
nor U10445 (N_10445,N_10269,N_10311);
nand U10446 (N_10446,N_10323,N_10261);
xnor U10447 (N_10447,N_10282,N_10339);
xor U10448 (N_10448,N_10248,N_10317);
xor U10449 (N_10449,N_10279,N_10254);
xnor U10450 (N_10450,N_10280,N_10385);
and U10451 (N_10451,N_10350,N_10299);
nor U10452 (N_10452,N_10315,N_10325);
and U10453 (N_10453,N_10308,N_10384);
xor U10454 (N_10454,N_10386,N_10343);
xor U10455 (N_10455,N_10348,N_10260);
xnor U10456 (N_10456,N_10329,N_10379);
and U10457 (N_10457,N_10262,N_10284);
and U10458 (N_10458,N_10246,N_10273);
and U10459 (N_10459,N_10395,N_10331);
and U10460 (N_10460,N_10272,N_10388);
or U10461 (N_10461,N_10346,N_10353);
nor U10462 (N_10462,N_10376,N_10333);
nand U10463 (N_10463,N_10358,N_10372);
xnor U10464 (N_10464,N_10296,N_10367);
or U10465 (N_10465,N_10253,N_10330);
xnor U10466 (N_10466,N_10247,N_10393);
nand U10467 (N_10467,N_10382,N_10275);
xnor U10468 (N_10468,N_10257,N_10281);
and U10469 (N_10469,N_10302,N_10249);
nor U10470 (N_10470,N_10306,N_10290);
or U10471 (N_10471,N_10259,N_10378);
xnor U10472 (N_10472,N_10392,N_10355);
and U10473 (N_10473,N_10271,N_10338);
and U10474 (N_10474,N_10293,N_10328);
nor U10475 (N_10475,N_10277,N_10335);
nor U10476 (N_10476,N_10332,N_10255);
or U10477 (N_10477,N_10359,N_10301);
xnor U10478 (N_10478,N_10304,N_10278);
nand U10479 (N_10479,N_10326,N_10396);
or U10480 (N_10480,N_10389,N_10292);
xnor U10481 (N_10481,N_10267,N_10335);
nor U10482 (N_10482,N_10390,N_10294);
nor U10483 (N_10483,N_10247,N_10323);
nand U10484 (N_10484,N_10354,N_10287);
or U10485 (N_10485,N_10301,N_10293);
nand U10486 (N_10486,N_10331,N_10340);
xnor U10487 (N_10487,N_10375,N_10381);
nand U10488 (N_10488,N_10252,N_10397);
and U10489 (N_10489,N_10250,N_10262);
or U10490 (N_10490,N_10383,N_10273);
or U10491 (N_10491,N_10335,N_10342);
nor U10492 (N_10492,N_10327,N_10329);
nor U10493 (N_10493,N_10363,N_10353);
xor U10494 (N_10494,N_10292,N_10355);
nand U10495 (N_10495,N_10343,N_10242);
xor U10496 (N_10496,N_10348,N_10364);
nor U10497 (N_10497,N_10368,N_10340);
nor U10498 (N_10498,N_10331,N_10343);
and U10499 (N_10499,N_10291,N_10385);
nand U10500 (N_10500,N_10368,N_10298);
nand U10501 (N_10501,N_10331,N_10339);
nor U10502 (N_10502,N_10333,N_10267);
xor U10503 (N_10503,N_10343,N_10282);
nor U10504 (N_10504,N_10349,N_10383);
or U10505 (N_10505,N_10321,N_10345);
or U10506 (N_10506,N_10309,N_10341);
and U10507 (N_10507,N_10313,N_10332);
nand U10508 (N_10508,N_10267,N_10372);
or U10509 (N_10509,N_10249,N_10282);
and U10510 (N_10510,N_10251,N_10249);
xor U10511 (N_10511,N_10302,N_10379);
or U10512 (N_10512,N_10240,N_10255);
xor U10513 (N_10513,N_10265,N_10312);
xnor U10514 (N_10514,N_10366,N_10268);
nand U10515 (N_10515,N_10341,N_10294);
and U10516 (N_10516,N_10247,N_10282);
nand U10517 (N_10517,N_10356,N_10398);
and U10518 (N_10518,N_10326,N_10320);
and U10519 (N_10519,N_10328,N_10344);
nand U10520 (N_10520,N_10311,N_10398);
or U10521 (N_10521,N_10312,N_10252);
and U10522 (N_10522,N_10243,N_10341);
nand U10523 (N_10523,N_10302,N_10385);
nand U10524 (N_10524,N_10376,N_10395);
nor U10525 (N_10525,N_10369,N_10277);
nor U10526 (N_10526,N_10346,N_10251);
nor U10527 (N_10527,N_10378,N_10363);
or U10528 (N_10528,N_10346,N_10303);
or U10529 (N_10529,N_10293,N_10247);
or U10530 (N_10530,N_10298,N_10330);
and U10531 (N_10531,N_10249,N_10279);
and U10532 (N_10532,N_10328,N_10241);
or U10533 (N_10533,N_10352,N_10341);
or U10534 (N_10534,N_10281,N_10368);
xnor U10535 (N_10535,N_10371,N_10330);
and U10536 (N_10536,N_10388,N_10301);
or U10537 (N_10537,N_10324,N_10277);
or U10538 (N_10538,N_10297,N_10259);
nor U10539 (N_10539,N_10244,N_10346);
xor U10540 (N_10540,N_10323,N_10370);
nor U10541 (N_10541,N_10260,N_10332);
xor U10542 (N_10542,N_10292,N_10388);
and U10543 (N_10543,N_10299,N_10252);
xor U10544 (N_10544,N_10280,N_10257);
nor U10545 (N_10545,N_10364,N_10316);
nand U10546 (N_10546,N_10383,N_10255);
and U10547 (N_10547,N_10322,N_10243);
and U10548 (N_10548,N_10281,N_10271);
nand U10549 (N_10549,N_10260,N_10322);
xor U10550 (N_10550,N_10326,N_10350);
nand U10551 (N_10551,N_10285,N_10342);
and U10552 (N_10552,N_10359,N_10331);
xnor U10553 (N_10553,N_10268,N_10295);
or U10554 (N_10554,N_10338,N_10348);
nor U10555 (N_10555,N_10316,N_10390);
and U10556 (N_10556,N_10342,N_10360);
nand U10557 (N_10557,N_10360,N_10387);
or U10558 (N_10558,N_10284,N_10393);
or U10559 (N_10559,N_10351,N_10252);
xor U10560 (N_10560,N_10507,N_10540);
nor U10561 (N_10561,N_10519,N_10413);
or U10562 (N_10562,N_10469,N_10483);
xnor U10563 (N_10563,N_10539,N_10553);
nor U10564 (N_10564,N_10550,N_10494);
and U10565 (N_10565,N_10537,N_10501);
or U10566 (N_10566,N_10411,N_10503);
nor U10567 (N_10567,N_10427,N_10541);
nor U10568 (N_10568,N_10451,N_10512);
nand U10569 (N_10569,N_10437,N_10468);
nor U10570 (N_10570,N_10429,N_10490);
or U10571 (N_10571,N_10405,N_10491);
or U10572 (N_10572,N_10525,N_10528);
xor U10573 (N_10573,N_10495,N_10461);
or U10574 (N_10574,N_10435,N_10425);
xnor U10575 (N_10575,N_10510,N_10544);
and U10576 (N_10576,N_10552,N_10459);
nand U10577 (N_10577,N_10477,N_10419);
and U10578 (N_10578,N_10422,N_10444);
and U10579 (N_10579,N_10516,N_10450);
or U10580 (N_10580,N_10443,N_10466);
and U10581 (N_10581,N_10445,N_10511);
nor U10582 (N_10582,N_10538,N_10484);
and U10583 (N_10583,N_10545,N_10497);
xor U10584 (N_10584,N_10471,N_10496);
or U10585 (N_10585,N_10489,N_10407);
xor U10586 (N_10586,N_10438,N_10558);
and U10587 (N_10587,N_10473,N_10474);
or U10588 (N_10588,N_10522,N_10487);
nand U10589 (N_10589,N_10408,N_10548);
or U10590 (N_10590,N_10559,N_10465);
xor U10591 (N_10591,N_10467,N_10480);
xor U10592 (N_10592,N_10527,N_10504);
nor U10593 (N_10593,N_10420,N_10448);
nor U10594 (N_10594,N_10442,N_10457);
nand U10595 (N_10595,N_10410,N_10488);
nor U10596 (N_10596,N_10547,N_10460);
nor U10597 (N_10597,N_10464,N_10499);
nand U10598 (N_10598,N_10421,N_10432);
nor U10599 (N_10599,N_10530,N_10482);
and U10600 (N_10600,N_10481,N_10533);
and U10601 (N_10601,N_10514,N_10426);
nor U10602 (N_10602,N_10400,N_10434);
xor U10603 (N_10603,N_10508,N_10518);
nor U10604 (N_10604,N_10406,N_10412);
and U10605 (N_10605,N_10416,N_10529);
xor U10606 (N_10606,N_10446,N_10555);
nor U10607 (N_10607,N_10431,N_10535);
nand U10608 (N_10608,N_10492,N_10418);
and U10609 (N_10609,N_10523,N_10470);
xor U10610 (N_10610,N_10458,N_10517);
nand U10611 (N_10611,N_10521,N_10462);
xor U10612 (N_10612,N_10509,N_10513);
and U10613 (N_10613,N_10531,N_10415);
xnor U10614 (N_10614,N_10500,N_10536);
or U10615 (N_10615,N_10506,N_10502);
nand U10616 (N_10616,N_10554,N_10551);
nand U10617 (N_10617,N_10433,N_10404);
nor U10618 (N_10618,N_10449,N_10439);
nor U10619 (N_10619,N_10549,N_10401);
xnor U10620 (N_10620,N_10557,N_10403);
nor U10621 (N_10621,N_10472,N_10453);
nor U10622 (N_10622,N_10428,N_10430);
or U10623 (N_10623,N_10456,N_10436);
nor U10624 (N_10624,N_10475,N_10505);
and U10625 (N_10625,N_10423,N_10534);
xor U10626 (N_10626,N_10414,N_10485);
and U10627 (N_10627,N_10463,N_10543);
or U10628 (N_10628,N_10441,N_10455);
or U10629 (N_10629,N_10520,N_10424);
and U10630 (N_10630,N_10454,N_10409);
nor U10631 (N_10631,N_10440,N_10526);
and U10632 (N_10632,N_10532,N_10479);
xnor U10633 (N_10633,N_10498,N_10417);
and U10634 (N_10634,N_10452,N_10447);
or U10635 (N_10635,N_10478,N_10515);
xnor U10636 (N_10636,N_10476,N_10524);
nand U10637 (N_10637,N_10493,N_10402);
and U10638 (N_10638,N_10486,N_10556);
or U10639 (N_10639,N_10546,N_10542);
and U10640 (N_10640,N_10529,N_10421);
or U10641 (N_10641,N_10551,N_10494);
and U10642 (N_10642,N_10452,N_10541);
or U10643 (N_10643,N_10427,N_10517);
or U10644 (N_10644,N_10404,N_10432);
xnor U10645 (N_10645,N_10405,N_10549);
xor U10646 (N_10646,N_10528,N_10480);
or U10647 (N_10647,N_10544,N_10412);
nand U10648 (N_10648,N_10431,N_10440);
or U10649 (N_10649,N_10534,N_10528);
nand U10650 (N_10650,N_10402,N_10518);
xor U10651 (N_10651,N_10471,N_10400);
or U10652 (N_10652,N_10448,N_10433);
and U10653 (N_10653,N_10439,N_10410);
nand U10654 (N_10654,N_10501,N_10402);
nand U10655 (N_10655,N_10551,N_10475);
and U10656 (N_10656,N_10406,N_10400);
or U10657 (N_10657,N_10416,N_10480);
xnor U10658 (N_10658,N_10470,N_10434);
and U10659 (N_10659,N_10554,N_10490);
or U10660 (N_10660,N_10472,N_10481);
nand U10661 (N_10661,N_10549,N_10516);
nor U10662 (N_10662,N_10419,N_10408);
xor U10663 (N_10663,N_10477,N_10553);
and U10664 (N_10664,N_10478,N_10519);
or U10665 (N_10665,N_10441,N_10485);
nor U10666 (N_10666,N_10466,N_10432);
nor U10667 (N_10667,N_10415,N_10463);
xor U10668 (N_10668,N_10520,N_10499);
xnor U10669 (N_10669,N_10472,N_10409);
or U10670 (N_10670,N_10559,N_10402);
and U10671 (N_10671,N_10417,N_10460);
nor U10672 (N_10672,N_10505,N_10530);
and U10673 (N_10673,N_10431,N_10423);
xnor U10674 (N_10674,N_10431,N_10426);
or U10675 (N_10675,N_10419,N_10559);
xnor U10676 (N_10676,N_10539,N_10436);
or U10677 (N_10677,N_10516,N_10518);
xnor U10678 (N_10678,N_10467,N_10549);
xor U10679 (N_10679,N_10405,N_10495);
and U10680 (N_10680,N_10481,N_10483);
xor U10681 (N_10681,N_10438,N_10462);
nand U10682 (N_10682,N_10516,N_10479);
nor U10683 (N_10683,N_10495,N_10499);
or U10684 (N_10684,N_10412,N_10547);
xnor U10685 (N_10685,N_10555,N_10501);
and U10686 (N_10686,N_10533,N_10497);
nand U10687 (N_10687,N_10405,N_10468);
nand U10688 (N_10688,N_10446,N_10519);
nor U10689 (N_10689,N_10444,N_10515);
nand U10690 (N_10690,N_10466,N_10423);
and U10691 (N_10691,N_10441,N_10525);
nor U10692 (N_10692,N_10435,N_10530);
and U10693 (N_10693,N_10518,N_10540);
xor U10694 (N_10694,N_10469,N_10508);
and U10695 (N_10695,N_10548,N_10487);
nand U10696 (N_10696,N_10531,N_10500);
nor U10697 (N_10697,N_10559,N_10459);
nand U10698 (N_10698,N_10505,N_10523);
xor U10699 (N_10699,N_10416,N_10439);
xnor U10700 (N_10700,N_10480,N_10432);
nand U10701 (N_10701,N_10481,N_10487);
nor U10702 (N_10702,N_10400,N_10423);
nor U10703 (N_10703,N_10521,N_10408);
xnor U10704 (N_10704,N_10528,N_10459);
and U10705 (N_10705,N_10525,N_10536);
and U10706 (N_10706,N_10410,N_10470);
or U10707 (N_10707,N_10404,N_10528);
or U10708 (N_10708,N_10409,N_10522);
xor U10709 (N_10709,N_10514,N_10530);
nand U10710 (N_10710,N_10482,N_10520);
or U10711 (N_10711,N_10513,N_10506);
nand U10712 (N_10712,N_10514,N_10430);
nor U10713 (N_10713,N_10548,N_10488);
nand U10714 (N_10714,N_10449,N_10413);
nand U10715 (N_10715,N_10488,N_10506);
xnor U10716 (N_10716,N_10497,N_10430);
or U10717 (N_10717,N_10408,N_10404);
nand U10718 (N_10718,N_10492,N_10442);
nor U10719 (N_10719,N_10454,N_10457);
nand U10720 (N_10720,N_10682,N_10582);
nor U10721 (N_10721,N_10708,N_10646);
nor U10722 (N_10722,N_10688,N_10683);
nor U10723 (N_10723,N_10679,N_10586);
and U10724 (N_10724,N_10633,N_10685);
xnor U10725 (N_10725,N_10605,N_10572);
nor U10726 (N_10726,N_10621,N_10623);
nand U10727 (N_10727,N_10600,N_10637);
nor U10728 (N_10728,N_10568,N_10567);
and U10729 (N_10729,N_10625,N_10664);
xnor U10730 (N_10730,N_10640,N_10676);
nand U10731 (N_10731,N_10581,N_10585);
nand U10732 (N_10732,N_10570,N_10649);
nand U10733 (N_10733,N_10593,N_10589);
and U10734 (N_10734,N_10716,N_10642);
nor U10735 (N_10735,N_10715,N_10561);
or U10736 (N_10736,N_10670,N_10632);
nand U10737 (N_10737,N_10699,N_10631);
and U10738 (N_10738,N_10604,N_10575);
nand U10739 (N_10739,N_10574,N_10647);
xor U10740 (N_10740,N_10563,N_10710);
nand U10741 (N_10741,N_10615,N_10610);
nand U10742 (N_10742,N_10587,N_10656);
and U10743 (N_10743,N_10571,N_10609);
nor U10744 (N_10744,N_10626,N_10620);
nor U10745 (N_10745,N_10598,N_10636);
or U10746 (N_10746,N_10564,N_10645);
nor U10747 (N_10747,N_10599,N_10662);
xnor U10748 (N_10748,N_10616,N_10680);
nor U10749 (N_10749,N_10692,N_10681);
or U10750 (N_10750,N_10591,N_10641);
or U10751 (N_10751,N_10566,N_10596);
nor U10752 (N_10752,N_10630,N_10562);
nor U10753 (N_10753,N_10659,N_10704);
nand U10754 (N_10754,N_10638,N_10660);
or U10755 (N_10755,N_10560,N_10628);
xor U10756 (N_10756,N_10677,N_10622);
or U10757 (N_10757,N_10653,N_10694);
and U10758 (N_10758,N_10652,N_10665);
and U10759 (N_10759,N_10655,N_10606);
and U10760 (N_10760,N_10675,N_10601);
and U10761 (N_10761,N_10577,N_10629);
or U10762 (N_10762,N_10617,N_10613);
and U10763 (N_10763,N_10657,N_10619);
and U10764 (N_10764,N_10717,N_10713);
and U10765 (N_10765,N_10594,N_10671);
or U10766 (N_10766,N_10707,N_10718);
xor U10767 (N_10767,N_10651,N_10608);
and U10768 (N_10768,N_10687,N_10611);
and U10769 (N_10769,N_10627,N_10666);
or U10770 (N_10770,N_10584,N_10573);
nor U10771 (N_10771,N_10706,N_10635);
and U10772 (N_10772,N_10648,N_10576);
nor U10773 (N_10773,N_10644,N_10719);
or U10774 (N_10774,N_10569,N_10588);
or U10775 (N_10775,N_10674,N_10689);
or U10776 (N_10776,N_10592,N_10669);
nor U10777 (N_10777,N_10612,N_10583);
xnor U10778 (N_10778,N_10691,N_10697);
and U10779 (N_10779,N_10668,N_10714);
and U10780 (N_10780,N_10678,N_10701);
and U10781 (N_10781,N_10673,N_10579);
nor U10782 (N_10782,N_10700,N_10684);
or U10783 (N_10783,N_10672,N_10590);
and U10784 (N_10784,N_10693,N_10667);
nor U10785 (N_10785,N_10686,N_10602);
or U10786 (N_10786,N_10711,N_10696);
or U10787 (N_10787,N_10634,N_10705);
and U10788 (N_10788,N_10658,N_10614);
and U10789 (N_10789,N_10618,N_10650);
xor U10790 (N_10790,N_10624,N_10690);
xor U10791 (N_10791,N_10698,N_10597);
and U10792 (N_10792,N_10702,N_10695);
nand U10793 (N_10793,N_10607,N_10712);
nor U10794 (N_10794,N_10603,N_10654);
nand U10795 (N_10795,N_10709,N_10580);
or U10796 (N_10796,N_10578,N_10643);
nor U10797 (N_10797,N_10639,N_10661);
and U10798 (N_10798,N_10703,N_10595);
or U10799 (N_10799,N_10663,N_10565);
and U10800 (N_10800,N_10680,N_10583);
nand U10801 (N_10801,N_10567,N_10639);
and U10802 (N_10802,N_10671,N_10699);
or U10803 (N_10803,N_10654,N_10652);
and U10804 (N_10804,N_10713,N_10600);
xnor U10805 (N_10805,N_10576,N_10715);
or U10806 (N_10806,N_10628,N_10600);
xnor U10807 (N_10807,N_10703,N_10596);
nor U10808 (N_10808,N_10709,N_10630);
nand U10809 (N_10809,N_10668,N_10701);
nor U10810 (N_10810,N_10656,N_10710);
and U10811 (N_10811,N_10672,N_10564);
and U10812 (N_10812,N_10654,N_10622);
nand U10813 (N_10813,N_10632,N_10675);
nor U10814 (N_10814,N_10639,N_10636);
nand U10815 (N_10815,N_10623,N_10606);
or U10816 (N_10816,N_10699,N_10646);
xnor U10817 (N_10817,N_10712,N_10628);
and U10818 (N_10818,N_10580,N_10695);
or U10819 (N_10819,N_10602,N_10624);
or U10820 (N_10820,N_10597,N_10560);
or U10821 (N_10821,N_10571,N_10675);
nand U10822 (N_10822,N_10577,N_10666);
nor U10823 (N_10823,N_10617,N_10597);
or U10824 (N_10824,N_10605,N_10690);
or U10825 (N_10825,N_10674,N_10680);
nor U10826 (N_10826,N_10690,N_10677);
and U10827 (N_10827,N_10663,N_10703);
nand U10828 (N_10828,N_10688,N_10566);
and U10829 (N_10829,N_10670,N_10678);
or U10830 (N_10830,N_10610,N_10596);
xor U10831 (N_10831,N_10613,N_10619);
nand U10832 (N_10832,N_10630,N_10587);
nand U10833 (N_10833,N_10655,N_10624);
and U10834 (N_10834,N_10678,N_10716);
or U10835 (N_10835,N_10633,N_10623);
nand U10836 (N_10836,N_10621,N_10596);
nand U10837 (N_10837,N_10613,N_10581);
nor U10838 (N_10838,N_10683,N_10673);
xor U10839 (N_10839,N_10621,N_10636);
nor U10840 (N_10840,N_10633,N_10715);
nand U10841 (N_10841,N_10578,N_10694);
or U10842 (N_10842,N_10589,N_10697);
nor U10843 (N_10843,N_10717,N_10610);
nor U10844 (N_10844,N_10652,N_10655);
nor U10845 (N_10845,N_10705,N_10581);
or U10846 (N_10846,N_10666,N_10692);
nand U10847 (N_10847,N_10714,N_10653);
xor U10848 (N_10848,N_10686,N_10625);
nor U10849 (N_10849,N_10614,N_10626);
xor U10850 (N_10850,N_10635,N_10717);
or U10851 (N_10851,N_10716,N_10666);
nor U10852 (N_10852,N_10565,N_10606);
or U10853 (N_10853,N_10645,N_10652);
and U10854 (N_10854,N_10612,N_10580);
xnor U10855 (N_10855,N_10675,N_10700);
and U10856 (N_10856,N_10691,N_10561);
or U10857 (N_10857,N_10649,N_10711);
and U10858 (N_10858,N_10644,N_10679);
nor U10859 (N_10859,N_10620,N_10715);
nand U10860 (N_10860,N_10685,N_10608);
and U10861 (N_10861,N_10585,N_10562);
nor U10862 (N_10862,N_10673,N_10677);
xor U10863 (N_10863,N_10699,N_10675);
nand U10864 (N_10864,N_10673,N_10582);
and U10865 (N_10865,N_10613,N_10664);
and U10866 (N_10866,N_10665,N_10715);
nand U10867 (N_10867,N_10679,N_10664);
nand U10868 (N_10868,N_10581,N_10580);
nor U10869 (N_10869,N_10632,N_10702);
nand U10870 (N_10870,N_10564,N_10655);
xnor U10871 (N_10871,N_10670,N_10714);
and U10872 (N_10872,N_10573,N_10603);
xor U10873 (N_10873,N_10704,N_10690);
nand U10874 (N_10874,N_10576,N_10656);
nor U10875 (N_10875,N_10679,N_10594);
xor U10876 (N_10876,N_10588,N_10700);
nor U10877 (N_10877,N_10647,N_10607);
or U10878 (N_10878,N_10578,N_10618);
nand U10879 (N_10879,N_10668,N_10633);
nor U10880 (N_10880,N_10857,N_10795);
nand U10881 (N_10881,N_10819,N_10731);
nand U10882 (N_10882,N_10786,N_10843);
nand U10883 (N_10883,N_10771,N_10826);
or U10884 (N_10884,N_10869,N_10764);
and U10885 (N_10885,N_10834,N_10746);
and U10886 (N_10886,N_10783,N_10745);
or U10887 (N_10887,N_10726,N_10847);
or U10888 (N_10888,N_10794,N_10809);
nand U10889 (N_10889,N_10808,N_10846);
and U10890 (N_10890,N_10866,N_10821);
nor U10891 (N_10891,N_10760,N_10828);
and U10892 (N_10892,N_10788,N_10790);
nand U10893 (N_10893,N_10729,N_10763);
nand U10894 (N_10894,N_10767,N_10782);
and U10895 (N_10895,N_10802,N_10738);
nor U10896 (N_10896,N_10751,N_10791);
nand U10897 (N_10897,N_10820,N_10836);
or U10898 (N_10898,N_10827,N_10770);
or U10899 (N_10899,N_10837,N_10854);
nor U10900 (N_10900,N_10733,N_10872);
or U10901 (N_10901,N_10728,N_10870);
and U10902 (N_10902,N_10750,N_10734);
nand U10903 (N_10903,N_10752,N_10784);
and U10904 (N_10904,N_10800,N_10725);
xnor U10905 (N_10905,N_10789,N_10863);
or U10906 (N_10906,N_10865,N_10798);
nand U10907 (N_10907,N_10864,N_10817);
and U10908 (N_10908,N_10811,N_10844);
and U10909 (N_10909,N_10851,N_10878);
or U10910 (N_10910,N_10774,N_10769);
or U10911 (N_10911,N_10829,N_10749);
and U10912 (N_10912,N_10754,N_10841);
or U10913 (N_10913,N_10858,N_10793);
nor U10914 (N_10914,N_10765,N_10761);
nor U10915 (N_10915,N_10768,N_10742);
nand U10916 (N_10916,N_10831,N_10812);
and U10917 (N_10917,N_10806,N_10839);
nand U10918 (N_10918,N_10842,N_10822);
xor U10919 (N_10919,N_10856,N_10735);
xnor U10920 (N_10920,N_10773,N_10830);
xnor U10921 (N_10921,N_10727,N_10780);
or U10922 (N_10922,N_10721,N_10823);
or U10923 (N_10923,N_10739,N_10720);
nor U10924 (N_10924,N_10840,N_10807);
nor U10925 (N_10925,N_10833,N_10804);
and U10926 (N_10926,N_10792,N_10813);
nand U10927 (N_10927,N_10785,N_10805);
or U10928 (N_10928,N_10776,N_10861);
nand U10929 (N_10929,N_10860,N_10759);
or U10930 (N_10930,N_10781,N_10815);
and U10931 (N_10931,N_10775,N_10801);
and U10932 (N_10932,N_10758,N_10777);
nand U10933 (N_10933,N_10873,N_10722);
and U10934 (N_10934,N_10816,N_10757);
and U10935 (N_10935,N_10744,N_10877);
nor U10936 (N_10936,N_10778,N_10879);
or U10937 (N_10937,N_10818,N_10845);
or U10938 (N_10938,N_10724,N_10772);
nand U10939 (N_10939,N_10838,N_10850);
nand U10940 (N_10940,N_10762,N_10859);
or U10941 (N_10941,N_10814,N_10832);
xor U10942 (N_10942,N_10747,N_10756);
nand U10943 (N_10943,N_10755,N_10787);
nand U10944 (N_10944,N_10853,N_10748);
or U10945 (N_10945,N_10743,N_10867);
nand U10946 (N_10946,N_10740,N_10737);
nand U10947 (N_10947,N_10835,N_10799);
nand U10948 (N_10948,N_10796,N_10871);
xor U10949 (N_10949,N_10824,N_10876);
nand U10950 (N_10950,N_10868,N_10875);
nand U10951 (N_10951,N_10732,N_10855);
xnor U10952 (N_10952,N_10779,N_10741);
and U10953 (N_10953,N_10862,N_10848);
or U10954 (N_10954,N_10736,N_10803);
nor U10955 (N_10955,N_10874,N_10852);
and U10956 (N_10956,N_10849,N_10825);
and U10957 (N_10957,N_10766,N_10730);
nand U10958 (N_10958,N_10723,N_10810);
xnor U10959 (N_10959,N_10753,N_10797);
and U10960 (N_10960,N_10815,N_10877);
nand U10961 (N_10961,N_10874,N_10838);
or U10962 (N_10962,N_10728,N_10744);
nor U10963 (N_10963,N_10815,N_10789);
or U10964 (N_10964,N_10756,N_10730);
xnor U10965 (N_10965,N_10762,N_10791);
or U10966 (N_10966,N_10824,N_10744);
or U10967 (N_10967,N_10814,N_10790);
nand U10968 (N_10968,N_10830,N_10874);
or U10969 (N_10969,N_10815,N_10850);
xor U10970 (N_10970,N_10830,N_10764);
and U10971 (N_10971,N_10808,N_10755);
nor U10972 (N_10972,N_10753,N_10806);
or U10973 (N_10973,N_10781,N_10831);
nor U10974 (N_10974,N_10846,N_10778);
xor U10975 (N_10975,N_10862,N_10805);
nand U10976 (N_10976,N_10724,N_10838);
and U10977 (N_10977,N_10748,N_10722);
and U10978 (N_10978,N_10757,N_10780);
xor U10979 (N_10979,N_10860,N_10867);
nand U10980 (N_10980,N_10775,N_10763);
or U10981 (N_10981,N_10785,N_10871);
nand U10982 (N_10982,N_10783,N_10742);
and U10983 (N_10983,N_10797,N_10790);
and U10984 (N_10984,N_10725,N_10813);
nand U10985 (N_10985,N_10725,N_10834);
xor U10986 (N_10986,N_10770,N_10751);
nand U10987 (N_10987,N_10767,N_10864);
nand U10988 (N_10988,N_10838,N_10734);
xnor U10989 (N_10989,N_10797,N_10737);
nor U10990 (N_10990,N_10874,N_10764);
and U10991 (N_10991,N_10808,N_10804);
and U10992 (N_10992,N_10721,N_10836);
and U10993 (N_10993,N_10857,N_10842);
or U10994 (N_10994,N_10817,N_10763);
xor U10995 (N_10995,N_10753,N_10732);
or U10996 (N_10996,N_10816,N_10872);
xor U10997 (N_10997,N_10721,N_10841);
and U10998 (N_10998,N_10771,N_10840);
or U10999 (N_10999,N_10848,N_10797);
xnor U11000 (N_11000,N_10805,N_10777);
xor U11001 (N_11001,N_10774,N_10861);
nand U11002 (N_11002,N_10837,N_10817);
nor U11003 (N_11003,N_10759,N_10743);
or U11004 (N_11004,N_10814,N_10726);
or U11005 (N_11005,N_10840,N_10774);
xor U11006 (N_11006,N_10777,N_10765);
or U11007 (N_11007,N_10744,N_10762);
nand U11008 (N_11008,N_10837,N_10831);
nor U11009 (N_11009,N_10826,N_10815);
nand U11010 (N_11010,N_10877,N_10764);
nand U11011 (N_11011,N_10817,N_10786);
or U11012 (N_11012,N_10834,N_10724);
or U11013 (N_11013,N_10737,N_10788);
nand U11014 (N_11014,N_10775,N_10810);
and U11015 (N_11015,N_10876,N_10844);
xnor U11016 (N_11016,N_10799,N_10794);
nand U11017 (N_11017,N_10727,N_10775);
and U11018 (N_11018,N_10746,N_10823);
xnor U11019 (N_11019,N_10777,N_10866);
nor U11020 (N_11020,N_10823,N_10779);
nor U11021 (N_11021,N_10874,N_10808);
nor U11022 (N_11022,N_10856,N_10725);
or U11023 (N_11023,N_10873,N_10819);
xor U11024 (N_11024,N_10864,N_10720);
nand U11025 (N_11025,N_10807,N_10736);
xnor U11026 (N_11026,N_10738,N_10808);
xnor U11027 (N_11027,N_10860,N_10794);
or U11028 (N_11028,N_10738,N_10758);
nand U11029 (N_11029,N_10818,N_10812);
nor U11030 (N_11030,N_10837,N_10824);
or U11031 (N_11031,N_10833,N_10849);
nand U11032 (N_11032,N_10845,N_10879);
nor U11033 (N_11033,N_10751,N_10788);
xnor U11034 (N_11034,N_10793,N_10822);
or U11035 (N_11035,N_10739,N_10810);
or U11036 (N_11036,N_10826,N_10745);
nand U11037 (N_11037,N_10829,N_10760);
nand U11038 (N_11038,N_10814,N_10779);
nor U11039 (N_11039,N_10747,N_10857);
xor U11040 (N_11040,N_10996,N_10889);
and U11041 (N_11041,N_11009,N_10928);
xnor U11042 (N_11042,N_10979,N_10957);
nor U11043 (N_11043,N_10927,N_11002);
and U11044 (N_11044,N_11036,N_10967);
xnor U11045 (N_11045,N_10906,N_10891);
and U11046 (N_11046,N_11027,N_10946);
xnor U11047 (N_11047,N_10915,N_11033);
and U11048 (N_11048,N_10969,N_10975);
xor U11049 (N_11049,N_10907,N_10948);
or U11050 (N_11050,N_10908,N_11032);
nor U11051 (N_11051,N_11035,N_10963);
or U11052 (N_11052,N_10960,N_10893);
or U11053 (N_11053,N_10880,N_10914);
or U11054 (N_11054,N_11013,N_10972);
and U11055 (N_11055,N_10993,N_10973);
nor U11056 (N_11056,N_10986,N_10929);
or U11057 (N_11057,N_10925,N_11001);
nor U11058 (N_11058,N_10989,N_10970);
or U11059 (N_11059,N_10899,N_11024);
nand U11060 (N_11060,N_11031,N_10951);
nor U11061 (N_11061,N_10949,N_10933);
and U11062 (N_11062,N_10981,N_11010);
nand U11063 (N_11063,N_11012,N_10945);
xnor U11064 (N_11064,N_10964,N_10994);
or U11065 (N_11065,N_10987,N_11015);
or U11066 (N_11066,N_10913,N_11017);
or U11067 (N_11067,N_11025,N_10898);
nand U11068 (N_11068,N_10953,N_11008);
nor U11069 (N_11069,N_11016,N_10944);
or U11070 (N_11070,N_10926,N_10980);
and U11071 (N_11071,N_10974,N_10905);
or U11072 (N_11072,N_11006,N_10930);
and U11073 (N_11073,N_10968,N_10937);
or U11074 (N_11074,N_11021,N_10942);
or U11075 (N_11075,N_10995,N_10954);
or U11076 (N_11076,N_10904,N_10940);
xor U11077 (N_11077,N_10901,N_11039);
nor U11078 (N_11078,N_10936,N_10971);
and U11079 (N_11079,N_10956,N_10982);
nor U11080 (N_11080,N_10999,N_10932);
and U11081 (N_11081,N_11029,N_11003);
or U11082 (N_11082,N_10884,N_10911);
xnor U11083 (N_11083,N_10881,N_10984);
xor U11084 (N_11084,N_10966,N_11028);
xnor U11085 (N_11085,N_10941,N_11026);
nand U11086 (N_11086,N_11037,N_10988);
and U11087 (N_11087,N_11034,N_10983);
or U11088 (N_11088,N_10958,N_10895);
xnor U11089 (N_11089,N_11022,N_10977);
or U11090 (N_11090,N_11038,N_10947);
nor U11091 (N_11091,N_10931,N_10950);
xor U11092 (N_11092,N_10902,N_11014);
nor U11093 (N_11093,N_10903,N_10919);
and U11094 (N_11094,N_10978,N_10961);
or U11095 (N_11095,N_10990,N_11020);
xnor U11096 (N_11096,N_10985,N_10943);
xor U11097 (N_11097,N_11000,N_10959);
xnor U11098 (N_11098,N_10955,N_11005);
xor U11099 (N_11099,N_10888,N_10886);
nand U11100 (N_11100,N_10917,N_11011);
or U11101 (N_11101,N_10887,N_10997);
xnor U11102 (N_11102,N_10912,N_11030);
and U11103 (N_11103,N_10976,N_10900);
xor U11104 (N_11104,N_11023,N_10885);
nand U11105 (N_11105,N_10924,N_11019);
nand U11106 (N_11106,N_10962,N_10935);
and U11107 (N_11107,N_11018,N_10882);
nor U11108 (N_11108,N_10923,N_10894);
or U11109 (N_11109,N_10921,N_10910);
or U11110 (N_11110,N_10909,N_10920);
nor U11111 (N_11111,N_10892,N_10952);
or U11112 (N_11112,N_10890,N_10896);
or U11113 (N_11113,N_10998,N_10916);
or U11114 (N_11114,N_10991,N_11007);
nor U11115 (N_11115,N_10992,N_10883);
xnor U11116 (N_11116,N_10922,N_10965);
or U11117 (N_11117,N_10934,N_11004);
and U11118 (N_11118,N_10939,N_10938);
nand U11119 (N_11119,N_10897,N_10918);
nand U11120 (N_11120,N_10972,N_11028);
and U11121 (N_11121,N_10962,N_11034);
nor U11122 (N_11122,N_10911,N_11028);
or U11123 (N_11123,N_10904,N_11010);
xnor U11124 (N_11124,N_10979,N_10983);
nor U11125 (N_11125,N_10970,N_10967);
nor U11126 (N_11126,N_11018,N_11034);
nand U11127 (N_11127,N_10950,N_10949);
nor U11128 (N_11128,N_11036,N_10885);
nand U11129 (N_11129,N_10940,N_10981);
or U11130 (N_11130,N_10880,N_10980);
or U11131 (N_11131,N_10898,N_10953);
xor U11132 (N_11132,N_10967,N_10950);
nand U11133 (N_11133,N_10891,N_11001);
and U11134 (N_11134,N_10980,N_10959);
xor U11135 (N_11135,N_10934,N_10944);
nor U11136 (N_11136,N_10888,N_10913);
xor U11137 (N_11137,N_10939,N_10941);
nor U11138 (N_11138,N_10960,N_10967);
nand U11139 (N_11139,N_10951,N_10999);
nor U11140 (N_11140,N_11027,N_10914);
or U11141 (N_11141,N_11010,N_10937);
nor U11142 (N_11142,N_11012,N_10999);
or U11143 (N_11143,N_10970,N_10918);
xor U11144 (N_11144,N_11039,N_10905);
xor U11145 (N_11145,N_10932,N_10915);
and U11146 (N_11146,N_10957,N_10940);
xor U11147 (N_11147,N_10918,N_10978);
nor U11148 (N_11148,N_10908,N_10883);
nand U11149 (N_11149,N_11002,N_10900);
nand U11150 (N_11150,N_10936,N_10996);
or U11151 (N_11151,N_10979,N_11019);
nand U11152 (N_11152,N_10946,N_10885);
xnor U11153 (N_11153,N_10889,N_10993);
and U11154 (N_11154,N_10968,N_10989);
and U11155 (N_11155,N_10939,N_11001);
or U11156 (N_11156,N_10885,N_10921);
nand U11157 (N_11157,N_10971,N_10933);
and U11158 (N_11158,N_10939,N_11006);
nand U11159 (N_11159,N_10983,N_10963);
xnor U11160 (N_11160,N_10994,N_11034);
and U11161 (N_11161,N_10951,N_10946);
xnor U11162 (N_11162,N_10897,N_10942);
xnor U11163 (N_11163,N_10956,N_10991);
xor U11164 (N_11164,N_10941,N_10928);
nor U11165 (N_11165,N_11015,N_10883);
or U11166 (N_11166,N_11023,N_10981);
nor U11167 (N_11167,N_10942,N_10985);
nand U11168 (N_11168,N_10920,N_10995);
or U11169 (N_11169,N_10887,N_10938);
nor U11170 (N_11170,N_11004,N_10988);
nand U11171 (N_11171,N_11025,N_11008);
xnor U11172 (N_11172,N_11004,N_11008);
or U11173 (N_11173,N_11015,N_11017);
or U11174 (N_11174,N_10892,N_10906);
and U11175 (N_11175,N_10996,N_10989);
nor U11176 (N_11176,N_11025,N_10965);
xnor U11177 (N_11177,N_10965,N_10886);
nand U11178 (N_11178,N_10907,N_10938);
nand U11179 (N_11179,N_10943,N_10958);
or U11180 (N_11180,N_10916,N_11033);
nor U11181 (N_11181,N_11034,N_10955);
and U11182 (N_11182,N_10938,N_10895);
or U11183 (N_11183,N_10957,N_11022);
nor U11184 (N_11184,N_10941,N_10969);
xor U11185 (N_11185,N_10887,N_10993);
xnor U11186 (N_11186,N_10936,N_10937);
nand U11187 (N_11187,N_10974,N_10887);
nand U11188 (N_11188,N_10970,N_10966);
xor U11189 (N_11189,N_11038,N_10979);
nand U11190 (N_11190,N_10910,N_10951);
or U11191 (N_11191,N_10911,N_10948);
or U11192 (N_11192,N_10995,N_11030);
nor U11193 (N_11193,N_10992,N_11028);
xor U11194 (N_11194,N_10967,N_10986);
nand U11195 (N_11195,N_10958,N_11033);
nor U11196 (N_11196,N_10887,N_11020);
nor U11197 (N_11197,N_10956,N_10960);
xnor U11198 (N_11198,N_10996,N_11004);
or U11199 (N_11199,N_11010,N_10920);
nor U11200 (N_11200,N_11091,N_11148);
xor U11201 (N_11201,N_11157,N_11102);
and U11202 (N_11202,N_11173,N_11099);
xnor U11203 (N_11203,N_11181,N_11196);
nand U11204 (N_11204,N_11087,N_11176);
or U11205 (N_11205,N_11083,N_11198);
xnor U11206 (N_11206,N_11060,N_11160);
and U11207 (N_11207,N_11130,N_11076);
nor U11208 (N_11208,N_11117,N_11104);
and U11209 (N_11209,N_11109,N_11180);
and U11210 (N_11210,N_11077,N_11186);
nor U11211 (N_11211,N_11053,N_11171);
or U11212 (N_11212,N_11151,N_11079);
or U11213 (N_11213,N_11161,N_11075);
nand U11214 (N_11214,N_11058,N_11155);
nand U11215 (N_11215,N_11068,N_11066);
nand U11216 (N_11216,N_11140,N_11044);
or U11217 (N_11217,N_11048,N_11191);
nand U11218 (N_11218,N_11074,N_11110);
nand U11219 (N_11219,N_11067,N_11197);
and U11220 (N_11220,N_11051,N_11065);
xnor U11221 (N_11221,N_11118,N_11111);
and U11222 (N_11222,N_11187,N_11081);
and U11223 (N_11223,N_11142,N_11199);
xor U11224 (N_11224,N_11159,N_11049);
or U11225 (N_11225,N_11092,N_11139);
xor U11226 (N_11226,N_11093,N_11095);
or U11227 (N_11227,N_11178,N_11073);
and U11228 (N_11228,N_11138,N_11125);
xor U11229 (N_11229,N_11047,N_11128);
and U11230 (N_11230,N_11040,N_11189);
and U11231 (N_11231,N_11041,N_11156);
or U11232 (N_11232,N_11094,N_11135);
xnor U11233 (N_11233,N_11175,N_11107);
or U11234 (N_11234,N_11165,N_11054);
nand U11235 (N_11235,N_11114,N_11120);
xor U11236 (N_11236,N_11063,N_11133);
or U11237 (N_11237,N_11174,N_11062);
xnor U11238 (N_11238,N_11136,N_11042);
xor U11239 (N_11239,N_11082,N_11069);
xnor U11240 (N_11240,N_11131,N_11134);
nand U11241 (N_11241,N_11106,N_11123);
nor U11242 (N_11242,N_11055,N_11192);
nand U11243 (N_11243,N_11097,N_11052);
or U11244 (N_11244,N_11124,N_11112);
and U11245 (N_11245,N_11177,N_11144);
xnor U11246 (N_11246,N_11085,N_11098);
xnor U11247 (N_11247,N_11183,N_11096);
xor U11248 (N_11248,N_11056,N_11050);
nand U11249 (N_11249,N_11129,N_11162);
and U11250 (N_11250,N_11149,N_11141);
nand U11251 (N_11251,N_11152,N_11184);
or U11252 (N_11252,N_11127,N_11119);
nand U11253 (N_11253,N_11170,N_11046);
and U11254 (N_11254,N_11057,N_11088);
nor U11255 (N_11255,N_11150,N_11145);
nor U11256 (N_11256,N_11147,N_11108);
or U11257 (N_11257,N_11121,N_11137);
and U11258 (N_11258,N_11070,N_11154);
nor U11259 (N_11259,N_11168,N_11193);
nand U11260 (N_11260,N_11061,N_11146);
xor U11261 (N_11261,N_11071,N_11080);
or U11262 (N_11262,N_11126,N_11143);
nor U11263 (N_11263,N_11169,N_11072);
or U11264 (N_11264,N_11166,N_11116);
or U11265 (N_11265,N_11194,N_11195);
and U11266 (N_11266,N_11172,N_11132);
or U11267 (N_11267,N_11043,N_11167);
xor U11268 (N_11268,N_11158,N_11078);
and U11269 (N_11269,N_11089,N_11101);
nand U11270 (N_11270,N_11084,N_11105);
and U11271 (N_11271,N_11103,N_11090);
or U11272 (N_11272,N_11100,N_11190);
xor U11273 (N_11273,N_11164,N_11045);
xnor U11274 (N_11274,N_11086,N_11122);
nand U11275 (N_11275,N_11182,N_11113);
nor U11276 (N_11276,N_11059,N_11064);
xnor U11277 (N_11277,N_11163,N_11188);
xor U11278 (N_11278,N_11185,N_11153);
or U11279 (N_11279,N_11115,N_11179);
nand U11280 (N_11280,N_11042,N_11094);
nand U11281 (N_11281,N_11130,N_11053);
xor U11282 (N_11282,N_11192,N_11193);
and U11283 (N_11283,N_11075,N_11109);
nor U11284 (N_11284,N_11194,N_11116);
nand U11285 (N_11285,N_11124,N_11117);
and U11286 (N_11286,N_11196,N_11135);
nor U11287 (N_11287,N_11113,N_11082);
nand U11288 (N_11288,N_11165,N_11113);
nor U11289 (N_11289,N_11084,N_11199);
and U11290 (N_11290,N_11139,N_11185);
and U11291 (N_11291,N_11123,N_11117);
nor U11292 (N_11292,N_11121,N_11199);
nand U11293 (N_11293,N_11047,N_11073);
or U11294 (N_11294,N_11051,N_11066);
nor U11295 (N_11295,N_11087,N_11082);
or U11296 (N_11296,N_11052,N_11135);
nand U11297 (N_11297,N_11079,N_11192);
or U11298 (N_11298,N_11057,N_11124);
nand U11299 (N_11299,N_11164,N_11079);
nor U11300 (N_11300,N_11133,N_11065);
and U11301 (N_11301,N_11158,N_11044);
or U11302 (N_11302,N_11075,N_11108);
and U11303 (N_11303,N_11118,N_11090);
xnor U11304 (N_11304,N_11174,N_11166);
xnor U11305 (N_11305,N_11187,N_11178);
nor U11306 (N_11306,N_11172,N_11089);
and U11307 (N_11307,N_11180,N_11077);
and U11308 (N_11308,N_11139,N_11084);
and U11309 (N_11309,N_11146,N_11063);
nor U11310 (N_11310,N_11064,N_11170);
or U11311 (N_11311,N_11091,N_11177);
or U11312 (N_11312,N_11086,N_11062);
nor U11313 (N_11313,N_11054,N_11162);
nor U11314 (N_11314,N_11139,N_11193);
xor U11315 (N_11315,N_11099,N_11102);
xnor U11316 (N_11316,N_11156,N_11123);
or U11317 (N_11317,N_11177,N_11088);
xor U11318 (N_11318,N_11058,N_11099);
nor U11319 (N_11319,N_11121,N_11075);
nand U11320 (N_11320,N_11094,N_11193);
and U11321 (N_11321,N_11050,N_11091);
nand U11322 (N_11322,N_11136,N_11109);
nor U11323 (N_11323,N_11167,N_11161);
or U11324 (N_11324,N_11194,N_11068);
xnor U11325 (N_11325,N_11085,N_11149);
and U11326 (N_11326,N_11186,N_11068);
or U11327 (N_11327,N_11191,N_11154);
nand U11328 (N_11328,N_11050,N_11185);
nand U11329 (N_11329,N_11079,N_11179);
and U11330 (N_11330,N_11076,N_11120);
or U11331 (N_11331,N_11127,N_11147);
xnor U11332 (N_11332,N_11146,N_11092);
and U11333 (N_11333,N_11148,N_11155);
nand U11334 (N_11334,N_11089,N_11134);
nand U11335 (N_11335,N_11058,N_11162);
and U11336 (N_11336,N_11134,N_11173);
and U11337 (N_11337,N_11120,N_11157);
and U11338 (N_11338,N_11072,N_11130);
and U11339 (N_11339,N_11105,N_11163);
nor U11340 (N_11340,N_11072,N_11193);
nor U11341 (N_11341,N_11167,N_11076);
nand U11342 (N_11342,N_11065,N_11110);
nand U11343 (N_11343,N_11074,N_11118);
and U11344 (N_11344,N_11100,N_11046);
nor U11345 (N_11345,N_11125,N_11111);
or U11346 (N_11346,N_11061,N_11180);
and U11347 (N_11347,N_11193,N_11129);
or U11348 (N_11348,N_11121,N_11176);
nor U11349 (N_11349,N_11099,N_11093);
nand U11350 (N_11350,N_11180,N_11184);
nor U11351 (N_11351,N_11071,N_11113);
nand U11352 (N_11352,N_11185,N_11049);
nor U11353 (N_11353,N_11150,N_11078);
and U11354 (N_11354,N_11069,N_11110);
or U11355 (N_11355,N_11167,N_11143);
nor U11356 (N_11356,N_11154,N_11040);
nor U11357 (N_11357,N_11056,N_11095);
or U11358 (N_11358,N_11168,N_11061);
and U11359 (N_11359,N_11054,N_11155);
or U11360 (N_11360,N_11243,N_11244);
or U11361 (N_11361,N_11258,N_11262);
xnor U11362 (N_11362,N_11304,N_11238);
or U11363 (N_11363,N_11303,N_11297);
and U11364 (N_11364,N_11336,N_11346);
nand U11365 (N_11365,N_11237,N_11224);
and U11366 (N_11366,N_11259,N_11285);
and U11367 (N_11367,N_11225,N_11327);
or U11368 (N_11368,N_11232,N_11354);
nand U11369 (N_11369,N_11350,N_11203);
nand U11370 (N_11370,N_11208,N_11226);
xnor U11371 (N_11371,N_11293,N_11311);
and U11372 (N_11372,N_11313,N_11269);
xor U11373 (N_11373,N_11248,N_11287);
or U11374 (N_11374,N_11256,N_11289);
or U11375 (N_11375,N_11318,N_11267);
xnor U11376 (N_11376,N_11266,N_11206);
xnor U11377 (N_11377,N_11321,N_11342);
xnor U11378 (N_11378,N_11337,N_11257);
or U11379 (N_11379,N_11273,N_11218);
and U11380 (N_11380,N_11331,N_11216);
nor U11381 (N_11381,N_11275,N_11341);
and U11382 (N_11382,N_11205,N_11290);
nor U11383 (N_11383,N_11295,N_11250);
or U11384 (N_11384,N_11357,N_11310);
nor U11385 (N_11385,N_11242,N_11358);
and U11386 (N_11386,N_11277,N_11325);
nand U11387 (N_11387,N_11333,N_11211);
nor U11388 (N_11388,N_11322,N_11316);
or U11389 (N_11389,N_11209,N_11200);
nand U11390 (N_11390,N_11235,N_11264);
nand U11391 (N_11391,N_11344,N_11340);
and U11392 (N_11392,N_11249,N_11260);
xnor U11393 (N_11393,N_11241,N_11219);
and U11394 (N_11394,N_11351,N_11312);
or U11395 (N_11395,N_11348,N_11320);
nand U11396 (N_11396,N_11306,N_11230);
or U11397 (N_11397,N_11272,N_11292);
xnor U11398 (N_11398,N_11246,N_11229);
xnor U11399 (N_11399,N_11210,N_11301);
and U11400 (N_11400,N_11314,N_11247);
xnor U11401 (N_11401,N_11296,N_11233);
or U11402 (N_11402,N_11339,N_11240);
nand U11403 (N_11403,N_11212,N_11239);
or U11404 (N_11404,N_11279,N_11352);
and U11405 (N_11405,N_11284,N_11234);
and U11406 (N_11406,N_11328,N_11265);
nor U11407 (N_11407,N_11245,N_11355);
and U11408 (N_11408,N_11270,N_11231);
nor U11409 (N_11409,N_11254,N_11345);
nand U11410 (N_11410,N_11326,N_11215);
xnor U11411 (N_11411,N_11323,N_11201);
nor U11412 (N_11412,N_11283,N_11222);
or U11413 (N_11413,N_11281,N_11299);
xor U11414 (N_11414,N_11288,N_11204);
and U11415 (N_11415,N_11338,N_11280);
or U11416 (N_11416,N_11319,N_11308);
or U11417 (N_11417,N_11347,N_11276);
nand U11418 (N_11418,N_11263,N_11307);
and U11419 (N_11419,N_11252,N_11291);
nand U11420 (N_11420,N_11220,N_11286);
nand U11421 (N_11421,N_11298,N_11282);
nand U11422 (N_11422,N_11300,N_11223);
nor U11423 (N_11423,N_11329,N_11334);
or U11424 (N_11424,N_11294,N_11317);
nand U11425 (N_11425,N_11202,N_11278);
and U11426 (N_11426,N_11255,N_11353);
nand U11427 (N_11427,N_11274,N_11302);
nand U11428 (N_11428,N_11268,N_11253);
nor U11429 (N_11429,N_11359,N_11213);
nor U11430 (N_11430,N_11356,N_11221);
xnor U11431 (N_11431,N_11330,N_11227);
or U11432 (N_11432,N_11217,N_11207);
nand U11433 (N_11433,N_11349,N_11261);
nor U11434 (N_11434,N_11251,N_11343);
xnor U11435 (N_11435,N_11335,N_11305);
nor U11436 (N_11436,N_11271,N_11309);
nand U11437 (N_11437,N_11214,N_11236);
nand U11438 (N_11438,N_11324,N_11332);
and U11439 (N_11439,N_11228,N_11315);
xor U11440 (N_11440,N_11279,N_11344);
and U11441 (N_11441,N_11284,N_11212);
and U11442 (N_11442,N_11307,N_11220);
nor U11443 (N_11443,N_11208,N_11347);
nand U11444 (N_11444,N_11277,N_11223);
nor U11445 (N_11445,N_11341,N_11203);
or U11446 (N_11446,N_11321,N_11215);
nand U11447 (N_11447,N_11322,N_11294);
nand U11448 (N_11448,N_11346,N_11330);
nand U11449 (N_11449,N_11291,N_11315);
xnor U11450 (N_11450,N_11220,N_11224);
or U11451 (N_11451,N_11202,N_11353);
and U11452 (N_11452,N_11287,N_11275);
xnor U11453 (N_11453,N_11208,N_11277);
xor U11454 (N_11454,N_11239,N_11358);
nand U11455 (N_11455,N_11234,N_11255);
and U11456 (N_11456,N_11277,N_11212);
nor U11457 (N_11457,N_11242,N_11216);
and U11458 (N_11458,N_11327,N_11347);
xnor U11459 (N_11459,N_11224,N_11357);
nor U11460 (N_11460,N_11285,N_11276);
nand U11461 (N_11461,N_11316,N_11312);
nand U11462 (N_11462,N_11335,N_11242);
and U11463 (N_11463,N_11276,N_11342);
xor U11464 (N_11464,N_11238,N_11340);
nor U11465 (N_11465,N_11313,N_11231);
or U11466 (N_11466,N_11346,N_11266);
nand U11467 (N_11467,N_11273,N_11325);
xor U11468 (N_11468,N_11257,N_11245);
nor U11469 (N_11469,N_11339,N_11306);
and U11470 (N_11470,N_11220,N_11314);
nor U11471 (N_11471,N_11333,N_11221);
or U11472 (N_11472,N_11237,N_11243);
and U11473 (N_11473,N_11246,N_11270);
xor U11474 (N_11474,N_11257,N_11332);
xor U11475 (N_11475,N_11286,N_11232);
or U11476 (N_11476,N_11292,N_11355);
nor U11477 (N_11477,N_11272,N_11241);
or U11478 (N_11478,N_11253,N_11350);
nor U11479 (N_11479,N_11317,N_11249);
nand U11480 (N_11480,N_11258,N_11353);
or U11481 (N_11481,N_11351,N_11356);
or U11482 (N_11482,N_11283,N_11225);
nand U11483 (N_11483,N_11259,N_11338);
or U11484 (N_11484,N_11200,N_11286);
xnor U11485 (N_11485,N_11318,N_11333);
nor U11486 (N_11486,N_11227,N_11221);
or U11487 (N_11487,N_11216,N_11293);
and U11488 (N_11488,N_11315,N_11335);
nor U11489 (N_11489,N_11310,N_11247);
or U11490 (N_11490,N_11305,N_11351);
and U11491 (N_11491,N_11335,N_11285);
xor U11492 (N_11492,N_11290,N_11317);
xnor U11493 (N_11493,N_11310,N_11216);
or U11494 (N_11494,N_11301,N_11351);
xor U11495 (N_11495,N_11338,N_11251);
and U11496 (N_11496,N_11300,N_11322);
nand U11497 (N_11497,N_11359,N_11229);
nor U11498 (N_11498,N_11301,N_11296);
nand U11499 (N_11499,N_11276,N_11270);
and U11500 (N_11500,N_11341,N_11244);
and U11501 (N_11501,N_11298,N_11284);
or U11502 (N_11502,N_11289,N_11299);
and U11503 (N_11503,N_11359,N_11257);
or U11504 (N_11504,N_11271,N_11330);
and U11505 (N_11505,N_11243,N_11320);
nor U11506 (N_11506,N_11202,N_11331);
xor U11507 (N_11507,N_11235,N_11276);
nand U11508 (N_11508,N_11321,N_11251);
nand U11509 (N_11509,N_11238,N_11205);
xnor U11510 (N_11510,N_11275,N_11264);
or U11511 (N_11511,N_11330,N_11209);
nand U11512 (N_11512,N_11256,N_11209);
or U11513 (N_11513,N_11293,N_11331);
and U11514 (N_11514,N_11311,N_11357);
nand U11515 (N_11515,N_11348,N_11218);
or U11516 (N_11516,N_11261,N_11303);
nand U11517 (N_11517,N_11201,N_11271);
or U11518 (N_11518,N_11286,N_11351);
or U11519 (N_11519,N_11242,N_11231);
nor U11520 (N_11520,N_11445,N_11449);
and U11521 (N_11521,N_11380,N_11406);
nand U11522 (N_11522,N_11407,N_11458);
nor U11523 (N_11523,N_11501,N_11383);
nand U11524 (N_11524,N_11486,N_11518);
xor U11525 (N_11525,N_11479,N_11370);
and U11526 (N_11526,N_11457,N_11361);
nand U11527 (N_11527,N_11425,N_11382);
xnor U11528 (N_11528,N_11469,N_11417);
or U11529 (N_11529,N_11442,N_11477);
xor U11530 (N_11530,N_11405,N_11426);
and U11531 (N_11531,N_11438,N_11395);
nand U11532 (N_11532,N_11429,N_11385);
xor U11533 (N_11533,N_11362,N_11456);
xor U11534 (N_11534,N_11419,N_11423);
xnor U11535 (N_11535,N_11388,N_11513);
nor U11536 (N_11536,N_11495,N_11399);
or U11537 (N_11537,N_11367,N_11428);
and U11538 (N_11538,N_11492,N_11500);
or U11539 (N_11539,N_11494,N_11448);
or U11540 (N_11540,N_11422,N_11483);
xor U11541 (N_11541,N_11424,N_11410);
nand U11542 (N_11542,N_11474,N_11489);
nor U11543 (N_11543,N_11390,N_11514);
nor U11544 (N_11544,N_11368,N_11439);
and U11545 (N_11545,N_11502,N_11369);
nor U11546 (N_11546,N_11432,N_11476);
xnor U11547 (N_11547,N_11508,N_11412);
nand U11548 (N_11548,N_11505,N_11499);
nor U11549 (N_11549,N_11487,N_11393);
or U11550 (N_11550,N_11462,N_11427);
or U11551 (N_11551,N_11365,N_11491);
xor U11552 (N_11552,N_11484,N_11481);
nand U11553 (N_11553,N_11416,N_11374);
or U11554 (N_11554,N_11467,N_11517);
or U11555 (N_11555,N_11409,N_11397);
or U11556 (N_11556,N_11459,N_11444);
nand U11557 (N_11557,N_11404,N_11435);
and U11558 (N_11558,N_11375,N_11391);
nand U11559 (N_11559,N_11377,N_11516);
and U11560 (N_11560,N_11387,N_11400);
and U11561 (N_11561,N_11381,N_11447);
nor U11562 (N_11562,N_11455,N_11446);
or U11563 (N_11563,N_11408,N_11394);
xor U11564 (N_11564,N_11401,N_11496);
and U11565 (N_11565,N_11434,N_11504);
and U11566 (N_11566,N_11403,N_11468);
and U11567 (N_11567,N_11515,N_11450);
nand U11568 (N_11568,N_11413,N_11473);
xnor U11569 (N_11569,N_11360,N_11437);
xnor U11570 (N_11570,N_11463,N_11414);
and U11571 (N_11571,N_11373,N_11480);
nor U11572 (N_11572,N_11436,N_11418);
and U11573 (N_11573,N_11415,N_11372);
nor U11574 (N_11574,N_11379,N_11493);
or U11575 (N_11575,N_11398,N_11512);
nand U11576 (N_11576,N_11460,N_11509);
or U11577 (N_11577,N_11490,N_11364);
nor U11578 (N_11578,N_11478,N_11511);
nand U11579 (N_11579,N_11396,N_11475);
nand U11580 (N_11580,N_11378,N_11366);
and U11581 (N_11581,N_11411,N_11466);
and U11582 (N_11582,N_11443,N_11441);
xnor U11583 (N_11583,N_11497,N_11498);
or U11584 (N_11584,N_11519,N_11451);
xor U11585 (N_11585,N_11421,N_11363);
xor U11586 (N_11586,N_11452,N_11371);
xor U11587 (N_11587,N_11389,N_11461);
xnor U11588 (N_11588,N_11453,N_11482);
nand U11589 (N_11589,N_11420,N_11464);
and U11590 (N_11590,N_11384,N_11440);
and U11591 (N_11591,N_11503,N_11488);
nor U11592 (N_11592,N_11471,N_11454);
nor U11593 (N_11593,N_11376,N_11507);
nor U11594 (N_11594,N_11472,N_11402);
nor U11595 (N_11595,N_11485,N_11465);
nor U11596 (N_11596,N_11510,N_11392);
or U11597 (N_11597,N_11470,N_11506);
xnor U11598 (N_11598,N_11430,N_11431);
and U11599 (N_11599,N_11433,N_11386);
nand U11600 (N_11600,N_11468,N_11491);
nor U11601 (N_11601,N_11368,N_11511);
nor U11602 (N_11602,N_11501,N_11408);
and U11603 (N_11603,N_11491,N_11487);
nor U11604 (N_11604,N_11452,N_11488);
nand U11605 (N_11605,N_11514,N_11494);
and U11606 (N_11606,N_11467,N_11515);
nor U11607 (N_11607,N_11462,N_11390);
and U11608 (N_11608,N_11511,N_11388);
and U11609 (N_11609,N_11361,N_11486);
nor U11610 (N_11610,N_11427,N_11450);
nor U11611 (N_11611,N_11494,N_11381);
xor U11612 (N_11612,N_11369,N_11504);
xnor U11613 (N_11613,N_11402,N_11498);
xor U11614 (N_11614,N_11463,N_11383);
nand U11615 (N_11615,N_11510,N_11518);
xor U11616 (N_11616,N_11424,N_11457);
nor U11617 (N_11617,N_11485,N_11412);
xor U11618 (N_11618,N_11490,N_11451);
nor U11619 (N_11619,N_11484,N_11399);
nand U11620 (N_11620,N_11373,N_11424);
or U11621 (N_11621,N_11395,N_11502);
xor U11622 (N_11622,N_11466,N_11425);
or U11623 (N_11623,N_11438,N_11378);
or U11624 (N_11624,N_11363,N_11370);
nand U11625 (N_11625,N_11503,N_11497);
xor U11626 (N_11626,N_11395,N_11375);
xnor U11627 (N_11627,N_11393,N_11365);
nor U11628 (N_11628,N_11405,N_11516);
nand U11629 (N_11629,N_11511,N_11463);
nand U11630 (N_11630,N_11488,N_11444);
nor U11631 (N_11631,N_11379,N_11519);
or U11632 (N_11632,N_11408,N_11461);
or U11633 (N_11633,N_11422,N_11397);
and U11634 (N_11634,N_11503,N_11432);
and U11635 (N_11635,N_11388,N_11449);
nor U11636 (N_11636,N_11463,N_11428);
xor U11637 (N_11637,N_11445,N_11472);
and U11638 (N_11638,N_11488,N_11406);
nor U11639 (N_11639,N_11421,N_11408);
and U11640 (N_11640,N_11400,N_11435);
and U11641 (N_11641,N_11433,N_11478);
and U11642 (N_11642,N_11385,N_11432);
xnor U11643 (N_11643,N_11376,N_11515);
xnor U11644 (N_11644,N_11459,N_11410);
or U11645 (N_11645,N_11487,N_11398);
and U11646 (N_11646,N_11465,N_11427);
nor U11647 (N_11647,N_11387,N_11502);
or U11648 (N_11648,N_11443,N_11509);
nand U11649 (N_11649,N_11492,N_11426);
and U11650 (N_11650,N_11415,N_11431);
nand U11651 (N_11651,N_11516,N_11457);
nand U11652 (N_11652,N_11423,N_11410);
nand U11653 (N_11653,N_11441,N_11497);
xor U11654 (N_11654,N_11454,N_11376);
nor U11655 (N_11655,N_11378,N_11420);
xnor U11656 (N_11656,N_11361,N_11493);
and U11657 (N_11657,N_11369,N_11511);
nand U11658 (N_11658,N_11475,N_11360);
or U11659 (N_11659,N_11378,N_11502);
or U11660 (N_11660,N_11490,N_11456);
xnor U11661 (N_11661,N_11376,N_11435);
or U11662 (N_11662,N_11501,N_11369);
nand U11663 (N_11663,N_11413,N_11410);
nand U11664 (N_11664,N_11439,N_11401);
and U11665 (N_11665,N_11483,N_11370);
nand U11666 (N_11666,N_11438,N_11461);
xor U11667 (N_11667,N_11449,N_11465);
and U11668 (N_11668,N_11486,N_11441);
and U11669 (N_11669,N_11390,N_11384);
and U11670 (N_11670,N_11399,N_11396);
and U11671 (N_11671,N_11494,N_11511);
nand U11672 (N_11672,N_11485,N_11476);
nor U11673 (N_11673,N_11468,N_11432);
nor U11674 (N_11674,N_11427,N_11417);
or U11675 (N_11675,N_11369,N_11363);
nand U11676 (N_11676,N_11451,N_11486);
xor U11677 (N_11677,N_11447,N_11390);
nand U11678 (N_11678,N_11406,N_11385);
and U11679 (N_11679,N_11457,N_11449);
nand U11680 (N_11680,N_11672,N_11544);
nand U11681 (N_11681,N_11556,N_11676);
nor U11682 (N_11682,N_11520,N_11615);
or U11683 (N_11683,N_11667,N_11578);
or U11684 (N_11684,N_11633,N_11576);
nand U11685 (N_11685,N_11524,N_11634);
xnor U11686 (N_11686,N_11564,N_11668);
nand U11687 (N_11687,N_11596,N_11553);
nor U11688 (N_11688,N_11612,N_11588);
or U11689 (N_11689,N_11525,N_11542);
or U11690 (N_11690,N_11572,N_11597);
or U11691 (N_11691,N_11539,N_11593);
nor U11692 (N_11692,N_11563,N_11577);
and U11693 (N_11693,N_11656,N_11650);
xor U11694 (N_11694,N_11534,N_11529);
xnor U11695 (N_11695,N_11671,N_11620);
or U11696 (N_11696,N_11674,N_11666);
nor U11697 (N_11697,N_11590,N_11624);
nand U11698 (N_11698,N_11603,N_11533);
or U11699 (N_11699,N_11579,N_11643);
nor U11700 (N_11700,N_11611,N_11554);
or U11701 (N_11701,N_11558,N_11653);
nor U11702 (N_11702,N_11561,N_11531);
nand U11703 (N_11703,N_11607,N_11616);
nor U11704 (N_11704,N_11655,N_11657);
nor U11705 (N_11705,N_11566,N_11550);
nor U11706 (N_11706,N_11568,N_11625);
and U11707 (N_11707,N_11573,N_11608);
and U11708 (N_11708,N_11582,N_11585);
or U11709 (N_11709,N_11548,N_11545);
and U11710 (N_11710,N_11673,N_11535);
nor U11711 (N_11711,N_11654,N_11532);
or U11712 (N_11712,N_11587,N_11583);
xor U11713 (N_11713,N_11647,N_11543);
xnor U11714 (N_11714,N_11557,N_11637);
nor U11715 (N_11715,N_11523,N_11559);
xnor U11716 (N_11716,N_11600,N_11640);
and U11717 (N_11717,N_11522,N_11549);
or U11718 (N_11718,N_11644,N_11575);
nor U11719 (N_11719,N_11599,N_11536);
nor U11720 (N_11720,N_11530,N_11677);
or U11721 (N_11721,N_11613,N_11630);
and U11722 (N_11722,N_11580,N_11661);
or U11723 (N_11723,N_11646,N_11649);
nor U11724 (N_11724,N_11628,N_11675);
nor U11725 (N_11725,N_11619,N_11632);
nor U11726 (N_11726,N_11614,N_11595);
xnor U11727 (N_11727,N_11598,N_11562);
or U11728 (N_11728,N_11669,N_11605);
nor U11729 (N_11729,N_11581,N_11629);
xnor U11730 (N_11730,N_11658,N_11670);
and U11731 (N_11731,N_11538,N_11665);
nor U11732 (N_11732,N_11592,N_11610);
xnor U11733 (N_11733,N_11622,N_11623);
nor U11734 (N_11734,N_11526,N_11567);
xor U11735 (N_11735,N_11636,N_11540);
or U11736 (N_11736,N_11546,N_11601);
and U11737 (N_11737,N_11541,N_11552);
xor U11738 (N_11738,N_11621,N_11638);
and U11739 (N_11739,N_11660,N_11589);
or U11740 (N_11740,N_11602,N_11662);
nor U11741 (N_11741,N_11547,N_11664);
nor U11742 (N_11742,N_11606,N_11635);
nand U11743 (N_11743,N_11570,N_11569);
xnor U11744 (N_11744,N_11642,N_11604);
or U11745 (N_11745,N_11586,N_11645);
nor U11746 (N_11746,N_11641,N_11651);
or U11747 (N_11747,N_11537,N_11594);
nand U11748 (N_11748,N_11527,N_11528);
xnor U11749 (N_11749,N_11631,N_11551);
and U11750 (N_11750,N_11571,N_11663);
and U11751 (N_11751,N_11565,N_11639);
nor U11752 (N_11752,N_11678,N_11652);
xnor U11753 (N_11753,N_11591,N_11648);
nand U11754 (N_11754,N_11627,N_11574);
or U11755 (N_11755,N_11626,N_11555);
nor U11756 (N_11756,N_11618,N_11679);
xnor U11757 (N_11757,N_11584,N_11617);
and U11758 (N_11758,N_11560,N_11659);
or U11759 (N_11759,N_11609,N_11521);
nor U11760 (N_11760,N_11672,N_11641);
xnor U11761 (N_11761,N_11596,N_11554);
and U11762 (N_11762,N_11590,N_11606);
nor U11763 (N_11763,N_11546,N_11559);
and U11764 (N_11764,N_11578,N_11535);
nand U11765 (N_11765,N_11540,N_11564);
nand U11766 (N_11766,N_11655,N_11667);
nand U11767 (N_11767,N_11552,N_11588);
nand U11768 (N_11768,N_11533,N_11527);
xor U11769 (N_11769,N_11653,N_11561);
xor U11770 (N_11770,N_11667,N_11535);
nand U11771 (N_11771,N_11603,N_11554);
nor U11772 (N_11772,N_11569,N_11561);
or U11773 (N_11773,N_11653,N_11542);
xor U11774 (N_11774,N_11558,N_11673);
nand U11775 (N_11775,N_11590,N_11651);
nor U11776 (N_11776,N_11658,N_11521);
nand U11777 (N_11777,N_11575,N_11591);
nand U11778 (N_11778,N_11596,N_11571);
nand U11779 (N_11779,N_11524,N_11576);
or U11780 (N_11780,N_11664,N_11534);
xnor U11781 (N_11781,N_11618,N_11547);
nand U11782 (N_11782,N_11670,N_11607);
or U11783 (N_11783,N_11546,N_11679);
or U11784 (N_11784,N_11641,N_11569);
and U11785 (N_11785,N_11629,N_11638);
and U11786 (N_11786,N_11612,N_11663);
and U11787 (N_11787,N_11535,N_11654);
nor U11788 (N_11788,N_11577,N_11522);
nor U11789 (N_11789,N_11534,N_11628);
and U11790 (N_11790,N_11571,N_11625);
nor U11791 (N_11791,N_11603,N_11615);
or U11792 (N_11792,N_11662,N_11594);
nor U11793 (N_11793,N_11560,N_11540);
nor U11794 (N_11794,N_11572,N_11590);
nor U11795 (N_11795,N_11586,N_11576);
nor U11796 (N_11796,N_11603,N_11571);
or U11797 (N_11797,N_11551,N_11561);
nand U11798 (N_11798,N_11558,N_11662);
nand U11799 (N_11799,N_11591,N_11521);
nand U11800 (N_11800,N_11535,N_11593);
nand U11801 (N_11801,N_11537,N_11622);
nor U11802 (N_11802,N_11593,N_11640);
and U11803 (N_11803,N_11638,N_11677);
xor U11804 (N_11804,N_11628,N_11666);
or U11805 (N_11805,N_11565,N_11647);
or U11806 (N_11806,N_11656,N_11547);
or U11807 (N_11807,N_11660,N_11538);
nor U11808 (N_11808,N_11548,N_11633);
nor U11809 (N_11809,N_11522,N_11606);
xor U11810 (N_11810,N_11639,N_11610);
xnor U11811 (N_11811,N_11622,N_11654);
nor U11812 (N_11812,N_11579,N_11592);
xor U11813 (N_11813,N_11561,N_11575);
or U11814 (N_11814,N_11556,N_11667);
nand U11815 (N_11815,N_11565,N_11676);
and U11816 (N_11816,N_11543,N_11544);
or U11817 (N_11817,N_11566,N_11526);
nor U11818 (N_11818,N_11535,N_11531);
and U11819 (N_11819,N_11647,N_11652);
nor U11820 (N_11820,N_11526,N_11626);
nor U11821 (N_11821,N_11587,N_11660);
xor U11822 (N_11822,N_11538,N_11661);
nand U11823 (N_11823,N_11520,N_11673);
or U11824 (N_11824,N_11561,N_11555);
nor U11825 (N_11825,N_11525,N_11600);
and U11826 (N_11826,N_11678,N_11661);
or U11827 (N_11827,N_11596,N_11599);
nand U11828 (N_11828,N_11611,N_11525);
nand U11829 (N_11829,N_11611,N_11614);
nand U11830 (N_11830,N_11642,N_11672);
and U11831 (N_11831,N_11524,N_11642);
xor U11832 (N_11832,N_11525,N_11628);
xnor U11833 (N_11833,N_11539,N_11670);
nor U11834 (N_11834,N_11670,N_11660);
and U11835 (N_11835,N_11535,N_11598);
nor U11836 (N_11836,N_11631,N_11621);
or U11837 (N_11837,N_11654,N_11599);
and U11838 (N_11838,N_11639,N_11528);
or U11839 (N_11839,N_11600,N_11578);
and U11840 (N_11840,N_11822,N_11752);
xor U11841 (N_11841,N_11806,N_11699);
nor U11842 (N_11842,N_11783,N_11813);
or U11843 (N_11843,N_11835,N_11803);
nand U11844 (N_11844,N_11839,N_11683);
or U11845 (N_11845,N_11834,N_11824);
or U11846 (N_11846,N_11777,N_11810);
nor U11847 (N_11847,N_11804,N_11761);
nor U11848 (N_11848,N_11749,N_11681);
nand U11849 (N_11849,N_11764,N_11735);
nand U11850 (N_11850,N_11780,N_11718);
and U11851 (N_11851,N_11809,N_11733);
nor U11852 (N_11852,N_11686,N_11708);
and U11853 (N_11853,N_11836,N_11812);
and U11854 (N_11854,N_11720,N_11744);
nand U11855 (N_11855,N_11741,N_11758);
xnor U11856 (N_11856,N_11730,N_11711);
and U11857 (N_11857,N_11696,N_11837);
xnor U11858 (N_11858,N_11693,N_11801);
nor U11859 (N_11859,N_11745,N_11760);
and U11860 (N_11860,N_11727,N_11717);
nor U11861 (N_11861,N_11721,N_11797);
or U11862 (N_11862,N_11759,N_11821);
xor U11863 (N_11863,N_11828,N_11784);
nand U11864 (N_11864,N_11808,N_11800);
nand U11865 (N_11865,N_11724,N_11737);
or U11866 (N_11866,N_11826,N_11782);
and U11867 (N_11867,N_11771,N_11689);
nor U11868 (N_11868,N_11767,N_11788);
xor U11869 (N_11869,N_11795,N_11705);
or U11870 (N_11870,N_11792,N_11714);
or U11871 (N_11871,N_11704,N_11713);
xnor U11872 (N_11872,N_11723,N_11710);
xnor U11873 (N_11873,N_11684,N_11774);
xnor U11874 (N_11874,N_11814,N_11831);
or U11875 (N_11875,N_11794,N_11755);
or U11876 (N_11876,N_11778,N_11793);
and U11877 (N_11877,N_11817,N_11682);
nor U11878 (N_11878,N_11748,N_11832);
and U11879 (N_11879,N_11743,N_11707);
or U11880 (N_11880,N_11786,N_11716);
or U11881 (N_11881,N_11754,N_11773);
nand U11882 (N_11882,N_11740,N_11747);
nor U11883 (N_11883,N_11739,N_11763);
and U11884 (N_11884,N_11818,N_11706);
nand U11885 (N_11885,N_11680,N_11688);
or U11886 (N_11886,N_11742,N_11732);
or U11887 (N_11887,N_11838,N_11805);
xor U11888 (N_11888,N_11796,N_11697);
and U11889 (N_11889,N_11779,N_11789);
or U11890 (N_11890,N_11750,N_11746);
xor U11891 (N_11891,N_11691,N_11702);
nand U11892 (N_11892,N_11791,N_11685);
nor U11893 (N_11893,N_11729,N_11715);
or U11894 (N_11894,N_11829,N_11719);
xnor U11895 (N_11895,N_11807,N_11785);
and U11896 (N_11896,N_11769,N_11725);
or U11897 (N_11897,N_11736,N_11772);
xnor U11898 (N_11898,N_11823,N_11833);
xnor U11899 (N_11899,N_11753,N_11731);
or U11900 (N_11900,N_11811,N_11815);
nand U11901 (N_11901,N_11798,N_11695);
nand U11902 (N_11902,N_11751,N_11766);
or U11903 (N_11903,N_11768,N_11722);
or U11904 (N_11904,N_11825,N_11734);
xor U11905 (N_11905,N_11694,N_11819);
xor U11906 (N_11906,N_11703,N_11756);
xor U11907 (N_11907,N_11799,N_11820);
and U11908 (N_11908,N_11762,N_11690);
nand U11909 (N_11909,N_11757,N_11790);
nor U11910 (N_11910,N_11709,N_11781);
or U11911 (N_11911,N_11698,N_11738);
xnor U11912 (N_11912,N_11692,N_11830);
nor U11913 (N_11913,N_11775,N_11712);
or U11914 (N_11914,N_11726,N_11827);
nand U11915 (N_11915,N_11728,N_11816);
and U11916 (N_11916,N_11802,N_11700);
xnor U11917 (N_11917,N_11787,N_11770);
nor U11918 (N_11918,N_11776,N_11701);
or U11919 (N_11919,N_11687,N_11765);
and U11920 (N_11920,N_11781,N_11766);
xor U11921 (N_11921,N_11686,N_11753);
nor U11922 (N_11922,N_11728,N_11790);
and U11923 (N_11923,N_11785,N_11731);
and U11924 (N_11924,N_11773,N_11682);
nor U11925 (N_11925,N_11701,N_11837);
xnor U11926 (N_11926,N_11690,N_11699);
nor U11927 (N_11927,N_11680,N_11806);
nor U11928 (N_11928,N_11788,N_11787);
or U11929 (N_11929,N_11752,N_11832);
and U11930 (N_11930,N_11680,N_11786);
and U11931 (N_11931,N_11837,N_11717);
xor U11932 (N_11932,N_11805,N_11742);
or U11933 (N_11933,N_11832,N_11757);
xor U11934 (N_11934,N_11747,N_11772);
or U11935 (N_11935,N_11702,N_11782);
and U11936 (N_11936,N_11699,N_11706);
or U11937 (N_11937,N_11768,N_11821);
or U11938 (N_11938,N_11834,N_11763);
nor U11939 (N_11939,N_11815,N_11819);
or U11940 (N_11940,N_11767,N_11751);
and U11941 (N_11941,N_11708,N_11775);
or U11942 (N_11942,N_11786,N_11685);
and U11943 (N_11943,N_11702,N_11819);
and U11944 (N_11944,N_11824,N_11750);
xnor U11945 (N_11945,N_11715,N_11821);
nand U11946 (N_11946,N_11786,N_11708);
or U11947 (N_11947,N_11681,N_11824);
or U11948 (N_11948,N_11814,N_11748);
nand U11949 (N_11949,N_11721,N_11825);
and U11950 (N_11950,N_11753,N_11701);
nor U11951 (N_11951,N_11729,N_11745);
nor U11952 (N_11952,N_11692,N_11726);
nand U11953 (N_11953,N_11705,N_11777);
nand U11954 (N_11954,N_11767,N_11705);
or U11955 (N_11955,N_11792,N_11770);
or U11956 (N_11956,N_11713,N_11723);
and U11957 (N_11957,N_11684,N_11680);
nand U11958 (N_11958,N_11752,N_11695);
and U11959 (N_11959,N_11820,N_11715);
or U11960 (N_11960,N_11749,N_11737);
xnor U11961 (N_11961,N_11806,N_11685);
and U11962 (N_11962,N_11808,N_11810);
xnor U11963 (N_11963,N_11791,N_11718);
or U11964 (N_11964,N_11812,N_11755);
nand U11965 (N_11965,N_11739,N_11778);
or U11966 (N_11966,N_11735,N_11783);
and U11967 (N_11967,N_11704,N_11821);
or U11968 (N_11968,N_11682,N_11721);
nand U11969 (N_11969,N_11696,N_11778);
xor U11970 (N_11970,N_11737,N_11694);
and U11971 (N_11971,N_11748,N_11778);
and U11972 (N_11972,N_11737,N_11703);
or U11973 (N_11973,N_11765,N_11779);
nand U11974 (N_11974,N_11819,N_11762);
or U11975 (N_11975,N_11833,N_11781);
or U11976 (N_11976,N_11714,N_11794);
and U11977 (N_11977,N_11772,N_11767);
and U11978 (N_11978,N_11770,N_11683);
nor U11979 (N_11979,N_11788,N_11792);
nor U11980 (N_11980,N_11760,N_11692);
or U11981 (N_11981,N_11774,N_11740);
and U11982 (N_11982,N_11778,N_11803);
nor U11983 (N_11983,N_11835,N_11704);
or U11984 (N_11984,N_11832,N_11795);
xnor U11985 (N_11985,N_11693,N_11709);
nand U11986 (N_11986,N_11686,N_11695);
nor U11987 (N_11987,N_11718,N_11828);
xnor U11988 (N_11988,N_11736,N_11759);
nand U11989 (N_11989,N_11766,N_11793);
nor U11990 (N_11990,N_11793,N_11745);
nand U11991 (N_11991,N_11720,N_11801);
nand U11992 (N_11992,N_11721,N_11836);
and U11993 (N_11993,N_11795,N_11756);
nand U11994 (N_11994,N_11833,N_11838);
nand U11995 (N_11995,N_11682,N_11748);
and U11996 (N_11996,N_11764,N_11779);
nor U11997 (N_11997,N_11699,N_11753);
nor U11998 (N_11998,N_11832,N_11721);
and U11999 (N_11999,N_11757,N_11806);
or U12000 (N_12000,N_11979,N_11936);
and U12001 (N_12001,N_11849,N_11908);
nand U12002 (N_12002,N_11848,N_11913);
xor U12003 (N_12003,N_11869,N_11945);
or U12004 (N_12004,N_11846,N_11991);
nand U12005 (N_12005,N_11922,N_11875);
or U12006 (N_12006,N_11890,N_11884);
nor U12007 (N_12007,N_11928,N_11910);
nand U12008 (N_12008,N_11864,N_11844);
or U12009 (N_12009,N_11932,N_11883);
or U12010 (N_12010,N_11924,N_11990);
xnor U12011 (N_12011,N_11964,N_11926);
and U12012 (N_12012,N_11987,N_11958);
nand U12013 (N_12013,N_11969,N_11904);
or U12014 (N_12014,N_11851,N_11903);
xnor U12015 (N_12015,N_11876,N_11856);
and U12016 (N_12016,N_11859,N_11885);
xnor U12017 (N_12017,N_11920,N_11940);
xnor U12018 (N_12018,N_11973,N_11914);
and U12019 (N_12019,N_11872,N_11947);
or U12020 (N_12020,N_11917,N_11967);
and U12021 (N_12021,N_11988,N_11935);
nor U12022 (N_12022,N_11850,N_11980);
or U12023 (N_12023,N_11986,N_11888);
or U12024 (N_12024,N_11965,N_11972);
and U12025 (N_12025,N_11882,N_11933);
nor U12026 (N_12026,N_11960,N_11898);
and U12027 (N_12027,N_11974,N_11897);
nor U12028 (N_12028,N_11954,N_11998);
xnor U12029 (N_12029,N_11927,N_11877);
nand U12030 (N_12030,N_11886,N_11997);
nor U12031 (N_12031,N_11867,N_11962);
and U12032 (N_12032,N_11871,N_11930);
nor U12033 (N_12033,N_11881,N_11915);
or U12034 (N_12034,N_11878,N_11946);
nor U12035 (N_12035,N_11906,N_11918);
xor U12036 (N_12036,N_11956,N_11843);
nand U12037 (N_12037,N_11842,N_11951);
nand U12038 (N_12038,N_11942,N_11845);
or U12039 (N_12039,N_11981,N_11978);
nor U12040 (N_12040,N_11992,N_11862);
xor U12041 (N_12041,N_11996,N_11925);
nand U12042 (N_12042,N_11853,N_11902);
or U12043 (N_12043,N_11982,N_11870);
and U12044 (N_12044,N_11880,N_11966);
nand U12045 (N_12045,N_11858,N_11873);
or U12046 (N_12046,N_11909,N_11953);
nand U12047 (N_12047,N_11985,N_11983);
nor U12048 (N_12048,N_11949,N_11912);
or U12049 (N_12049,N_11984,N_11855);
xnor U12050 (N_12050,N_11923,N_11937);
nor U12051 (N_12051,N_11999,N_11916);
nand U12052 (N_12052,N_11968,N_11975);
and U12053 (N_12053,N_11866,N_11874);
or U12054 (N_12054,N_11847,N_11941);
or U12055 (N_12055,N_11959,N_11895);
nor U12056 (N_12056,N_11901,N_11970);
xnor U12057 (N_12057,N_11929,N_11852);
and U12058 (N_12058,N_11868,N_11943);
or U12059 (N_12059,N_11934,N_11994);
nor U12060 (N_12060,N_11963,N_11919);
and U12061 (N_12061,N_11948,N_11889);
nor U12062 (N_12062,N_11894,N_11976);
or U12063 (N_12063,N_11887,N_11840);
nand U12064 (N_12064,N_11944,N_11993);
xnor U12065 (N_12065,N_11891,N_11931);
xnor U12066 (N_12066,N_11961,N_11971);
nand U12067 (N_12067,N_11863,N_11892);
nor U12068 (N_12068,N_11955,N_11950);
nor U12069 (N_12069,N_11841,N_11854);
or U12070 (N_12070,N_11861,N_11899);
xor U12071 (N_12071,N_11900,N_11989);
nor U12072 (N_12072,N_11907,N_11860);
nor U12073 (N_12073,N_11905,N_11938);
xnor U12074 (N_12074,N_11921,N_11911);
or U12075 (N_12075,N_11977,N_11952);
and U12076 (N_12076,N_11865,N_11896);
or U12077 (N_12077,N_11893,N_11957);
nor U12078 (N_12078,N_11939,N_11879);
nand U12079 (N_12079,N_11995,N_11857);
and U12080 (N_12080,N_11978,N_11954);
or U12081 (N_12081,N_11885,N_11955);
nor U12082 (N_12082,N_11936,N_11934);
or U12083 (N_12083,N_11994,N_11951);
nand U12084 (N_12084,N_11968,N_11893);
nand U12085 (N_12085,N_11973,N_11913);
and U12086 (N_12086,N_11920,N_11906);
or U12087 (N_12087,N_11924,N_11988);
xor U12088 (N_12088,N_11877,N_11918);
nand U12089 (N_12089,N_11949,N_11942);
nand U12090 (N_12090,N_11844,N_11886);
and U12091 (N_12091,N_11848,N_11852);
nand U12092 (N_12092,N_11849,N_11916);
or U12093 (N_12093,N_11949,N_11842);
xor U12094 (N_12094,N_11976,N_11889);
nand U12095 (N_12095,N_11852,N_11856);
xor U12096 (N_12096,N_11997,N_11949);
xnor U12097 (N_12097,N_11866,N_11998);
xnor U12098 (N_12098,N_11932,N_11998);
or U12099 (N_12099,N_11887,N_11960);
and U12100 (N_12100,N_11852,N_11841);
nand U12101 (N_12101,N_11929,N_11902);
nor U12102 (N_12102,N_11854,N_11945);
nand U12103 (N_12103,N_11894,N_11912);
and U12104 (N_12104,N_11852,N_11887);
xor U12105 (N_12105,N_11996,N_11886);
and U12106 (N_12106,N_11927,N_11925);
xnor U12107 (N_12107,N_11912,N_11988);
nor U12108 (N_12108,N_11847,N_11894);
and U12109 (N_12109,N_11872,N_11987);
or U12110 (N_12110,N_11969,N_11854);
nand U12111 (N_12111,N_11855,N_11938);
nand U12112 (N_12112,N_11947,N_11898);
xnor U12113 (N_12113,N_11851,N_11979);
xnor U12114 (N_12114,N_11949,N_11887);
and U12115 (N_12115,N_11958,N_11992);
xnor U12116 (N_12116,N_11912,N_11979);
nor U12117 (N_12117,N_11871,N_11858);
and U12118 (N_12118,N_11868,N_11957);
nor U12119 (N_12119,N_11919,N_11847);
xnor U12120 (N_12120,N_11995,N_11986);
xor U12121 (N_12121,N_11996,N_11935);
xor U12122 (N_12122,N_11972,N_11926);
nand U12123 (N_12123,N_11937,N_11887);
nand U12124 (N_12124,N_11881,N_11856);
xnor U12125 (N_12125,N_11870,N_11913);
nand U12126 (N_12126,N_11999,N_11985);
xor U12127 (N_12127,N_11854,N_11903);
xnor U12128 (N_12128,N_11947,N_11983);
nand U12129 (N_12129,N_11907,N_11993);
and U12130 (N_12130,N_11935,N_11842);
nand U12131 (N_12131,N_11941,N_11962);
nand U12132 (N_12132,N_11892,N_11984);
nor U12133 (N_12133,N_11881,N_11861);
nor U12134 (N_12134,N_11943,N_11862);
nor U12135 (N_12135,N_11964,N_11899);
and U12136 (N_12136,N_11992,N_11935);
xor U12137 (N_12137,N_11932,N_11874);
or U12138 (N_12138,N_11915,N_11845);
or U12139 (N_12139,N_11912,N_11992);
xnor U12140 (N_12140,N_11984,N_11990);
nor U12141 (N_12141,N_11850,N_11875);
nand U12142 (N_12142,N_11850,N_11951);
nand U12143 (N_12143,N_11847,N_11875);
and U12144 (N_12144,N_11986,N_11957);
xnor U12145 (N_12145,N_11988,N_11946);
nand U12146 (N_12146,N_11883,N_11943);
and U12147 (N_12147,N_11999,N_11939);
xor U12148 (N_12148,N_11923,N_11949);
and U12149 (N_12149,N_11922,N_11954);
nor U12150 (N_12150,N_11925,N_11988);
nand U12151 (N_12151,N_11859,N_11985);
xnor U12152 (N_12152,N_11858,N_11894);
xnor U12153 (N_12153,N_11844,N_11962);
nor U12154 (N_12154,N_11990,N_11969);
or U12155 (N_12155,N_11845,N_11847);
nor U12156 (N_12156,N_11987,N_11923);
nor U12157 (N_12157,N_11939,N_11848);
nand U12158 (N_12158,N_11946,N_11970);
nor U12159 (N_12159,N_11858,N_11930);
nand U12160 (N_12160,N_12053,N_12077);
xnor U12161 (N_12161,N_12092,N_12025);
or U12162 (N_12162,N_12125,N_12149);
or U12163 (N_12163,N_12098,N_12080);
or U12164 (N_12164,N_12020,N_12007);
and U12165 (N_12165,N_12128,N_12017);
nand U12166 (N_12166,N_12045,N_12134);
or U12167 (N_12167,N_12066,N_12078);
or U12168 (N_12168,N_12099,N_12148);
nor U12169 (N_12169,N_12144,N_12024);
and U12170 (N_12170,N_12062,N_12143);
nand U12171 (N_12171,N_12088,N_12038);
nor U12172 (N_12172,N_12104,N_12159);
or U12173 (N_12173,N_12087,N_12133);
and U12174 (N_12174,N_12093,N_12030);
nand U12175 (N_12175,N_12055,N_12137);
and U12176 (N_12176,N_12082,N_12076);
xor U12177 (N_12177,N_12052,N_12131);
and U12178 (N_12178,N_12006,N_12027);
and U12179 (N_12179,N_12111,N_12047);
nor U12180 (N_12180,N_12158,N_12127);
and U12181 (N_12181,N_12130,N_12152);
nor U12182 (N_12182,N_12058,N_12145);
and U12183 (N_12183,N_12153,N_12147);
and U12184 (N_12184,N_12032,N_12132);
xor U12185 (N_12185,N_12083,N_12108);
nor U12186 (N_12186,N_12067,N_12000);
nand U12187 (N_12187,N_12035,N_12079);
and U12188 (N_12188,N_12016,N_12011);
or U12189 (N_12189,N_12106,N_12065);
and U12190 (N_12190,N_12061,N_12094);
or U12191 (N_12191,N_12095,N_12064);
or U12192 (N_12192,N_12048,N_12155);
nor U12193 (N_12193,N_12049,N_12150);
xor U12194 (N_12194,N_12001,N_12063);
or U12195 (N_12195,N_12115,N_12085);
nand U12196 (N_12196,N_12086,N_12039);
xor U12197 (N_12197,N_12101,N_12028);
nor U12198 (N_12198,N_12113,N_12084);
xnor U12199 (N_12199,N_12042,N_12021);
or U12200 (N_12200,N_12117,N_12105);
nand U12201 (N_12201,N_12043,N_12072);
nand U12202 (N_12202,N_12118,N_12068);
nor U12203 (N_12203,N_12151,N_12100);
nand U12204 (N_12204,N_12119,N_12012);
or U12205 (N_12205,N_12069,N_12116);
xnor U12206 (N_12206,N_12026,N_12057);
and U12207 (N_12207,N_12097,N_12121);
nand U12208 (N_12208,N_12090,N_12123);
nor U12209 (N_12209,N_12122,N_12091);
and U12210 (N_12210,N_12029,N_12010);
or U12211 (N_12211,N_12014,N_12013);
and U12212 (N_12212,N_12036,N_12075);
and U12213 (N_12213,N_12142,N_12018);
nor U12214 (N_12214,N_12050,N_12139);
and U12215 (N_12215,N_12073,N_12138);
nor U12216 (N_12216,N_12056,N_12154);
and U12217 (N_12217,N_12051,N_12040);
and U12218 (N_12218,N_12110,N_12074);
or U12219 (N_12219,N_12124,N_12003);
nand U12220 (N_12220,N_12009,N_12041);
and U12221 (N_12221,N_12002,N_12022);
nand U12222 (N_12222,N_12107,N_12109);
nand U12223 (N_12223,N_12136,N_12015);
nor U12224 (N_12224,N_12141,N_12008);
and U12225 (N_12225,N_12081,N_12146);
and U12226 (N_12226,N_12135,N_12156);
or U12227 (N_12227,N_12005,N_12033);
xor U12228 (N_12228,N_12059,N_12103);
nor U12229 (N_12229,N_12112,N_12023);
nor U12230 (N_12230,N_12004,N_12070);
and U12231 (N_12231,N_12031,N_12140);
nand U12232 (N_12232,N_12060,N_12129);
and U12233 (N_12233,N_12157,N_12096);
and U12234 (N_12234,N_12044,N_12126);
or U12235 (N_12235,N_12089,N_12054);
and U12236 (N_12236,N_12120,N_12037);
nor U12237 (N_12237,N_12102,N_12019);
or U12238 (N_12238,N_12071,N_12114);
xor U12239 (N_12239,N_12046,N_12034);
nor U12240 (N_12240,N_12112,N_12140);
nand U12241 (N_12241,N_12156,N_12051);
or U12242 (N_12242,N_12032,N_12135);
and U12243 (N_12243,N_12115,N_12079);
nor U12244 (N_12244,N_12053,N_12024);
nor U12245 (N_12245,N_12070,N_12115);
or U12246 (N_12246,N_12020,N_12010);
nand U12247 (N_12247,N_12096,N_12158);
nor U12248 (N_12248,N_12084,N_12034);
and U12249 (N_12249,N_12145,N_12073);
nand U12250 (N_12250,N_12043,N_12140);
nand U12251 (N_12251,N_12065,N_12151);
xnor U12252 (N_12252,N_12139,N_12062);
nand U12253 (N_12253,N_12038,N_12068);
nor U12254 (N_12254,N_12061,N_12053);
and U12255 (N_12255,N_12094,N_12154);
nor U12256 (N_12256,N_12087,N_12017);
xnor U12257 (N_12257,N_12031,N_12126);
nand U12258 (N_12258,N_12069,N_12111);
or U12259 (N_12259,N_12139,N_12052);
nor U12260 (N_12260,N_12015,N_12026);
nor U12261 (N_12261,N_12154,N_12022);
xnor U12262 (N_12262,N_12143,N_12109);
nand U12263 (N_12263,N_12143,N_12099);
or U12264 (N_12264,N_12017,N_12091);
nor U12265 (N_12265,N_12149,N_12001);
and U12266 (N_12266,N_12124,N_12033);
xor U12267 (N_12267,N_12034,N_12127);
nand U12268 (N_12268,N_12098,N_12103);
nor U12269 (N_12269,N_12052,N_12153);
nor U12270 (N_12270,N_12060,N_12036);
and U12271 (N_12271,N_12012,N_12055);
or U12272 (N_12272,N_12022,N_12028);
nor U12273 (N_12273,N_12039,N_12053);
and U12274 (N_12274,N_12125,N_12126);
nand U12275 (N_12275,N_12099,N_12119);
and U12276 (N_12276,N_12111,N_12057);
nor U12277 (N_12277,N_12004,N_12039);
xnor U12278 (N_12278,N_12095,N_12105);
xor U12279 (N_12279,N_12137,N_12082);
and U12280 (N_12280,N_12159,N_12038);
or U12281 (N_12281,N_12132,N_12044);
and U12282 (N_12282,N_12037,N_12016);
xor U12283 (N_12283,N_12007,N_12047);
nor U12284 (N_12284,N_12135,N_12036);
xor U12285 (N_12285,N_12146,N_12051);
nor U12286 (N_12286,N_12048,N_12134);
and U12287 (N_12287,N_12033,N_12034);
nor U12288 (N_12288,N_12075,N_12081);
xnor U12289 (N_12289,N_12077,N_12115);
nor U12290 (N_12290,N_12057,N_12010);
and U12291 (N_12291,N_12044,N_12031);
or U12292 (N_12292,N_12111,N_12048);
nand U12293 (N_12293,N_12062,N_12136);
and U12294 (N_12294,N_12056,N_12060);
xor U12295 (N_12295,N_12071,N_12003);
or U12296 (N_12296,N_12044,N_12001);
xor U12297 (N_12297,N_12155,N_12088);
nor U12298 (N_12298,N_12015,N_12123);
nor U12299 (N_12299,N_12069,N_12145);
nand U12300 (N_12300,N_12081,N_12106);
nor U12301 (N_12301,N_12076,N_12092);
or U12302 (N_12302,N_12104,N_12067);
or U12303 (N_12303,N_12156,N_12145);
nand U12304 (N_12304,N_12063,N_12070);
nor U12305 (N_12305,N_12096,N_12143);
nand U12306 (N_12306,N_12114,N_12034);
nor U12307 (N_12307,N_12133,N_12100);
and U12308 (N_12308,N_12069,N_12121);
xnor U12309 (N_12309,N_12060,N_12110);
and U12310 (N_12310,N_12022,N_12093);
nand U12311 (N_12311,N_12130,N_12016);
nor U12312 (N_12312,N_12049,N_12099);
nor U12313 (N_12313,N_12032,N_12098);
or U12314 (N_12314,N_12089,N_12037);
nand U12315 (N_12315,N_12134,N_12115);
nor U12316 (N_12316,N_12133,N_12037);
xnor U12317 (N_12317,N_12008,N_12070);
nor U12318 (N_12318,N_12128,N_12092);
nor U12319 (N_12319,N_12094,N_12129);
and U12320 (N_12320,N_12284,N_12182);
or U12321 (N_12321,N_12198,N_12194);
nor U12322 (N_12322,N_12200,N_12163);
or U12323 (N_12323,N_12220,N_12219);
and U12324 (N_12324,N_12275,N_12201);
nor U12325 (N_12325,N_12302,N_12312);
nand U12326 (N_12326,N_12185,N_12184);
nand U12327 (N_12327,N_12271,N_12167);
or U12328 (N_12328,N_12304,N_12295);
and U12329 (N_12329,N_12172,N_12171);
xnor U12330 (N_12330,N_12301,N_12269);
xnor U12331 (N_12331,N_12170,N_12223);
and U12332 (N_12332,N_12204,N_12226);
and U12333 (N_12333,N_12168,N_12266);
nand U12334 (N_12334,N_12288,N_12319);
or U12335 (N_12335,N_12208,N_12303);
or U12336 (N_12336,N_12270,N_12217);
and U12337 (N_12337,N_12293,N_12289);
nand U12338 (N_12338,N_12309,N_12178);
and U12339 (N_12339,N_12209,N_12202);
nand U12340 (N_12340,N_12297,N_12294);
and U12341 (N_12341,N_12177,N_12256);
and U12342 (N_12342,N_12286,N_12274);
xor U12343 (N_12343,N_12212,N_12285);
xnor U12344 (N_12344,N_12227,N_12290);
or U12345 (N_12345,N_12317,N_12180);
and U12346 (N_12346,N_12310,N_12243);
or U12347 (N_12347,N_12193,N_12251);
nand U12348 (N_12348,N_12232,N_12165);
or U12349 (N_12349,N_12189,N_12233);
nor U12350 (N_12350,N_12166,N_12252);
nor U12351 (N_12351,N_12257,N_12300);
and U12352 (N_12352,N_12173,N_12305);
or U12353 (N_12353,N_12282,N_12192);
nand U12354 (N_12354,N_12179,N_12176);
and U12355 (N_12355,N_12277,N_12273);
nand U12356 (N_12356,N_12196,N_12203);
nand U12357 (N_12357,N_12237,N_12246);
and U12358 (N_12358,N_12258,N_12186);
nor U12359 (N_12359,N_12287,N_12272);
nor U12360 (N_12360,N_12169,N_12239);
xnor U12361 (N_12361,N_12238,N_12162);
xnor U12362 (N_12362,N_12183,N_12164);
nor U12363 (N_12363,N_12240,N_12281);
xnor U12364 (N_12364,N_12315,N_12236);
and U12365 (N_12365,N_12260,N_12313);
nand U12366 (N_12366,N_12175,N_12191);
nand U12367 (N_12367,N_12299,N_12210);
and U12368 (N_12368,N_12306,N_12318);
nor U12369 (N_12369,N_12213,N_12283);
nor U12370 (N_12370,N_12161,N_12264);
xor U12371 (N_12371,N_12199,N_12263);
nor U12372 (N_12372,N_12268,N_12279);
xnor U12373 (N_12373,N_12298,N_12195);
nand U12374 (N_12374,N_12259,N_12276);
and U12375 (N_12375,N_12228,N_12216);
xnor U12376 (N_12376,N_12160,N_12314);
or U12377 (N_12377,N_12247,N_12253);
nor U12378 (N_12378,N_12215,N_12244);
and U12379 (N_12379,N_12311,N_12174);
nand U12380 (N_12380,N_12206,N_12218);
nand U12381 (N_12381,N_12197,N_12280);
nand U12382 (N_12382,N_12278,N_12230);
nor U12383 (N_12383,N_12242,N_12316);
nand U12384 (N_12384,N_12248,N_12292);
nand U12385 (N_12385,N_12214,N_12308);
xor U12386 (N_12386,N_12254,N_12207);
or U12387 (N_12387,N_12291,N_12235);
xor U12388 (N_12388,N_12307,N_12224);
nor U12389 (N_12389,N_12249,N_12181);
nor U12390 (N_12390,N_12190,N_12296);
nand U12391 (N_12391,N_12265,N_12261);
nor U12392 (N_12392,N_12234,N_12245);
nand U12393 (N_12393,N_12221,N_12250);
nor U12394 (N_12394,N_12225,N_12255);
and U12395 (N_12395,N_12262,N_12229);
xor U12396 (N_12396,N_12187,N_12241);
and U12397 (N_12397,N_12267,N_12205);
and U12398 (N_12398,N_12231,N_12211);
nand U12399 (N_12399,N_12222,N_12188);
xor U12400 (N_12400,N_12220,N_12266);
and U12401 (N_12401,N_12212,N_12276);
and U12402 (N_12402,N_12306,N_12314);
nand U12403 (N_12403,N_12162,N_12222);
and U12404 (N_12404,N_12242,N_12202);
xor U12405 (N_12405,N_12247,N_12212);
and U12406 (N_12406,N_12250,N_12217);
nor U12407 (N_12407,N_12275,N_12209);
nand U12408 (N_12408,N_12235,N_12238);
xnor U12409 (N_12409,N_12252,N_12232);
and U12410 (N_12410,N_12238,N_12180);
or U12411 (N_12411,N_12254,N_12311);
nor U12412 (N_12412,N_12261,N_12225);
xor U12413 (N_12413,N_12269,N_12264);
xnor U12414 (N_12414,N_12223,N_12260);
nor U12415 (N_12415,N_12249,N_12316);
nor U12416 (N_12416,N_12279,N_12248);
or U12417 (N_12417,N_12208,N_12251);
nand U12418 (N_12418,N_12211,N_12198);
nand U12419 (N_12419,N_12302,N_12290);
or U12420 (N_12420,N_12238,N_12178);
nor U12421 (N_12421,N_12174,N_12178);
nand U12422 (N_12422,N_12194,N_12262);
and U12423 (N_12423,N_12212,N_12241);
nand U12424 (N_12424,N_12228,N_12262);
and U12425 (N_12425,N_12213,N_12229);
nand U12426 (N_12426,N_12260,N_12249);
nand U12427 (N_12427,N_12244,N_12206);
nand U12428 (N_12428,N_12242,N_12231);
nor U12429 (N_12429,N_12239,N_12215);
nand U12430 (N_12430,N_12312,N_12275);
xnor U12431 (N_12431,N_12184,N_12198);
xor U12432 (N_12432,N_12168,N_12308);
and U12433 (N_12433,N_12244,N_12234);
or U12434 (N_12434,N_12214,N_12278);
nand U12435 (N_12435,N_12271,N_12299);
nor U12436 (N_12436,N_12306,N_12206);
nor U12437 (N_12437,N_12199,N_12214);
xnor U12438 (N_12438,N_12293,N_12283);
nor U12439 (N_12439,N_12236,N_12287);
or U12440 (N_12440,N_12209,N_12277);
nor U12441 (N_12441,N_12301,N_12297);
nor U12442 (N_12442,N_12287,N_12215);
or U12443 (N_12443,N_12237,N_12263);
xor U12444 (N_12444,N_12256,N_12232);
xnor U12445 (N_12445,N_12162,N_12264);
nand U12446 (N_12446,N_12244,N_12216);
xnor U12447 (N_12447,N_12270,N_12237);
and U12448 (N_12448,N_12204,N_12269);
nand U12449 (N_12449,N_12293,N_12278);
xor U12450 (N_12450,N_12186,N_12305);
xnor U12451 (N_12451,N_12175,N_12195);
xor U12452 (N_12452,N_12193,N_12316);
xnor U12453 (N_12453,N_12244,N_12288);
nor U12454 (N_12454,N_12223,N_12229);
nand U12455 (N_12455,N_12188,N_12303);
nand U12456 (N_12456,N_12316,N_12314);
xnor U12457 (N_12457,N_12301,N_12194);
and U12458 (N_12458,N_12217,N_12304);
nand U12459 (N_12459,N_12318,N_12301);
xor U12460 (N_12460,N_12190,N_12291);
xor U12461 (N_12461,N_12273,N_12274);
nor U12462 (N_12462,N_12194,N_12251);
xor U12463 (N_12463,N_12272,N_12267);
and U12464 (N_12464,N_12238,N_12239);
or U12465 (N_12465,N_12282,N_12275);
xnor U12466 (N_12466,N_12249,N_12285);
nand U12467 (N_12467,N_12246,N_12302);
nor U12468 (N_12468,N_12242,N_12160);
and U12469 (N_12469,N_12160,N_12187);
xnor U12470 (N_12470,N_12169,N_12212);
xor U12471 (N_12471,N_12198,N_12248);
xnor U12472 (N_12472,N_12289,N_12168);
xor U12473 (N_12473,N_12227,N_12198);
xnor U12474 (N_12474,N_12288,N_12277);
nand U12475 (N_12475,N_12193,N_12221);
and U12476 (N_12476,N_12267,N_12187);
nand U12477 (N_12477,N_12263,N_12256);
nor U12478 (N_12478,N_12244,N_12306);
or U12479 (N_12479,N_12230,N_12174);
xnor U12480 (N_12480,N_12454,N_12443);
xor U12481 (N_12481,N_12373,N_12368);
or U12482 (N_12482,N_12463,N_12320);
or U12483 (N_12483,N_12335,N_12460);
xnor U12484 (N_12484,N_12392,N_12396);
xor U12485 (N_12485,N_12438,N_12372);
nor U12486 (N_12486,N_12324,N_12439);
or U12487 (N_12487,N_12337,N_12367);
nand U12488 (N_12488,N_12475,N_12338);
or U12489 (N_12489,N_12321,N_12461);
and U12490 (N_12490,N_12447,N_12331);
xor U12491 (N_12491,N_12459,N_12325);
nand U12492 (N_12492,N_12474,N_12382);
and U12493 (N_12493,N_12430,N_12424);
nand U12494 (N_12494,N_12355,N_12332);
nor U12495 (N_12495,N_12413,N_12334);
or U12496 (N_12496,N_12383,N_12477);
and U12497 (N_12497,N_12440,N_12339);
and U12498 (N_12498,N_12351,N_12434);
nand U12499 (N_12499,N_12344,N_12445);
nand U12500 (N_12500,N_12455,N_12346);
and U12501 (N_12501,N_12336,N_12411);
xor U12502 (N_12502,N_12386,N_12416);
or U12503 (N_12503,N_12352,N_12410);
and U12504 (N_12504,N_12387,N_12436);
nor U12505 (N_12505,N_12348,N_12343);
or U12506 (N_12506,N_12465,N_12391);
xnor U12507 (N_12507,N_12400,N_12423);
or U12508 (N_12508,N_12379,N_12366);
xnor U12509 (N_12509,N_12422,N_12361);
or U12510 (N_12510,N_12452,N_12425);
nand U12511 (N_12511,N_12435,N_12406);
or U12512 (N_12512,N_12453,N_12329);
or U12513 (N_12513,N_12398,N_12376);
xnor U12514 (N_12514,N_12380,N_12441);
or U12515 (N_12515,N_12417,N_12472);
nand U12516 (N_12516,N_12328,N_12415);
and U12517 (N_12517,N_12420,N_12356);
nand U12518 (N_12518,N_12421,N_12405);
and U12519 (N_12519,N_12437,N_12450);
xnor U12520 (N_12520,N_12479,N_12458);
nor U12521 (N_12521,N_12412,N_12374);
and U12522 (N_12522,N_12384,N_12381);
xnor U12523 (N_12523,N_12370,N_12470);
and U12524 (N_12524,N_12468,N_12402);
or U12525 (N_12525,N_12389,N_12466);
xnor U12526 (N_12526,N_12467,N_12326);
xnor U12527 (N_12527,N_12446,N_12362);
and U12528 (N_12528,N_12444,N_12464);
and U12529 (N_12529,N_12451,N_12364);
nand U12530 (N_12530,N_12418,N_12350);
nand U12531 (N_12531,N_12327,N_12365);
xor U12532 (N_12532,N_12401,N_12442);
and U12533 (N_12533,N_12347,N_12385);
nor U12534 (N_12534,N_12340,N_12377);
or U12535 (N_12535,N_12426,N_12395);
nor U12536 (N_12536,N_12345,N_12323);
nand U12537 (N_12537,N_12378,N_12419);
nand U12538 (N_12538,N_12360,N_12414);
or U12539 (N_12539,N_12469,N_12462);
xor U12540 (N_12540,N_12449,N_12322);
nor U12541 (N_12541,N_12342,N_12333);
nor U12542 (N_12542,N_12375,N_12428);
or U12543 (N_12543,N_12357,N_12359);
xnor U12544 (N_12544,N_12397,N_12394);
xor U12545 (N_12545,N_12358,N_12404);
xnor U12546 (N_12546,N_12363,N_12471);
and U12547 (N_12547,N_12448,N_12388);
nor U12548 (N_12548,N_12432,N_12427);
or U12549 (N_12549,N_12431,N_12393);
xor U12550 (N_12550,N_12371,N_12457);
xor U12551 (N_12551,N_12369,N_12349);
and U12552 (N_12552,N_12476,N_12407);
xnor U12553 (N_12553,N_12433,N_12399);
xnor U12554 (N_12554,N_12473,N_12408);
xnor U12555 (N_12555,N_12456,N_12390);
or U12556 (N_12556,N_12478,N_12409);
and U12557 (N_12557,N_12354,N_12429);
nor U12558 (N_12558,N_12353,N_12330);
nand U12559 (N_12559,N_12403,N_12341);
or U12560 (N_12560,N_12429,N_12449);
and U12561 (N_12561,N_12352,N_12362);
nand U12562 (N_12562,N_12329,N_12333);
nand U12563 (N_12563,N_12438,N_12380);
and U12564 (N_12564,N_12409,N_12443);
or U12565 (N_12565,N_12438,N_12341);
and U12566 (N_12566,N_12471,N_12323);
or U12567 (N_12567,N_12430,N_12381);
nor U12568 (N_12568,N_12442,N_12334);
or U12569 (N_12569,N_12430,N_12470);
nand U12570 (N_12570,N_12465,N_12324);
and U12571 (N_12571,N_12475,N_12458);
and U12572 (N_12572,N_12349,N_12346);
xor U12573 (N_12573,N_12348,N_12414);
or U12574 (N_12574,N_12374,N_12420);
nand U12575 (N_12575,N_12447,N_12443);
nand U12576 (N_12576,N_12359,N_12400);
or U12577 (N_12577,N_12411,N_12456);
and U12578 (N_12578,N_12386,N_12453);
nor U12579 (N_12579,N_12354,N_12343);
nand U12580 (N_12580,N_12397,N_12327);
and U12581 (N_12581,N_12444,N_12334);
or U12582 (N_12582,N_12352,N_12348);
or U12583 (N_12583,N_12444,N_12335);
or U12584 (N_12584,N_12335,N_12435);
nor U12585 (N_12585,N_12380,N_12440);
xor U12586 (N_12586,N_12436,N_12452);
or U12587 (N_12587,N_12408,N_12398);
or U12588 (N_12588,N_12372,N_12385);
xor U12589 (N_12589,N_12325,N_12411);
nand U12590 (N_12590,N_12476,N_12343);
nor U12591 (N_12591,N_12459,N_12465);
and U12592 (N_12592,N_12355,N_12433);
xor U12593 (N_12593,N_12465,N_12419);
nor U12594 (N_12594,N_12420,N_12348);
or U12595 (N_12595,N_12466,N_12341);
nor U12596 (N_12596,N_12381,N_12383);
or U12597 (N_12597,N_12364,N_12466);
and U12598 (N_12598,N_12337,N_12455);
and U12599 (N_12599,N_12364,N_12408);
or U12600 (N_12600,N_12352,N_12450);
xnor U12601 (N_12601,N_12449,N_12444);
or U12602 (N_12602,N_12341,N_12411);
xnor U12603 (N_12603,N_12323,N_12339);
xnor U12604 (N_12604,N_12396,N_12382);
xnor U12605 (N_12605,N_12326,N_12384);
nor U12606 (N_12606,N_12361,N_12469);
or U12607 (N_12607,N_12322,N_12432);
nor U12608 (N_12608,N_12458,N_12373);
or U12609 (N_12609,N_12399,N_12336);
xor U12610 (N_12610,N_12428,N_12429);
and U12611 (N_12611,N_12344,N_12462);
xnor U12612 (N_12612,N_12325,N_12320);
and U12613 (N_12613,N_12455,N_12380);
or U12614 (N_12614,N_12435,N_12470);
nor U12615 (N_12615,N_12371,N_12460);
and U12616 (N_12616,N_12444,N_12412);
or U12617 (N_12617,N_12431,N_12379);
xnor U12618 (N_12618,N_12333,N_12434);
nor U12619 (N_12619,N_12346,N_12335);
xnor U12620 (N_12620,N_12351,N_12383);
nor U12621 (N_12621,N_12359,N_12425);
and U12622 (N_12622,N_12408,N_12440);
nand U12623 (N_12623,N_12326,N_12419);
nand U12624 (N_12624,N_12373,N_12335);
or U12625 (N_12625,N_12356,N_12464);
nor U12626 (N_12626,N_12449,N_12385);
and U12627 (N_12627,N_12346,N_12399);
and U12628 (N_12628,N_12327,N_12478);
xor U12629 (N_12629,N_12453,N_12455);
and U12630 (N_12630,N_12419,N_12441);
or U12631 (N_12631,N_12414,N_12478);
or U12632 (N_12632,N_12464,N_12427);
xor U12633 (N_12633,N_12327,N_12393);
nand U12634 (N_12634,N_12423,N_12476);
xor U12635 (N_12635,N_12403,N_12471);
or U12636 (N_12636,N_12382,N_12377);
nand U12637 (N_12637,N_12355,N_12327);
and U12638 (N_12638,N_12472,N_12343);
nand U12639 (N_12639,N_12445,N_12401);
xnor U12640 (N_12640,N_12627,N_12583);
xor U12641 (N_12641,N_12534,N_12531);
or U12642 (N_12642,N_12537,N_12570);
nand U12643 (N_12643,N_12555,N_12608);
nor U12644 (N_12644,N_12607,N_12597);
and U12645 (N_12645,N_12571,N_12572);
nand U12646 (N_12646,N_12566,N_12510);
or U12647 (N_12647,N_12581,N_12529);
or U12648 (N_12648,N_12545,N_12511);
nor U12649 (N_12649,N_12500,N_12502);
nand U12650 (N_12650,N_12574,N_12549);
and U12651 (N_12651,N_12526,N_12538);
xnor U12652 (N_12652,N_12576,N_12519);
xor U12653 (N_12653,N_12635,N_12498);
xnor U12654 (N_12654,N_12505,N_12616);
nor U12655 (N_12655,N_12614,N_12528);
xnor U12656 (N_12656,N_12551,N_12518);
xor U12657 (N_12657,N_12630,N_12596);
nand U12658 (N_12658,N_12560,N_12497);
xor U12659 (N_12659,N_12515,N_12632);
or U12660 (N_12660,N_12604,N_12599);
nand U12661 (N_12661,N_12564,N_12554);
nand U12662 (N_12662,N_12633,N_12508);
and U12663 (N_12663,N_12580,N_12568);
and U12664 (N_12664,N_12569,N_12486);
xnor U12665 (N_12665,N_12530,N_12595);
nand U12666 (N_12666,N_12621,N_12586);
nand U12667 (N_12667,N_12482,N_12557);
nand U12668 (N_12668,N_12490,N_12619);
xor U12669 (N_12669,N_12584,N_12638);
and U12670 (N_12670,N_12634,N_12567);
nor U12671 (N_12671,N_12626,N_12598);
nor U12672 (N_12672,N_12600,N_12481);
and U12673 (N_12673,N_12588,N_12577);
nand U12674 (N_12674,N_12590,N_12575);
xnor U12675 (N_12675,N_12629,N_12593);
and U12676 (N_12676,N_12524,N_12532);
xnor U12677 (N_12677,N_12624,N_12506);
and U12678 (N_12678,N_12520,N_12527);
and U12679 (N_12679,N_12546,N_12533);
nand U12680 (N_12680,N_12536,N_12544);
xnor U12681 (N_12681,N_12615,N_12605);
nand U12682 (N_12682,N_12561,N_12503);
nor U12683 (N_12683,N_12541,N_12494);
and U12684 (N_12684,N_12585,N_12514);
or U12685 (N_12685,N_12578,N_12525);
nand U12686 (N_12686,N_12550,N_12542);
and U12687 (N_12687,N_12556,N_12613);
or U12688 (N_12688,N_12573,N_12522);
or U12689 (N_12689,N_12602,N_12483);
nand U12690 (N_12690,N_12507,N_12489);
xor U12691 (N_12691,N_12637,N_12639);
or U12692 (N_12692,N_12558,N_12636);
nor U12693 (N_12693,N_12628,N_12618);
or U12694 (N_12694,N_12487,N_12562);
or U12695 (N_12695,N_12623,N_12543);
nand U12696 (N_12696,N_12540,N_12488);
xnor U12697 (N_12697,N_12587,N_12548);
and U12698 (N_12698,N_12579,N_12603);
xnor U12699 (N_12699,N_12594,N_12601);
and U12700 (N_12700,N_12493,N_12591);
and U12701 (N_12701,N_12492,N_12559);
nand U12702 (N_12702,N_12611,N_12504);
nand U12703 (N_12703,N_12509,N_12631);
nand U12704 (N_12704,N_12499,N_12484);
and U12705 (N_12705,N_12547,N_12609);
and U12706 (N_12706,N_12539,N_12582);
and U12707 (N_12707,N_12617,N_12610);
xnor U12708 (N_12708,N_12523,N_12485);
nor U12709 (N_12709,N_12625,N_12622);
nor U12710 (N_12710,N_12553,N_12512);
nand U12711 (N_12711,N_12565,N_12521);
nor U12712 (N_12712,N_12513,N_12620);
or U12713 (N_12713,N_12491,N_12516);
xor U12714 (N_12714,N_12612,N_12496);
nand U12715 (N_12715,N_12606,N_12517);
nor U12716 (N_12716,N_12592,N_12535);
or U12717 (N_12717,N_12501,N_12480);
or U12718 (N_12718,N_12563,N_12589);
nor U12719 (N_12719,N_12552,N_12495);
and U12720 (N_12720,N_12603,N_12573);
nor U12721 (N_12721,N_12547,N_12573);
nor U12722 (N_12722,N_12578,N_12490);
xnor U12723 (N_12723,N_12630,N_12591);
or U12724 (N_12724,N_12637,N_12503);
and U12725 (N_12725,N_12569,N_12571);
xnor U12726 (N_12726,N_12579,N_12549);
nand U12727 (N_12727,N_12591,N_12609);
nor U12728 (N_12728,N_12524,N_12481);
nor U12729 (N_12729,N_12631,N_12482);
nor U12730 (N_12730,N_12492,N_12484);
or U12731 (N_12731,N_12501,N_12556);
xnor U12732 (N_12732,N_12521,N_12567);
or U12733 (N_12733,N_12489,N_12579);
nand U12734 (N_12734,N_12535,N_12615);
or U12735 (N_12735,N_12609,N_12633);
xor U12736 (N_12736,N_12594,N_12570);
xnor U12737 (N_12737,N_12554,N_12502);
or U12738 (N_12738,N_12606,N_12550);
nand U12739 (N_12739,N_12612,N_12629);
nor U12740 (N_12740,N_12544,N_12541);
and U12741 (N_12741,N_12504,N_12484);
nand U12742 (N_12742,N_12579,N_12627);
or U12743 (N_12743,N_12600,N_12504);
nor U12744 (N_12744,N_12588,N_12571);
nor U12745 (N_12745,N_12568,N_12560);
and U12746 (N_12746,N_12522,N_12607);
nand U12747 (N_12747,N_12513,N_12532);
and U12748 (N_12748,N_12627,N_12562);
xor U12749 (N_12749,N_12517,N_12487);
nand U12750 (N_12750,N_12595,N_12624);
and U12751 (N_12751,N_12543,N_12496);
nand U12752 (N_12752,N_12545,N_12578);
or U12753 (N_12753,N_12607,N_12571);
nand U12754 (N_12754,N_12538,N_12576);
nand U12755 (N_12755,N_12595,N_12574);
nand U12756 (N_12756,N_12511,N_12572);
nor U12757 (N_12757,N_12618,N_12481);
xor U12758 (N_12758,N_12541,N_12556);
and U12759 (N_12759,N_12551,N_12623);
xnor U12760 (N_12760,N_12619,N_12527);
and U12761 (N_12761,N_12638,N_12513);
xnor U12762 (N_12762,N_12621,N_12495);
nand U12763 (N_12763,N_12596,N_12611);
nand U12764 (N_12764,N_12508,N_12507);
xor U12765 (N_12765,N_12615,N_12482);
xor U12766 (N_12766,N_12556,N_12639);
nand U12767 (N_12767,N_12618,N_12489);
xnor U12768 (N_12768,N_12601,N_12489);
or U12769 (N_12769,N_12542,N_12583);
or U12770 (N_12770,N_12522,N_12589);
xnor U12771 (N_12771,N_12541,N_12573);
xnor U12772 (N_12772,N_12594,N_12628);
and U12773 (N_12773,N_12570,N_12529);
or U12774 (N_12774,N_12627,N_12567);
nor U12775 (N_12775,N_12578,N_12615);
and U12776 (N_12776,N_12563,N_12576);
and U12777 (N_12777,N_12527,N_12588);
nor U12778 (N_12778,N_12526,N_12544);
and U12779 (N_12779,N_12506,N_12576);
nand U12780 (N_12780,N_12637,N_12560);
nand U12781 (N_12781,N_12570,N_12606);
and U12782 (N_12782,N_12583,N_12616);
or U12783 (N_12783,N_12581,N_12602);
and U12784 (N_12784,N_12598,N_12633);
xnor U12785 (N_12785,N_12533,N_12629);
and U12786 (N_12786,N_12490,N_12488);
and U12787 (N_12787,N_12618,N_12515);
nand U12788 (N_12788,N_12511,N_12601);
and U12789 (N_12789,N_12483,N_12612);
and U12790 (N_12790,N_12513,N_12510);
xor U12791 (N_12791,N_12638,N_12495);
nor U12792 (N_12792,N_12608,N_12508);
and U12793 (N_12793,N_12548,N_12607);
or U12794 (N_12794,N_12549,N_12538);
and U12795 (N_12795,N_12589,N_12602);
nand U12796 (N_12796,N_12569,N_12492);
nor U12797 (N_12797,N_12571,N_12635);
xnor U12798 (N_12798,N_12573,N_12564);
xnor U12799 (N_12799,N_12549,N_12566);
xor U12800 (N_12800,N_12758,N_12666);
or U12801 (N_12801,N_12659,N_12789);
and U12802 (N_12802,N_12676,N_12646);
or U12803 (N_12803,N_12675,N_12694);
nor U12804 (N_12804,N_12774,N_12660);
nor U12805 (N_12805,N_12664,N_12743);
or U12806 (N_12806,N_12671,N_12641);
xor U12807 (N_12807,N_12689,N_12711);
or U12808 (N_12808,N_12715,N_12765);
and U12809 (N_12809,N_12750,N_12658);
or U12810 (N_12810,N_12643,N_12795);
or U12811 (N_12811,N_12754,N_12681);
nand U12812 (N_12812,N_12776,N_12709);
nor U12813 (N_12813,N_12787,N_12678);
nor U12814 (N_12814,N_12724,N_12642);
nand U12815 (N_12815,N_12751,N_12661);
nor U12816 (N_12816,N_12733,N_12772);
xnor U12817 (N_12817,N_12704,N_12718);
or U12818 (N_12818,N_12712,N_12738);
nand U12819 (N_12819,N_12691,N_12687);
and U12820 (N_12820,N_12727,N_12648);
or U12821 (N_12821,N_12667,N_12730);
or U12822 (N_12822,N_12794,N_12720);
and U12823 (N_12823,N_12753,N_12662);
xnor U12824 (N_12824,N_12645,N_12708);
nor U12825 (N_12825,N_12763,N_12721);
nor U12826 (N_12826,N_12699,N_12655);
nand U12827 (N_12827,N_12663,N_12784);
and U12828 (N_12828,N_12756,N_12732);
nor U12829 (N_12829,N_12734,N_12656);
or U12830 (N_12830,N_12683,N_12652);
xnor U12831 (N_12831,N_12785,N_12755);
or U12832 (N_12832,N_12702,N_12741);
nand U12833 (N_12833,N_12728,N_12697);
and U12834 (N_12834,N_12701,N_12647);
xnor U12835 (N_12835,N_12749,N_12747);
xor U12836 (N_12836,N_12799,N_12792);
xor U12837 (N_12837,N_12767,N_12722);
nor U12838 (N_12838,N_12696,N_12651);
and U12839 (N_12839,N_12737,N_12686);
nor U12840 (N_12840,N_12759,N_12713);
xor U12841 (N_12841,N_12669,N_12672);
xnor U12842 (N_12842,N_12752,N_12716);
or U12843 (N_12843,N_12757,N_12719);
nand U12844 (N_12844,N_12793,N_12698);
xor U12845 (N_12845,N_12788,N_12773);
nand U12846 (N_12846,N_12786,N_12769);
nand U12847 (N_12847,N_12706,N_12726);
nand U12848 (N_12848,N_12778,N_12717);
xor U12849 (N_12849,N_12674,N_12640);
xor U12850 (N_12850,N_12700,N_12770);
or U12851 (N_12851,N_12710,N_12771);
nor U12852 (N_12852,N_12653,N_12690);
nand U12853 (N_12853,N_12791,N_12644);
and U12854 (N_12854,N_12682,N_12766);
nand U12855 (N_12855,N_12725,N_12779);
or U12856 (N_12856,N_12775,N_12739);
and U12857 (N_12857,N_12740,N_12695);
nor U12858 (N_12858,N_12680,N_12692);
nand U12859 (N_12859,N_12729,N_12744);
nor U12860 (N_12860,N_12764,N_12777);
nor U12861 (N_12861,N_12705,N_12670);
and U12862 (N_12862,N_12761,N_12668);
or U12863 (N_12863,N_12745,N_12798);
nand U12864 (N_12864,N_12768,N_12684);
nor U12865 (N_12865,N_12677,N_12782);
nand U12866 (N_12866,N_12703,N_12707);
nor U12867 (N_12867,N_12783,N_12746);
or U12868 (N_12868,N_12796,N_12781);
or U12869 (N_12869,N_12780,N_12762);
nor U12870 (N_12870,N_12797,N_12688);
xnor U12871 (N_12871,N_12735,N_12679);
or U12872 (N_12872,N_12736,N_12790);
and U12873 (N_12873,N_12760,N_12731);
and U12874 (N_12874,N_12673,N_12685);
xor U12875 (N_12875,N_12649,N_12748);
and U12876 (N_12876,N_12654,N_12650);
and U12877 (N_12877,N_12723,N_12657);
nor U12878 (N_12878,N_12742,N_12714);
and U12879 (N_12879,N_12665,N_12693);
nor U12880 (N_12880,N_12774,N_12781);
xor U12881 (N_12881,N_12789,N_12750);
xnor U12882 (N_12882,N_12694,N_12695);
nor U12883 (N_12883,N_12796,N_12726);
and U12884 (N_12884,N_12795,N_12678);
and U12885 (N_12885,N_12754,N_12698);
nor U12886 (N_12886,N_12752,N_12676);
or U12887 (N_12887,N_12703,N_12777);
or U12888 (N_12888,N_12685,N_12717);
nand U12889 (N_12889,N_12737,N_12799);
nor U12890 (N_12890,N_12694,N_12775);
and U12891 (N_12891,N_12766,N_12778);
and U12892 (N_12892,N_12776,N_12753);
xor U12893 (N_12893,N_12784,N_12749);
and U12894 (N_12894,N_12755,N_12778);
or U12895 (N_12895,N_12706,N_12731);
xnor U12896 (N_12896,N_12657,N_12693);
xnor U12897 (N_12897,N_12728,N_12716);
nor U12898 (N_12898,N_12710,N_12686);
xnor U12899 (N_12899,N_12762,N_12655);
or U12900 (N_12900,N_12711,N_12687);
and U12901 (N_12901,N_12695,N_12668);
or U12902 (N_12902,N_12744,N_12695);
nor U12903 (N_12903,N_12707,N_12640);
nand U12904 (N_12904,N_12788,N_12761);
or U12905 (N_12905,N_12759,N_12701);
nand U12906 (N_12906,N_12713,N_12722);
or U12907 (N_12907,N_12666,N_12702);
nor U12908 (N_12908,N_12701,N_12768);
and U12909 (N_12909,N_12739,N_12672);
nor U12910 (N_12910,N_12698,N_12708);
and U12911 (N_12911,N_12736,N_12688);
nand U12912 (N_12912,N_12656,N_12749);
nor U12913 (N_12913,N_12767,N_12671);
nand U12914 (N_12914,N_12654,N_12778);
nand U12915 (N_12915,N_12684,N_12645);
xnor U12916 (N_12916,N_12719,N_12783);
xor U12917 (N_12917,N_12697,N_12734);
or U12918 (N_12918,N_12733,N_12656);
nor U12919 (N_12919,N_12751,N_12651);
or U12920 (N_12920,N_12712,N_12727);
and U12921 (N_12921,N_12642,N_12666);
and U12922 (N_12922,N_12778,N_12747);
nand U12923 (N_12923,N_12669,N_12643);
and U12924 (N_12924,N_12662,N_12729);
and U12925 (N_12925,N_12786,N_12779);
nand U12926 (N_12926,N_12718,N_12728);
nor U12927 (N_12927,N_12653,N_12799);
nor U12928 (N_12928,N_12752,N_12781);
xor U12929 (N_12929,N_12760,N_12655);
and U12930 (N_12930,N_12749,N_12709);
nand U12931 (N_12931,N_12796,N_12732);
and U12932 (N_12932,N_12774,N_12790);
and U12933 (N_12933,N_12663,N_12670);
or U12934 (N_12934,N_12705,N_12750);
nand U12935 (N_12935,N_12670,N_12643);
nor U12936 (N_12936,N_12678,N_12727);
nor U12937 (N_12937,N_12757,N_12717);
and U12938 (N_12938,N_12733,N_12659);
nand U12939 (N_12939,N_12702,N_12791);
and U12940 (N_12940,N_12694,N_12790);
nand U12941 (N_12941,N_12722,N_12665);
nor U12942 (N_12942,N_12723,N_12731);
and U12943 (N_12943,N_12740,N_12746);
xor U12944 (N_12944,N_12675,N_12688);
or U12945 (N_12945,N_12760,N_12642);
nand U12946 (N_12946,N_12763,N_12742);
nor U12947 (N_12947,N_12796,N_12656);
or U12948 (N_12948,N_12641,N_12643);
xor U12949 (N_12949,N_12699,N_12677);
and U12950 (N_12950,N_12716,N_12647);
or U12951 (N_12951,N_12795,N_12791);
or U12952 (N_12952,N_12726,N_12780);
nand U12953 (N_12953,N_12751,N_12741);
nor U12954 (N_12954,N_12677,N_12724);
or U12955 (N_12955,N_12737,N_12684);
nand U12956 (N_12956,N_12640,N_12720);
or U12957 (N_12957,N_12750,N_12691);
or U12958 (N_12958,N_12715,N_12794);
nand U12959 (N_12959,N_12649,N_12792);
or U12960 (N_12960,N_12900,N_12927);
nor U12961 (N_12961,N_12824,N_12953);
xnor U12962 (N_12962,N_12882,N_12856);
xnor U12963 (N_12963,N_12901,N_12846);
xor U12964 (N_12964,N_12865,N_12845);
xnor U12965 (N_12965,N_12866,N_12903);
and U12966 (N_12966,N_12832,N_12844);
and U12967 (N_12967,N_12841,N_12908);
nand U12968 (N_12968,N_12802,N_12848);
and U12969 (N_12969,N_12909,N_12890);
nand U12970 (N_12970,N_12859,N_12835);
or U12971 (N_12971,N_12899,N_12852);
xnor U12972 (N_12972,N_12923,N_12884);
xnor U12973 (N_12973,N_12810,N_12888);
nand U12974 (N_12974,N_12956,N_12877);
nand U12975 (N_12975,N_12922,N_12941);
or U12976 (N_12976,N_12860,N_12915);
nor U12977 (N_12977,N_12934,N_12834);
and U12978 (N_12978,N_12878,N_12943);
nand U12979 (N_12979,N_12838,N_12914);
and U12980 (N_12980,N_12849,N_12818);
xnor U12981 (N_12981,N_12843,N_12812);
nor U12982 (N_12982,N_12942,N_12836);
nor U12983 (N_12983,N_12898,N_12958);
nor U12984 (N_12984,N_12921,N_12815);
nor U12985 (N_12985,N_12930,N_12938);
or U12986 (N_12986,N_12857,N_12875);
nand U12987 (N_12987,N_12807,N_12946);
and U12988 (N_12988,N_12891,N_12904);
or U12989 (N_12989,N_12868,N_12840);
nand U12990 (N_12990,N_12851,N_12804);
nor U12991 (N_12991,N_12842,N_12881);
xnor U12992 (N_12992,N_12825,N_12952);
nand U12993 (N_12993,N_12855,N_12907);
or U12994 (N_12994,N_12826,N_12803);
or U12995 (N_12995,N_12918,N_12885);
and U12996 (N_12996,N_12853,N_12837);
nand U12997 (N_12997,N_12831,N_12910);
or U12998 (N_12998,N_12827,N_12811);
nor U12999 (N_12999,N_12896,N_12945);
or U13000 (N_13000,N_12872,N_12912);
xor U13001 (N_13001,N_12905,N_12933);
or U13002 (N_13002,N_12949,N_12948);
nor U13003 (N_13003,N_12839,N_12954);
nand U13004 (N_13004,N_12847,N_12821);
nor U13005 (N_13005,N_12830,N_12957);
nand U13006 (N_13006,N_12858,N_12928);
or U13007 (N_13007,N_12816,N_12886);
xor U13008 (N_13008,N_12864,N_12808);
xor U13009 (N_13009,N_12913,N_12889);
nand U13010 (N_13010,N_12919,N_12820);
or U13011 (N_13011,N_12880,N_12873);
and U13012 (N_13012,N_12959,N_12828);
and U13013 (N_13013,N_12926,N_12876);
and U13014 (N_13014,N_12937,N_12863);
or U13015 (N_13015,N_12813,N_12944);
or U13016 (N_13016,N_12939,N_12822);
or U13017 (N_13017,N_12879,N_12809);
nor U13018 (N_13018,N_12906,N_12870);
xor U13019 (N_13019,N_12867,N_12801);
nand U13020 (N_13020,N_12911,N_12947);
xnor U13021 (N_13021,N_12819,N_12924);
or U13022 (N_13022,N_12929,N_12823);
nand U13023 (N_13023,N_12861,N_12833);
or U13024 (N_13024,N_12869,N_12883);
or U13025 (N_13025,N_12925,N_12916);
nor U13026 (N_13026,N_12955,N_12874);
or U13027 (N_13027,N_12814,N_12892);
xnor U13028 (N_13028,N_12806,N_12817);
and U13029 (N_13029,N_12950,N_12854);
xnor U13030 (N_13030,N_12887,N_12917);
xor U13031 (N_13031,N_12894,N_12871);
nand U13032 (N_13032,N_12936,N_12951);
xor U13033 (N_13033,N_12893,N_12897);
or U13034 (N_13034,N_12940,N_12829);
nand U13035 (N_13035,N_12920,N_12805);
nand U13036 (N_13036,N_12902,N_12931);
nand U13037 (N_13037,N_12932,N_12850);
or U13038 (N_13038,N_12935,N_12895);
and U13039 (N_13039,N_12800,N_12862);
xnor U13040 (N_13040,N_12888,N_12925);
nor U13041 (N_13041,N_12878,N_12888);
and U13042 (N_13042,N_12935,N_12957);
nand U13043 (N_13043,N_12878,N_12898);
or U13044 (N_13044,N_12828,N_12951);
nor U13045 (N_13045,N_12803,N_12808);
nor U13046 (N_13046,N_12806,N_12946);
xnor U13047 (N_13047,N_12903,N_12842);
nand U13048 (N_13048,N_12808,N_12908);
nand U13049 (N_13049,N_12864,N_12869);
xnor U13050 (N_13050,N_12953,N_12803);
xnor U13051 (N_13051,N_12949,N_12862);
xor U13052 (N_13052,N_12805,N_12880);
and U13053 (N_13053,N_12807,N_12940);
nor U13054 (N_13054,N_12922,N_12932);
and U13055 (N_13055,N_12895,N_12884);
nand U13056 (N_13056,N_12928,N_12905);
nor U13057 (N_13057,N_12955,N_12800);
and U13058 (N_13058,N_12894,N_12887);
and U13059 (N_13059,N_12823,N_12904);
or U13060 (N_13060,N_12883,N_12909);
and U13061 (N_13061,N_12902,N_12873);
xnor U13062 (N_13062,N_12918,N_12934);
and U13063 (N_13063,N_12826,N_12821);
or U13064 (N_13064,N_12820,N_12896);
or U13065 (N_13065,N_12946,N_12920);
nand U13066 (N_13066,N_12921,N_12939);
or U13067 (N_13067,N_12896,N_12898);
nor U13068 (N_13068,N_12955,N_12887);
nor U13069 (N_13069,N_12883,N_12898);
and U13070 (N_13070,N_12856,N_12848);
nand U13071 (N_13071,N_12934,N_12926);
nand U13072 (N_13072,N_12946,N_12814);
or U13073 (N_13073,N_12947,N_12897);
xnor U13074 (N_13074,N_12829,N_12866);
nand U13075 (N_13075,N_12959,N_12934);
nand U13076 (N_13076,N_12870,N_12840);
or U13077 (N_13077,N_12952,N_12959);
xnor U13078 (N_13078,N_12897,N_12880);
nand U13079 (N_13079,N_12877,N_12954);
nor U13080 (N_13080,N_12820,N_12818);
xnor U13081 (N_13081,N_12925,N_12851);
xor U13082 (N_13082,N_12900,N_12902);
or U13083 (N_13083,N_12903,N_12870);
or U13084 (N_13084,N_12947,N_12887);
and U13085 (N_13085,N_12811,N_12822);
nor U13086 (N_13086,N_12839,N_12921);
xnor U13087 (N_13087,N_12855,N_12868);
and U13088 (N_13088,N_12815,N_12829);
or U13089 (N_13089,N_12923,N_12947);
xor U13090 (N_13090,N_12917,N_12838);
xnor U13091 (N_13091,N_12884,N_12846);
nor U13092 (N_13092,N_12954,N_12956);
xnor U13093 (N_13093,N_12833,N_12915);
nor U13094 (N_13094,N_12881,N_12914);
nand U13095 (N_13095,N_12863,N_12870);
nor U13096 (N_13096,N_12911,N_12856);
nand U13097 (N_13097,N_12854,N_12922);
xor U13098 (N_13098,N_12849,N_12901);
or U13099 (N_13099,N_12808,N_12853);
nand U13100 (N_13100,N_12912,N_12842);
or U13101 (N_13101,N_12889,N_12872);
xnor U13102 (N_13102,N_12917,N_12918);
xor U13103 (N_13103,N_12894,N_12888);
xnor U13104 (N_13104,N_12829,N_12819);
xor U13105 (N_13105,N_12843,N_12850);
and U13106 (N_13106,N_12858,N_12872);
and U13107 (N_13107,N_12857,N_12891);
or U13108 (N_13108,N_12896,N_12821);
and U13109 (N_13109,N_12926,N_12941);
nor U13110 (N_13110,N_12921,N_12908);
and U13111 (N_13111,N_12925,N_12828);
xnor U13112 (N_13112,N_12933,N_12953);
nand U13113 (N_13113,N_12885,N_12814);
xnor U13114 (N_13114,N_12851,N_12875);
xor U13115 (N_13115,N_12878,N_12931);
and U13116 (N_13116,N_12942,N_12852);
and U13117 (N_13117,N_12852,N_12844);
and U13118 (N_13118,N_12911,N_12909);
nor U13119 (N_13119,N_12957,N_12842);
xnor U13120 (N_13120,N_13111,N_13010);
or U13121 (N_13121,N_13069,N_13113);
and U13122 (N_13122,N_13104,N_13102);
nor U13123 (N_13123,N_13107,N_13086);
and U13124 (N_13124,N_13071,N_13022);
nor U13125 (N_13125,N_13060,N_13002);
and U13126 (N_13126,N_13096,N_12970);
nand U13127 (N_13127,N_13003,N_13036);
nand U13128 (N_13128,N_12987,N_13074);
nand U13129 (N_13129,N_13065,N_13034);
or U13130 (N_13130,N_12991,N_13118);
nor U13131 (N_13131,N_13042,N_12977);
and U13132 (N_13132,N_13011,N_12992);
nor U13133 (N_13133,N_12981,N_12961);
nand U13134 (N_13134,N_13035,N_13017);
nor U13135 (N_13135,N_13047,N_12986);
and U13136 (N_13136,N_13117,N_13044);
xor U13137 (N_13137,N_13062,N_12976);
or U13138 (N_13138,N_13066,N_13025);
nand U13139 (N_13139,N_13038,N_13080);
nor U13140 (N_13140,N_13006,N_13112);
xnor U13141 (N_13141,N_12985,N_13001);
and U13142 (N_13142,N_13109,N_13051);
or U13143 (N_13143,N_12975,N_13054);
and U13144 (N_13144,N_13043,N_12969);
or U13145 (N_13145,N_13018,N_13024);
nor U13146 (N_13146,N_13082,N_13059);
nand U13147 (N_13147,N_13081,N_13068);
nor U13148 (N_13148,N_13108,N_12965);
or U13149 (N_13149,N_13105,N_13037);
or U13150 (N_13150,N_13028,N_13005);
nor U13151 (N_13151,N_13046,N_13067);
nand U13152 (N_13152,N_13099,N_12999);
nor U13153 (N_13153,N_13097,N_13100);
or U13154 (N_13154,N_12998,N_13088);
nor U13155 (N_13155,N_13052,N_13033);
nand U13156 (N_13156,N_13106,N_13076);
xor U13157 (N_13157,N_13084,N_13055);
nor U13158 (N_13158,N_13009,N_13029);
nand U13159 (N_13159,N_12994,N_12982);
and U13160 (N_13160,N_13061,N_12974);
nor U13161 (N_13161,N_13089,N_13072);
nand U13162 (N_13162,N_13053,N_12997);
xnor U13163 (N_13163,N_13023,N_12990);
and U13164 (N_13164,N_13016,N_13083);
xor U13165 (N_13165,N_13116,N_12960);
nor U13166 (N_13166,N_12962,N_12993);
and U13167 (N_13167,N_13098,N_12979);
xor U13168 (N_13168,N_13090,N_12984);
xor U13169 (N_13169,N_13114,N_13073);
nor U13170 (N_13170,N_13040,N_13075);
xnor U13171 (N_13171,N_13004,N_13103);
nand U13172 (N_13172,N_13048,N_13115);
xnor U13173 (N_13173,N_13019,N_13058);
nand U13174 (N_13174,N_13027,N_13026);
xnor U13175 (N_13175,N_13056,N_13078);
and U13176 (N_13176,N_12980,N_13077);
and U13177 (N_13177,N_13039,N_13057);
and U13178 (N_13178,N_12967,N_12971);
or U13179 (N_13179,N_12968,N_13021);
nor U13180 (N_13180,N_13012,N_13091);
and U13181 (N_13181,N_13014,N_12963);
nand U13182 (N_13182,N_13110,N_13101);
and U13183 (N_13183,N_13000,N_12973);
and U13184 (N_13184,N_13093,N_13095);
and U13185 (N_13185,N_13049,N_13041);
or U13186 (N_13186,N_13013,N_13031);
xor U13187 (N_13187,N_12966,N_12983);
and U13188 (N_13188,N_13094,N_13008);
xnor U13189 (N_13189,N_13063,N_13015);
and U13190 (N_13190,N_13030,N_13087);
nand U13191 (N_13191,N_13119,N_12972);
and U13192 (N_13192,N_13045,N_12988);
nand U13193 (N_13193,N_12989,N_12964);
nor U13194 (N_13194,N_13085,N_12995);
nor U13195 (N_13195,N_13032,N_13092);
nor U13196 (N_13196,N_13079,N_12978);
nor U13197 (N_13197,N_13020,N_13050);
nand U13198 (N_13198,N_12996,N_13007);
nand U13199 (N_13199,N_13064,N_13070);
and U13200 (N_13200,N_13078,N_13036);
nand U13201 (N_13201,N_13096,N_13056);
nand U13202 (N_13202,N_13115,N_12995);
nand U13203 (N_13203,N_12962,N_13084);
nand U13204 (N_13204,N_13102,N_13081);
xor U13205 (N_13205,N_13007,N_12962);
nand U13206 (N_13206,N_13110,N_12997);
nor U13207 (N_13207,N_12970,N_13117);
nand U13208 (N_13208,N_12966,N_13062);
and U13209 (N_13209,N_13026,N_13111);
nand U13210 (N_13210,N_13006,N_12991);
xor U13211 (N_13211,N_12977,N_13032);
nor U13212 (N_13212,N_13078,N_13067);
xor U13213 (N_13213,N_13112,N_13034);
and U13214 (N_13214,N_13049,N_12981);
or U13215 (N_13215,N_13092,N_13065);
xnor U13216 (N_13216,N_12991,N_13094);
nor U13217 (N_13217,N_13063,N_13087);
xor U13218 (N_13218,N_12967,N_13063);
nor U13219 (N_13219,N_13107,N_13044);
nand U13220 (N_13220,N_13050,N_12975);
and U13221 (N_13221,N_13056,N_13119);
and U13222 (N_13222,N_13069,N_13052);
nor U13223 (N_13223,N_13061,N_12995);
or U13224 (N_13224,N_13080,N_13014);
xor U13225 (N_13225,N_13001,N_13017);
nand U13226 (N_13226,N_13007,N_13054);
xor U13227 (N_13227,N_13034,N_13045);
nor U13228 (N_13228,N_13105,N_12981);
xor U13229 (N_13229,N_13020,N_13003);
nand U13230 (N_13230,N_12972,N_13066);
nor U13231 (N_13231,N_12985,N_12988);
and U13232 (N_13232,N_13081,N_13049);
nor U13233 (N_13233,N_13112,N_13081);
nor U13234 (N_13234,N_13113,N_13020);
xor U13235 (N_13235,N_13100,N_13010);
xor U13236 (N_13236,N_13043,N_13031);
xnor U13237 (N_13237,N_13055,N_12961);
and U13238 (N_13238,N_13104,N_13065);
and U13239 (N_13239,N_13047,N_12988);
or U13240 (N_13240,N_13009,N_13024);
and U13241 (N_13241,N_13109,N_13119);
nand U13242 (N_13242,N_13005,N_13044);
or U13243 (N_13243,N_13068,N_13049);
xnor U13244 (N_13244,N_13118,N_13100);
xnor U13245 (N_13245,N_13004,N_13080);
xor U13246 (N_13246,N_12985,N_13111);
and U13247 (N_13247,N_13018,N_13080);
xor U13248 (N_13248,N_13041,N_13092);
xor U13249 (N_13249,N_13119,N_13012);
xor U13250 (N_13250,N_13035,N_13039);
nor U13251 (N_13251,N_13052,N_13064);
nor U13252 (N_13252,N_12978,N_13030);
nand U13253 (N_13253,N_12988,N_13095);
nand U13254 (N_13254,N_13070,N_13119);
xor U13255 (N_13255,N_13114,N_13012);
or U13256 (N_13256,N_13037,N_13073);
xnor U13257 (N_13257,N_13036,N_13070);
nor U13258 (N_13258,N_13067,N_13033);
and U13259 (N_13259,N_13059,N_13043);
or U13260 (N_13260,N_13007,N_13052);
xor U13261 (N_13261,N_13068,N_12967);
nor U13262 (N_13262,N_13091,N_13054);
or U13263 (N_13263,N_13101,N_13027);
and U13264 (N_13264,N_12985,N_13073);
nor U13265 (N_13265,N_13113,N_13077);
nor U13266 (N_13266,N_13004,N_12979);
or U13267 (N_13267,N_12984,N_12995);
xnor U13268 (N_13268,N_12984,N_13059);
or U13269 (N_13269,N_12965,N_13081);
nor U13270 (N_13270,N_13054,N_13036);
xnor U13271 (N_13271,N_13087,N_13015);
or U13272 (N_13272,N_13085,N_13037);
or U13273 (N_13273,N_13055,N_13105);
and U13274 (N_13274,N_12963,N_13069);
nand U13275 (N_13275,N_12972,N_13077);
nand U13276 (N_13276,N_13066,N_12988);
or U13277 (N_13277,N_13116,N_13013);
nand U13278 (N_13278,N_13086,N_12987);
nor U13279 (N_13279,N_13014,N_13059);
and U13280 (N_13280,N_13167,N_13155);
or U13281 (N_13281,N_13274,N_13189);
nand U13282 (N_13282,N_13158,N_13163);
nand U13283 (N_13283,N_13276,N_13252);
nand U13284 (N_13284,N_13211,N_13132);
xor U13285 (N_13285,N_13157,N_13187);
nand U13286 (N_13286,N_13168,N_13150);
nor U13287 (N_13287,N_13166,N_13208);
or U13288 (N_13288,N_13230,N_13193);
nor U13289 (N_13289,N_13121,N_13268);
xor U13290 (N_13290,N_13179,N_13220);
xnor U13291 (N_13291,N_13237,N_13260);
or U13292 (N_13292,N_13266,N_13241);
and U13293 (N_13293,N_13156,N_13209);
xor U13294 (N_13294,N_13272,N_13191);
nand U13295 (N_13295,N_13217,N_13178);
or U13296 (N_13296,N_13173,N_13122);
nand U13297 (N_13297,N_13257,N_13259);
nor U13298 (N_13298,N_13131,N_13232);
xor U13299 (N_13299,N_13176,N_13244);
nor U13300 (N_13300,N_13123,N_13261);
nor U13301 (N_13301,N_13127,N_13222);
and U13302 (N_13302,N_13223,N_13231);
xor U13303 (N_13303,N_13253,N_13125);
nand U13304 (N_13304,N_13174,N_13200);
or U13305 (N_13305,N_13201,N_13198);
nor U13306 (N_13306,N_13169,N_13188);
xnor U13307 (N_13307,N_13250,N_13145);
and U13308 (N_13308,N_13172,N_13271);
or U13309 (N_13309,N_13204,N_13182);
and U13310 (N_13310,N_13219,N_13248);
or U13311 (N_13311,N_13228,N_13210);
nand U13312 (N_13312,N_13245,N_13240);
and U13313 (N_13313,N_13161,N_13226);
or U13314 (N_13314,N_13148,N_13141);
nor U13315 (N_13315,N_13277,N_13196);
and U13316 (N_13316,N_13243,N_13153);
and U13317 (N_13317,N_13258,N_13267);
nor U13318 (N_13318,N_13236,N_13207);
and U13319 (N_13319,N_13235,N_13275);
and U13320 (N_13320,N_13190,N_13137);
nand U13321 (N_13321,N_13227,N_13130);
nand U13322 (N_13322,N_13213,N_13262);
nand U13323 (N_13323,N_13264,N_13170);
xnor U13324 (N_13324,N_13234,N_13133);
nor U13325 (N_13325,N_13256,N_13184);
xnor U13326 (N_13326,N_13181,N_13195);
nor U13327 (N_13327,N_13238,N_13194);
or U13328 (N_13328,N_13147,N_13242);
nand U13329 (N_13329,N_13151,N_13254);
nand U13330 (N_13330,N_13136,N_13139);
xor U13331 (N_13331,N_13177,N_13216);
or U13332 (N_13332,N_13214,N_13159);
or U13333 (N_13333,N_13185,N_13206);
nand U13334 (N_13334,N_13229,N_13263);
or U13335 (N_13335,N_13203,N_13225);
and U13336 (N_13336,N_13205,N_13140);
xnor U13337 (N_13337,N_13197,N_13154);
and U13338 (N_13338,N_13249,N_13162);
nand U13339 (N_13339,N_13134,N_13124);
xnor U13340 (N_13340,N_13143,N_13164);
nand U13341 (N_13341,N_13233,N_13224);
nor U13342 (N_13342,N_13192,N_13215);
nor U13343 (N_13343,N_13183,N_13212);
xnor U13344 (N_13344,N_13165,N_13239);
and U13345 (N_13345,N_13138,N_13269);
or U13346 (N_13346,N_13270,N_13128);
or U13347 (N_13347,N_13202,N_13126);
nor U13348 (N_13348,N_13255,N_13120);
nand U13349 (N_13349,N_13218,N_13247);
nor U13350 (N_13350,N_13142,N_13199);
nor U13351 (N_13351,N_13246,N_13129);
or U13352 (N_13352,N_13144,N_13180);
or U13353 (N_13353,N_13149,N_13273);
and U13354 (N_13354,N_13175,N_13186);
and U13355 (N_13355,N_13171,N_13265);
nor U13356 (N_13356,N_13152,N_13160);
and U13357 (N_13357,N_13135,N_13251);
or U13358 (N_13358,N_13278,N_13279);
xnor U13359 (N_13359,N_13146,N_13221);
or U13360 (N_13360,N_13259,N_13228);
or U13361 (N_13361,N_13271,N_13269);
nor U13362 (N_13362,N_13130,N_13125);
nand U13363 (N_13363,N_13159,N_13153);
xnor U13364 (N_13364,N_13274,N_13278);
or U13365 (N_13365,N_13172,N_13265);
and U13366 (N_13366,N_13122,N_13166);
nor U13367 (N_13367,N_13157,N_13244);
nor U13368 (N_13368,N_13255,N_13129);
or U13369 (N_13369,N_13181,N_13144);
and U13370 (N_13370,N_13184,N_13273);
and U13371 (N_13371,N_13120,N_13223);
xor U13372 (N_13372,N_13220,N_13214);
and U13373 (N_13373,N_13152,N_13128);
and U13374 (N_13374,N_13170,N_13150);
and U13375 (N_13375,N_13151,N_13156);
xnor U13376 (N_13376,N_13128,N_13229);
nand U13377 (N_13377,N_13277,N_13126);
xor U13378 (N_13378,N_13142,N_13183);
or U13379 (N_13379,N_13249,N_13128);
xnor U13380 (N_13380,N_13152,N_13220);
or U13381 (N_13381,N_13261,N_13208);
or U13382 (N_13382,N_13231,N_13237);
xnor U13383 (N_13383,N_13257,N_13156);
and U13384 (N_13384,N_13153,N_13219);
or U13385 (N_13385,N_13279,N_13168);
or U13386 (N_13386,N_13146,N_13177);
nand U13387 (N_13387,N_13194,N_13153);
nand U13388 (N_13388,N_13134,N_13155);
xor U13389 (N_13389,N_13129,N_13131);
and U13390 (N_13390,N_13197,N_13249);
nand U13391 (N_13391,N_13172,N_13181);
and U13392 (N_13392,N_13218,N_13141);
xor U13393 (N_13393,N_13269,N_13207);
xor U13394 (N_13394,N_13263,N_13214);
xnor U13395 (N_13395,N_13247,N_13158);
nand U13396 (N_13396,N_13122,N_13124);
and U13397 (N_13397,N_13129,N_13189);
xor U13398 (N_13398,N_13225,N_13218);
xor U13399 (N_13399,N_13271,N_13202);
nand U13400 (N_13400,N_13272,N_13270);
xor U13401 (N_13401,N_13233,N_13207);
and U13402 (N_13402,N_13228,N_13220);
xnor U13403 (N_13403,N_13130,N_13173);
nand U13404 (N_13404,N_13120,N_13162);
xor U13405 (N_13405,N_13186,N_13147);
nand U13406 (N_13406,N_13229,N_13204);
xnor U13407 (N_13407,N_13203,N_13256);
nor U13408 (N_13408,N_13240,N_13144);
nand U13409 (N_13409,N_13191,N_13231);
nor U13410 (N_13410,N_13178,N_13244);
xnor U13411 (N_13411,N_13251,N_13196);
and U13412 (N_13412,N_13209,N_13271);
nand U13413 (N_13413,N_13122,N_13156);
nand U13414 (N_13414,N_13254,N_13259);
or U13415 (N_13415,N_13139,N_13186);
xor U13416 (N_13416,N_13185,N_13232);
xnor U13417 (N_13417,N_13126,N_13241);
nand U13418 (N_13418,N_13157,N_13202);
or U13419 (N_13419,N_13172,N_13167);
or U13420 (N_13420,N_13276,N_13162);
or U13421 (N_13421,N_13256,N_13183);
nand U13422 (N_13422,N_13229,N_13217);
or U13423 (N_13423,N_13167,N_13144);
nand U13424 (N_13424,N_13245,N_13183);
xnor U13425 (N_13425,N_13129,N_13181);
nor U13426 (N_13426,N_13260,N_13194);
xor U13427 (N_13427,N_13273,N_13277);
nor U13428 (N_13428,N_13126,N_13235);
or U13429 (N_13429,N_13239,N_13151);
or U13430 (N_13430,N_13262,N_13221);
and U13431 (N_13431,N_13198,N_13167);
nor U13432 (N_13432,N_13126,N_13210);
xor U13433 (N_13433,N_13227,N_13171);
xnor U13434 (N_13434,N_13276,N_13232);
nand U13435 (N_13435,N_13137,N_13161);
or U13436 (N_13436,N_13274,N_13133);
xnor U13437 (N_13437,N_13270,N_13208);
and U13438 (N_13438,N_13279,N_13126);
xnor U13439 (N_13439,N_13157,N_13150);
nand U13440 (N_13440,N_13292,N_13390);
and U13441 (N_13441,N_13321,N_13367);
nand U13442 (N_13442,N_13378,N_13432);
nand U13443 (N_13443,N_13335,N_13424);
xnor U13444 (N_13444,N_13293,N_13286);
nor U13445 (N_13445,N_13309,N_13403);
or U13446 (N_13446,N_13434,N_13338);
nand U13447 (N_13447,N_13337,N_13412);
nor U13448 (N_13448,N_13359,N_13428);
or U13449 (N_13449,N_13426,N_13388);
nand U13450 (N_13450,N_13304,N_13352);
xnor U13451 (N_13451,N_13281,N_13384);
and U13452 (N_13452,N_13353,N_13336);
nand U13453 (N_13453,N_13316,N_13408);
nor U13454 (N_13454,N_13413,N_13411);
xor U13455 (N_13455,N_13333,N_13297);
nor U13456 (N_13456,N_13416,N_13280);
and U13457 (N_13457,N_13393,N_13398);
xnor U13458 (N_13458,N_13318,N_13366);
nor U13459 (N_13459,N_13394,N_13389);
xnor U13460 (N_13460,N_13294,N_13395);
xnor U13461 (N_13461,N_13298,N_13377);
and U13462 (N_13462,N_13355,N_13375);
xor U13463 (N_13463,N_13414,N_13332);
nor U13464 (N_13464,N_13427,N_13320);
and U13465 (N_13465,N_13420,N_13369);
nand U13466 (N_13466,N_13307,N_13419);
or U13467 (N_13467,N_13402,N_13284);
nor U13468 (N_13468,N_13439,N_13285);
or U13469 (N_13469,N_13331,N_13317);
nand U13470 (N_13470,N_13396,N_13409);
or U13471 (N_13471,N_13404,N_13370);
nor U13472 (N_13472,N_13374,N_13417);
xor U13473 (N_13473,N_13334,N_13382);
nand U13474 (N_13474,N_13422,N_13385);
nand U13475 (N_13475,N_13328,N_13364);
or U13476 (N_13476,N_13310,N_13347);
nor U13477 (N_13477,N_13387,N_13429);
nor U13478 (N_13478,N_13344,N_13392);
nor U13479 (N_13479,N_13324,N_13283);
and U13480 (N_13480,N_13350,N_13348);
xor U13481 (N_13481,N_13365,N_13372);
and U13482 (N_13482,N_13421,N_13371);
nand U13483 (N_13483,N_13399,N_13343);
nor U13484 (N_13484,N_13308,N_13291);
and U13485 (N_13485,N_13360,N_13368);
or U13486 (N_13486,N_13325,N_13289);
nand U13487 (N_13487,N_13322,N_13423);
nor U13488 (N_13488,N_13376,N_13300);
nand U13489 (N_13489,N_13379,N_13357);
and U13490 (N_13490,N_13341,N_13346);
xnor U13491 (N_13491,N_13288,N_13386);
and U13492 (N_13492,N_13430,N_13407);
or U13493 (N_13493,N_13342,N_13349);
xor U13494 (N_13494,N_13391,N_13330);
xor U13495 (N_13495,N_13299,N_13438);
nand U13496 (N_13496,N_13305,N_13358);
nand U13497 (N_13497,N_13356,N_13361);
or U13498 (N_13498,N_13296,N_13362);
xnor U13499 (N_13499,N_13351,N_13415);
nand U13500 (N_13500,N_13381,N_13400);
nand U13501 (N_13501,N_13437,N_13418);
or U13502 (N_13502,N_13397,N_13436);
and U13503 (N_13503,N_13340,N_13287);
and U13504 (N_13504,N_13302,N_13319);
nand U13505 (N_13505,N_13301,N_13311);
or U13506 (N_13506,N_13313,N_13323);
nor U13507 (N_13507,N_13306,N_13425);
nor U13508 (N_13508,N_13380,N_13312);
xor U13509 (N_13509,N_13326,N_13345);
nand U13510 (N_13510,N_13295,N_13431);
or U13511 (N_13511,N_13303,N_13282);
nor U13512 (N_13512,N_13406,N_13314);
nand U13513 (N_13513,N_13363,N_13354);
or U13514 (N_13514,N_13373,N_13401);
and U13515 (N_13515,N_13435,N_13410);
or U13516 (N_13516,N_13433,N_13327);
nor U13517 (N_13517,N_13315,N_13383);
nand U13518 (N_13518,N_13290,N_13339);
or U13519 (N_13519,N_13329,N_13405);
or U13520 (N_13520,N_13347,N_13367);
and U13521 (N_13521,N_13328,N_13309);
xnor U13522 (N_13522,N_13386,N_13349);
or U13523 (N_13523,N_13396,N_13435);
or U13524 (N_13524,N_13286,N_13315);
nor U13525 (N_13525,N_13410,N_13393);
nor U13526 (N_13526,N_13361,N_13303);
nand U13527 (N_13527,N_13384,N_13285);
nand U13528 (N_13528,N_13380,N_13360);
nand U13529 (N_13529,N_13346,N_13439);
or U13530 (N_13530,N_13418,N_13334);
xor U13531 (N_13531,N_13371,N_13404);
nand U13532 (N_13532,N_13321,N_13427);
nand U13533 (N_13533,N_13414,N_13281);
nand U13534 (N_13534,N_13382,N_13357);
or U13535 (N_13535,N_13404,N_13365);
nand U13536 (N_13536,N_13282,N_13358);
and U13537 (N_13537,N_13297,N_13334);
xnor U13538 (N_13538,N_13350,N_13431);
and U13539 (N_13539,N_13332,N_13394);
nand U13540 (N_13540,N_13372,N_13282);
and U13541 (N_13541,N_13395,N_13352);
and U13542 (N_13542,N_13286,N_13337);
nand U13543 (N_13543,N_13322,N_13343);
nand U13544 (N_13544,N_13419,N_13404);
or U13545 (N_13545,N_13308,N_13303);
nor U13546 (N_13546,N_13383,N_13282);
nand U13547 (N_13547,N_13293,N_13364);
nor U13548 (N_13548,N_13280,N_13307);
and U13549 (N_13549,N_13291,N_13342);
nor U13550 (N_13550,N_13417,N_13320);
nor U13551 (N_13551,N_13348,N_13424);
nor U13552 (N_13552,N_13349,N_13429);
or U13553 (N_13553,N_13295,N_13353);
nor U13554 (N_13554,N_13380,N_13436);
xor U13555 (N_13555,N_13294,N_13379);
and U13556 (N_13556,N_13415,N_13406);
or U13557 (N_13557,N_13349,N_13355);
or U13558 (N_13558,N_13319,N_13305);
xnor U13559 (N_13559,N_13353,N_13349);
and U13560 (N_13560,N_13332,N_13309);
nor U13561 (N_13561,N_13282,N_13360);
and U13562 (N_13562,N_13293,N_13438);
xor U13563 (N_13563,N_13317,N_13346);
nand U13564 (N_13564,N_13363,N_13396);
and U13565 (N_13565,N_13387,N_13363);
and U13566 (N_13566,N_13333,N_13358);
nand U13567 (N_13567,N_13383,N_13425);
nand U13568 (N_13568,N_13373,N_13294);
xnor U13569 (N_13569,N_13363,N_13349);
nor U13570 (N_13570,N_13422,N_13315);
or U13571 (N_13571,N_13435,N_13312);
nand U13572 (N_13572,N_13430,N_13307);
or U13573 (N_13573,N_13434,N_13310);
xor U13574 (N_13574,N_13429,N_13379);
and U13575 (N_13575,N_13411,N_13408);
nor U13576 (N_13576,N_13400,N_13369);
xnor U13577 (N_13577,N_13429,N_13336);
xor U13578 (N_13578,N_13378,N_13371);
or U13579 (N_13579,N_13280,N_13319);
nor U13580 (N_13580,N_13436,N_13377);
and U13581 (N_13581,N_13363,N_13282);
or U13582 (N_13582,N_13415,N_13365);
nand U13583 (N_13583,N_13415,N_13323);
or U13584 (N_13584,N_13329,N_13412);
and U13585 (N_13585,N_13280,N_13369);
or U13586 (N_13586,N_13402,N_13407);
and U13587 (N_13587,N_13307,N_13410);
and U13588 (N_13588,N_13281,N_13386);
nor U13589 (N_13589,N_13314,N_13383);
or U13590 (N_13590,N_13326,N_13299);
and U13591 (N_13591,N_13413,N_13390);
or U13592 (N_13592,N_13404,N_13381);
nand U13593 (N_13593,N_13399,N_13323);
xnor U13594 (N_13594,N_13411,N_13401);
and U13595 (N_13595,N_13325,N_13424);
and U13596 (N_13596,N_13326,N_13351);
xnor U13597 (N_13597,N_13437,N_13433);
or U13598 (N_13598,N_13318,N_13356);
nand U13599 (N_13599,N_13313,N_13395);
nor U13600 (N_13600,N_13509,N_13484);
nor U13601 (N_13601,N_13536,N_13599);
nand U13602 (N_13602,N_13452,N_13445);
and U13603 (N_13603,N_13505,N_13517);
nor U13604 (N_13604,N_13469,N_13463);
or U13605 (N_13605,N_13557,N_13454);
nor U13606 (N_13606,N_13561,N_13527);
or U13607 (N_13607,N_13443,N_13476);
or U13608 (N_13608,N_13472,N_13524);
or U13609 (N_13609,N_13512,N_13528);
or U13610 (N_13610,N_13507,N_13532);
nor U13611 (N_13611,N_13578,N_13508);
and U13612 (N_13612,N_13568,N_13579);
nand U13613 (N_13613,N_13464,N_13598);
nor U13614 (N_13614,N_13471,N_13529);
and U13615 (N_13615,N_13550,N_13547);
or U13616 (N_13616,N_13496,N_13582);
nand U13617 (N_13617,N_13516,N_13467);
nor U13618 (N_13618,N_13573,N_13447);
or U13619 (N_13619,N_13566,N_13590);
or U13620 (N_13620,N_13560,N_13595);
nor U13621 (N_13621,N_13450,N_13585);
nor U13622 (N_13622,N_13518,N_13474);
or U13623 (N_13623,N_13548,N_13537);
nand U13624 (N_13624,N_13570,N_13580);
or U13625 (N_13625,N_13549,N_13481);
nand U13626 (N_13626,N_13554,N_13564);
nor U13627 (N_13627,N_13441,N_13543);
and U13628 (N_13628,N_13501,N_13456);
or U13629 (N_13629,N_13540,N_13470);
or U13630 (N_13630,N_13577,N_13588);
xnor U13631 (N_13631,N_13519,N_13572);
xor U13632 (N_13632,N_13515,N_13446);
and U13633 (N_13633,N_13499,N_13592);
and U13634 (N_13634,N_13493,N_13525);
xnor U13635 (N_13635,N_13576,N_13571);
nand U13636 (N_13636,N_13535,N_13460);
xor U13637 (N_13637,N_13495,N_13565);
xnor U13638 (N_13638,N_13486,N_13526);
xor U13639 (N_13639,N_13596,N_13475);
or U13640 (N_13640,N_13523,N_13492);
xor U13641 (N_13641,N_13468,N_13538);
xnor U13642 (N_13642,N_13531,N_13551);
and U13643 (N_13643,N_13544,N_13491);
nand U13644 (N_13644,N_13442,N_13506);
and U13645 (N_13645,N_13479,N_13466);
and U13646 (N_13646,N_13457,N_13589);
xor U13647 (N_13647,N_13489,N_13478);
nor U13648 (N_13648,N_13597,N_13511);
or U13649 (N_13649,N_13533,N_13584);
or U13650 (N_13650,N_13465,N_13574);
nor U13651 (N_13651,N_13510,N_13562);
nand U13652 (N_13652,N_13594,N_13483);
xnor U13653 (N_13653,N_13448,N_13502);
and U13654 (N_13654,N_13453,N_13497);
nand U13655 (N_13655,N_13461,N_13513);
xnor U13656 (N_13656,N_13586,N_13451);
or U13657 (N_13657,N_13559,N_13514);
nor U13658 (N_13658,N_13556,N_13520);
nand U13659 (N_13659,N_13563,N_13462);
nand U13660 (N_13660,N_13440,N_13449);
nand U13661 (N_13661,N_13487,N_13552);
and U13662 (N_13662,N_13444,N_13553);
nor U13663 (N_13663,N_13593,N_13555);
nor U13664 (N_13664,N_13488,N_13459);
or U13665 (N_13665,N_13587,N_13482);
nand U13666 (N_13666,N_13473,N_13583);
and U13667 (N_13667,N_13541,N_13500);
xor U13668 (N_13668,N_13545,N_13558);
nand U13669 (N_13669,N_13485,N_13534);
nor U13670 (N_13670,N_13521,N_13458);
nand U13671 (N_13671,N_13477,N_13530);
xor U13672 (N_13672,N_13542,N_13480);
nand U13673 (N_13673,N_13539,N_13504);
or U13674 (N_13674,N_13569,N_13567);
nor U13675 (N_13675,N_13591,N_13503);
or U13676 (N_13676,N_13498,N_13546);
nand U13677 (N_13677,N_13455,N_13490);
and U13678 (N_13678,N_13581,N_13522);
nand U13679 (N_13679,N_13575,N_13494);
nand U13680 (N_13680,N_13534,N_13472);
xnor U13681 (N_13681,N_13512,N_13572);
nor U13682 (N_13682,N_13598,N_13593);
nor U13683 (N_13683,N_13542,N_13527);
or U13684 (N_13684,N_13481,N_13506);
nor U13685 (N_13685,N_13523,N_13590);
and U13686 (N_13686,N_13507,N_13562);
and U13687 (N_13687,N_13539,N_13533);
and U13688 (N_13688,N_13442,N_13556);
and U13689 (N_13689,N_13504,N_13488);
nor U13690 (N_13690,N_13483,N_13516);
xnor U13691 (N_13691,N_13494,N_13568);
nor U13692 (N_13692,N_13441,N_13453);
xor U13693 (N_13693,N_13502,N_13503);
nand U13694 (N_13694,N_13566,N_13443);
or U13695 (N_13695,N_13593,N_13572);
xnor U13696 (N_13696,N_13583,N_13459);
or U13697 (N_13697,N_13566,N_13479);
xor U13698 (N_13698,N_13529,N_13592);
xor U13699 (N_13699,N_13582,N_13485);
and U13700 (N_13700,N_13504,N_13531);
nand U13701 (N_13701,N_13568,N_13463);
nor U13702 (N_13702,N_13470,N_13453);
xor U13703 (N_13703,N_13573,N_13558);
nand U13704 (N_13704,N_13481,N_13504);
nor U13705 (N_13705,N_13456,N_13443);
xor U13706 (N_13706,N_13454,N_13545);
xor U13707 (N_13707,N_13566,N_13555);
or U13708 (N_13708,N_13447,N_13575);
nand U13709 (N_13709,N_13523,N_13583);
or U13710 (N_13710,N_13462,N_13522);
and U13711 (N_13711,N_13485,N_13553);
xor U13712 (N_13712,N_13539,N_13482);
or U13713 (N_13713,N_13497,N_13451);
nor U13714 (N_13714,N_13464,N_13475);
and U13715 (N_13715,N_13448,N_13518);
and U13716 (N_13716,N_13555,N_13469);
or U13717 (N_13717,N_13474,N_13471);
nor U13718 (N_13718,N_13516,N_13590);
nand U13719 (N_13719,N_13447,N_13568);
nor U13720 (N_13720,N_13541,N_13486);
and U13721 (N_13721,N_13490,N_13574);
xor U13722 (N_13722,N_13530,N_13459);
xnor U13723 (N_13723,N_13578,N_13456);
or U13724 (N_13724,N_13567,N_13577);
or U13725 (N_13725,N_13553,N_13519);
nand U13726 (N_13726,N_13589,N_13585);
nand U13727 (N_13727,N_13488,N_13496);
nor U13728 (N_13728,N_13479,N_13453);
nor U13729 (N_13729,N_13531,N_13492);
and U13730 (N_13730,N_13442,N_13542);
nor U13731 (N_13731,N_13555,N_13565);
nor U13732 (N_13732,N_13490,N_13580);
or U13733 (N_13733,N_13548,N_13474);
or U13734 (N_13734,N_13510,N_13462);
or U13735 (N_13735,N_13598,N_13508);
nor U13736 (N_13736,N_13524,N_13473);
and U13737 (N_13737,N_13464,N_13528);
nor U13738 (N_13738,N_13524,N_13453);
nor U13739 (N_13739,N_13441,N_13536);
and U13740 (N_13740,N_13583,N_13470);
nor U13741 (N_13741,N_13501,N_13509);
or U13742 (N_13742,N_13471,N_13588);
nand U13743 (N_13743,N_13445,N_13581);
or U13744 (N_13744,N_13587,N_13480);
nor U13745 (N_13745,N_13504,N_13533);
and U13746 (N_13746,N_13551,N_13535);
nor U13747 (N_13747,N_13552,N_13513);
xor U13748 (N_13748,N_13583,N_13540);
xor U13749 (N_13749,N_13478,N_13545);
xnor U13750 (N_13750,N_13460,N_13506);
xnor U13751 (N_13751,N_13554,N_13544);
or U13752 (N_13752,N_13489,N_13515);
nor U13753 (N_13753,N_13537,N_13472);
nor U13754 (N_13754,N_13442,N_13470);
or U13755 (N_13755,N_13550,N_13526);
xnor U13756 (N_13756,N_13463,N_13577);
xnor U13757 (N_13757,N_13471,N_13509);
nand U13758 (N_13758,N_13503,N_13506);
nor U13759 (N_13759,N_13507,N_13460);
or U13760 (N_13760,N_13631,N_13713);
nor U13761 (N_13761,N_13751,N_13673);
and U13762 (N_13762,N_13648,N_13750);
or U13763 (N_13763,N_13661,N_13682);
or U13764 (N_13764,N_13743,N_13641);
and U13765 (N_13765,N_13611,N_13703);
nand U13766 (N_13766,N_13671,N_13714);
xor U13767 (N_13767,N_13635,N_13685);
and U13768 (N_13768,N_13670,N_13659);
and U13769 (N_13769,N_13606,N_13607);
and U13770 (N_13770,N_13731,N_13689);
nor U13771 (N_13771,N_13701,N_13727);
and U13772 (N_13772,N_13640,N_13675);
nor U13773 (N_13773,N_13752,N_13663);
or U13774 (N_13774,N_13711,N_13694);
or U13775 (N_13775,N_13696,N_13706);
or U13776 (N_13776,N_13748,N_13683);
xnor U13777 (N_13777,N_13744,N_13721);
nand U13778 (N_13778,N_13742,N_13600);
xor U13779 (N_13779,N_13643,N_13680);
nor U13780 (N_13780,N_13738,N_13686);
xnor U13781 (N_13781,N_13616,N_13617);
nand U13782 (N_13782,N_13665,N_13737);
nand U13783 (N_13783,N_13627,N_13649);
xor U13784 (N_13784,N_13759,N_13695);
nand U13785 (N_13785,N_13603,N_13735);
and U13786 (N_13786,N_13740,N_13757);
nor U13787 (N_13787,N_13693,N_13669);
nor U13788 (N_13788,N_13656,N_13630);
nor U13789 (N_13789,N_13609,N_13700);
nand U13790 (N_13790,N_13653,N_13712);
and U13791 (N_13791,N_13645,N_13647);
nand U13792 (N_13792,N_13687,N_13749);
nor U13793 (N_13793,N_13602,N_13612);
nand U13794 (N_13794,N_13732,N_13632);
nor U13795 (N_13795,N_13739,N_13716);
nand U13796 (N_13796,N_13610,N_13741);
xnor U13797 (N_13797,N_13668,N_13676);
xnor U13798 (N_13798,N_13646,N_13681);
xor U13799 (N_13799,N_13664,N_13718);
nor U13800 (N_13800,N_13708,N_13726);
nand U13801 (N_13801,N_13746,N_13704);
xor U13802 (N_13802,N_13722,N_13754);
and U13803 (N_13803,N_13725,N_13644);
or U13804 (N_13804,N_13658,N_13639);
or U13805 (N_13805,N_13719,N_13699);
and U13806 (N_13806,N_13715,N_13628);
nor U13807 (N_13807,N_13672,N_13690);
nor U13808 (N_13808,N_13626,N_13604);
and U13809 (N_13809,N_13698,N_13650);
nor U13810 (N_13810,N_13705,N_13657);
xor U13811 (N_13811,N_13623,N_13614);
xor U13812 (N_13812,N_13755,N_13636);
nand U13813 (N_13813,N_13660,N_13723);
or U13814 (N_13814,N_13625,N_13720);
or U13815 (N_13815,N_13654,N_13709);
and U13816 (N_13816,N_13674,N_13613);
nor U13817 (N_13817,N_13666,N_13634);
xor U13818 (N_13818,N_13638,N_13692);
nand U13819 (N_13819,N_13707,N_13618);
and U13820 (N_13820,N_13667,N_13608);
xor U13821 (N_13821,N_13745,N_13697);
nand U13822 (N_13822,N_13605,N_13601);
and U13823 (N_13823,N_13729,N_13651);
nor U13824 (N_13824,N_13688,N_13734);
or U13825 (N_13825,N_13622,N_13637);
and U13826 (N_13826,N_13629,N_13678);
nor U13827 (N_13827,N_13710,N_13702);
and U13828 (N_13828,N_13652,N_13619);
or U13829 (N_13829,N_13756,N_13633);
or U13830 (N_13830,N_13655,N_13621);
nor U13831 (N_13831,N_13758,N_13724);
xnor U13832 (N_13832,N_13662,N_13728);
nor U13833 (N_13833,N_13691,N_13642);
xnor U13834 (N_13834,N_13615,N_13747);
and U13835 (N_13835,N_13684,N_13624);
nor U13836 (N_13836,N_13717,N_13620);
nand U13837 (N_13837,N_13753,N_13733);
nor U13838 (N_13838,N_13730,N_13677);
nor U13839 (N_13839,N_13679,N_13736);
and U13840 (N_13840,N_13719,N_13715);
nand U13841 (N_13841,N_13616,N_13704);
and U13842 (N_13842,N_13709,N_13637);
nand U13843 (N_13843,N_13716,N_13682);
xor U13844 (N_13844,N_13665,N_13603);
nand U13845 (N_13845,N_13660,N_13693);
xnor U13846 (N_13846,N_13616,N_13751);
and U13847 (N_13847,N_13706,N_13739);
nor U13848 (N_13848,N_13692,N_13722);
nand U13849 (N_13849,N_13658,N_13741);
and U13850 (N_13850,N_13643,N_13714);
or U13851 (N_13851,N_13754,N_13608);
nor U13852 (N_13852,N_13609,N_13717);
and U13853 (N_13853,N_13750,N_13669);
and U13854 (N_13854,N_13684,N_13610);
and U13855 (N_13855,N_13681,N_13625);
nand U13856 (N_13856,N_13709,N_13741);
and U13857 (N_13857,N_13627,N_13705);
nand U13858 (N_13858,N_13742,N_13662);
and U13859 (N_13859,N_13715,N_13729);
xnor U13860 (N_13860,N_13684,N_13628);
nand U13861 (N_13861,N_13642,N_13746);
xnor U13862 (N_13862,N_13746,N_13662);
xor U13863 (N_13863,N_13740,N_13713);
and U13864 (N_13864,N_13620,N_13721);
and U13865 (N_13865,N_13691,N_13686);
or U13866 (N_13866,N_13670,N_13600);
nor U13867 (N_13867,N_13644,N_13687);
and U13868 (N_13868,N_13698,N_13629);
or U13869 (N_13869,N_13685,N_13723);
xor U13870 (N_13870,N_13622,N_13740);
nand U13871 (N_13871,N_13735,N_13692);
nand U13872 (N_13872,N_13759,N_13735);
nor U13873 (N_13873,N_13657,N_13608);
and U13874 (N_13874,N_13735,N_13652);
or U13875 (N_13875,N_13715,N_13759);
xnor U13876 (N_13876,N_13687,N_13632);
or U13877 (N_13877,N_13609,N_13649);
or U13878 (N_13878,N_13611,N_13623);
nand U13879 (N_13879,N_13648,N_13701);
and U13880 (N_13880,N_13680,N_13621);
nand U13881 (N_13881,N_13737,N_13609);
or U13882 (N_13882,N_13612,N_13748);
xnor U13883 (N_13883,N_13737,N_13743);
xor U13884 (N_13884,N_13650,N_13682);
or U13885 (N_13885,N_13748,N_13709);
nand U13886 (N_13886,N_13667,N_13676);
and U13887 (N_13887,N_13605,N_13680);
nor U13888 (N_13888,N_13691,N_13613);
xnor U13889 (N_13889,N_13600,N_13692);
nor U13890 (N_13890,N_13622,N_13746);
nor U13891 (N_13891,N_13743,N_13677);
xnor U13892 (N_13892,N_13673,N_13602);
nand U13893 (N_13893,N_13691,N_13629);
xnor U13894 (N_13894,N_13637,N_13743);
xor U13895 (N_13895,N_13619,N_13739);
nand U13896 (N_13896,N_13670,N_13732);
xor U13897 (N_13897,N_13717,N_13656);
xor U13898 (N_13898,N_13689,N_13628);
or U13899 (N_13899,N_13653,N_13755);
nor U13900 (N_13900,N_13755,N_13702);
nor U13901 (N_13901,N_13709,N_13613);
nor U13902 (N_13902,N_13714,N_13606);
xnor U13903 (N_13903,N_13633,N_13702);
nor U13904 (N_13904,N_13759,N_13679);
nand U13905 (N_13905,N_13639,N_13740);
or U13906 (N_13906,N_13645,N_13701);
nand U13907 (N_13907,N_13723,N_13724);
and U13908 (N_13908,N_13609,N_13675);
nor U13909 (N_13909,N_13670,N_13668);
xnor U13910 (N_13910,N_13664,N_13693);
xor U13911 (N_13911,N_13731,N_13658);
nor U13912 (N_13912,N_13639,N_13711);
and U13913 (N_13913,N_13722,N_13613);
nor U13914 (N_13914,N_13669,N_13717);
nand U13915 (N_13915,N_13740,N_13666);
nand U13916 (N_13916,N_13643,N_13755);
nand U13917 (N_13917,N_13643,N_13692);
and U13918 (N_13918,N_13630,N_13625);
and U13919 (N_13919,N_13644,N_13667);
nor U13920 (N_13920,N_13832,N_13813);
or U13921 (N_13921,N_13844,N_13766);
and U13922 (N_13922,N_13816,N_13880);
xnor U13923 (N_13923,N_13918,N_13871);
nand U13924 (N_13924,N_13897,N_13812);
nand U13925 (N_13925,N_13796,N_13849);
or U13926 (N_13926,N_13857,N_13896);
and U13927 (N_13927,N_13868,N_13835);
xor U13928 (N_13928,N_13775,N_13895);
nand U13929 (N_13929,N_13799,N_13807);
nor U13930 (N_13930,N_13908,N_13772);
or U13931 (N_13931,N_13904,N_13768);
nor U13932 (N_13932,N_13767,N_13782);
and U13933 (N_13933,N_13874,N_13803);
and U13934 (N_13934,N_13792,N_13777);
nor U13935 (N_13935,N_13906,N_13811);
or U13936 (N_13936,N_13876,N_13909);
nor U13937 (N_13937,N_13824,N_13826);
and U13938 (N_13938,N_13900,N_13855);
and U13939 (N_13939,N_13847,N_13825);
or U13940 (N_13940,N_13852,N_13914);
nor U13941 (N_13941,N_13860,N_13804);
and U13942 (N_13942,N_13787,N_13911);
nor U13943 (N_13943,N_13762,N_13886);
and U13944 (N_13944,N_13821,N_13850);
nand U13945 (N_13945,N_13838,N_13862);
nor U13946 (N_13946,N_13873,N_13810);
xor U13947 (N_13947,N_13848,N_13823);
xnor U13948 (N_13948,N_13890,N_13892);
nand U13949 (N_13949,N_13845,N_13903);
nor U13950 (N_13950,N_13919,N_13814);
nand U13951 (N_13951,N_13834,N_13801);
or U13952 (N_13952,N_13789,N_13798);
or U13953 (N_13953,N_13770,N_13776);
xnor U13954 (N_13954,N_13875,N_13843);
or U13955 (N_13955,N_13894,N_13902);
xnor U13956 (N_13956,N_13869,N_13800);
xnor U13957 (N_13957,N_13831,N_13783);
nand U13958 (N_13958,N_13881,N_13888);
nand U13959 (N_13959,N_13889,N_13828);
xor U13960 (N_13960,N_13917,N_13794);
xnor U13961 (N_13961,N_13865,N_13829);
and U13962 (N_13962,N_13859,N_13887);
xnor U13963 (N_13963,N_13915,N_13820);
and U13964 (N_13964,N_13830,N_13879);
xor U13965 (N_13965,N_13806,N_13842);
xnor U13966 (N_13966,N_13819,N_13785);
and U13967 (N_13967,N_13905,N_13893);
xor U13968 (N_13968,N_13822,N_13872);
xnor U13969 (N_13969,N_13765,N_13907);
nor U13970 (N_13970,N_13779,N_13884);
nand U13971 (N_13971,N_13809,N_13856);
nor U13972 (N_13972,N_13778,N_13836);
nor U13973 (N_13973,N_13861,N_13771);
or U13974 (N_13974,N_13795,N_13781);
nor U13975 (N_13975,N_13817,N_13764);
nand U13976 (N_13976,N_13870,N_13790);
and U13977 (N_13977,N_13833,N_13910);
nand U13978 (N_13978,N_13839,N_13898);
or U13979 (N_13979,N_13916,N_13793);
nor U13980 (N_13980,N_13840,N_13786);
or U13981 (N_13981,N_13773,N_13841);
xor U13982 (N_13982,N_13858,N_13818);
nor U13983 (N_13983,N_13837,N_13864);
and U13984 (N_13984,N_13878,N_13815);
nand U13985 (N_13985,N_13853,N_13867);
nor U13986 (N_13986,N_13797,N_13882);
and U13987 (N_13987,N_13885,N_13846);
and U13988 (N_13988,N_13769,N_13899);
nand U13989 (N_13989,N_13913,N_13827);
nand U13990 (N_13990,N_13791,N_13891);
nor U13991 (N_13991,N_13761,N_13760);
or U13992 (N_13992,N_13780,N_13866);
nor U13993 (N_13993,N_13863,N_13851);
nand U13994 (N_13994,N_13901,N_13854);
xor U13995 (N_13995,N_13763,N_13883);
nor U13996 (N_13996,N_13784,N_13808);
and U13997 (N_13997,N_13802,N_13788);
or U13998 (N_13998,N_13805,N_13912);
and U13999 (N_13999,N_13877,N_13774);
and U14000 (N_14000,N_13793,N_13840);
and U14001 (N_14001,N_13885,N_13881);
nand U14002 (N_14002,N_13829,N_13784);
and U14003 (N_14003,N_13835,N_13882);
nand U14004 (N_14004,N_13903,N_13766);
nand U14005 (N_14005,N_13808,N_13838);
or U14006 (N_14006,N_13803,N_13767);
nand U14007 (N_14007,N_13788,N_13883);
nand U14008 (N_14008,N_13797,N_13842);
nand U14009 (N_14009,N_13793,N_13826);
nor U14010 (N_14010,N_13829,N_13884);
or U14011 (N_14011,N_13900,N_13895);
nor U14012 (N_14012,N_13905,N_13837);
or U14013 (N_14013,N_13916,N_13898);
nand U14014 (N_14014,N_13869,N_13857);
or U14015 (N_14015,N_13826,N_13855);
or U14016 (N_14016,N_13830,N_13824);
nand U14017 (N_14017,N_13785,N_13880);
and U14018 (N_14018,N_13854,N_13887);
and U14019 (N_14019,N_13914,N_13862);
nand U14020 (N_14020,N_13803,N_13898);
or U14021 (N_14021,N_13850,N_13849);
nand U14022 (N_14022,N_13841,N_13911);
nor U14023 (N_14023,N_13834,N_13862);
or U14024 (N_14024,N_13895,N_13831);
and U14025 (N_14025,N_13806,N_13876);
or U14026 (N_14026,N_13899,N_13900);
nor U14027 (N_14027,N_13795,N_13801);
nand U14028 (N_14028,N_13822,N_13912);
xnor U14029 (N_14029,N_13765,N_13852);
nor U14030 (N_14030,N_13760,N_13857);
or U14031 (N_14031,N_13841,N_13788);
xnor U14032 (N_14032,N_13874,N_13768);
nand U14033 (N_14033,N_13768,N_13833);
nor U14034 (N_14034,N_13881,N_13901);
nor U14035 (N_14035,N_13848,N_13912);
or U14036 (N_14036,N_13915,N_13877);
xor U14037 (N_14037,N_13837,N_13821);
nor U14038 (N_14038,N_13778,N_13784);
nand U14039 (N_14039,N_13765,N_13891);
nor U14040 (N_14040,N_13855,N_13806);
nor U14041 (N_14041,N_13913,N_13917);
xor U14042 (N_14042,N_13782,N_13818);
nand U14043 (N_14043,N_13857,N_13853);
and U14044 (N_14044,N_13887,N_13760);
xnor U14045 (N_14045,N_13887,N_13844);
xnor U14046 (N_14046,N_13794,N_13839);
nand U14047 (N_14047,N_13839,N_13854);
nor U14048 (N_14048,N_13889,N_13914);
and U14049 (N_14049,N_13766,N_13819);
and U14050 (N_14050,N_13895,N_13870);
nor U14051 (N_14051,N_13849,N_13889);
or U14052 (N_14052,N_13881,N_13835);
xnor U14053 (N_14053,N_13785,N_13837);
and U14054 (N_14054,N_13813,N_13907);
nand U14055 (N_14055,N_13776,N_13912);
nand U14056 (N_14056,N_13850,N_13799);
nor U14057 (N_14057,N_13867,N_13807);
nor U14058 (N_14058,N_13888,N_13804);
xnor U14059 (N_14059,N_13851,N_13834);
and U14060 (N_14060,N_13837,N_13826);
or U14061 (N_14061,N_13848,N_13800);
and U14062 (N_14062,N_13785,N_13822);
xnor U14063 (N_14063,N_13879,N_13848);
xnor U14064 (N_14064,N_13762,N_13854);
and U14065 (N_14065,N_13780,N_13864);
xnor U14066 (N_14066,N_13782,N_13881);
nand U14067 (N_14067,N_13766,N_13874);
or U14068 (N_14068,N_13898,N_13874);
xnor U14069 (N_14069,N_13807,N_13837);
nand U14070 (N_14070,N_13893,N_13788);
xor U14071 (N_14071,N_13762,N_13814);
xnor U14072 (N_14072,N_13882,N_13917);
nand U14073 (N_14073,N_13792,N_13849);
xor U14074 (N_14074,N_13879,N_13865);
nand U14075 (N_14075,N_13890,N_13834);
or U14076 (N_14076,N_13780,N_13872);
and U14077 (N_14077,N_13899,N_13885);
xor U14078 (N_14078,N_13787,N_13838);
and U14079 (N_14079,N_13850,N_13828);
or U14080 (N_14080,N_14003,N_13942);
xor U14081 (N_14081,N_14031,N_14056);
and U14082 (N_14082,N_14064,N_13939);
xor U14083 (N_14083,N_13936,N_13986);
xnor U14084 (N_14084,N_13991,N_14041);
or U14085 (N_14085,N_14062,N_13985);
xor U14086 (N_14086,N_13979,N_14009);
or U14087 (N_14087,N_14004,N_13965);
nor U14088 (N_14088,N_13967,N_13990);
or U14089 (N_14089,N_14047,N_14068);
nand U14090 (N_14090,N_14018,N_14079);
or U14091 (N_14091,N_13953,N_13929);
nand U14092 (N_14092,N_14051,N_13964);
and U14093 (N_14093,N_14033,N_13970);
nand U14094 (N_14094,N_14048,N_13937);
nand U14095 (N_14095,N_13971,N_13928);
nor U14096 (N_14096,N_14052,N_13963);
and U14097 (N_14097,N_13994,N_13961);
and U14098 (N_14098,N_14019,N_13968);
nand U14099 (N_14099,N_14058,N_14021);
xnor U14100 (N_14100,N_14049,N_13972);
xnor U14101 (N_14101,N_14029,N_13959);
nand U14102 (N_14102,N_14013,N_14043);
nor U14103 (N_14103,N_13940,N_14026);
nand U14104 (N_14104,N_13999,N_13945);
and U14105 (N_14105,N_14008,N_13938);
nor U14106 (N_14106,N_13949,N_13933);
or U14107 (N_14107,N_13998,N_13930);
or U14108 (N_14108,N_14061,N_14017);
or U14109 (N_14109,N_13973,N_14046);
xor U14110 (N_14110,N_14059,N_13952);
nor U14111 (N_14111,N_13993,N_13982);
or U14112 (N_14112,N_13974,N_14039);
nand U14113 (N_14113,N_13955,N_14044);
nand U14114 (N_14114,N_14032,N_14075);
and U14115 (N_14115,N_14054,N_13954);
and U14116 (N_14116,N_13922,N_14050);
nand U14117 (N_14117,N_13957,N_13977);
nand U14118 (N_14118,N_13981,N_13931);
or U14119 (N_14119,N_14028,N_14067);
or U14120 (N_14120,N_13924,N_14060);
nor U14121 (N_14121,N_14035,N_14077);
or U14122 (N_14122,N_13947,N_13978);
xor U14123 (N_14123,N_13926,N_14007);
and U14124 (N_14124,N_13960,N_14078);
or U14125 (N_14125,N_14027,N_14037);
xor U14126 (N_14126,N_14066,N_13980);
or U14127 (N_14127,N_13997,N_13925);
nor U14128 (N_14128,N_13966,N_14016);
and U14129 (N_14129,N_14057,N_14074);
xnor U14130 (N_14130,N_14015,N_14076);
nor U14131 (N_14131,N_13975,N_14070);
nor U14132 (N_14132,N_14053,N_14023);
xnor U14133 (N_14133,N_14014,N_14071);
or U14134 (N_14134,N_14030,N_14012);
and U14135 (N_14135,N_14010,N_14073);
nand U14136 (N_14136,N_14005,N_13941);
and U14137 (N_14137,N_13921,N_14069);
nor U14138 (N_14138,N_14011,N_14006);
and U14139 (N_14139,N_13987,N_13976);
xnor U14140 (N_14140,N_14042,N_14045);
nor U14141 (N_14141,N_14022,N_13969);
xnor U14142 (N_14142,N_13950,N_13956);
and U14143 (N_14143,N_13989,N_13951);
nand U14144 (N_14144,N_13958,N_13943);
or U14145 (N_14145,N_14002,N_14024);
or U14146 (N_14146,N_13962,N_13995);
or U14147 (N_14147,N_13934,N_13935);
nand U14148 (N_14148,N_14025,N_14036);
and U14149 (N_14149,N_13923,N_13932);
xor U14150 (N_14150,N_13946,N_13984);
nand U14151 (N_14151,N_14038,N_13983);
nor U14152 (N_14152,N_14034,N_13996);
nor U14153 (N_14153,N_14001,N_14055);
nor U14154 (N_14154,N_14020,N_13948);
and U14155 (N_14155,N_14063,N_14065);
or U14156 (N_14156,N_13992,N_13920);
and U14157 (N_14157,N_14040,N_13944);
nor U14158 (N_14158,N_13927,N_14072);
or U14159 (N_14159,N_14000,N_13988);
or U14160 (N_14160,N_14049,N_14050);
or U14161 (N_14161,N_14077,N_14054);
nand U14162 (N_14162,N_14043,N_13985);
nor U14163 (N_14163,N_14034,N_13938);
nand U14164 (N_14164,N_13941,N_13946);
nor U14165 (N_14165,N_14012,N_13953);
or U14166 (N_14166,N_14010,N_14037);
nor U14167 (N_14167,N_13973,N_14075);
nand U14168 (N_14168,N_14066,N_14041);
nor U14169 (N_14169,N_14042,N_13997);
xnor U14170 (N_14170,N_13998,N_13988);
nor U14171 (N_14171,N_14028,N_13983);
nor U14172 (N_14172,N_14061,N_13986);
nor U14173 (N_14173,N_13937,N_13960);
nor U14174 (N_14174,N_14012,N_13996);
or U14175 (N_14175,N_14077,N_13988);
or U14176 (N_14176,N_14053,N_14063);
nand U14177 (N_14177,N_14071,N_13980);
xnor U14178 (N_14178,N_14033,N_14012);
or U14179 (N_14179,N_13955,N_13976);
and U14180 (N_14180,N_14063,N_14028);
nor U14181 (N_14181,N_13956,N_13957);
and U14182 (N_14182,N_14049,N_14074);
nor U14183 (N_14183,N_14031,N_14023);
and U14184 (N_14184,N_14074,N_14037);
and U14185 (N_14185,N_14004,N_14062);
and U14186 (N_14186,N_13933,N_14011);
or U14187 (N_14187,N_14036,N_14026);
and U14188 (N_14188,N_14012,N_13976);
or U14189 (N_14189,N_14015,N_13940);
and U14190 (N_14190,N_14026,N_14050);
xnor U14191 (N_14191,N_14024,N_14035);
or U14192 (N_14192,N_13924,N_13970);
nand U14193 (N_14193,N_13938,N_13965);
xnor U14194 (N_14194,N_14047,N_13956);
and U14195 (N_14195,N_14012,N_14040);
and U14196 (N_14196,N_13995,N_14075);
nand U14197 (N_14197,N_13925,N_14012);
nand U14198 (N_14198,N_13973,N_14054);
or U14199 (N_14199,N_14022,N_13954);
and U14200 (N_14200,N_13968,N_14006);
or U14201 (N_14201,N_14066,N_13922);
xnor U14202 (N_14202,N_13933,N_14042);
or U14203 (N_14203,N_14058,N_13972);
and U14204 (N_14204,N_14042,N_13996);
or U14205 (N_14205,N_13947,N_14017);
or U14206 (N_14206,N_14034,N_14040);
or U14207 (N_14207,N_14077,N_13938);
nor U14208 (N_14208,N_14016,N_13975);
and U14209 (N_14209,N_13932,N_14009);
nor U14210 (N_14210,N_13980,N_13997);
and U14211 (N_14211,N_14022,N_14004);
or U14212 (N_14212,N_13999,N_14040);
nand U14213 (N_14213,N_14017,N_13978);
and U14214 (N_14214,N_13930,N_14006);
or U14215 (N_14215,N_14034,N_14070);
nand U14216 (N_14216,N_14071,N_13961);
and U14217 (N_14217,N_13933,N_14047);
and U14218 (N_14218,N_14056,N_13987);
nand U14219 (N_14219,N_14009,N_14077);
and U14220 (N_14220,N_13946,N_14051);
or U14221 (N_14221,N_14061,N_14068);
or U14222 (N_14222,N_13926,N_14016);
xor U14223 (N_14223,N_13948,N_14071);
nor U14224 (N_14224,N_13944,N_13994);
xnor U14225 (N_14225,N_13935,N_13930);
xnor U14226 (N_14226,N_13923,N_14046);
nand U14227 (N_14227,N_13927,N_13968);
nand U14228 (N_14228,N_14060,N_14040);
and U14229 (N_14229,N_13993,N_13920);
xnor U14230 (N_14230,N_14058,N_14075);
or U14231 (N_14231,N_14068,N_13937);
xnor U14232 (N_14232,N_14038,N_13963);
and U14233 (N_14233,N_13957,N_13963);
nor U14234 (N_14234,N_13958,N_14003);
nand U14235 (N_14235,N_13970,N_14058);
nor U14236 (N_14236,N_13924,N_14027);
xnor U14237 (N_14237,N_14066,N_13924);
nand U14238 (N_14238,N_13948,N_13961);
and U14239 (N_14239,N_14008,N_13968);
nor U14240 (N_14240,N_14161,N_14203);
or U14241 (N_14241,N_14134,N_14080);
nor U14242 (N_14242,N_14147,N_14223);
or U14243 (N_14243,N_14105,N_14138);
nand U14244 (N_14244,N_14196,N_14207);
nand U14245 (N_14245,N_14179,N_14213);
or U14246 (N_14246,N_14093,N_14173);
nor U14247 (N_14247,N_14238,N_14231);
or U14248 (N_14248,N_14234,N_14136);
xnor U14249 (N_14249,N_14108,N_14191);
and U14250 (N_14250,N_14091,N_14230);
nand U14251 (N_14251,N_14205,N_14126);
xor U14252 (N_14252,N_14183,N_14117);
or U14253 (N_14253,N_14225,N_14184);
nand U14254 (N_14254,N_14082,N_14192);
xor U14255 (N_14255,N_14085,N_14104);
nor U14256 (N_14256,N_14120,N_14190);
nand U14257 (N_14257,N_14174,N_14089);
or U14258 (N_14258,N_14124,N_14233);
and U14259 (N_14259,N_14197,N_14155);
or U14260 (N_14260,N_14135,N_14111);
nor U14261 (N_14261,N_14101,N_14185);
and U14262 (N_14262,N_14095,N_14209);
nand U14263 (N_14263,N_14220,N_14235);
xor U14264 (N_14264,N_14216,N_14211);
or U14265 (N_14265,N_14171,N_14215);
and U14266 (N_14266,N_14123,N_14169);
nor U14267 (N_14267,N_14218,N_14236);
or U14268 (N_14268,N_14226,N_14160);
xnor U14269 (N_14269,N_14081,N_14088);
nand U14270 (N_14270,N_14102,N_14114);
and U14271 (N_14271,N_14178,N_14163);
nor U14272 (N_14272,N_14150,N_14151);
xor U14273 (N_14273,N_14144,N_14159);
nor U14274 (N_14274,N_14212,N_14121);
and U14275 (N_14275,N_14129,N_14127);
xnor U14276 (N_14276,N_14164,N_14090);
and U14277 (N_14277,N_14199,N_14156);
or U14278 (N_14278,N_14176,N_14224);
and U14279 (N_14279,N_14146,N_14172);
xnor U14280 (N_14280,N_14200,N_14142);
nor U14281 (N_14281,N_14098,N_14113);
nand U14282 (N_14282,N_14137,N_14193);
nand U14283 (N_14283,N_14112,N_14219);
nand U14284 (N_14284,N_14096,N_14186);
or U14285 (N_14285,N_14100,N_14103);
or U14286 (N_14286,N_14157,N_14170);
or U14287 (N_14287,N_14115,N_14167);
and U14288 (N_14288,N_14162,N_14106);
nor U14289 (N_14289,N_14217,N_14141);
nand U14290 (N_14290,N_14118,N_14208);
or U14291 (N_14291,N_14086,N_14194);
or U14292 (N_14292,N_14154,N_14110);
or U14293 (N_14293,N_14229,N_14149);
nand U14294 (N_14294,N_14109,N_14168);
xor U14295 (N_14295,N_14092,N_14214);
nor U14296 (N_14296,N_14195,N_14228);
nand U14297 (N_14297,N_14140,N_14119);
xnor U14298 (N_14298,N_14187,N_14189);
nand U14299 (N_14299,N_14227,N_14094);
nor U14300 (N_14300,N_14130,N_14177);
xnor U14301 (N_14301,N_14182,N_14181);
and U14302 (N_14302,N_14083,N_14166);
nor U14303 (N_14303,N_14232,N_14221);
nor U14304 (N_14304,N_14133,N_14204);
xor U14305 (N_14305,N_14143,N_14122);
or U14306 (N_14306,N_14239,N_14180);
and U14307 (N_14307,N_14084,N_14165);
and U14308 (N_14308,N_14202,N_14139);
nand U14309 (N_14309,N_14222,N_14153);
or U14310 (N_14310,N_14097,N_14131);
nor U14311 (N_14311,N_14125,N_14201);
nand U14312 (N_14312,N_14132,N_14145);
and U14313 (N_14313,N_14116,N_14237);
and U14314 (N_14314,N_14188,N_14148);
and U14315 (N_14315,N_14175,N_14158);
nand U14316 (N_14316,N_14152,N_14128);
xor U14317 (N_14317,N_14210,N_14206);
nor U14318 (N_14318,N_14099,N_14087);
nor U14319 (N_14319,N_14198,N_14107);
or U14320 (N_14320,N_14201,N_14176);
xor U14321 (N_14321,N_14181,N_14104);
nand U14322 (N_14322,N_14093,N_14098);
nor U14323 (N_14323,N_14107,N_14191);
and U14324 (N_14324,N_14122,N_14199);
nor U14325 (N_14325,N_14176,N_14119);
nor U14326 (N_14326,N_14141,N_14198);
nor U14327 (N_14327,N_14195,N_14214);
nor U14328 (N_14328,N_14118,N_14102);
and U14329 (N_14329,N_14145,N_14201);
and U14330 (N_14330,N_14142,N_14192);
or U14331 (N_14331,N_14134,N_14145);
nand U14332 (N_14332,N_14128,N_14114);
or U14333 (N_14333,N_14134,N_14120);
nand U14334 (N_14334,N_14170,N_14123);
and U14335 (N_14335,N_14237,N_14190);
nand U14336 (N_14336,N_14112,N_14233);
nand U14337 (N_14337,N_14159,N_14210);
and U14338 (N_14338,N_14169,N_14215);
or U14339 (N_14339,N_14217,N_14185);
nor U14340 (N_14340,N_14230,N_14205);
or U14341 (N_14341,N_14115,N_14192);
or U14342 (N_14342,N_14196,N_14097);
xor U14343 (N_14343,N_14186,N_14137);
and U14344 (N_14344,N_14150,N_14230);
nor U14345 (N_14345,N_14186,N_14169);
nor U14346 (N_14346,N_14090,N_14176);
xor U14347 (N_14347,N_14177,N_14156);
xnor U14348 (N_14348,N_14222,N_14095);
nand U14349 (N_14349,N_14163,N_14095);
nand U14350 (N_14350,N_14212,N_14116);
or U14351 (N_14351,N_14088,N_14190);
nor U14352 (N_14352,N_14166,N_14159);
xnor U14353 (N_14353,N_14167,N_14094);
nand U14354 (N_14354,N_14163,N_14188);
nor U14355 (N_14355,N_14133,N_14212);
nand U14356 (N_14356,N_14171,N_14157);
nand U14357 (N_14357,N_14168,N_14166);
xnor U14358 (N_14358,N_14185,N_14111);
nand U14359 (N_14359,N_14167,N_14110);
and U14360 (N_14360,N_14234,N_14209);
nand U14361 (N_14361,N_14114,N_14150);
nor U14362 (N_14362,N_14214,N_14131);
and U14363 (N_14363,N_14163,N_14176);
nor U14364 (N_14364,N_14085,N_14111);
nor U14365 (N_14365,N_14156,N_14136);
xor U14366 (N_14366,N_14167,N_14208);
or U14367 (N_14367,N_14124,N_14086);
nand U14368 (N_14368,N_14097,N_14101);
or U14369 (N_14369,N_14108,N_14083);
nand U14370 (N_14370,N_14082,N_14189);
nor U14371 (N_14371,N_14239,N_14186);
xor U14372 (N_14372,N_14169,N_14192);
xor U14373 (N_14373,N_14085,N_14160);
and U14374 (N_14374,N_14085,N_14148);
or U14375 (N_14375,N_14217,N_14219);
and U14376 (N_14376,N_14130,N_14149);
or U14377 (N_14377,N_14174,N_14099);
or U14378 (N_14378,N_14100,N_14224);
and U14379 (N_14379,N_14103,N_14096);
nand U14380 (N_14380,N_14140,N_14147);
nor U14381 (N_14381,N_14141,N_14124);
or U14382 (N_14382,N_14231,N_14147);
and U14383 (N_14383,N_14130,N_14225);
and U14384 (N_14384,N_14179,N_14147);
xor U14385 (N_14385,N_14220,N_14226);
and U14386 (N_14386,N_14159,N_14167);
xor U14387 (N_14387,N_14200,N_14085);
xnor U14388 (N_14388,N_14188,N_14108);
nand U14389 (N_14389,N_14111,N_14199);
or U14390 (N_14390,N_14084,N_14080);
or U14391 (N_14391,N_14158,N_14104);
nand U14392 (N_14392,N_14096,N_14224);
xnor U14393 (N_14393,N_14184,N_14089);
and U14394 (N_14394,N_14204,N_14083);
nor U14395 (N_14395,N_14096,N_14111);
nand U14396 (N_14396,N_14093,N_14176);
xor U14397 (N_14397,N_14237,N_14137);
xnor U14398 (N_14398,N_14151,N_14125);
or U14399 (N_14399,N_14239,N_14195);
xor U14400 (N_14400,N_14360,N_14310);
nor U14401 (N_14401,N_14265,N_14293);
nand U14402 (N_14402,N_14289,N_14317);
or U14403 (N_14403,N_14267,N_14359);
nand U14404 (N_14404,N_14398,N_14271);
nor U14405 (N_14405,N_14258,N_14288);
xnor U14406 (N_14406,N_14295,N_14263);
nor U14407 (N_14407,N_14326,N_14299);
or U14408 (N_14408,N_14361,N_14277);
or U14409 (N_14409,N_14322,N_14268);
nor U14410 (N_14410,N_14335,N_14357);
or U14411 (N_14411,N_14314,N_14308);
nand U14412 (N_14412,N_14246,N_14375);
xor U14413 (N_14413,N_14391,N_14249);
and U14414 (N_14414,N_14351,N_14254);
nor U14415 (N_14415,N_14383,N_14396);
nor U14416 (N_14416,N_14393,N_14388);
or U14417 (N_14417,N_14387,N_14294);
or U14418 (N_14418,N_14259,N_14284);
and U14419 (N_14419,N_14346,N_14342);
and U14420 (N_14420,N_14307,N_14313);
nor U14421 (N_14421,N_14324,N_14376);
xnor U14422 (N_14422,N_14377,N_14287);
nand U14423 (N_14423,N_14290,N_14353);
xor U14424 (N_14424,N_14339,N_14392);
and U14425 (N_14425,N_14261,N_14372);
nand U14426 (N_14426,N_14241,N_14275);
nand U14427 (N_14427,N_14382,N_14337);
or U14428 (N_14428,N_14363,N_14251);
and U14429 (N_14429,N_14368,N_14330);
or U14430 (N_14430,N_14381,N_14384);
or U14431 (N_14431,N_14319,N_14243);
and U14432 (N_14432,N_14292,N_14305);
or U14433 (N_14433,N_14250,N_14352);
or U14434 (N_14434,N_14374,N_14399);
or U14435 (N_14435,N_14276,N_14338);
xnor U14436 (N_14436,N_14390,N_14323);
and U14437 (N_14437,N_14345,N_14266);
or U14438 (N_14438,N_14344,N_14343);
xor U14439 (N_14439,N_14298,N_14242);
nor U14440 (N_14440,N_14260,N_14311);
and U14441 (N_14441,N_14362,N_14272);
or U14442 (N_14442,N_14350,N_14328);
and U14443 (N_14443,N_14312,N_14331);
or U14444 (N_14444,N_14325,N_14301);
xnor U14445 (N_14445,N_14253,N_14296);
nand U14446 (N_14446,N_14355,N_14282);
or U14447 (N_14447,N_14378,N_14245);
nor U14448 (N_14448,N_14248,N_14385);
xnor U14449 (N_14449,N_14395,N_14332);
and U14450 (N_14450,N_14367,N_14302);
nand U14451 (N_14451,N_14257,N_14386);
or U14452 (N_14452,N_14274,N_14394);
and U14453 (N_14453,N_14291,N_14364);
nor U14454 (N_14454,N_14269,N_14279);
nor U14455 (N_14455,N_14341,N_14283);
and U14456 (N_14456,N_14329,N_14304);
and U14457 (N_14457,N_14252,N_14309);
and U14458 (N_14458,N_14278,N_14247);
nand U14459 (N_14459,N_14358,N_14370);
nor U14460 (N_14460,N_14369,N_14262);
nand U14461 (N_14461,N_14315,N_14356);
xor U14462 (N_14462,N_14244,N_14334);
nor U14463 (N_14463,N_14336,N_14316);
and U14464 (N_14464,N_14306,N_14397);
or U14465 (N_14465,N_14347,N_14389);
nor U14466 (N_14466,N_14303,N_14281);
or U14467 (N_14467,N_14327,N_14255);
xor U14468 (N_14468,N_14366,N_14373);
nand U14469 (N_14469,N_14300,N_14286);
xnor U14470 (N_14470,N_14365,N_14349);
nand U14471 (N_14471,N_14297,N_14371);
nand U14472 (N_14472,N_14256,N_14264);
xor U14473 (N_14473,N_14280,N_14348);
nand U14474 (N_14474,N_14273,N_14380);
or U14475 (N_14475,N_14321,N_14240);
or U14476 (N_14476,N_14379,N_14333);
or U14477 (N_14477,N_14285,N_14320);
xor U14478 (N_14478,N_14318,N_14340);
nand U14479 (N_14479,N_14354,N_14270);
xnor U14480 (N_14480,N_14301,N_14385);
nand U14481 (N_14481,N_14338,N_14308);
nor U14482 (N_14482,N_14368,N_14350);
nand U14483 (N_14483,N_14284,N_14311);
and U14484 (N_14484,N_14390,N_14266);
or U14485 (N_14485,N_14393,N_14392);
or U14486 (N_14486,N_14349,N_14339);
xnor U14487 (N_14487,N_14352,N_14358);
and U14488 (N_14488,N_14391,N_14278);
or U14489 (N_14489,N_14299,N_14321);
or U14490 (N_14490,N_14332,N_14379);
nand U14491 (N_14491,N_14362,N_14292);
or U14492 (N_14492,N_14349,N_14331);
xnor U14493 (N_14493,N_14281,N_14337);
or U14494 (N_14494,N_14276,N_14372);
xnor U14495 (N_14495,N_14370,N_14396);
or U14496 (N_14496,N_14330,N_14285);
nand U14497 (N_14497,N_14359,N_14255);
nand U14498 (N_14498,N_14300,N_14348);
nand U14499 (N_14499,N_14382,N_14244);
xor U14500 (N_14500,N_14262,N_14251);
and U14501 (N_14501,N_14304,N_14382);
xor U14502 (N_14502,N_14385,N_14244);
nor U14503 (N_14503,N_14246,N_14358);
nor U14504 (N_14504,N_14388,N_14312);
xor U14505 (N_14505,N_14390,N_14355);
nor U14506 (N_14506,N_14374,N_14342);
nand U14507 (N_14507,N_14250,N_14325);
or U14508 (N_14508,N_14397,N_14255);
xnor U14509 (N_14509,N_14314,N_14390);
or U14510 (N_14510,N_14385,N_14319);
nor U14511 (N_14511,N_14329,N_14340);
nor U14512 (N_14512,N_14394,N_14289);
and U14513 (N_14513,N_14272,N_14264);
xnor U14514 (N_14514,N_14300,N_14342);
and U14515 (N_14515,N_14353,N_14278);
xnor U14516 (N_14516,N_14382,N_14334);
and U14517 (N_14517,N_14392,N_14347);
or U14518 (N_14518,N_14392,N_14294);
nor U14519 (N_14519,N_14397,N_14367);
and U14520 (N_14520,N_14386,N_14272);
nand U14521 (N_14521,N_14350,N_14284);
xor U14522 (N_14522,N_14293,N_14339);
nand U14523 (N_14523,N_14344,N_14352);
and U14524 (N_14524,N_14325,N_14381);
nand U14525 (N_14525,N_14251,N_14289);
xor U14526 (N_14526,N_14342,N_14269);
xor U14527 (N_14527,N_14257,N_14351);
nand U14528 (N_14528,N_14368,N_14243);
nand U14529 (N_14529,N_14286,N_14315);
or U14530 (N_14530,N_14331,N_14385);
nand U14531 (N_14531,N_14255,N_14283);
xor U14532 (N_14532,N_14387,N_14345);
nand U14533 (N_14533,N_14324,N_14336);
and U14534 (N_14534,N_14366,N_14265);
nand U14535 (N_14535,N_14394,N_14297);
nor U14536 (N_14536,N_14365,N_14390);
xnor U14537 (N_14537,N_14242,N_14324);
nand U14538 (N_14538,N_14254,N_14390);
nand U14539 (N_14539,N_14311,N_14334);
and U14540 (N_14540,N_14358,N_14283);
xor U14541 (N_14541,N_14363,N_14366);
xor U14542 (N_14542,N_14277,N_14267);
and U14543 (N_14543,N_14324,N_14315);
nor U14544 (N_14544,N_14321,N_14341);
and U14545 (N_14545,N_14320,N_14276);
nand U14546 (N_14546,N_14291,N_14242);
xnor U14547 (N_14547,N_14385,N_14390);
xnor U14548 (N_14548,N_14321,N_14323);
nor U14549 (N_14549,N_14300,N_14390);
nor U14550 (N_14550,N_14298,N_14300);
or U14551 (N_14551,N_14398,N_14340);
xor U14552 (N_14552,N_14345,N_14359);
xor U14553 (N_14553,N_14399,N_14342);
or U14554 (N_14554,N_14367,N_14324);
nor U14555 (N_14555,N_14367,N_14370);
nor U14556 (N_14556,N_14302,N_14310);
nor U14557 (N_14557,N_14296,N_14280);
or U14558 (N_14558,N_14390,N_14324);
nand U14559 (N_14559,N_14263,N_14347);
or U14560 (N_14560,N_14513,N_14536);
nand U14561 (N_14561,N_14414,N_14527);
or U14562 (N_14562,N_14486,N_14495);
xnor U14563 (N_14563,N_14440,N_14556);
nand U14564 (N_14564,N_14433,N_14485);
and U14565 (N_14565,N_14450,N_14411);
nand U14566 (N_14566,N_14553,N_14468);
xnor U14567 (N_14567,N_14533,N_14424);
and U14568 (N_14568,N_14464,N_14451);
nand U14569 (N_14569,N_14415,N_14554);
or U14570 (N_14570,N_14490,N_14518);
or U14571 (N_14571,N_14413,N_14478);
or U14572 (N_14572,N_14500,N_14430);
nand U14573 (N_14573,N_14474,N_14448);
nand U14574 (N_14574,N_14425,N_14503);
and U14575 (N_14575,N_14452,N_14479);
nor U14576 (N_14576,N_14548,N_14416);
xnor U14577 (N_14577,N_14405,N_14489);
and U14578 (N_14578,N_14487,N_14447);
nand U14579 (N_14579,N_14537,N_14459);
and U14580 (N_14580,N_14473,N_14545);
and U14581 (N_14581,N_14484,N_14494);
nor U14582 (N_14582,N_14531,N_14491);
xnor U14583 (N_14583,N_14454,N_14516);
or U14584 (N_14584,N_14535,N_14492);
or U14585 (N_14585,N_14539,N_14442);
nor U14586 (N_14586,N_14552,N_14463);
nor U14587 (N_14587,N_14543,N_14434);
nand U14588 (N_14588,N_14488,N_14446);
or U14589 (N_14589,N_14432,N_14462);
nor U14590 (N_14590,N_14444,N_14481);
xor U14591 (N_14591,N_14505,N_14520);
or U14592 (N_14592,N_14529,N_14512);
or U14593 (N_14593,N_14508,N_14557);
nor U14594 (N_14594,N_14404,N_14412);
nand U14595 (N_14595,N_14426,N_14402);
xnor U14596 (N_14596,N_14437,N_14528);
or U14597 (N_14597,N_14538,N_14403);
xnor U14598 (N_14598,N_14517,N_14534);
nor U14599 (N_14599,N_14524,N_14496);
or U14600 (N_14600,N_14507,N_14458);
xnor U14601 (N_14601,N_14441,N_14455);
xnor U14602 (N_14602,N_14559,N_14525);
and U14603 (N_14603,N_14429,N_14502);
xnor U14604 (N_14604,N_14497,N_14476);
nand U14605 (N_14605,N_14445,N_14438);
and U14606 (N_14606,N_14428,N_14523);
xor U14607 (N_14607,N_14470,N_14421);
and U14608 (N_14608,N_14427,N_14435);
nor U14609 (N_14609,N_14465,N_14400);
nand U14610 (N_14610,N_14514,N_14483);
nand U14611 (N_14611,N_14469,N_14546);
xnor U14612 (N_14612,N_14555,N_14558);
nor U14613 (N_14613,N_14510,N_14453);
and U14614 (N_14614,N_14449,N_14519);
xnor U14615 (N_14615,N_14540,N_14509);
nand U14616 (N_14616,N_14477,N_14475);
and U14617 (N_14617,N_14504,N_14472);
or U14618 (N_14618,N_14501,N_14408);
nor U14619 (N_14619,N_14550,N_14542);
or U14620 (N_14620,N_14522,N_14544);
nand U14621 (N_14621,N_14407,N_14532);
and U14622 (N_14622,N_14541,N_14436);
or U14623 (N_14623,N_14401,N_14530);
xor U14624 (N_14624,N_14521,N_14511);
and U14625 (N_14625,N_14439,N_14506);
or U14626 (N_14626,N_14409,N_14420);
nand U14627 (N_14627,N_14493,N_14443);
xor U14628 (N_14628,N_14547,N_14480);
nand U14629 (N_14629,N_14406,N_14422);
and U14630 (N_14630,N_14515,N_14431);
xnor U14631 (N_14631,N_14526,N_14423);
nand U14632 (N_14632,N_14551,N_14471);
nand U14633 (N_14633,N_14461,N_14410);
or U14634 (N_14634,N_14457,N_14417);
and U14635 (N_14635,N_14498,N_14466);
and U14636 (N_14636,N_14549,N_14467);
xnor U14637 (N_14637,N_14419,N_14499);
and U14638 (N_14638,N_14460,N_14418);
xor U14639 (N_14639,N_14456,N_14482);
and U14640 (N_14640,N_14513,N_14542);
nor U14641 (N_14641,N_14529,N_14531);
xor U14642 (N_14642,N_14404,N_14403);
nand U14643 (N_14643,N_14411,N_14465);
xor U14644 (N_14644,N_14527,N_14551);
or U14645 (N_14645,N_14511,N_14417);
nor U14646 (N_14646,N_14426,N_14554);
and U14647 (N_14647,N_14419,N_14555);
or U14648 (N_14648,N_14461,N_14523);
or U14649 (N_14649,N_14467,N_14518);
or U14650 (N_14650,N_14445,N_14480);
and U14651 (N_14651,N_14511,N_14406);
xor U14652 (N_14652,N_14539,N_14432);
and U14653 (N_14653,N_14447,N_14559);
nand U14654 (N_14654,N_14469,N_14467);
and U14655 (N_14655,N_14525,N_14504);
xor U14656 (N_14656,N_14489,N_14488);
and U14657 (N_14657,N_14420,N_14513);
and U14658 (N_14658,N_14546,N_14530);
xor U14659 (N_14659,N_14418,N_14405);
nand U14660 (N_14660,N_14412,N_14540);
or U14661 (N_14661,N_14506,N_14442);
or U14662 (N_14662,N_14480,N_14433);
or U14663 (N_14663,N_14551,N_14435);
xnor U14664 (N_14664,N_14463,N_14438);
nor U14665 (N_14665,N_14400,N_14506);
and U14666 (N_14666,N_14453,N_14484);
xor U14667 (N_14667,N_14520,N_14458);
or U14668 (N_14668,N_14410,N_14413);
and U14669 (N_14669,N_14539,N_14471);
or U14670 (N_14670,N_14501,N_14522);
and U14671 (N_14671,N_14423,N_14549);
or U14672 (N_14672,N_14515,N_14547);
or U14673 (N_14673,N_14476,N_14496);
nor U14674 (N_14674,N_14537,N_14534);
xnor U14675 (N_14675,N_14443,N_14506);
or U14676 (N_14676,N_14409,N_14505);
nand U14677 (N_14677,N_14490,N_14487);
nand U14678 (N_14678,N_14540,N_14529);
nor U14679 (N_14679,N_14525,N_14500);
nand U14680 (N_14680,N_14425,N_14519);
nand U14681 (N_14681,N_14505,N_14499);
or U14682 (N_14682,N_14414,N_14439);
xor U14683 (N_14683,N_14488,N_14425);
and U14684 (N_14684,N_14441,N_14462);
xnor U14685 (N_14685,N_14500,N_14551);
or U14686 (N_14686,N_14518,N_14511);
nor U14687 (N_14687,N_14425,N_14554);
xnor U14688 (N_14688,N_14483,N_14546);
and U14689 (N_14689,N_14548,N_14545);
nor U14690 (N_14690,N_14490,N_14420);
or U14691 (N_14691,N_14521,N_14483);
or U14692 (N_14692,N_14504,N_14493);
and U14693 (N_14693,N_14445,N_14433);
or U14694 (N_14694,N_14464,N_14493);
nand U14695 (N_14695,N_14467,N_14520);
nor U14696 (N_14696,N_14524,N_14429);
nand U14697 (N_14697,N_14516,N_14477);
or U14698 (N_14698,N_14412,N_14559);
or U14699 (N_14699,N_14502,N_14513);
nor U14700 (N_14700,N_14439,N_14436);
nor U14701 (N_14701,N_14451,N_14416);
xor U14702 (N_14702,N_14446,N_14426);
nor U14703 (N_14703,N_14456,N_14559);
and U14704 (N_14704,N_14556,N_14544);
nor U14705 (N_14705,N_14437,N_14462);
xnor U14706 (N_14706,N_14423,N_14533);
xnor U14707 (N_14707,N_14461,N_14433);
nand U14708 (N_14708,N_14434,N_14426);
and U14709 (N_14709,N_14432,N_14524);
xnor U14710 (N_14710,N_14438,N_14497);
nor U14711 (N_14711,N_14407,N_14444);
nand U14712 (N_14712,N_14511,N_14514);
and U14713 (N_14713,N_14427,N_14501);
or U14714 (N_14714,N_14463,N_14465);
or U14715 (N_14715,N_14550,N_14557);
xnor U14716 (N_14716,N_14494,N_14533);
nand U14717 (N_14717,N_14522,N_14490);
xor U14718 (N_14718,N_14421,N_14468);
nor U14719 (N_14719,N_14464,N_14415);
xor U14720 (N_14720,N_14601,N_14711);
nand U14721 (N_14721,N_14580,N_14603);
nand U14722 (N_14722,N_14642,N_14609);
or U14723 (N_14723,N_14612,N_14617);
or U14724 (N_14724,N_14599,N_14573);
or U14725 (N_14725,N_14588,N_14687);
and U14726 (N_14726,N_14679,N_14566);
nor U14727 (N_14727,N_14598,N_14641);
nand U14728 (N_14728,N_14637,N_14686);
nand U14729 (N_14729,N_14657,N_14632);
nand U14730 (N_14730,N_14633,N_14688);
nand U14731 (N_14731,N_14690,N_14593);
nor U14732 (N_14732,N_14674,N_14715);
xnor U14733 (N_14733,N_14619,N_14705);
and U14734 (N_14734,N_14704,N_14636);
nand U14735 (N_14735,N_14639,N_14663);
nor U14736 (N_14736,N_14570,N_14654);
and U14737 (N_14737,N_14596,N_14615);
or U14738 (N_14738,N_14635,N_14565);
xor U14739 (N_14739,N_14613,N_14577);
nand U14740 (N_14740,N_14594,N_14622);
xnor U14741 (N_14741,N_14600,N_14666);
nand U14742 (N_14742,N_14714,N_14591);
and U14743 (N_14743,N_14651,N_14578);
nor U14744 (N_14744,N_14579,N_14698);
or U14745 (N_14745,N_14648,N_14629);
or U14746 (N_14746,N_14586,N_14621);
nand U14747 (N_14747,N_14631,N_14630);
xnor U14748 (N_14748,N_14569,N_14667);
and U14749 (N_14749,N_14712,N_14575);
xor U14750 (N_14750,N_14655,N_14634);
and U14751 (N_14751,N_14645,N_14713);
nor U14752 (N_14752,N_14656,N_14644);
nor U14753 (N_14753,N_14691,N_14652);
nand U14754 (N_14754,N_14627,N_14626);
nand U14755 (N_14755,N_14659,N_14673);
and U14756 (N_14756,N_14563,N_14694);
or U14757 (N_14757,N_14590,N_14562);
or U14758 (N_14758,N_14692,N_14697);
nor U14759 (N_14759,N_14611,N_14669);
nor U14760 (N_14760,N_14571,N_14574);
xnor U14761 (N_14761,N_14606,N_14682);
and U14762 (N_14762,N_14683,N_14620);
xor U14763 (N_14763,N_14701,N_14581);
and U14764 (N_14764,N_14681,N_14680);
or U14765 (N_14765,N_14605,N_14592);
nand U14766 (N_14766,N_14561,N_14589);
xnor U14767 (N_14767,N_14707,N_14678);
nor U14768 (N_14768,N_14567,N_14647);
nor U14769 (N_14769,N_14582,N_14676);
and U14770 (N_14770,N_14709,N_14608);
nor U14771 (N_14771,N_14672,N_14628);
nand U14772 (N_14772,N_14660,N_14584);
xnor U14773 (N_14773,N_14703,N_14618);
or U14774 (N_14774,N_14675,N_14710);
nand U14775 (N_14775,N_14595,N_14668);
nand U14776 (N_14776,N_14706,N_14695);
and U14777 (N_14777,N_14610,N_14719);
xnor U14778 (N_14778,N_14576,N_14587);
and U14779 (N_14779,N_14699,N_14717);
xor U14780 (N_14780,N_14670,N_14602);
xor U14781 (N_14781,N_14649,N_14685);
or U14782 (N_14782,N_14708,N_14623);
xor U14783 (N_14783,N_14604,N_14696);
or U14784 (N_14784,N_14702,N_14585);
xnor U14785 (N_14785,N_14560,N_14718);
xor U14786 (N_14786,N_14662,N_14646);
and U14787 (N_14787,N_14661,N_14564);
nand U14788 (N_14788,N_14664,N_14650);
or U14789 (N_14789,N_14607,N_14614);
and U14790 (N_14790,N_14572,N_14640);
nand U14791 (N_14791,N_14716,N_14653);
and U14792 (N_14792,N_14689,N_14597);
nand U14793 (N_14793,N_14693,N_14671);
nor U14794 (N_14794,N_14643,N_14568);
and U14795 (N_14795,N_14583,N_14625);
nand U14796 (N_14796,N_14677,N_14665);
nand U14797 (N_14797,N_14658,N_14616);
xnor U14798 (N_14798,N_14638,N_14684);
nand U14799 (N_14799,N_14624,N_14700);
and U14800 (N_14800,N_14650,N_14707);
or U14801 (N_14801,N_14573,N_14716);
nand U14802 (N_14802,N_14653,N_14586);
and U14803 (N_14803,N_14588,N_14650);
and U14804 (N_14804,N_14579,N_14648);
or U14805 (N_14805,N_14682,N_14586);
nor U14806 (N_14806,N_14621,N_14567);
nand U14807 (N_14807,N_14662,N_14592);
xnor U14808 (N_14808,N_14560,N_14694);
xor U14809 (N_14809,N_14583,N_14699);
or U14810 (N_14810,N_14568,N_14621);
and U14811 (N_14811,N_14691,N_14616);
xnor U14812 (N_14812,N_14664,N_14649);
xnor U14813 (N_14813,N_14638,N_14576);
or U14814 (N_14814,N_14654,N_14704);
nor U14815 (N_14815,N_14711,N_14602);
xor U14816 (N_14816,N_14585,N_14680);
or U14817 (N_14817,N_14710,N_14719);
nor U14818 (N_14818,N_14657,N_14606);
xor U14819 (N_14819,N_14561,N_14679);
nand U14820 (N_14820,N_14580,N_14596);
or U14821 (N_14821,N_14678,N_14709);
and U14822 (N_14822,N_14716,N_14561);
or U14823 (N_14823,N_14668,N_14628);
xnor U14824 (N_14824,N_14598,N_14708);
xor U14825 (N_14825,N_14577,N_14702);
and U14826 (N_14826,N_14647,N_14668);
nand U14827 (N_14827,N_14652,N_14593);
and U14828 (N_14828,N_14604,N_14584);
or U14829 (N_14829,N_14561,N_14689);
nand U14830 (N_14830,N_14577,N_14635);
and U14831 (N_14831,N_14704,N_14708);
xnor U14832 (N_14832,N_14561,N_14696);
and U14833 (N_14833,N_14562,N_14710);
nor U14834 (N_14834,N_14646,N_14712);
nor U14835 (N_14835,N_14608,N_14674);
nand U14836 (N_14836,N_14586,N_14693);
nand U14837 (N_14837,N_14603,N_14717);
and U14838 (N_14838,N_14695,N_14678);
nand U14839 (N_14839,N_14566,N_14631);
nand U14840 (N_14840,N_14590,N_14683);
xor U14841 (N_14841,N_14596,N_14684);
nand U14842 (N_14842,N_14645,N_14636);
or U14843 (N_14843,N_14641,N_14584);
nand U14844 (N_14844,N_14562,N_14647);
or U14845 (N_14845,N_14607,N_14563);
or U14846 (N_14846,N_14660,N_14661);
or U14847 (N_14847,N_14584,N_14597);
nand U14848 (N_14848,N_14662,N_14615);
and U14849 (N_14849,N_14683,N_14645);
nor U14850 (N_14850,N_14685,N_14719);
nor U14851 (N_14851,N_14688,N_14707);
xor U14852 (N_14852,N_14648,N_14698);
nor U14853 (N_14853,N_14562,N_14662);
and U14854 (N_14854,N_14592,N_14624);
and U14855 (N_14855,N_14661,N_14628);
xor U14856 (N_14856,N_14585,N_14621);
nand U14857 (N_14857,N_14636,N_14581);
or U14858 (N_14858,N_14706,N_14714);
nand U14859 (N_14859,N_14711,N_14700);
nor U14860 (N_14860,N_14571,N_14641);
xor U14861 (N_14861,N_14566,N_14628);
or U14862 (N_14862,N_14606,N_14709);
or U14863 (N_14863,N_14609,N_14629);
and U14864 (N_14864,N_14642,N_14584);
or U14865 (N_14865,N_14629,N_14561);
or U14866 (N_14866,N_14579,N_14568);
or U14867 (N_14867,N_14675,N_14699);
and U14868 (N_14868,N_14613,N_14706);
or U14869 (N_14869,N_14664,N_14594);
or U14870 (N_14870,N_14667,N_14624);
nor U14871 (N_14871,N_14594,N_14712);
or U14872 (N_14872,N_14582,N_14668);
nand U14873 (N_14873,N_14683,N_14588);
or U14874 (N_14874,N_14578,N_14703);
nand U14875 (N_14875,N_14612,N_14638);
or U14876 (N_14876,N_14697,N_14688);
xor U14877 (N_14877,N_14716,N_14659);
nor U14878 (N_14878,N_14624,N_14588);
nor U14879 (N_14879,N_14648,N_14627);
and U14880 (N_14880,N_14823,N_14809);
and U14881 (N_14881,N_14792,N_14816);
nand U14882 (N_14882,N_14822,N_14732);
nand U14883 (N_14883,N_14742,N_14785);
xnor U14884 (N_14884,N_14782,N_14807);
xor U14885 (N_14885,N_14865,N_14875);
nand U14886 (N_14886,N_14866,N_14727);
nor U14887 (N_14887,N_14850,N_14802);
nand U14888 (N_14888,N_14847,N_14759);
nor U14889 (N_14889,N_14749,N_14805);
and U14890 (N_14890,N_14838,N_14728);
nand U14891 (N_14891,N_14818,N_14862);
nor U14892 (N_14892,N_14870,N_14832);
and U14893 (N_14893,N_14817,N_14801);
xnor U14894 (N_14894,N_14783,N_14828);
and U14895 (N_14895,N_14798,N_14754);
nor U14896 (N_14896,N_14824,N_14833);
nor U14897 (N_14897,N_14762,N_14840);
nor U14898 (N_14898,N_14836,N_14763);
or U14899 (N_14899,N_14812,N_14819);
and U14900 (N_14900,N_14835,N_14748);
or U14901 (N_14901,N_14874,N_14808);
and U14902 (N_14902,N_14803,N_14730);
nand U14903 (N_14903,N_14753,N_14741);
and U14904 (N_14904,N_14829,N_14804);
nor U14905 (N_14905,N_14767,N_14859);
xnor U14906 (N_14906,N_14839,N_14806);
nor U14907 (N_14907,N_14872,N_14733);
nand U14908 (N_14908,N_14775,N_14744);
nor U14909 (N_14909,N_14745,N_14857);
xor U14910 (N_14910,N_14820,N_14723);
and U14911 (N_14911,N_14821,N_14858);
or U14912 (N_14912,N_14793,N_14796);
and U14913 (N_14913,N_14771,N_14769);
xor U14914 (N_14914,N_14845,N_14867);
nand U14915 (N_14915,N_14811,N_14787);
nand U14916 (N_14916,N_14766,N_14747);
nor U14917 (N_14917,N_14722,N_14720);
nand U14918 (N_14918,N_14831,N_14764);
nand U14919 (N_14919,N_14735,N_14813);
nand U14920 (N_14920,N_14842,N_14871);
xor U14921 (N_14921,N_14757,N_14810);
nand U14922 (N_14922,N_14837,N_14770);
and U14923 (N_14923,N_14815,N_14786);
xor U14924 (N_14924,N_14799,N_14740);
or U14925 (N_14925,N_14751,N_14860);
nand U14926 (N_14926,N_14724,N_14774);
xor U14927 (N_14927,N_14868,N_14876);
xnor U14928 (N_14928,N_14841,N_14773);
nor U14929 (N_14929,N_14873,N_14765);
xor U14930 (N_14930,N_14848,N_14794);
nor U14931 (N_14931,N_14746,N_14852);
xor U14932 (N_14932,N_14800,N_14755);
nand U14933 (N_14933,N_14846,N_14855);
and U14934 (N_14934,N_14750,N_14779);
nand U14935 (N_14935,N_14778,N_14736);
nor U14936 (N_14936,N_14758,N_14791);
and U14937 (N_14937,N_14739,N_14869);
nand U14938 (N_14938,N_14789,N_14856);
nand U14939 (N_14939,N_14826,N_14843);
xor U14940 (N_14940,N_14737,N_14760);
or U14941 (N_14941,N_14861,N_14795);
or U14942 (N_14942,N_14761,N_14776);
and U14943 (N_14943,N_14731,N_14777);
nor U14944 (N_14944,N_14878,N_14879);
or U14945 (N_14945,N_14734,N_14827);
nand U14946 (N_14946,N_14877,N_14756);
and U14947 (N_14947,N_14780,N_14725);
or U14948 (N_14948,N_14788,N_14849);
and U14949 (N_14949,N_14830,N_14738);
nor U14950 (N_14950,N_14853,N_14790);
or U14951 (N_14951,N_14772,N_14851);
nor U14952 (N_14952,N_14721,N_14864);
nand U14953 (N_14953,N_14752,N_14863);
nor U14954 (N_14954,N_14814,N_14844);
and U14955 (N_14955,N_14781,N_14825);
xor U14956 (N_14956,N_14784,N_14797);
nor U14957 (N_14957,N_14768,N_14834);
or U14958 (N_14958,N_14729,N_14854);
xor U14959 (N_14959,N_14743,N_14726);
xnor U14960 (N_14960,N_14726,N_14772);
and U14961 (N_14961,N_14850,N_14810);
nand U14962 (N_14962,N_14778,N_14794);
nor U14963 (N_14963,N_14855,N_14867);
or U14964 (N_14964,N_14813,N_14859);
or U14965 (N_14965,N_14858,N_14764);
and U14966 (N_14966,N_14828,N_14771);
and U14967 (N_14967,N_14805,N_14773);
nand U14968 (N_14968,N_14825,N_14782);
or U14969 (N_14969,N_14731,N_14720);
or U14970 (N_14970,N_14789,N_14728);
or U14971 (N_14971,N_14827,N_14819);
and U14972 (N_14972,N_14806,N_14741);
nor U14973 (N_14973,N_14747,N_14836);
xnor U14974 (N_14974,N_14722,N_14796);
nand U14975 (N_14975,N_14812,N_14754);
or U14976 (N_14976,N_14746,N_14826);
nor U14977 (N_14977,N_14772,N_14752);
or U14978 (N_14978,N_14831,N_14794);
xnor U14979 (N_14979,N_14750,N_14866);
xor U14980 (N_14980,N_14787,N_14755);
or U14981 (N_14981,N_14768,N_14778);
or U14982 (N_14982,N_14813,N_14784);
and U14983 (N_14983,N_14755,N_14845);
nor U14984 (N_14984,N_14731,N_14875);
nor U14985 (N_14985,N_14808,N_14729);
nand U14986 (N_14986,N_14782,N_14795);
xor U14987 (N_14987,N_14738,N_14749);
nand U14988 (N_14988,N_14759,N_14736);
nand U14989 (N_14989,N_14868,N_14848);
nor U14990 (N_14990,N_14721,N_14873);
nand U14991 (N_14991,N_14813,N_14733);
and U14992 (N_14992,N_14795,N_14739);
nor U14993 (N_14993,N_14818,N_14843);
xor U14994 (N_14994,N_14724,N_14862);
nor U14995 (N_14995,N_14776,N_14809);
xor U14996 (N_14996,N_14865,N_14829);
xor U14997 (N_14997,N_14825,N_14779);
and U14998 (N_14998,N_14726,N_14829);
nand U14999 (N_14999,N_14722,N_14752);
nor U15000 (N_15000,N_14776,N_14879);
nor U15001 (N_15001,N_14762,N_14828);
and U15002 (N_15002,N_14870,N_14815);
nand U15003 (N_15003,N_14780,N_14795);
xor U15004 (N_15004,N_14846,N_14733);
or U15005 (N_15005,N_14755,N_14830);
and U15006 (N_15006,N_14731,N_14826);
nand U15007 (N_15007,N_14838,N_14863);
nand U15008 (N_15008,N_14744,N_14793);
xnor U15009 (N_15009,N_14739,N_14877);
xor U15010 (N_15010,N_14849,N_14721);
nor U15011 (N_15011,N_14827,N_14740);
nand U15012 (N_15012,N_14801,N_14807);
nor U15013 (N_15013,N_14840,N_14835);
and U15014 (N_15014,N_14830,N_14790);
or U15015 (N_15015,N_14735,N_14761);
xnor U15016 (N_15016,N_14761,N_14802);
nor U15017 (N_15017,N_14771,N_14825);
and U15018 (N_15018,N_14744,N_14721);
nand U15019 (N_15019,N_14830,N_14857);
or U15020 (N_15020,N_14867,N_14861);
or U15021 (N_15021,N_14738,N_14767);
xnor U15022 (N_15022,N_14828,N_14798);
nor U15023 (N_15023,N_14803,N_14770);
or U15024 (N_15024,N_14792,N_14724);
and U15025 (N_15025,N_14729,N_14867);
xor U15026 (N_15026,N_14831,N_14747);
nor U15027 (N_15027,N_14836,N_14835);
nand U15028 (N_15028,N_14871,N_14788);
xor U15029 (N_15029,N_14790,N_14812);
xnor U15030 (N_15030,N_14833,N_14781);
xnor U15031 (N_15031,N_14873,N_14785);
and U15032 (N_15032,N_14859,N_14736);
nor U15033 (N_15033,N_14758,N_14721);
or U15034 (N_15034,N_14761,N_14729);
xor U15035 (N_15035,N_14822,N_14733);
or U15036 (N_15036,N_14810,N_14775);
xor U15037 (N_15037,N_14769,N_14752);
nand U15038 (N_15038,N_14823,N_14828);
nand U15039 (N_15039,N_14820,N_14756);
nand U15040 (N_15040,N_15027,N_15011);
and U15041 (N_15041,N_14910,N_14989);
nand U15042 (N_15042,N_15015,N_15030);
and U15043 (N_15043,N_14924,N_15032);
nand U15044 (N_15044,N_14883,N_14917);
nand U15045 (N_15045,N_15033,N_14888);
and U15046 (N_15046,N_15029,N_14896);
nor U15047 (N_15047,N_15019,N_14885);
xnor U15048 (N_15048,N_14937,N_14939);
or U15049 (N_15049,N_15009,N_15003);
or U15050 (N_15050,N_14908,N_14987);
and U15051 (N_15051,N_14988,N_15036);
nand U15052 (N_15052,N_14884,N_15022);
or U15053 (N_15053,N_14956,N_15026);
xor U15054 (N_15054,N_15010,N_14902);
nor U15055 (N_15055,N_14925,N_14999);
or U15056 (N_15056,N_14930,N_14991);
or U15057 (N_15057,N_14949,N_14997);
nor U15058 (N_15058,N_15013,N_14998);
nand U15059 (N_15059,N_14945,N_15017);
and U15060 (N_15060,N_14955,N_14996);
or U15061 (N_15061,N_14976,N_14882);
nand U15062 (N_15062,N_14951,N_14899);
nor U15063 (N_15063,N_15035,N_14895);
nor U15064 (N_15064,N_14957,N_14960);
or U15065 (N_15065,N_14978,N_14948);
nand U15066 (N_15066,N_14915,N_14913);
and U15067 (N_15067,N_14942,N_14894);
and U15068 (N_15068,N_15037,N_15001);
nor U15069 (N_15069,N_14932,N_14938);
or U15070 (N_15070,N_15038,N_14995);
and U15071 (N_15071,N_15023,N_14912);
nor U15072 (N_15072,N_14905,N_14892);
xnor U15073 (N_15073,N_14952,N_14903);
xnor U15074 (N_15074,N_14934,N_15028);
and U15075 (N_15075,N_15016,N_14972);
or U15076 (N_15076,N_14909,N_14964);
nor U15077 (N_15077,N_14940,N_14966);
xnor U15078 (N_15078,N_14943,N_14977);
nand U15079 (N_15079,N_14907,N_14979);
nand U15080 (N_15080,N_14981,N_15034);
and U15081 (N_15081,N_14967,N_14953);
xnor U15082 (N_15082,N_15039,N_14887);
xor U15083 (N_15083,N_14946,N_14904);
or U15084 (N_15084,N_14900,N_14984);
and U15085 (N_15085,N_14993,N_15021);
and U15086 (N_15086,N_14897,N_15025);
and U15087 (N_15087,N_14886,N_14901);
and U15088 (N_15088,N_14947,N_14926);
nor U15089 (N_15089,N_15018,N_14963);
xor U15090 (N_15090,N_14922,N_14959);
and U15091 (N_15091,N_14890,N_14880);
and U15092 (N_15092,N_14994,N_15004);
nand U15093 (N_15093,N_14931,N_14980);
and U15094 (N_15094,N_14920,N_14954);
or U15095 (N_15095,N_14970,N_14893);
and U15096 (N_15096,N_14928,N_14962);
nand U15097 (N_15097,N_15008,N_14918);
xor U15098 (N_15098,N_14983,N_14969);
or U15099 (N_15099,N_14973,N_15024);
xor U15100 (N_15100,N_14916,N_15012);
nor U15101 (N_15101,N_14914,N_14971);
nand U15102 (N_15102,N_14921,N_14982);
nor U15103 (N_15103,N_14929,N_15014);
and U15104 (N_15104,N_14992,N_14950);
xor U15105 (N_15105,N_14958,N_15031);
and U15106 (N_15106,N_14936,N_15005);
and U15107 (N_15107,N_14898,N_15002);
and U15108 (N_15108,N_14933,N_14927);
nand U15109 (N_15109,N_15007,N_14889);
and U15110 (N_15110,N_14965,N_15020);
and U15111 (N_15111,N_14986,N_14974);
nor U15112 (N_15112,N_14935,N_14923);
nor U15113 (N_15113,N_15006,N_14944);
xor U15114 (N_15114,N_14919,N_15000);
and U15115 (N_15115,N_14911,N_14985);
or U15116 (N_15116,N_14975,N_14968);
and U15117 (N_15117,N_14891,N_14881);
and U15118 (N_15118,N_14961,N_14906);
and U15119 (N_15119,N_14941,N_14990);
nor U15120 (N_15120,N_14893,N_14883);
nor U15121 (N_15121,N_15007,N_14898);
xor U15122 (N_15122,N_14981,N_14968);
and U15123 (N_15123,N_14937,N_14911);
or U15124 (N_15124,N_14945,N_14944);
nand U15125 (N_15125,N_15018,N_15021);
nor U15126 (N_15126,N_14962,N_14963);
and U15127 (N_15127,N_14977,N_14947);
nor U15128 (N_15128,N_14940,N_14887);
or U15129 (N_15129,N_15025,N_14920);
nor U15130 (N_15130,N_14906,N_14996);
nor U15131 (N_15131,N_15036,N_14965);
and U15132 (N_15132,N_14942,N_15020);
or U15133 (N_15133,N_14982,N_15020);
xor U15134 (N_15134,N_15001,N_14902);
xor U15135 (N_15135,N_14947,N_14918);
nor U15136 (N_15136,N_14989,N_14923);
or U15137 (N_15137,N_14910,N_15016);
or U15138 (N_15138,N_14948,N_14912);
or U15139 (N_15139,N_14958,N_14909);
or U15140 (N_15140,N_14964,N_14899);
xor U15141 (N_15141,N_14886,N_14915);
nand U15142 (N_15142,N_14965,N_14938);
and U15143 (N_15143,N_14911,N_14982);
xnor U15144 (N_15144,N_14918,N_14919);
xor U15145 (N_15145,N_14935,N_14962);
and U15146 (N_15146,N_14885,N_14917);
or U15147 (N_15147,N_14993,N_14986);
xor U15148 (N_15148,N_14964,N_14998);
and U15149 (N_15149,N_14941,N_14984);
xnor U15150 (N_15150,N_14896,N_14990);
or U15151 (N_15151,N_15015,N_14940);
and U15152 (N_15152,N_15030,N_14957);
nor U15153 (N_15153,N_14925,N_14941);
xnor U15154 (N_15154,N_14972,N_14973);
or U15155 (N_15155,N_14932,N_15037);
nor U15156 (N_15156,N_15007,N_15036);
nor U15157 (N_15157,N_14926,N_14895);
xnor U15158 (N_15158,N_14883,N_14881);
or U15159 (N_15159,N_15007,N_15014);
nor U15160 (N_15160,N_15034,N_14978);
nor U15161 (N_15161,N_14947,N_14911);
nand U15162 (N_15162,N_14903,N_15035);
nor U15163 (N_15163,N_14916,N_14989);
xnor U15164 (N_15164,N_14976,N_14898);
nand U15165 (N_15165,N_14995,N_15022);
xnor U15166 (N_15166,N_15008,N_15003);
nand U15167 (N_15167,N_14919,N_14938);
nor U15168 (N_15168,N_14896,N_15024);
xor U15169 (N_15169,N_15006,N_14997);
nor U15170 (N_15170,N_14946,N_14981);
and U15171 (N_15171,N_14910,N_15004);
and U15172 (N_15172,N_14915,N_14984);
and U15173 (N_15173,N_15007,N_15039);
nand U15174 (N_15174,N_14971,N_14892);
nand U15175 (N_15175,N_14915,N_14992);
nand U15176 (N_15176,N_14963,N_14970);
nor U15177 (N_15177,N_15032,N_14974);
xor U15178 (N_15178,N_14881,N_14941);
and U15179 (N_15179,N_14920,N_14950);
nor U15180 (N_15180,N_14937,N_14961);
xnor U15181 (N_15181,N_14882,N_14968);
nor U15182 (N_15182,N_14924,N_15000);
or U15183 (N_15183,N_14958,N_15009);
nand U15184 (N_15184,N_14943,N_14939);
nand U15185 (N_15185,N_14927,N_15008);
xnor U15186 (N_15186,N_14893,N_14889);
nor U15187 (N_15187,N_14975,N_14894);
nand U15188 (N_15188,N_14994,N_14944);
and U15189 (N_15189,N_14963,N_14921);
and U15190 (N_15190,N_14937,N_14934);
and U15191 (N_15191,N_15039,N_15027);
nor U15192 (N_15192,N_14891,N_14996);
xor U15193 (N_15193,N_14976,N_15015);
xnor U15194 (N_15194,N_14983,N_15018);
nor U15195 (N_15195,N_14968,N_14934);
nor U15196 (N_15196,N_14908,N_14918);
nor U15197 (N_15197,N_14909,N_15036);
or U15198 (N_15198,N_14894,N_14890);
nor U15199 (N_15199,N_14979,N_14981);
and U15200 (N_15200,N_15190,N_15082);
nor U15201 (N_15201,N_15046,N_15067);
xor U15202 (N_15202,N_15066,N_15105);
nand U15203 (N_15203,N_15120,N_15103);
nand U15204 (N_15204,N_15130,N_15172);
xor U15205 (N_15205,N_15176,N_15171);
nand U15206 (N_15206,N_15166,N_15064);
xnor U15207 (N_15207,N_15041,N_15148);
xor U15208 (N_15208,N_15068,N_15052);
and U15209 (N_15209,N_15090,N_15075);
or U15210 (N_15210,N_15179,N_15054);
xnor U15211 (N_15211,N_15069,N_15085);
nand U15212 (N_15212,N_15157,N_15086);
or U15213 (N_15213,N_15196,N_15057);
xnor U15214 (N_15214,N_15113,N_15106);
xnor U15215 (N_15215,N_15073,N_15117);
xor U15216 (N_15216,N_15127,N_15189);
and U15217 (N_15217,N_15142,N_15059);
nand U15218 (N_15218,N_15154,N_15193);
and U15219 (N_15219,N_15123,N_15124);
nor U15220 (N_15220,N_15074,N_15131);
xor U15221 (N_15221,N_15173,N_15164);
or U15222 (N_15222,N_15182,N_15165);
xor U15223 (N_15223,N_15137,N_15099);
or U15224 (N_15224,N_15092,N_15144);
and U15225 (N_15225,N_15167,N_15198);
nand U15226 (N_15226,N_15135,N_15048);
and U15227 (N_15227,N_15134,N_15097);
nor U15228 (N_15228,N_15118,N_15102);
and U15229 (N_15229,N_15070,N_15186);
or U15230 (N_15230,N_15043,N_15191);
nor U15231 (N_15231,N_15168,N_15056);
and U15232 (N_15232,N_15040,N_15177);
xnor U15233 (N_15233,N_15096,N_15141);
xor U15234 (N_15234,N_15170,N_15169);
nor U15235 (N_15235,N_15108,N_15119);
xor U15236 (N_15236,N_15091,N_15079);
xnor U15237 (N_15237,N_15049,N_15116);
nor U15238 (N_15238,N_15093,N_15051);
nor U15239 (N_15239,N_15072,N_15163);
nor U15240 (N_15240,N_15149,N_15161);
nand U15241 (N_15241,N_15076,N_15151);
nand U15242 (N_15242,N_15050,N_15044);
xnor U15243 (N_15243,N_15194,N_15143);
or U15244 (N_15244,N_15089,N_15178);
nor U15245 (N_15245,N_15109,N_15195);
nor U15246 (N_15246,N_15133,N_15114);
xnor U15247 (N_15247,N_15175,N_15063);
and U15248 (N_15248,N_15184,N_15139);
and U15249 (N_15249,N_15045,N_15162);
nor U15250 (N_15250,N_15145,N_15192);
nand U15251 (N_15251,N_15188,N_15047);
nand U15252 (N_15252,N_15053,N_15183);
and U15253 (N_15253,N_15065,N_15125);
or U15254 (N_15254,N_15174,N_15110);
or U15255 (N_15255,N_15155,N_15095);
or U15256 (N_15256,N_15080,N_15078);
or U15257 (N_15257,N_15129,N_15060);
xor U15258 (N_15258,N_15147,N_15150);
or U15259 (N_15259,N_15126,N_15122);
nand U15260 (N_15260,N_15197,N_15107);
or U15261 (N_15261,N_15152,N_15132);
nor U15262 (N_15262,N_15087,N_15084);
nor U15263 (N_15263,N_15098,N_15058);
or U15264 (N_15264,N_15160,N_15062);
and U15265 (N_15265,N_15180,N_15156);
xor U15266 (N_15266,N_15146,N_15199);
or U15267 (N_15267,N_15159,N_15181);
or U15268 (N_15268,N_15185,N_15138);
xor U15269 (N_15269,N_15128,N_15104);
and U15270 (N_15270,N_15100,N_15055);
nand U15271 (N_15271,N_15111,N_15077);
or U15272 (N_15272,N_15187,N_15153);
and U15273 (N_15273,N_15088,N_15121);
nand U15274 (N_15274,N_15061,N_15071);
nand U15275 (N_15275,N_15083,N_15136);
nor U15276 (N_15276,N_15158,N_15112);
nand U15277 (N_15277,N_15115,N_15101);
or U15278 (N_15278,N_15081,N_15140);
nor U15279 (N_15279,N_15094,N_15042);
or U15280 (N_15280,N_15136,N_15183);
or U15281 (N_15281,N_15096,N_15080);
or U15282 (N_15282,N_15124,N_15135);
xnor U15283 (N_15283,N_15112,N_15106);
nand U15284 (N_15284,N_15178,N_15087);
nand U15285 (N_15285,N_15189,N_15135);
nor U15286 (N_15286,N_15077,N_15108);
and U15287 (N_15287,N_15170,N_15070);
or U15288 (N_15288,N_15042,N_15167);
xnor U15289 (N_15289,N_15080,N_15068);
and U15290 (N_15290,N_15196,N_15178);
and U15291 (N_15291,N_15141,N_15167);
or U15292 (N_15292,N_15091,N_15074);
or U15293 (N_15293,N_15196,N_15076);
nor U15294 (N_15294,N_15042,N_15151);
or U15295 (N_15295,N_15109,N_15060);
nand U15296 (N_15296,N_15075,N_15197);
and U15297 (N_15297,N_15077,N_15098);
nand U15298 (N_15298,N_15196,N_15138);
nand U15299 (N_15299,N_15080,N_15127);
nand U15300 (N_15300,N_15157,N_15067);
nand U15301 (N_15301,N_15185,N_15147);
xor U15302 (N_15302,N_15188,N_15079);
nand U15303 (N_15303,N_15050,N_15155);
nand U15304 (N_15304,N_15068,N_15074);
and U15305 (N_15305,N_15109,N_15133);
xor U15306 (N_15306,N_15148,N_15140);
nand U15307 (N_15307,N_15102,N_15180);
and U15308 (N_15308,N_15147,N_15199);
nor U15309 (N_15309,N_15180,N_15078);
and U15310 (N_15310,N_15125,N_15189);
and U15311 (N_15311,N_15188,N_15128);
nand U15312 (N_15312,N_15111,N_15194);
and U15313 (N_15313,N_15120,N_15150);
nor U15314 (N_15314,N_15163,N_15183);
xnor U15315 (N_15315,N_15144,N_15069);
and U15316 (N_15316,N_15061,N_15084);
or U15317 (N_15317,N_15088,N_15147);
nand U15318 (N_15318,N_15107,N_15159);
and U15319 (N_15319,N_15049,N_15068);
nand U15320 (N_15320,N_15198,N_15147);
and U15321 (N_15321,N_15116,N_15163);
or U15322 (N_15322,N_15075,N_15125);
nand U15323 (N_15323,N_15118,N_15107);
nand U15324 (N_15324,N_15057,N_15139);
or U15325 (N_15325,N_15189,N_15118);
nand U15326 (N_15326,N_15087,N_15101);
nand U15327 (N_15327,N_15060,N_15162);
or U15328 (N_15328,N_15065,N_15083);
nor U15329 (N_15329,N_15154,N_15134);
and U15330 (N_15330,N_15163,N_15127);
or U15331 (N_15331,N_15169,N_15177);
or U15332 (N_15332,N_15144,N_15119);
or U15333 (N_15333,N_15071,N_15161);
or U15334 (N_15334,N_15138,N_15109);
or U15335 (N_15335,N_15040,N_15140);
nand U15336 (N_15336,N_15080,N_15165);
or U15337 (N_15337,N_15132,N_15169);
or U15338 (N_15338,N_15059,N_15086);
nor U15339 (N_15339,N_15188,N_15094);
or U15340 (N_15340,N_15184,N_15170);
xnor U15341 (N_15341,N_15081,N_15064);
nand U15342 (N_15342,N_15042,N_15054);
or U15343 (N_15343,N_15182,N_15088);
xnor U15344 (N_15344,N_15179,N_15155);
xnor U15345 (N_15345,N_15087,N_15171);
xnor U15346 (N_15346,N_15106,N_15045);
and U15347 (N_15347,N_15163,N_15171);
xnor U15348 (N_15348,N_15111,N_15174);
xor U15349 (N_15349,N_15162,N_15101);
and U15350 (N_15350,N_15067,N_15124);
xnor U15351 (N_15351,N_15193,N_15133);
nor U15352 (N_15352,N_15137,N_15156);
or U15353 (N_15353,N_15170,N_15156);
nand U15354 (N_15354,N_15173,N_15179);
and U15355 (N_15355,N_15123,N_15072);
and U15356 (N_15356,N_15197,N_15170);
nand U15357 (N_15357,N_15181,N_15184);
and U15358 (N_15358,N_15130,N_15154);
or U15359 (N_15359,N_15190,N_15162);
or U15360 (N_15360,N_15262,N_15256);
or U15361 (N_15361,N_15215,N_15313);
and U15362 (N_15362,N_15292,N_15250);
and U15363 (N_15363,N_15279,N_15304);
and U15364 (N_15364,N_15217,N_15223);
xnor U15365 (N_15365,N_15239,N_15246);
and U15366 (N_15366,N_15259,N_15240);
nand U15367 (N_15367,N_15346,N_15334);
or U15368 (N_15368,N_15283,N_15245);
or U15369 (N_15369,N_15332,N_15309);
xor U15370 (N_15370,N_15322,N_15298);
and U15371 (N_15371,N_15242,N_15236);
xor U15372 (N_15372,N_15280,N_15335);
and U15373 (N_15373,N_15251,N_15340);
and U15374 (N_15374,N_15229,N_15318);
nand U15375 (N_15375,N_15349,N_15237);
nor U15376 (N_15376,N_15290,N_15354);
nor U15377 (N_15377,N_15352,N_15338);
xnor U15378 (N_15378,N_15202,N_15265);
xor U15379 (N_15379,N_15268,N_15303);
xor U15380 (N_15380,N_15296,N_15226);
nor U15381 (N_15381,N_15281,N_15321);
and U15382 (N_15382,N_15337,N_15289);
nand U15383 (N_15383,N_15254,N_15211);
nor U15384 (N_15384,N_15266,N_15232);
and U15385 (N_15385,N_15287,N_15359);
nand U15386 (N_15386,N_15231,N_15221);
and U15387 (N_15387,N_15306,N_15307);
nor U15388 (N_15388,N_15234,N_15210);
and U15389 (N_15389,N_15312,N_15314);
nor U15390 (N_15390,N_15324,N_15227);
xnor U15391 (N_15391,N_15285,N_15331);
nand U15392 (N_15392,N_15228,N_15209);
and U15393 (N_15393,N_15342,N_15213);
xor U15394 (N_15394,N_15272,N_15358);
and U15395 (N_15395,N_15276,N_15257);
nor U15396 (N_15396,N_15328,N_15297);
and U15397 (N_15397,N_15219,N_15264);
xnor U15398 (N_15398,N_15244,N_15238);
nor U15399 (N_15399,N_15282,N_15235);
nor U15400 (N_15400,N_15201,N_15295);
nand U15401 (N_15401,N_15300,N_15225);
nor U15402 (N_15402,N_15325,N_15305);
nor U15403 (N_15403,N_15327,N_15208);
and U15404 (N_15404,N_15243,N_15205);
nand U15405 (N_15405,N_15315,N_15271);
and U15406 (N_15406,N_15348,N_15316);
or U15407 (N_15407,N_15347,N_15293);
or U15408 (N_15408,N_15206,N_15339);
and U15409 (N_15409,N_15267,N_15357);
nor U15410 (N_15410,N_15253,N_15356);
and U15411 (N_15411,N_15353,N_15274);
nor U15412 (N_15412,N_15273,N_15269);
and U15413 (N_15413,N_15286,N_15323);
and U15414 (N_15414,N_15222,N_15230);
and U15415 (N_15415,N_15326,N_15345);
or U15416 (N_15416,N_15355,N_15320);
nand U15417 (N_15417,N_15301,N_15329);
and U15418 (N_15418,N_15341,N_15319);
or U15419 (N_15419,N_15220,N_15247);
nand U15420 (N_15420,N_15277,N_15212);
nand U15421 (N_15421,N_15308,N_15233);
nor U15422 (N_15422,N_15311,N_15330);
nor U15423 (N_15423,N_15255,N_15224);
and U15424 (N_15424,N_15284,N_15248);
nand U15425 (N_15425,N_15207,N_15252);
nand U15426 (N_15426,N_15203,N_15263);
and U15427 (N_15427,N_15351,N_15214);
xor U15428 (N_15428,N_15302,N_15275);
xnor U15429 (N_15429,N_15350,N_15249);
and U15430 (N_15430,N_15241,N_15344);
nor U15431 (N_15431,N_15291,N_15333);
and U15432 (N_15432,N_15260,N_15299);
and U15433 (N_15433,N_15294,N_15317);
nand U15434 (N_15434,N_15278,N_15218);
nor U15435 (N_15435,N_15200,N_15288);
and U15436 (N_15436,N_15204,N_15343);
nand U15437 (N_15437,N_15310,N_15270);
nor U15438 (N_15438,N_15216,N_15261);
nand U15439 (N_15439,N_15336,N_15258);
and U15440 (N_15440,N_15250,N_15305);
xnor U15441 (N_15441,N_15261,N_15206);
xnor U15442 (N_15442,N_15282,N_15332);
and U15443 (N_15443,N_15313,N_15201);
xor U15444 (N_15444,N_15230,N_15327);
xnor U15445 (N_15445,N_15280,N_15275);
or U15446 (N_15446,N_15281,N_15332);
nor U15447 (N_15447,N_15208,N_15262);
and U15448 (N_15448,N_15205,N_15253);
nand U15449 (N_15449,N_15323,N_15342);
nand U15450 (N_15450,N_15225,N_15233);
and U15451 (N_15451,N_15333,N_15253);
or U15452 (N_15452,N_15217,N_15312);
or U15453 (N_15453,N_15285,N_15335);
xnor U15454 (N_15454,N_15267,N_15284);
nand U15455 (N_15455,N_15272,N_15277);
nor U15456 (N_15456,N_15317,N_15347);
or U15457 (N_15457,N_15299,N_15342);
and U15458 (N_15458,N_15242,N_15264);
and U15459 (N_15459,N_15296,N_15307);
nand U15460 (N_15460,N_15266,N_15307);
xnor U15461 (N_15461,N_15222,N_15301);
nand U15462 (N_15462,N_15329,N_15230);
nand U15463 (N_15463,N_15300,N_15310);
and U15464 (N_15464,N_15262,N_15316);
nand U15465 (N_15465,N_15205,N_15282);
nand U15466 (N_15466,N_15240,N_15321);
nand U15467 (N_15467,N_15220,N_15286);
and U15468 (N_15468,N_15346,N_15283);
xnor U15469 (N_15469,N_15257,N_15286);
xnor U15470 (N_15470,N_15272,N_15286);
and U15471 (N_15471,N_15255,N_15318);
nor U15472 (N_15472,N_15299,N_15208);
nand U15473 (N_15473,N_15344,N_15231);
nor U15474 (N_15474,N_15209,N_15225);
xor U15475 (N_15475,N_15315,N_15331);
xor U15476 (N_15476,N_15308,N_15247);
xor U15477 (N_15477,N_15244,N_15303);
or U15478 (N_15478,N_15227,N_15213);
and U15479 (N_15479,N_15333,N_15320);
nor U15480 (N_15480,N_15321,N_15216);
and U15481 (N_15481,N_15346,N_15302);
or U15482 (N_15482,N_15279,N_15203);
nor U15483 (N_15483,N_15345,N_15224);
nand U15484 (N_15484,N_15356,N_15282);
xor U15485 (N_15485,N_15280,N_15291);
and U15486 (N_15486,N_15321,N_15244);
and U15487 (N_15487,N_15253,N_15336);
or U15488 (N_15488,N_15282,N_15277);
nand U15489 (N_15489,N_15203,N_15359);
and U15490 (N_15490,N_15321,N_15231);
or U15491 (N_15491,N_15300,N_15343);
and U15492 (N_15492,N_15326,N_15242);
or U15493 (N_15493,N_15235,N_15241);
nand U15494 (N_15494,N_15342,N_15326);
nand U15495 (N_15495,N_15297,N_15220);
and U15496 (N_15496,N_15333,N_15332);
nand U15497 (N_15497,N_15226,N_15340);
xor U15498 (N_15498,N_15344,N_15358);
nand U15499 (N_15499,N_15326,N_15260);
xnor U15500 (N_15500,N_15222,N_15288);
or U15501 (N_15501,N_15342,N_15263);
and U15502 (N_15502,N_15301,N_15247);
nor U15503 (N_15503,N_15325,N_15230);
or U15504 (N_15504,N_15232,N_15252);
and U15505 (N_15505,N_15265,N_15264);
nand U15506 (N_15506,N_15273,N_15282);
or U15507 (N_15507,N_15262,N_15319);
or U15508 (N_15508,N_15270,N_15246);
nor U15509 (N_15509,N_15315,N_15329);
or U15510 (N_15510,N_15259,N_15232);
nor U15511 (N_15511,N_15285,N_15332);
or U15512 (N_15512,N_15298,N_15276);
and U15513 (N_15513,N_15282,N_15227);
and U15514 (N_15514,N_15241,N_15282);
xnor U15515 (N_15515,N_15234,N_15265);
or U15516 (N_15516,N_15220,N_15335);
nor U15517 (N_15517,N_15318,N_15253);
and U15518 (N_15518,N_15290,N_15233);
xnor U15519 (N_15519,N_15336,N_15234);
nor U15520 (N_15520,N_15517,N_15463);
or U15521 (N_15521,N_15475,N_15454);
nor U15522 (N_15522,N_15455,N_15369);
nand U15523 (N_15523,N_15400,N_15484);
xor U15524 (N_15524,N_15456,N_15501);
or U15525 (N_15525,N_15437,N_15424);
and U15526 (N_15526,N_15417,N_15502);
nor U15527 (N_15527,N_15361,N_15490);
and U15528 (N_15528,N_15381,N_15518);
nand U15529 (N_15529,N_15445,N_15494);
nor U15530 (N_15530,N_15393,N_15458);
nand U15531 (N_15531,N_15507,N_15465);
nand U15532 (N_15532,N_15370,N_15396);
or U15533 (N_15533,N_15485,N_15371);
nor U15534 (N_15534,N_15491,N_15479);
or U15535 (N_15535,N_15380,N_15363);
nor U15536 (N_15536,N_15420,N_15449);
nor U15537 (N_15537,N_15433,N_15505);
nand U15538 (N_15538,N_15444,N_15403);
xor U15539 (N_15539,N_15384,N_15441);
nor U15540 (N_15540,N_15476,N_15410);
and U15541 (N_15541,N_15397,N_15429);
xnor U15542 (N_15542,N_15431,N_15452);
nor U15543 (N_15543,N_15503,N_15447);
nand U15544 (N_15544,N_15495,N_15432);
and U15545 (N_15545,N_15385,N_15499);
nand U15546 (N_15546,N_15504,N_15377);
nor U15547 (N_15547,N_15480,N_15478);
xnor U15548 (N_15548,N_15442,N_15440);
nor U15549 (N_15549,N_15481,N_15435);
nand U15550 (N_15550,N_15466,N_15422);
or U15551 (N_15551,N_15434,N_15468);
and U15552 (N_15552,N_15461,N_15487);
or U15553 (N_15553,N_15399,N_15492);
or U15554 (N_15554,N_15473,N_15411);
nand U15555 (N_15555,N_15388,N_15368);
xor U15556 (N_15556,N_15383,N_15394);
or U15557 (N_15557,N_15365,N_15443);
nand U15558 (N_15558,N_15459,N_15419);
or U15559 (N_15559,N_15418,N_15406);
or U15560 (N_15560,N_15413,N_15448);
or U15561 (N_15561,N_15372,N_15460);
and U15562 (N_15562,N_15412,N_15398);
nor U15563 (N_15563,N_15471,N_15438);
nand U15564 (N_15564,N_15405,N_15426);
and U15565 (N_15565,N_15391,N_15428);
or U15566 (N_15566,N_15427,N_15367);
xor U15567 (N_15567,N_15386,N_15477);
xnor U15568 (N_15568,N_15379,N_15416);
or U15569 (N_15569,N_15488,N_15514);
xor U15570 (N_15570,N_15423,N_15404);
nand U15571 (N_15571,N_15390,N_15408);
xor U15572 (N_15572,N_15401,N_15446);
nand U15573 (N_15573,N_15470,N_15414);
xor U15574 (N_15574,N_15421,N_15451);
or U15575 (N_15575,N_15472,N_15506);
or U15576 (N_15576,N_15512,N_15425);
nor U15577 (N_15577,N_15497,N_15374);
xnor U15578 (N_15578,N_15430,N_15389);
nand U15579 (N_15579,N_15469,N_15483);
nor U15580 (N_15580,N_15387,N_15409);
nor U15581 (N_15581,N_15496,N_15407);
nand U15582 (N_15582,N_15415,N_15366);
xnor U15583 (N_15583,N_15515,N_15486);
xor U15584 (N_15584,N_15402,N_15382);
xor U15585 (N_15585,N_15453,N_15464);
nand U15586 (N_15586,N_15519,N_15509);
or U15587 (N_15587,N_15457,N_15436);
or U15588 (N_15588,N_15362,N_15508);
xnor U15589 (N_15589,N_15395,N_15439);
and U15590 (N_15590,N_15500,N_15376);
or U15591 (N_15591,N_15364,N_15467);
or U15592 (N_15592,N_15489,N_15493);
and U15593 (N_15593,N_15513,N_15375);
or U15594 (N_15594,N_15373,N_15450);
and U15595 (N_15595,N_15498,N_15510);
nor U15596 (N_15596,N_15378,N_15360);
xnor U15597 (N_15597,N_15392,N_15474);
or U15598 (N_15598,N_15482,N_15462);
nor U15599 (N_15599,N_15511,N_15516);
nor U15600 (N_15600,N_15394,N_15380);
xnor U15601 (N_15601,N_15495,N_15374);
nand U15602 (N_15602,N_15377,N_15364);
xnor U15603 (N_15603,N_15502,N_15410);
and U15604 (N_15604,N_15470,N_15475);
nand U15605 (N_15605,N_15509,N_15393);
xnor U15606 (N_15606,N_15424,N_15377);
xnor U15607 (N_15607,N_15431,N_15480);
and U15608 (N_15608,N_15512,N_15456);
nor U15609 (N_15609,N_15468,N_15395);
nand U15610 (N_15610,N_15495,N_15491);
nor U15611 (N_15611,N_15404,N_15431);
nand U15612 (N_15612,N_15400,N_15469);
xnor U15613 (N_15613,N_15502,N_15464);
nand U15614 (N_15614,N_15400,N_15428);
or U15615 (N_15615,N_15492,N_15388);
xor U15616 (N_15616,N_15374,N_15506);
xnor U15617 (N_15617,N_15425,N_15459);
nand U15618 (N_15618,N_15404,N_15506);
nor U15619 (N_15619,N_15365,N_15471);
xor U15620 (N_15620,N_15452,N_15511);
nor U15621 (N_15621,N_15480,N_15500);
or U15622 (N_15622,N_15433,N_15517);
xnor U15623 (N_15623,N_15390,N_15436);
nor U15624 (N_15624,N_15366,N_15488);
or U15625 (N_15625,N_15496,N_15458);
nand U15626 (N_15626,N_15412,N_15467);
nor U15627 (N_15627,N_15434,N_15507);
nor U15628 (N_15628,N_15377,N_15510);
nand U15629 (N_15629,N_15511,N_15486);
or U15630 (N_15630,N_15519,N_15388);
nand U15631 (N_15631,N_15476,N_15370);
nand U15632 (N_15632,N_15457,N_15508);
xnor U15633 (N_15633,N_15457,N_15500);
or U15634 (N_15634,N_15462,N_15505);
xnor U15635 (N_15635,N_15512,N_15488);
nor U15636 (N_15636,N_15383,N_15411);
and U15637 (N_15637,N_15405,N_15486);
xor U15638 (N_15638,N_15442,N_15368);
or U15639 (N_15639,N_15367,N_15360);
and U15640 (N_15640,N_15400,N_15361);
or U15641 (N_15641,N_15400,N_15480);
and U15642 (N_15642,N_15508,N_15444);
or U15643 (N_15643,N_15467,N_15450);
xnor U15644 (N_15644,N_15513,N_15509);
nand U15645 (N_15645,N_15503,N_15470);
xor U15646 (N_15646,N_15370,N_15428);
or U15647 (N_15647,N_15463,N_15381);
and U15648 (N_15648,N_15400,N_15451);
nand U15649 (N_15649,N_15439,N_15385);
and U15650 (N_15650,N_15487,N_15374);
and U15651 (N_15651,N_15448,N_15441);
nand U15652 (N_15652,N_15404,N_15500);
or U15653 (N_15653,N_15414,N_15399);
or U15654 (N_15654,N_15417,N_15485);
nor U15655 (N_15655,N_15495,N_15510);
nand U15656 (N_15656,N_15509,N_15421);
nand U15657 (N_15657,N_15430,N_15455);
or U15658 (N_15658,N_15497,N_15380);
nor U15659 (N_15659,N_15481,N_15510);
xnor U15660 (N_15660,N_15425,N_15489);
and U15661 (N_15661,N_15425,N_15430);
xor U15662 (N_15662,N_15410,N_15499);
xnor U15663 (N_15663,N_15498,N_15387);
nor U15664 (N_15664,N_15502,N_15375);
nor U15665 (N_15665,N_15493,N_15492);
and U15666 (N_15666,N_15377,N_15410);
nor U15667 (N_15667,N_15449,N_15372);
nor U15668 (N_15668,N_15498,N_15379);
and U15669 (N_15669,N_15446,N_15501);
or U15670 (N_15670,N_15427,N_15447);
or U15671 (N_15671,N_15381,N_15435);
nor U15672 (N_15672,N_15425,N_15422);
xnor U15673 (N_15673,N_15437,N_15447);
xnor U15674 (N_15674,N_15461,N_15399);
and U15675 (N_15675,N_15438,N_15364);
xnor U15676 (N_15676,N_15381,N_15493);
xnor U15677 (N_15677,N_15498,N_15469);
nor U15678 (N_15678,N_15463,N_15441);
or U15679 (N_15679,N_15425,N_15409);
or U15680 (N_15680,N_15621,N_15678);
xor U15681 (N_15681,N_15565,N_15661);
nand U15682 (N_15682,N_15617,N_15526);
or U15683 (N_15683,N_15559,N_15638);
xnor U15684 (N_15684,N_15572,N_15564);
nor U15685 (N_15685,N_15532,N_15555);
nor U15686 (N_15686,N_15580,N_15541);
nand U15687 (N_15687,N_15651,N_15607);
nor U15688 (N_15688,N_15569,N_15627);
or U15689 (N_15689,N_15533,N_15552);
xnor U15690 (N_15690,N_15535,N_15579);
xnor U15691 (N_15691,N_15608,N_15528);
xor U15692 (N_15692,N_15645,N_15657);
or U15693 (N_15693,N_15522,N_15563);
nor U15694 (N_15694,N_15566,N_15647);
nor U15695 (N_15695,N_15521,N_15643);
or U15696 (N_15696,N_15656,N_15570);
xnor U15697 (N_15697,N_15574,N_15663);
nand U15698 (N_15698,N_15641,N_15586);
nand U15699 (N_15699,N_15665,N_15612);
xor U15700 (N_15700,N_15644,N_15675);
nand U15701 (N_15701,N_15615,N_15666);
xnor U15702 (N_15702,N_15536,N_15640);
xor U15703 (N_15703,N_15662,N_15573);
xor U15704 (N_15704,N_15576,N_15674);
and U15705 (N_15705,N_15525,N_15589);
and U15706 (N_15706,N_15670,N_15567);
and U15707 (N_15707,N_15628,N_15537);
and U15708 (N_15708,N_15629,N_15613);
nor U15709 (N_15709,N_15568,N_15637);
nor U15710 (N_15710,N_15530,N_15591);
and U15711 (N_15711,N_15616,N_15560);
nand U15712 (N_15712,N_15543,N_15545);
nor U15713 (N_15713,N_15550,N_15600);
nor U15714 (N_15714,N_15659,N_15658);
and U15715 (N_15715,N_15578,N_15587);
and U15716 (N_15716,N_15588,N_15634);
or U15717 (N_15717,N_15646,N_15603);
xor U15718 (N_15718,N_15606,N_15624);
xor U15719 (N_15719,N_15581,N_15648);
xor U15720 (N_15720,N_15632,N_15553);
xnor U15721 (N_15721,N_15664,N_15677);
and U15722 (N_15722,N_15575,N_15676);
xnor U15723 (N_15723,N_15554,N_15672);
and U15724 (N_15724,N_15660,N_15626);
nand U15725 (N_15725,N_15538,N_15642);
and U15726 (N_15726,N_15625,N_15611);
and U15727 (N_15727,N_15601,N_15679);
xor U15728 (N_15728,N_15546,N_15618);
or U15729 (N_15729,N_15653,N_15619);
nor U15730 (N_15730,N_15620,N_15649);
nor U15731 (N_15731,N_15597,N_15549);
nor U15732 (N_15732,N_15585,N_15520);
or U15733 (N_15733,N_15547,N_15594);
or U15734 (N_15734,N_15650,N_15595);
or U15735 (N_15735,N_15584,N_15668);
nand U15736 (N_15736,N_15652,N_15605);
and U15737 (N_15737,N_15673,N_15635);
xnor U15738 (N_15738,N_15654,N_15639);
or U15739 (N_15739,N_15540,N_15599);
nand U15740 (N_15740,N_15557,N_15614);
or U15741 (N_15741,N_15582,N_15539);
or U15742 (N_15742,N_15669,N_15523);
and U15743 (N_15743,N_15542,N_15630);
or U15744 (N_15744,N_15577,N_15610);
xnor U15745 (N_15745,N_15527,N_15531);
nor U15746 (N_15746,N_15529,N_15556);
nand U15747 (N_15747,N_15623,N_15604);
and U15748 (N_15748,N_15562,N_15524);
xnor U15749 (N_15749,N_15667,N_15534);
and U15750 (N_15750,N_15622,N_15655);
or U15751 (N_15751,N_15590,N_15583);
nand U15752 (N_15752,N_15592,N_15631);
or U15753 (N_15753,N_15544,N_15551);
nor U15754 (N_15754,N_15602,N_15593);
and U15755 (N_15755,N_15633,N_15596);
nor U15756 (N_15756,N_15636,N_15561);
nor U15757 (N_15757,N_15548,N_15558);
or U15758 (N_15758,N_15609,N_15571);
nor U15759 (N_15759,N_15598,N_15671);
and U15760 (N_15760,N_15582,N_15547);
nand U15761 (N_15761,N_15616,N_15569);
or U15762 (N_15762,N_15545,N_15523);
nand U15763 (N_15763,N_15641,N_15564);
and U15764 (N_15764,N_15619,N_15522);
nand U15765 (N_15765,N_15652,N_15574);
nand U15766 (N_15766,N_15532,N_15542);
or U15767 (N_15767,N_15548,N_15619);
xnor U15768 (N_15768,N_15623,N_15597);
nand U15769 (N_15769,N_15561,N_15584);
nand U15770 (N_15770,N_15539,N_15558);
or U15771 (N_15771,N_15542,N_15565);
nor U15772 (N_15772,N_15601,N_15540);
and U15773 (N_15773,N_15664,N_15536);
and U15774 (N_15774,N_15592,N_15563);
or U15775 (N_15775,N_15673,N_15611);
nor U15776 (N_15776,N_15581,N_15591);
nand U15777 (N_15777,N_15618,N_15641);
nor U15778 (N_15778,N_15594,N_15584);
and U15779 (N_15779,N_15542,N_15535);
nand U15780 (N_15780,N_15524,N_15560);
and U15781 (N_15781,N_15556,N_15563);
nor U15782 (N_15782,N_15543,N_15567);
xnor U15783 (N_15783,N_15546,N_15572);
xor U15784 (N_15784,N_15658,N_15534);
xor U15785 (N_15785,N_15538,N_15639);
nor U15786 (N_15786,N_15533,N_15565);
nor U15787 (N_15787,N_15584,N_15537);
nand U15788 (N_15788,N_15665,N_15557);
nand U15789 (N_15789,N_15662,N_15611);
xnor U15790 (N_15790,N_15615,N_15550);
and U15791 (N_15791,N_15531,N_15538);
nor U15792 (N_15792,N_15571,N_15561);
or U15793 (N_15793,N_15660,N_15553);
or U15794 (N_15794,N_15595,N_15549);
and U15795 (N_15795,N_15528,N_15606);
and U15796 (N_15796,N_15654,N_15595);
nor U15797 (N_15797,N_15597,N_15578);
and U15798 (N_15798,N_15556,N_15655);
xor U15799 (N_15799,N_15674,N_15616);
or U15800 (N_15800,N_15523,N_15636);
or U15801 (N_15801,N_15543,N_15523);
or U15802 (N_15802,N_15662,N_15560);
and U15803 (N_15803,N_15591,N_15656);
nor U15804 (N_15804,N_15561,N_15580);
nor U15805 (N_15805,N_15581,N_15547);
xnor U15806 (N_15806,N_15596,N_15557);
and U15807 (N_15807,N_15576,N_15548);
xor U15808 (N_15808,N_15529,N_15543);
xnor U15809 (N_15809,N_15639,N_15602);
nor U15810 (N_15810,N_15598,N_15674);
and U15811 (N_15811,N_15669,N_15633);
and U15812 (N_15812,N_15565,N_15600);
and U15813 (N_15813,N_15643,N_15564);
nand U15814 (N_15814,N_15538,N_15615);
xnor U15815 (N_15815,N_15532,N_15585);
or U15816 (N_15816,N_15654,N_15619);
or U15817 (N_15817,N_15558,N_15643);
nand U15818 (N_15818,N_15567,N_15557);
or U15819 (N_15819,N_15671,N_15584);
or U15820 (N_15820,N_15654,N_15588);
and U15821 (N_15821,N_15653,N_15548);
xnor U15822 (N_15822,N_15582,N_15524);
and U15823 (N_15823,N_15534,N_15574);
xnor U15824 (N_15824,N_15550,N_15575);
and U15825 (N_15825,N_15678,N_15578);
and U15826 (N_15826,N_15621,N_15666);
xor U15827 (N_15827,N_15538,N_15590);
xor U15828 (N_15828,N_15559,N_15587);
nor U15829 (N_15829,N_15598,N_15544);
or U15830 (N_15830,N_15615,N_15654);
nand U15831 (N_15831,N_15539,N_15670);
and U15832 (N_15832,N_15544,N_15646);
nor U15833 (N_15833,N_15525,N_15532);
and U15834 (N_15834,N_15559,N_15660);
or U15835 (N_15835,N_15667,N_15604);
xor U15836 (N_15836,N_15659,N_15590);
and U15837 (N_15837,N_15619,N_15671);
nor U15838 (N_15838,N_15580,N_15556);
xor U15839 (N_15839,N_15578,N_15533);
or U15840 (N_15840,N_15726,N_15757);
and U15841 (N_15841,N_15728,N_15836);
nand U15842 (N_15842,N_15704,N_15787);
or U15843 (N_15843,N_15750,N_15753);
nand U15844 (N_15844,N_15737,N_15703);
nor U15845 (N_15845,N_15797,N_15738);
nand U15846 (N_15846,N_15803,N_15721);
nor U15847 (N_15847,N_15835,N_15762);
nand U15848 (N_15848,N_15786,N_15814);
xnor U15849 (N_15849,N_15820,N_15724);
or U15850 (N_15850,N_15832,N_15815);
nand U15851 (N_15851,N_15816,N_15794);
and U15852 (N_15852,N_15740,N_15791);
or U15853 (N_15853,N_15772,N_15811);
and U15854 (N_15854,N_15729,N_15717);
xnor U15855 (N_15855,N_15807,N_15690);
nand U15856 (N_15856,N_15756,N_15776);
nor U15857 (N_15857,N_15681,N_15779);
xor U15858 (N_15858,N_15693,N_15705);
and U15859 (N_15859,N_15793,N_15680);
nand U15860 (N_15860,N_15831,N_15801);
or U15861 (N_15861,N_15698,N_15798);
nand U15862 (N_15862,N_15769,N_15819);
nor U15863 (N_15863,N_15701,N_15829);
nor U15864 (N_15864,N_15833,N_15805);
nand U15865 (N_15865,N_15684,N_15800);
xnor U15866 (N_15866,N_15700,N_15747);
nor U15867 (N_15867,N_15808,N_15763);
and U15868 (N_15868,N_15768,N_15839);
or U15869 (N_15869,N_15742,N_15720);
xor U15870 (N_15870,N_15727,N_15773);
or U15871 (N_15871,N_15716,N_15739);
nor U15872 (N_15872,N_15696,N_15709);
xnor U15873 (N_15873,N_15743,N_15688);
and U15874 (N_15874,N_15777,N_15706);
and U15875 (N_15875,N_15837,N_15691);
or U15876 (N_15876,N_15695,N_15802);
nand U15877 (N_15877,N_15766,N_15722);
nand U15878 (N_15878,N_15780,N_15751);
nand U15879 (N_15879,N_15785,N_15817);
and U15880 (N_15880,N_15775,N_15749);
nand U15881 (N_15881,N_15760,N_15730);
and U15882 (N_15882,N_15710,N_15697);
nand U15883 (N_15883,N_15685,N_15744);
xor U15884 (N_15884,N_15723,N_15838);
nand U15885 (N_15885,N_15788,N_15782);
nand U15886 (N_15886,N_15699,N_15795);
nor U15887 (N_15887,N_15790,N_15733);
nor U15888 (N_15888,N_15748,N_15821);
nor U15889 (N_15889,N_15799,N_15809);
xnor U15890 (N_15890,N_15810,N_15687);
nor U15891 (N_15891,N_15765,N_15735);
or U15892 (N_15892,N_15824,N_15746);
and U15893 (N_15893,N_15764,N_15731);
and U15894 (N_15894,N_15745,N_15796);
nand U15895 (N_15895,N_15767,N_15774);
or U15896 (N_15896,N_15758,N_15683);
nor U15897 (N_15897,N_15686,N_15713);
nor U15898 (N_15898,N_15718,N_15781);
and U15899 (N_15899,N_15812,N_15759);
or U15900 (N_15900,N_15828,N_15792);
nor U15901 (N_15901,N_15830,N_15725);
and U15902 (N_15902,N_15694,N_15714);
nor U15903 (N_15903,N_15754,N_15778);
or U15904 (N_15904,N_15818,N_15827);
nand U15905 (N_15905,N_15719,N_15804);
nor U15906 (N_15906,N_15692,N_15736);
nand U15907 (N_15907,N_15682,N_15732);
or U15908 (N_15908,N_15823,N_15771);
and U15909 (N_15909,N_15755,N_15834);
nand U15910 (N_15910,N_15813,N_15789);
xnor U15911 (N_15911,N_15734,N_15825);
and U15912 (N_15912,N_15711,N_15712);
nand U15913 (N_15913,N_15741,N_15708);
nor U15914 (N_15914,N_15806,N_15702);
nand U15915 (N_15915,N_15784,N_15689);
nor U15916 (N_15916,N_15761,N_15783);
nor U15917 (N_15917,N_15707,N_15752);
or U15918 (N_15918,N_15770,N_15826);
nand U15919 (N_15919,N_15822,N_15715);
xnor U15920 (N_15920,N_15773,N_15726);
and U15921 (N_15921,N_15811,N_15733);
or U15922 (N_15922,N_15826,N_15716);
xor U15923 (N_15923,N_15754,N_15796);
nor U15924 (N_15924,N_15782,N_15743);
xnor U15925 (N_15925,N_15694,N_15826);
xnor U15926 (N_15926,N_15821,N_15722);
xnor U15927 (N_15927,N_15759,N_15696);
xor U15928 (N_15928,N_15813,N_15827);
or U15929 (N_15929,N_15800,N_15802);
nor U15930 (N_15930,N_15756,N_15780);
xnor U15931 (N_15931,N_15765,N_15734);
xnor U15932 (N_15932,N_15760,N_15805);
and U15933 (N_15933,N_15682,N_15683);
nand U15934 (N_15934,N_15836,N_15734);
nand U15935 (N_15935,N_15707,N_15768);
nand U15936 (N_15936,N_15731,N_15692);
or U15937 (N_15937,N_15696,N_15745);
and U15938 (N_15938,N_15700,N_15838);
and U15939 (N_15939,N_15727,N_15787);
xnor U15940 (N_15940,N_15690,N_15687);
nand U15941 (N_15941,N_15759,N_15684);
and U15942 (N_15942,N_15820,N_15803);
xnor U15943 (N_15943,N_15752,N_15787);
and U15944 (N_15944,N_15763,N_15735);
nand U15945 (N_15945,N_15680,N_15697);
nand U15946 (N_15946,N_15794,N_15724);
nor U15947 (N_15947,N_15757,N_15833);
and U15948 (N_15948,N_15745,N_15819);
or U15949 (N_15949,N_15729,N_15715);
or U15950 (N_15950,N_15781,N_15711);
or U15951 (N_15951,N_15768,N_15752);
nor U15952 (N_15952,N_15764,N_15797);
nand U15953 (N_15953,N_15806,N_15696);
xor U15954 (N_15954,N_15740,N_15821);
xor U15955 (N_15955,N_15681,N_15796);
nor U15956 (N_15956,N_15802,N_15764);
or U15957 (N_15957,N_15738,N_15707);
and U15958 (N_15958,N_15709,N_15839);
and U15959 (N_15959,N_15696,N_15747);
nand U15960 (N_15960,N_15710,N_15824);
nand U15961 (N_15961,N_15796,N_15763);
nor U15962 (N_15962,N_15705,N_15740);
or U15963 (N_15963,N_15696,N_15804);
nor U15964 (N_15964,N_15777,N_15753);
nand U15965 (N_15965,N_15792,N_15736);
and U15966 (N_15966,N_15813,N_15791);
or U15967 (N_15967,N_15752,N_15749);
nand U15968 (N_15968,N_15782,N_15756);
nand U15969 (N_15969,N_15825,N_15839);
or U15970 (N_15970,N_15695,N_15826);
or U15971 (N_15971,N_15755,N_15734);
nand U15972 (N_15972,N_15697,N_15797);
nor U15973 (N_15973,N_15690,N_15781);
xor U15974 (N_15974,N_15785,N_15686);
or U15975 (N_15975,N_15715,N_15821);
nand U15976 (N_15976,N_15732,N_15822);
xor U15977 (N_15977,N_15775,N_15709);
nand U15978 (N_15978,N_15808,N_15742);
nor U15979 (N_15979,N_15721,N_15766);
xnor U15980 (N_15980,N_15746,N_15779);
and U15981 (N_15981,N_15793,N_15694);
nand U15982 (N_15982,N_15741,N_15709);
nor U15983 (N_15983,N_15696,N_15760);
xor U15984 (N_15984,N_15686,N_15720);
nand U15985 (N_15985,N_15729,N_15838);
or U15986 (N_15986,N_15728,N_15839);
and U15987 (N_15987,N_15729,N_15692);
and U15988 (N_15988,N_15751,N_15826);
or U15989 (N_15989,N_15686,N_15784);
xnor U15990 (N_15990,N_15725,N_15702);
or U15991 (N_15991,N_15761,N_15682);
nor U15992 (N_15992,N_15685,N_15727);
nand U15993 (N_15993,N_15783,N_15833);
xnor U15994 (N_15994,N_15725,N_15752);
nand U15995 (N_15995,N_15714,N_15808);
and U15996 (N_15996,N_15732,N_15685);
and U15997 (N_15997,N_15730,N_15778);
and U15998 (N_15998,N_15809,N_15725);
and U15999 (N_15999,N_15818,N_15725);
nand U16000 (N_16000,N_15971,N_15859);
xor U16001 (N_16001,N_15878,N_15979);
or U16002 (N_16002,N_15886,N_15923);
nand U16003 (N_16003,N_15911,N_15938);
and U16004 (N_16004,N_15847,N_15933);
xnor U16005 (N_16005,N_15887,N_15898);
nor U16006 (N_16006,N_15922,N_15928);
and U16007 (N_16007,N_15927,N_15947);
nand U16008 (N_16008,N_15858,N_15953);
xor U16009 (N_16009,N_15891,N_15934);
xor U16010 (N_16010,N_15875,N_15966);
and U16011 (N_16011,N_15910,N_15957);
xnor U16012 (N_16012,N_15991,N_15860);
nand U16013 (N_16013,N_15980,N_15985);
nand U16014 (N_16014,N_15855,N_15944);
xor U16015 (N_16015,N_15879,N_15972);
or U16016 (N_16016,N_15975,N_15955);
and U16017 (N_16017,N_15941,N_15948);
and U16018 (N_16018,N_15899,N_15998);
xor U16019 (N_16019,N_15849,N_15988);
or U16020 (N_16020,N_15907,N_15930);
nor U16021 (N_16021,N_15962,N_15937);
and U16022 (N_16022,N_15864,N_15936);
and U16023 (N_16023,N_15963,N_15908);
xnor U16024 (N_16024,N_15973,N_15935);
xnor U16025 (N_16025,N_15882,N_15968);
nand U16026 (N_16026,N_15904,N_15909);
and U16027 (N_16027,N_15854,N_15977);
nor U16028 (N_16028,N_15892,N_15844);
and U16029 (N_16029,N_15964,N_15919);
xor U16030 (N_16030,N_15984,N_15969);
or U16031 (N_16031,N_15913,N_15895);
or U16032 (N_16032,N_15863,N_15999);
and U16033 (N_16033,N_15992,N_15850);
and U16034 (N_16034,N_15884,N_15869);
nor U16035 (N_16035,N_15874,N_15906);
or U16036 (N_16036,N_15961,N_15918);
nand U16037 (N_16037,N_15921,N_15896);
xor U16038 (N_16038,N_15959,N_15940);
nand U16039 (N_16039,N_15877,N_15945);
nor U16040 (N_16040,N_15856,N_15853);
or U16041 (N_16041,N_15981,N_15926);
and U16042 (N_16042,N_15932,N_15956);
or U16043 (N_16043,N_15931,N_15846);
nor U16044 (N_16044,N_15916,N_15986);
xnor U16045 (N_16045,N_15840,N_15857);
nand U16046 (N_16046,N_15870,N_15845);
xnor U16047 (N_16047,N_15867,N_15917);
xor U16048 (N_16048,N_15897,N_15866);
and U16049 (N_16049,N_15880,N_15996);
and U16050 (N_16050,N_15976,N_15946);
and U16051 (N_16051,N_15894,N_15842);
and U16052 (N_16052,N_15861,N_15920);
xnor U16053 (N_16053,N_15905,N_15997);
or U16054 (N_16054,N_15943,N_15868);
nand U16055 (N_16055,N_15862,N_15843);
xnor U16056 (N_16056,N_15983,N_15974);
or U16057 (N_16057,N_15889,N_15924);
and U16058 (N_16058,N_15939,N_15888);
xnor U16059 (N_16059,N_15912,N_15967);
nand U16060 (N_16060,N_15987,N_15851);
nor U16061 (N_16061,N_15970,N_15965);
nor U16062 (N_16062,N_15990,N_15978);
nand U16063 (N_16063,N_15883,N_15929);
nand U16064 (N_16064,N_15942,N_15901);
xnor U16065 (N_16065,N_15841,N_15865);
or U16066 (N_16066,N_15951,N_15993);
or U16067 (N_16067,N_15925,N_15989);
and U16068 (N_16068,N_15994,N_15995);
or U16069 (N_16069,N_15873,N_15890);
nor U16070 (N_16070,N_15902,N_15954);
nor U16071 (N_16071,N_15893,N_15982);
and U16072 (N_16072,N_15952,N_15871);
or U16073 (N_16073,N_15900,N_15960);
or U16074 (N_16074,N_15848,N_15958);
xor U16075 (N_16075,N_15872,N_15949);
nor U16076 (N_16076,N_15950,N_15914);
nand U16077 (N_16077,N_15903,N_15915);
xor U16078 (N_16078,N_15881,N_15876);
or U16079 (N_16079,N_15852,N_15885);
or U16080 (N_16080,N_15851,N_15877);
and U16081 (N_16081,N_15956,N_15928);
xor U16082 (N_16082,N_15895,N_15925);
and U16083 (N_16083,N_15851,N_15938);
and U16084 (N_16084,N_15984,N_15891);
and U16085 (N_16085,N_15845,N_15862);
or U16086 (N_16086,N_15893,N_15937);
and U16087 (N_16087,N_15845,N_15877);
or U16088 (N_16088,N_15981,N_15955);
xor U16089 (N_16089,N_15850,N_15883);
nand U16090 (N_16090,N_15871,N_15969);
and U16091 (N_16091,N_15935,N_15862);
xor U16092 (N_16092,N_15992,N_15971);
nor U16093 (N_16093,N_15870,N_15923);
or U16094 (N_16094,N_15857,N_15916);
xnor U16095 (N_16095,N_15911,N_15883);
xor U16096 (N_16096,N_15939,N_15949);
xnor U16097 (N_16097,N_15981,N_15903);
and U16098 (N_16098,N_15884,N_15982);
xnor U16099 (N_16099,N_15954,N_15844);
nor U16100 (N_16100,N_15991,N_15908);
or U16101 (N_16101,N_15947,N_15890);
nor U16102 (N_16102,N_15846,N_15938);
nand U16103 (N_16103,N_15927,N_15940);
nor U16104 (N_16104,N_15957,N_15893);
xnor U16105 (N_16105,N_15946,N_15874);
nand U16106 (N_16106,N_15887,N_15980);
xnor U16107 (N_16107,N_15895,N_15926);
xor U16108 (N_16108,N_15859,N_15946);
or U16109 (N_16109,N_15976,N_15989);
and U16110 (N_16110,N_15967,N_15930);
nand U16111 (N_16111,N_15922,N_15997);
and U16112 (N_16112,N_15962,N_15952);
nor U16113 (N_16113,N_15979,N_15946);
nor U16114 (N_16114,N_15876,N_15918);
xnor U16115 (N_16115,N_15846,N_15890);
nand U16116 (N_16116,N_15892,N_15942);
and U16117 (N_16117,N_15893,N_15967);
or U16118 (N_16118,N_15924,N_15941);
nor U16119 (N_16119,N_15862,N_15983);
xnor U16120 (N_16120,N_15994,N_15899);
nand U16121 (N_16121,N_15850,N_15948);
nor U16122 (N_16122,N_15865,N_15848);
xor U16123 (N_16123,N_15997,N_15902);
nand U16124 (N_16124,N_15917,N_15986);
nand U16125 (N_16125,N_15942,N_15957);
or U16126 (N_16126,N_15942,N_15927);
or U16127 (N_16127,N_15864,N_15861);
and U16128 (N_16128,N_15916,N_15977);
nor U16129 (N_16129,N_15974,N_15958);
nand U16130 (N_16130,N_15971,N_15878);
xnor U16131 (N_16131,N_15947,N_15939);
nor U16132 (N_16132,N_15917,N_15909);
xor U16133 (N_16133,N_15941,N_15896);
or U16134 (N_16134,N_15842,N_15923);
or U16135 (N_16135,N_15922,N_15906);
and U16136 (N_16136,N_15969,N_15950);
or U16137 (N_16137,N_15864,N_15955);
xnor U16138 (N_16138,N_15981,N_15927);
nor U16139 (N_16139,N_15847,N_15870);
nor U16140 (N_16140,N_15960,N_15987);
xor U16141 (N_16141,N_15890,N_15877);
nor U16142 (N_16142,N_15877,N_15924);
xor U16143 (N_16143,N_15861,N_15992);
nor U16144 (N_16144,N_15934,N_15995);
xnor U16145 (N_16145,N_15849,N_15923);
xor U16146 (N_16146,N_15866,N_15965);
nor U16147 (N_16147,N_15866,N_15893);
nor U16148 (N_16148,N_15973,N_15840);
nor U16149 (N_16149,N_15871,N_15981);
or U16150 (N_16150,N_15939,N_15883);
xor U16151 (N_16151,N_15967,N_15868);
and U16152 (N_16152,N_15918,N_15962);
xor U16153 (N_16153,N_15970,N_15987);
and U16154 (N_16154,N_15878,N_15955);
and U16155 (N_16155,N_15848,N_15920);
xor U16156 (N_16156,N_15899,N_15960);
or U16157 (N_16157,N_15916,N_15979);
nand U16158 (N_16158,N_15881,N_15979);
nor U16159 (N_16159,N_15999,N_15851);
and U16160 (N_16160,N_16018,N_16121);
nand U16161 (N_16161,N_16142,N_16074);
nand U16162 (N_16162,N_16109,N_16032);
xnor U16163 (N_16163,N_16051,N_16122);
nand U16164 (N_16164,N_16103,N_16105);
and U16165 (N_16165,N_16143,N_16148);
or U16166 (N_16166,N_16128,N_16083);
xnor U16167 (N_16167,N_16067,N_16155);
xor U16168 (N_16168,N_16088,N_16002);
nor U16169 (N_16169,N_16138,N_16078);
and U16170 (N_16170,N_16059,N_16035);
xor U16171 (N_16171,N_16039,N_16118);
or U16172 (N_16172,N_16011,N_16094);
xor U16173 (N_16173,N_16098,N_16144);
or U16174 (N_16174,N_16130,N_16045);
nand U16175 (N_16175,N_16093,N_16038);
xor U16176 (N_16176,N_16071,N_16006);
xor U16177 (N_16177,N_16020,N_16111);
nor U16178 (N_16178,N_16022,N_16120);
or U16179 (N_16179,N_16115,N_16087);
nand U16180 (N_16180,N_16086,N_16021);
and U16181 (N_16181,N_16063,N_16053);
nor U16182 (N_16182,N_16146,N_16081);
nor U16183 (N_16183,N_16136,N_16040);
nand U16184 (N_16184,N_16084,N_16131);
and U16185 (N_16185,N_16129,N_16091);
xnor U16186 (N_16186,N_16116,N_16052);
xnor U16187 (N_16187,N_16057,N_16092);
or U16188 (N_16188,N_16062,N_16037);
nand U16189 (N_16189,N_16140,N_16099);
nand U16190 (N_16190,N_16069,N_16080);
xor U16191 (N_16191,N_16077,N_16061);
nand U16192 (N_16192,N_16012,N_16114);
xnor U16193 (N_16193,N_16149,N_16030);
or U16194 (N_16194,N_16075,N_16101);
nand U16195 (N_16195,N_16124,N_16119);
and U16196 (N_16196,N_16023,N_16041);
xor U16197 (N_16197,N_16150,N_16072);
xnor U16198 (N_16198,N_16153,N_16010);
xor U16199 (N_16199,N_16024,N_16090);
nor U16200 (N_16200,N_16089,N_16123);
nor U16201 (N_16201,N_16007,N_16108);
nor U16202 (N_16202,N_16154,N_16019);
and U16203 (N_16203,N_16141,N_16043);
nand U16204 (N_16204,N_16033,N_16147);
nor U16205 (N_16205,N_16009,N_16125);
xor U16206 (N_16206,N_16016,N_16157);
nor U16207 (N_16207,N_16042,N_16046);
xor U16208 (N_16208,N_16017,N_16055);
or U16209 (N_16209,N_16135,N_16049);
or U16210 (N_16210,N_16104,N_16132);
nor U16211 (N_16211,N_16100,N_16028);
nand U16212 (N_16212,N_16003,N_16048);
nor U16213 (N_16213,N_16000,N_16004);
or U16214 (N_16214,N_16079,N_16102);
or U16215 (N_16215,N_16068,N_16076);
xnor U16216 (N_16216,N_16065,N_16034);
or U16217 (N_16217,N_16085,N_16029);
or U16218 (N_16218,N_16073,N_16156);
nand U16219 (N_16219,N_16126,N_16106);
nand U16220 (N_16220,N_16127,N_16152);
nor U16221 (N_16221,N_16133,N_16047);
and U16222 (N_16222,N_16137,N_16064);
nor U16223 (N_16223,N_16096,N_16005);
nor U16224 (N_16224,N_16050,N_16110);
nand U16225 (N_16225,N_16060,N_16014);
and U16226 (N_16226,N_16054,N_16031);
or U16227 (N_16227,N_16015,N_16008);
xnor U16228 (N_16228,N_16058,N_16056);
and U16229 (N_16229,N_16066,N_16112);
nand U16230 (N_16230,N_16113,N_16070);
nor U16231 (N_16231,N_16036,N_16107);
and U16232 (N_16232,N_16044,N_16117);
xor U16233 (N_16233,N_16013,N_16159);
or U16234 (N_16234,N_16151,N_16095);
or U16235 (N_16235,N_16001,N_16145);
xor U16236 (N_16236,N_16097,N_16082);
xnor U16237 (N_16237,N_16134,N_16139);
xor U16238 (N_16238,N_16026,N_16027);
xnor U16239 (N_16239,N_16025,N_16158);
xor U16240 (N_16240,N_16133,N_16018);
xnor U16241 (N_16241,N_16130,N_16099);
nand U16242 (N_16242,N_16041,N_16087);
nor U16243 (N_16243,N_16029,N_16092);
or U16244 (N_16244,N_16149,N_16107);
or U16245 (N_16245,N_16082,N_16137);
and U16246 (N_16246,N_16050,N_16071);
or U16247 (N_16247,N_16122,N_16050);
or U16248 (N_16248,N_16021,N_16074);
xor U16249 (N_16249,N_16022,N_16086);
nor U16250 (N_16250,N_16071,N_16009);
xnor U16251 (N_16251,N_16145,N_16081);
xor U16252 (N_16252,N_16143,N_16067);
xnor U16253 (N_16253,N_16096,N_16136);
or U16254 (N_16254,N_16146,N_16036);
nor U16255 (N_16255,N_16029,N_16025);
nand U16256 (N_16256,N_16146,N_16106);
nand U16257 (N_16257,N_16036,N_16104);
or U16258 (N_16258,N_16159,N_16151);
nand U16259 (N_16259,N_16119,N_16056);
nor U16260 (N_16260,N_16055,N_16073);
or U16261 (N_16261,N_16124,N_16070);
nor U16262 (N_16262,N_16033,N_16140);
and U16263 (N_16263,N_16071,N_16124);
xor U16264 (N_16264,N_16124,N_16004);
nand U16265 (N_16265,N_16114,N_16105);
or U16266 (N_16266,N_16043,N_16089);
or U16267 (N_16267,N_16071,N_16033);
nor U16268 (N_16268,N_16005,N_16021);
xor U16269 (N_16269,N_16003,N_16058);
or U16270 (N_16270,N_16040,N_16127);
and U16271 (N_16271,N_16108,N_16054);
or U16272 (N_16272,N_16004,N_16040);
or U16273 (N_16273,N_16083,N_16013);
nor U16274 (N_16274,N_16067,N_16068);
xor U16275 (N_16275,N_16017,N_16027);
nor U16276 (N_16276,N_16126,N_16031);
nor U16277 (N_16277,N_16002,N_16094);
nand U16278 (N_16278,N_16025,N_16121);
nand U16279 (N_16279,N_16001,N_16156);
or U16280 (N_16280,N_16085,N_16058);
nor U16281 (N_16281,N_16046,N_16018);
nand U16282 (N_16282,N_16071,N_16119);
and U16283 (N_16283,N_16028,N_16149);
nor U16284 (N_16284,N_16074,N_16147);
xor U16285 (N_16285,N_16053,N_16052);
nand U16286 (N_16286,N_16133,N_16041);
and U16287 (N_16287,N_16137,N_16123);
xnor U16288 (N_16288,N_16017,N_16049);
nand U16289 (N_16289,N_16085,N_16010);
nor U16290 (N_16290,N_16136,N_16094);
xnor U16291 (N_16291,N_16112,N_16080);
nand U16292 (N_16292,N_16052,N_16056);
xnor U16293 (N_16293,N_16065,N_16135);
xnor U16294 (N_16294,N_16073,N_16144);
xor U16295 (N_16295,N_16146,N_16128);
nor U16296 (N_16296,N_16034,N_16030);
and U16297 (N_16297,N_16113,N_16065);
or U16298 (N_16298,N_16106,N_16155);
nor U16299 (N_16299,N_16125,N_16035);
or U16300 (N_16300,N_16057,N_16051);
or U16301 (N_16301,N_16158,N_16095);
nor U16302 (N_16302,N_16013,N_16023);
and U16303 (N_16303,N_16142,N_16056);
xnor U16304 (N_16304,N_16036,N_16004);
xor U16305 (N_16305,N_16013,N_16031);
nor U16306 (N_16306,N_16002,N_16068);
or U16307 (N_16307,N_16158,N_16109);
nand U16308 (N_16308,N_16146,N_16100);
and U16309 (N_16309,N_16040,N_16078);
nor U16310 (N_16310,N_16045,N_16108);
nand U16311 (N_16311,N_16027,N_16036);
nand U16312 (N_16312,N_16092,N_16082);
or U16313 (N_16313,N_16023,N_16147);
or U16314 (N_16314,N_16103,N_16009);
and U16315 (N_16315,N_16099,N_16035);
nand U16316 (N_16316,N_16118,N_16123);
and U16317 (N_16317,N_16068,N_16042);
and U16318 (N_16318,N_16151,N_16064);
and U16319 (N_16319,N_16159,N_16148);
xnor U16320 (N_16320,N_16178,N_16312);
xnor U16321 (N_16321,N_16171,N_16295);
or U16322 (N_16322,N_16278,N_16188);
nand U16323 (N_16323,N_16199,N_16283);
xnor U16324 (N_16324,N_16164,N_16166);
nor U16325 (N_16325,N_16204,N_16318);
nand U16326 (N_16326,N_16241,N_16269);
xor U16327 (N_16327,N_16249,N_16177);
or U16328 (N_16328,N_16225,N_16270);
and U16329 (N_16329,N_16265,N_16232);
xor U16330 (N_16330,N_16207,N_16293);
xnor U16331 (N_16331,N_16182,N_16203);
or U16332 (N_16332,N_16253,N_16161);
xor U16333 (N_16333,N_16294,N_16314);
nor U16334 (N_16334,N_16266,N_16217);
and U16335 (N_16335,N_16309,N_16288);
nor U16336 (N_16336,N_16172,N_16272);
nor U16337 (N_16337,N_16317,N_16306);
nor U16338 (N_16338,N_16302,N_16284);
or U16339 (N_16339,N_16206,N_16251);
or U16340 (N_16340,N_16274,N_16300);
or U16341 (N_16341,N_16224,N_16221);
nor U16342 (N_16342,N_16202,N_16313);
or U16343 (N_16343,N_16226,N_16311);
xor U16344 (N_16344,N_16259,N_16299);
nor U16345 (N_16345,N_16303,N_16165);
or U16346 (N_16346,N_16304,N_16200);
or U16347 (N_16347,N_16276,N_16185);
or U16348 (N_16348,N_16210,N_16256);
nor U16349 (N_16349,N_16229,N_16233);
nor U16350 (N_16350,N_16262,N_16192);
and U16351 (N_16351,N_16255,N_16254);
xor U16352 (N_16352,N_16220,N_16286);
and U16353 (N_16353,N_16163,N_16292);
nor U16354 (N_16354,N_16297,N_16277);
nor U16355 (N_16355,N_16205,N_16236);
xor U16356 (N_16356,N_16195,N_16267);
xnor U16357 (N_16357,N_16308,N_16234);
nand U16358 (N_16358,N_16271,N_16168);
xnor U16359 (N_16359,N_16243,N_16216);
and U16360 (N_16360,N_16189,N_16246);
xnor U16361 (N_16361,N_16201,N_16235);
or U16362 (N_16362,N_16307,N_16209);
and U16363 (N_16363,N_16231,N_16175);
nor U16364 (N_16364,N_16298,N_16190);
nand U16365 (N_16365,N_16174,N_16218);
or U16366 (N_16366,N_16227,N_16222);
nand U16367 (N_16367,N_16183,N_16242);
xor U16368 (N_16368,N_16223,N_16211);
and U16369 (N_16369,N_16181,N_16261);
nand U16370 (N_16370,N_16239,N_16310);
nor U16371 (N_16371,N_16169,N_16187);
nand U16372 (N_16372,N_16230,N_16180);
or U16373 (N_16373,N_16287,N_16296);
xnor U16374 (N_16374,N_16252,N_16291);
nand U16375 (N_16375,N_16173,N_16214);
nand U16376 (N_16376,N_16247,N_16319);
and U16377 (N_16377,N_16237,N_16281);
nor U16378 (N_16378,N_16245,N_16279);
or U16379 (N_16379,N_16316,N_16176);
or U16380 (N_16380,N_16264,N_16160);
nand U16381 (N_16381,N_16167,N_16305);
xor U16382 (N_16382,N_16257,N_16250);
nand U16383 (N_16383,N_16198,N_16301);
nand U16384 (N_16384,N_16289,N_16240);
or U16385 (N_16385,N_16248,N_16275);
and U16386 (N_16386,N_16197,N_16258);
nor U16387 (N_16387,N_16282,N_16215);
and U16388 (N_16388,N_16194,N_16170);
and U16389 (N_16389,N_16238,N_16228);
nor U16390 (N_16390,N_16213,N_16179);
nand U16391 (N_16391,N_16244,N_16268);
or U16392 (N_16392,N_16260,N_16193);
and U16393 (N_16393,N_16219,N_16280);
or U16394 (N_16394,N_16285,N_16263);
nor U16395 (N_16395,N_16186,N_16191);
or U16396 (N_16396,N_16208,N_16212);
or U16397 (N_16397,N_16196,N_16315);
xor U16398 (N_16398,N_16184,N_16273);
or U16399 (N_16399,N_16290,N_16162);
nor U16400 (N_16400,N_16254,N_16164);
or U16401 (N_16401,N_16197,N_16216);
nor U16402 (N_16402,N_16302,N_16163);
or U16403 (N_16403,N_16276,N_16190);
xnor U16404 (N_16404,N_16183,N_16307);
nor U16405 (N_16405,N_16200,N_16315);
nor U16406 (N_16406,N_16178,N_16241);
or U16407 (N_16407,N_16178,N_16264);
or U16408 (N_16408,N_16252,N_16225);
or U16409 (N_16409,N_16254,N_16261);
nand U16410 (N_16410,N_16174,N_16318);
nand U16411 (N_16411,N_16314,N_16161);
nand U16412 (N_16412,N_16259,N_16290);
xor U16413 (N_16413,N_16256,N_16204);
xnor U16414 (N_16414,N_16206,N_16196);
xor U16415 (N_16415,N_16238,N_16301);
nor U16416 (N_16416,N_16251,N_16277);
or U16417 (N_16417,N_16271,N_16233);
or U16418 (N_16418,N_16216,N_16303);
xor U16419 (N_16419,N_16175,N_16301);
and U16420 (N_16420,N_16230,N_16266);
and U16421 (N_16421,N_16192,N_16271);
xnor U16422 (N_16422,N_16171,N_16309);
nand U16423 (N_16423,N_16233,N_16269);
nand U16424 (N_16424,N_16227,N_16288);
nor U16425 (N_16425,N_16230,N_16198);
and U16426 (N_16426,N_16179,N_16196);
nand U16427 (N_16427,N_16254,N_16175);
nand U16428 (N_16428,N_16241,N_16167);
nand U16429 (N_16429,N_16299,N_16286);
nand U16430 (N_16430,N_16249,N_16243);
or U16431 (N_16431,N_16190,N_16283);
nand U16432 (N_16432,N_16312,N_16301);
or U16433 (N_16433,N_16237,N_16234);
nand U16434 (N_16434,N_16260,N_16294);
nor U16435 (N_16435,N_16223,N_16183);
or U16436 (N_16436,N_16273,N_16277);
xnor U16437 (N_16437,N_16205,N_16180);
nand U16438 (N_16438,N_16193,N_16187);
nand U16439 (N_16439,N_16302,N_16213);
nor U16440 (N_16440,N_16276,N_16166);
and U16441 (N_16441,N_16200,N_16234);
and U16442 (N_16442,N_16162,N_16217);
nor U16443 (N_16443,N_16254,N_16245);
or U16444 (N_16444,N_16182,N_16318);
xnor U16445 (N_16445,N_16262,N_16309);
nor U16446 (N_16446,N_16270,N_16218);
xor U16447 (N_16447,N_16309,N_16273);
and U16448 (N_16448,N_16270,N_16220);
xnor U16449 (N_16449,N_16206,N_16276);
xor U16450 (N_16450,N_16216,N_16280);
or U16451 (N_16451,N_16292,N_16265);
nor U16452 (N_16452,N_16220,N_16240);
or U16453 (N_16453,N_16188,N_16310);
xnor U16454 (N_16454,N_16161,N_16280);
and U16455 (N_16455,N_16179,N_16278);
or U16456 (N_16456,N_16218,N_16178);
xor U16457 (N_16457,N_16279,N_16210);
or U16458 (N_16458,N_16318,N_16306);
nand U16459 (N_16459,N_16256,N_16207);
xor U16460 (N_16460,N_16192,N_16207);
nand U16461 (N_16461,N_16284,N_16191);
and U16462 (N_16462,N_16276,N_16289);
nor U16463 (N_16463,N_16211,N_16201);
xor U16464 (N_16464,N_16239,N_16164);
or U16465 (N_16465,N_16300,N_16264);
and U16466 (N_16466,N_16238,N_16179);
or U16467 (N_16467,N_16214,N_16250);
xor U16468 (N_16468,N_16218,N_16167);
nor U16469 (N_16469,N_16168,N_16215);
xor U16470 (N_16470,N_16167,N_16273);
or U16471 (N_16471,N_16197,N_16315);
or U16472 (N_16472,N_16179,N_16276);
xor U16473 (N_16473,N_16215,N_16256);
nand U16474 (N_16474,N_16212,N_16292);
or U16475 (N_16475,N_16307,N_16163);
and U16476 (N_16476,N_16201,N_16205);
nand U16477 (N_16477,N_16221,N_16255);
or U16478 (N_16478,N_16226,N_16220);
nor U16479 (N_16479,N_16161,N_16261);
nand U16480 (N_16480,N_16441,N_16370);
xor U16481 (N_16481,N_16390,N_16386);
nand U16482 (N_16482,N_16472,N_16389);
and U16483 (N_16483,N_16430,N_16347);
xnor U16484 (N_16484,N_16443,N_16329);
or U16485 (N_16485,N_16433,N_16331);
xor U16486 (N_16486,N_16341,N_16456);
xnor U16487 (N_16487,N_16431,N_16469);
nor U16488 (N_16488,N_16477,N_16466);
and U16489 (N_16489,N_16320,N_16434);
xnor U16490 (N_16490,N_16412,N_16420);
nor U16491 (N_16491,N_16382,N_16408);
or U16492 (N_16492,N_16337,N_16454);
nor U16493 (N_16493,N_16413,N_16335);
and U16494 (N_16494,N_16416,N_16342);
or U16495 (N_16495,N_16368,N_16395);
and U16496 (N_16496,N_16340,N_16375);
nand U16497 (N_16497,N_16476,N_16378);
or U16498 (N_16498,N_16338,N_16376);
and U16499 (N_16499,N_16424,N_16421);
nand U16500 (N_16500,N_16427,N_16371);
and U16501 (N_16501,N_16381,N_16369);
or U16502 (N_16502,N_16323,N_16377);
nand U16503 (N_16503,N_16478,N_16440);
nor U16504 (N_16504,N_16445,N_16429);
or U16505 (N_16505,N_16460,N_16453);
nand U16506 (N_16506,N_16326,N_16464);
and U16507 (N_16507,N_16438,N_16447);
and U16508 (N_16508,N_16365,N_16327);
or U16509 (N_16509,N_16356,N_16334);
and U16510 (N_16510,N_16388,N_16398);
or U16511 (N_16511,N_16394,N_16468);
nand U16512 (N_16512,N_16372,N_16448);
or U16513 (N_16513,N_16405,N_16392);
and U16514 (N_16514,N_16407,N_16401);
or U16515 (N_16515,N_16459,N_16393);
and U16516 (N_16516,N_16415,N_16345);
nor U16517 (N_16517,N_16364,N_16399);
nor U16518 (N_16518,N_16474,N_16351);
xnor U16519 (N_16519,N_16436,N_16346);
or U16520 (N_16520,N_16452,N_16361);
xnor U16521 (N_16521,N_16339,N_16357);
or U16522 (N_16522,N_16411,N_16348);
and U16523 (N_16523,N_16450,N_16475);
nand U16524 (N_16524,N_16358,N_16462);
nor U16525 (N_16525,N_16330,N_16322);
and U16526 (N_16526,N_16410,N_16359);
xnor U16527 (N_16527,N_16353,N_16402);
and U16528 (N_16528,N_16374,N_16451);
xor U16529 (N_16529,N_16360,N_16373);
xor U16530 (N_16530,N_16355,N_16343);
xnor U16531 (N_16531,N_16344,N_16458);
nor U16532 (N_16532,N_16479,N_16328);
nand U16533 (N_16533,N_16467,N_16414);
nand U16534 (N_16534,N_16422,N_16465);
and U16535 (N_16535,N_16446,N_16367);
or U16536 (N_16536,N_16366,N_16333);
nor U16537 (N_16537,N_16324,N_16417);
and U16538 (N_16538,N_16385,N_16380);
xnor U16539 (N_16539,N_16336,N_16425);
and U16540 (N_16540,N_16432,N_16461);
and U16541 (N_16541,N_16379,N_16406);
nand U16542 (N_16542,N_16349,N_16423);
nand U16543 (N_16543,N_16362,N_16442);
and U16544 (N_16544,N_16384,N_16387);
nor U16545 (N_16545,N_16437,N_16409);
or U16546 (N_16546,N_16473,N_16363);
and U16547 (N_16547,N_16457,N_16400);
nor U16548 (N_16548,N_16396,N_16418);
or U16549 (N_16549,N_16403,N_16428);
nand U16550 (N_16550,N_16444,N_16352);
nor U16551 (N_16551,N_16471,N_16383);
nand U16552 (N_16552,N_16455,N_16350);
xor U16553 (N_16553,N_16419,N_16439);
nand U16554 (N_16554,N_16332,N_16321);
or U16555 (N_16555,N_16391,N_16354);
or U16556 (N_16556,N_16470,N_16397);
or U16557 (N_16557,N_16426,N_16435);
xnor U16558 (N_16558,N_16325,N_16463);
nand U16559 (N_16559,N_16404,N_16449);
nand U16560 (N_16560,N_16420,N_16455);
or U16561 (N_16561,N_16330,N_16339);
or U16562 (N_16562,N_16441,N_16432);
nor U16563 (N_16563,N_16328,N_16437);
and U16564 (N_16564,N_16340,N_16346);
or U16565 (N_16565,N_16473,N_16403);
and U16566 (N_16566,N_16373,N_16362);
nor U16567 (N_16567,N_16332,N_16468);
nand U16568 (N_16568,N_16344,N_16459);
and U16569 (N_16569,N_16428,N_16451);
nor U16570 (N_16570,N_16322,N_16467);
nor U16571 (N_16571,N_16391,N_16392);
nor U16572 (N_16572,N_16475,N_16350);
nand U16573 (N_16573,N_16336,N_16453);
nand U16574 (N_16574,N_16399,N_16458);
and U16575 (N_16575,N_16407,N_16405);
nand U16576 (N_16576,N_16434,N_16360);
and U16577 (N_16577,N_16341,N_16426);
or U16578 (N_16578,N_16423,N_16391);
and U16579 (N_16579,N_16479,N_16385);
and U16580 (N_16580,N_16333,N_16423);
nor U16581 (N_16581,N_16459,N_16366);
nor U16582 (N_16582,N_16431,N_16453);
or U16583 (N_16583,N_16428,N_16463);
xor U16584 (N_16584,N_16459,N_16368);
and U16585 (N_16585,N_16422,N_16472);
or U16586 (N_16586,N_16381,N_16443);
nand U16587 (N_16587,N_16322,N_16394);
xnor U16588 (N_16588,N_16337,N_16347);
nand U16589 (N_16589,N_16452,N_16460);
nor U16590 (N_16590,N_16327,N_16342);
xnor U16591 (N_16591,N_16355,N_16471);
xor U16592 (N_16592,N_16429,N_16418);
or U16593 (N_16593,N_16429,N_16450);
nor U16594 (N_16594,N_16422,N_16448);
nand U16595 (N_16595,N_16475,N_16420);
nand U16596 (N_16596,N_16479,N_16339);
and U16597 (N_16597,N_16356,N_16427);
or U16598 (N_16598,N_16422,N_16434);
and U16599 (N_16599,N_16460,N_16464);
or U16600 (N_16600,N_16463,N_16339);
or U16601 (N_16601,N_16433,N_16458);
or U16602 (N_16602,N_16391,N_16444);
and U16603 (N_16603,N_16435,N_16354);
xor U16604 (N_16604,N_16444,N_16461);
or U16605 (N_16605,N_16417,N_16361);
or U16606 (N_16606,N_16405,N_16360);
or U16607 (N_16607,N_16448,N_16338);
or U16608 (N_16608,N_16422,N_16322);
or U16609 (N_16609,N_16355,N_16403);
and U16610 (N_16610,N_16466,N_16436);
xnor U16611 (N_16611,N_16426,N_16398);
or U16612 (N_16612,N_16390,N_16339);
xor U16613 (N_16613,N_16395,N_16459);
xnor U16614 (N_16614,N_16470,N_16383);
and U16615 (N_16615,N_16320,N_16444);
xnor U16616 (N_16616,N_16421,N_16479);
and U16617 (N_16617,N_16361,N_16458);
xor U16618 (N_16618,N_16367,N_16388);
and U16619 (N_16619,N_16429,N_16374);
or U16620 (N_16620,N_16455,N_16392);
and U16621 (N_16621,N_16425,N_16324);
nor U16622 (N_16622,N_16463,N_16326);
xnor U16623 (N_16623,N_16386,N_16389);
and U16624 (N_16624,N_16329,N_16409);
or U16625 (N_16625,N_16445,N_16405);
nor U16626 (N_16626,N_16323,N_16397);
xnor U16627 (N_16627,N_16390,N_16415);
nand U16628 (N_16628,N_16367,N_16404);
nor U16629 (N_16629,N_16321,N_16422);
nor U16630 (N_16630,N_16453,N_16344);
xnor U16631 (N_16631,N_16344,N_16462);
and U16632 (N_16632,N_16347,N_16387);
nor U16633 (N_16633,N_16410,N_16357);
nand U16634 (N_16634,N_16414,N_16410);
nand U16635 (N_16635,N_16426,N_16446);
xor U16636 (N_16636,N_16344,N_16390);
xnor U16637 (N_16637,N_16387,N_16391);
xor U16638 (N_16638,N_16401,N_16369);
nor U16639 (N_16639,N_16425,N_16390);
xor U16640 (N_16640,N_16518,N_16500);
nor U16641 (N_16641,N_16556,N_16526);
nor U16642 (N_16642,N_16637,N_16546);
nor U16643 (N_16643,N_16602,N_16555);
or U16644 (N_16644,N_16521,N_16600);
or U16645 (N_16645,N_16510,N_16560);
nor U16646 (N_16646,N_16497,N_16488);
or U16647 (N_16647,N_16634,N_16534);
nand U16648 (N_16648,N_16545,N_16525);
and U16649 (N_16649,N_16530,N_16570);
or U16650 (N_16650,N_16508,N_16568);
xor U16651 (N_16651,N_16553,N_16586);
xnor U16652 (N_16652,N_16612,N_16496);
nand U16653 (N_16653,N_16481,N_16520);
nor U16654 (N_16654,N_16566,N_16561);
and U16655 (N_16655,N_16613,N_16494);
nor U16656 (N_16656,N_16551,N_16621);
or U16657 (N_16657,N_16523,N_16541);
or U16658 (N_16658,N_16605,N_16611);
nor U16659 (N_16659,N_16626,N_16597);
xnor U16660 (N_16660,N_16584,N_16486);
nor U16661 (N_16661,N_16573,N_16574);
nor U16662 (N_16662,N_16599,N_16615);
xor U16663 (N_16663,N_16569,N_16628);
nand U16664 (N_16664,N_16578,N_16544);
or U16665 (N_16665,N_16601,N_16583);
and U16666 (N_16666,N_16504,N_16515);
nand U16667 (N_16667,N_16483,N_16581);
xor U16668 (N_16668,N_16623,N_16639);
nand U16669 (N_16669,N_16577,N_16502);
nand U16670 (N_16670,N_16506,N_16572);
or U16671 (N_16671,N_16576,N_16625);
nor U16672 (N_16672,N_16490,N_16607);
xnor U16673 (N_16673,N_16565,N_16527);
or U16674 (N_16674,N_16616,N_16606);
nor U16675 (N_16675,N_16617,N_16563);
or U16676 (N_16676,N_16524,N_16498);
or U16677 (N_16677,N_16622,N_16575);
xnor U16678 (N_16678,N_16614,N_16608);
nor U16679 (N_16679,N_16509,N_16633);
and U16680 (N_16680,N_16540,N_16624);
and U16681 (N_16681,N_16550,N_16579);
xnor U16682 (N_16682,N_16604,N_16585);
and U16683 (N_16683,N_16491,N_16632);
nor U16684 (N_16684,N_16482,N_16595);
nand U16685 (N_16685,N_16594,N_16587);
or U16686 (N_16686,N_16591,N_16532);
nor U16687 (N_16687,N_16485,N_16517);
nand U16688 (N_16688,N_16516,N_16593);
or U16689 (N_16689,N_16582,N_16507);
and U16690 (N_16690,N_16596,N_16559);
or U16691 (N_16691,N_16480,N_16513);
nor U16692 (N_16692,N_16543,N_16535);
or U16693 (N_16693,N_16620,N_16598);
nor U16694 (N_16694,N_16489,N_16492);
or U16695 (N_16695,N_16564,N_16609);
nor U16696 (N_16696,N_16542,N_16501);
nor U16697 (N_16697,N_16592,N_16590);
or U16698 (N_16698,N_16484,N_16512);
or U16699 (N_16699,N_16511,N_16635);
nand U16700 (N_16700,N_16610,N_16538);
nor U16701 (N_16701,N_16547,N_16537);
nor U16702 (N_16702,N_16629,N_16514);
nor U16703 (N_16703,N_16533,N_16554);
nor U16704 (N_16704,N_16548,N_16631);
and U16705 (N_16705,N_16539,N_16562);
xnor U16706 (N_16706,N_16638,N_16495);
nand U16707 (N_16707,N_16536,N_16571);
and U16708 (N_16708,N_16529,N_16627);
or U16709 (N_16709,N_16531,N_16589);
or U16710 (N_16710,N_16567,N_16557);
nor U16711 (N_16711,N_16588,N_16503);
nor U16712 (N_16712,N_16505,N_16552);
nor U16713 (N_16713,N_16528,N_16630);
or U16714 (N_16714,N_16618,N_16487);
nand U16715 (N_16715,N_16619,N_16580);
nand U16716 (N_16716,N_16519,N_16522);
xor U16717 (N_16717,N_16558,N_16636);
and U16718 (N_16718,N_16499,N_16549);
or U16719 (N_16719,N_16493,N_16603);
and U16720 (N_16720,N_16613,N_16530);
nor U16721 (N_16721,N_16496,N_16598);
xnor U16722 (N_16722,N_16555,N_16567);
xor U16723 (N_16723,N_16529,N_16609);
and U16724 (N_16724,N_16537,N_16567);
or U16725 (N_16725,N_16494,N_16586);
and U16726 (N_16726,N_16481,N_16595);
nor U16727 (N_16727,N_16550,N_16597);
and U16728 (N_16728,N_16579,N_16589);
xnor U16729 (N_16729,N_16552,N_16557);
nor U16730 (N_16730,N_16556,N_16630);
and U16731 (N_16731,N_16621,N_16537);
nor U16732 (N_16732,N_16574,N_16638);
and U16733 (N_16733,N_16570,N_16519);
nand U16734 (N_16734,N_16619,N_16633);
xnor U16735 (N_16735,N_16617,N_16628);
nand U16736 (N_16736,N_16637,N_16538);
nor U16737 (N_16737,N_16597,N_16624);
nor U16738 (N_16738,N_16580,N_16635);
and U16739 (N_16739,N_16533,N_16493);
nand U16740 (N_16740,N_16610,N_16577);
or U16741 (N_16741,N_16544,N_16595);
nand U16742 (N_16742,N_16480,N_16512);
xnor U16743 (N_16743,N_16573,N_16566);
and U16744 (N_16744,N_16623,N_16491);
xnor U16745 (N_16745,N_16551,N_16618);
nand U16746 (N_16746,N_16593,N_16519);
xor U16747 (N_16747,N_16535,N_16612);
nor U16748 (N_16748,N_16502,N_16581);
nor U16749 (N_16749,N_16597,N_16520);
or U16750 (N_16750,N_16561,N_16588);
nor U16751 (N_16751,N_16497,N_16556);
and U16752 (N_16752,N_16501,N_16597);
xnor U16753 (N_16753,N_16526,N_16525);
and U16754 (N_16754,N_16628,N_16605);
and U16755 (N_16755,N_16626,N_16558);
nor U16756 (N_16756,N_16603,N_16500);
nor U16757 (N_16757,N_16527,N_16632);
xnor U16758 (N_16758,N_16615,N_16523);
and U16759 (N_16759,N_16605,N_16492);
and U16760 (N_16760,N_16505,N_16625);
xnor U16761 (N_16761,N_16522,N_16632);
xnor U16762 (N_16762,N_16586,N_16517);
and U16763 (N_16763,N_16500,N_16525);
nand U16764 (N_16764,N_16548,N_16598);
xor U16765 (N_16765,N_16593,N_16517);
and U16766 (N_16766,N_16618,N_16637);
xor U16767 (N_16767,N_16521,N_16529);
nor U16768 (N_16768,N_16494,N_16541);
or U16769 (N_16769,N_16558,N_16580);
or U16770 (N_16770,N_16606,N_16573);
and U16771 (N_16771,N_16619,N_16578);
and U16772 (N_16772,N_16608,N_16520);
nor U16773 (N_16773,N_16592,N_16581);
or U16774 (N_16774,N_16577,N_16538);
or U16775 (N_16775,N_16586,N_16489);
nor U16776 (N_16776,N_16608,N_16575);
or U16777 (N_16777,N_16502,N_16487);
nand U16778 (N_16778,N_16589,N_16532);
and U16779 (N_16779,N_16555,N_16510);
nand U16780 (N_16780,N_16588,N_16487);
or U16781 (N_16781,N_16638,N_16480);
xnor U16782 (N_16782,N_16504,N_16583);
nor U16783 (N_16783,N_16611,N_16531);
nand U16784 (N_16784,N_16524,N_16610);
and U16785 (N_16785,N_16572,N_16621);
and U16786 (N_16786,N_16585,N_16490);
xor U16787 (N_16787,N_16598,N_16607);
or U16788 (N_16788,N_16572,N_16517);
nand U16789 (N_16789,N_16591,N_16609);
xor U16790 (N_16790,N_16623,N_16590);
nand U16791 (N_16791,N_16616,N_16584);
xnor U16792 (N_16792,N_16498,N_16536);
nor U16793 (N_16793,N_16504,N_16586);
and U16794 (N_16794,N_16622,N_16547);
or U16795 (N_16795,N_16587,N_16556);
and U16796 (N_16796,N_16529,N_16610);
nor U16797 (N_16797,N_16487,N_16637);
nor U16798 (N_16798,N_16630,N_16626);
and U16799 (N_16799,N_16570,N_16608);
and U16800 (N_16800,N_16681,N_16745);
nand U16801 (N_16801,N_16722,N_16674);
xor U16802 (N_16802,N_16668,N_16784);
xor U16803 (N_16803,N_16795,N_16700);
nand U16804 (N_16804,N_16724,N_16673);
xor U16805 (N_16805,N_16780,N_16701);
nand U16806 (N_16806,N_16685,N_16758);
nand U16807 (N_16807,N_16676,N_16739);
xor U16808 (N_16808,N_16688,N_16647);
nand U16809 (N_16809,N_16680,N_16672);
and U16810 (N_16810,N_16648,N_16663);
or U16811 (N_16811,N_16798,N_16665);
xor U16812 (N_16812,N_16705,N_16693);
nand U16813 (N_16813,N_16746,N_16690);
nand U16814 (N_16814,N_16656,N_16651);
nand U16815 (N_16815,N_16742,N_16695);
nand U16816 (N_16816,N_16664,N_16706);
nor U16817 (N_16817,N_16738,N_16779);
nor U16818 (N_16818,N_16670,N_16642);
nand U16819 (N_16819,N_16692,N_16789);
nand U16820 (N_16820,N_16744,N_16749);
or U16821 (N_16821,N_16791,N_16752);
xor U16822 (N_16822,N_16734,N_16737);
or U16823 (N_16823,N_16707,N_16773);
nor U16824 (N_16824,N_16760,N_16759);
xor U16825 (N_16825,N_16644,N_16794);
and U16826 (N_16826,N_16708,N_16774);
or U16827 (N_16827,N_16640,N_16698);
nor U16828 (N_16828,N_16661,N_16709);
and U16829 (N_16829,N_16652,N_16653);
nor U16830 (N_16830,N_16799,N_16719);
nor U16831 (N_16831,N_16770,N_16776);
xnor U16832 (N_16832,N_16792,N_16777);
xor U16833 (N_16833,N_16753,N_16669);
nor U16834 (N_16834,N_16755,N_16743);
or U16835 (N_16835,N_16768,N_16714);
or U16836 (N_16836,N_16691,N_16733);
and U16837 (N_16837,N_16679,N_16713);
nor U16838 (N_16838,N_16730,N_16699);
or U16839 (N_16839,N_16741,N_16729);
or U16840 (N_16840,N_16717,N_16731);
nor U16841 (N_16841,N_16727,N_16715);
or U16842 (N_16842,N_16682,N_16694);
nor U16843 (N_16843,N_16797,N_16790);
and U16844 (N_16844,N_16787,N_16763);
xnor U16845 (N_16845,N_16660,N_16754);
xor U16846 (N_16846,N_16786,N_16783);
and U16847 (N_16847,N_16721,N_16767);
xor U16848 (N_16848,N_16646,N_16778);
nand U16849 (N_16849,N_16785,N_16726);
nor U16850 (N_16850,N_16765,N_16696);
nand U16851 (N_16851,N_16756,N_16728);
and U16852 (N_16852,N_16655,N_16750);
xnor U16853 (N_16853,N_16747,N_16736);
nor U16854 (N_16854,N_16761,N_16697);
and U16855 (N_16855,N_16748,N_16678);
xor U16856 (N_16856,N_16686,N_16764);
and U16857 (N_16857,N_16643,N_16772);
nand U16858 (N_16858,N_16684,N_16666);
and U16859 (N_16859,N_16732,N_16654);
and U16860 (N_16860,N_16771,N_16702);
and U16861 (N_16861,N_16704,N_16796);
and U16862 (N_16862,N_16650,N_16718);
nand U16863 (N_16863,N_16658,N_16769);
and U16864 (N_16864,N_16782,N_16689);
or U16865 (N_16865,N_16716,N_16677);
or U16866 (N_16866,N_16687,N_16703);
xnor U16867 (N_16867,N_16657,N_16725);
or U16868 (N_16868,N_16675,N_16641);
nor U16869 (N_16869,N_16762,N_16671);
or U16870 (N_16870,N_16723,N_16662);
xor U16871 (N_16871,N_16781,N_16757);
or U16872 (N_16872,N_16766,N_16740);
xnor U16873 (N_16873,N_16710,N_16659);
nor U16874 (N_16874,N_16649,N_16645);
nor U16875 (N_16875,N_16711,N_16683);
nor U16876 (N_16876,N_16793,N_16788);
or U16877 (N_16877,N_16712,N_16735);
or U16878 (N_16878,N_16667,N_16775);
and U16879 (N_16879,N_16720,N_16751);
nand U16880 (N_16880,N_16783,N_16748);
nand U16881 (N_16881,N_16684,N_16721);
nand U16882 (N_16882,N_16656,N_16665);
nand U16883 (N_16883,N_16792,N_16749);
and U16884 (N_16884,N_16642,N_16737);
nor U16885 (N_16885,N_16684,N_16679);
xor U16886 (N_16886,N_16740,N_16694);
nor U16887 (N_16887,N_16741,N_16687);
xnor U16888 (N_16888,N_16723,N_16702);
xor U16889 (N_16889,N_16749,N_16740);
xnor U16890 (N_16890,N_16723,N_16686);
nand U16891 (N_16891,N_16780,N_16682);
and U16892 (N_16892,N_16672,N_16704);
nand U16893 (N_16893,N_16647,N_16759);
and U16894 (N_16894,N_16763,N_16704);
nand U16895 (N_16895,N_16646,N_16758);
xor U16896 (N_16896,N_16647,N_16684);
nor U16897 (N_16897,N_16682,N_16753);
nand U16898 (N_16898,N_16686,N_16797);
and U16899 (N_16899,N_16710,N_16778);
and U16900 (N_16900,N_16646,N_16676);
nand U16901 (N_16901,N_16726,N_16675);
nand U16902 (N_16902,N_16754,N_16751);
nand U16903 (N_16903,N_16772,N_16767);
and U16904 (N_16904,N_16695,N_16782);
and U16905 (N_16905,N_16781,N_16773);
xor U16906 (N_16906,N_16706,N_16745);
nand U16907 (N_16907,N_16697,N_16744);
or U16908 (N_16908,N_16678,N_16717);
nand U16909 (N_16909,N_16646,N_16694);
nor U16910 (N_16910,N_16698,N_16682);
or U16911 (N_16911,N_16715,N_16642);
xnor U16912 (N_16912,N_16688,N_16691);
nand U16913 (N_16913,N_16710,N_16729);
xor U16914 (N_16914,N_16699,N_16661);
nor U16915 (N_16915,N_16755,N_16645);
or U16916 (N_16916,N_16730,N_16784);
nand U16917 (N_16917,N_16671,N_16659);
xnor U16918 (N_16918,N_16649,N_16673);
nand U16919 (N_16919,N_16698,N_16646);
nor U16920 (N_16920,N_16706,N_16709);
xor U16921 (N_16921,N_16673,N_16646);
and U16922 (N_16922,N_16786,N_16778);
nor U16923 (N_16923,N_16713,N_16702);
and U16924 (N_16924,N_16701,N_16685);
nand U16925 (N_16925,N_16685,N_16689);
nor U16926 (N_16926,N_16720,N_16739);
nand U16927 (N_16927,N_16756,N_16732);
nand U16928 (N_16928,N_16690,N_16714);
and U16929 (N_16929,N_16642,N_16753);
and U16930 (N_16930,N_16786,N_16764);
nor U16931 (N_16931,N_16741,N_16751);
or U16932 (N_16932,N_16770,N_16749);
nand U16933 (N_16933,N_16730,N_16693);
xor U16934 (N_16934,N_16748,N_16666);
and U16935 (N_16935,N_16770,N_16653);
xnor U16936 (N_16936,N_16780,N_16648);
or U16937 (N_16937,N_16678,N_16786);
or U16938 (N_16938,N_16796,N_16720);
nand U16939 (N_16939,N_16685,N_16658);
nand U16940 (N_16940,N_16733,N_16799);
nand U16941 (N_16941,N_16644,N_16762);
nor U16942 (N_16942,N_16732,N_16797);
and U16943 (N_16943,N_16798,N_16693);
nand U16944 (N_16944,N_16720,N_16724);
and U16945 (N_16945,N_16760,N_16736);
xor U16946 (N_16946,N_16713,N_16674);
or U16947 (N_16947,N_16713,N_16749);
or U16948 (N_16948,N_16736,N_16772);
nor U16949 (N_16949,N_16671,N_16748);
or U16950 (N_16950,N_16748,N_16759);
nand U16951 (N_16951,N_16653,N_16658);
nor U16952 (N_16952,N_16778,N_16785);
or U16953 (N_16953,N_16687,N_16777);
or U16954 (N_16954,N_16704,N_16748);
and U16955 (N_16955,N_16668,N_16686);
and U16956 (N_16956,N_16668,N_16676);
nand U16957 (N_16957,N_16763,N_16782);
nor U16958 (N_16958,N_16742,N_16770);
or U16959 (N_16959,N_16746,N_16751);
or U16960 (N_16960,N_16939,N_16947);
nand U16961 (N_16961,N_16917,N_16806);
xor U16962 (N_16962,N_16875,N_16814);
nor U16963 (N_16963,N_16863,N_16955);
or U16964 (N_16964,N_16893,N_16871);
or U16965 (N_16965,N_16802,N_16951);
or U16966 (N_16966,N_16923,N_16889);
and U16967 (N_16967,N_16852,N_16830);
nand U16968 (N_16968,N_16948,N_16847);
xor U16969 (N_16969,N_16815,N_16942);
nand U16970 (N_16970,N_16808,N_16884);
nor U16971 (N_16971,N_16858,N_16868);
or U16972 (N_16972,N_16899,N_16865);
and U16973 (N_16973,N_16914,N_16813);
xor U16974 (N_16974,N_16918,N_16901);
and U16975 (N_16975,N_16898,N_16861);
nand U16976 (N_16976,N_16824,N_16828);
nand U16977 (N_16977,N_16932,N_16856);
nor U16978 (N_16978,N_16800,N_16953);
and U16979 (N_16979,N_16897,N_16931);
nand U16980 (N_16980,N_16878,N_16869);
xor U16981 (N_16981,N_16834,N_16864);
or U16982 (N_16982,N_16925,N_16823);
nor U16983 (N_16983,N_16936,N_16900);
nor U16984 (N_16984,N_16816,N_16891);
nor U16985 (N_16985,N_16920,N_16850);
xor U16986 (N_16986,N_16956,N_16952);
nor U16987 (N_16987,N_16819,N_16810);
nor U16988 (N_16988,N_16831,N_16945);
nand U16989 (N_16989,N_16836,N_16921);
nand U16990 (N_16990,N_16853,N_16881);
or U16991 (N_16991,N_16801,N_16804);
and U16992 (N_16992,N_16912,N_16872);
xor U16993 (N_16993,N_16820,N_16957);
xnor U16994 (N_16994,N_16906,N_16840);
or U16995 (N_16995,N_16887,N_16911);
and U16996 (N_16996,N_16913,N_16894);
and U16997 (N_16997,N_16880,N_16924);
and U16998 (N_16998,N_16903,N_16922);
or U16999 (N_16999,N_16822,N_16905);
and U17000 (N_17000,N_16904,N_16859);
or U17001 (N_17001,N_16886,N_16907);
or U17002 (N_17002,N_16950,N_16832);
or U17003 (N_17003,N_16895,N_16896);
nor U17004 (N_17004,N_16848,N_16873);
or U17005 (N_17005,N_16844,N_16916);
and U17006 (N_17006,N_16902,N_16915);
and U17007 (N_17007,N_16937,N_16877);
nor U17008 (N_17008,N_16826,N_16882);
xnor U17009 (N_17009,N_16927,N_16857);
nor U17010 (N_17010,N_16829,N_16938);
nand U17011 (N_17011,N_16946,N_16944);
nor U17012 (N_17012,N_16940,N_16959);
and U17013 (N_17013,N_16890,N_16949);
or U17014 (N_17014,N_16837,N_16821);
or U17015 (N_17015,N_16805,N_16803);
nand U17016 (N_17016,N_16879,N_16811);
nor U17017 (N_17017,N_16817,N_16851);
xor U17018 (N_17018,N_16843,N_16909);
nand U17019 (N_17019,N_16827,N_16926);
nand U17020 (N_17020,N_16842,N_16825);
or U17021 (N_17021,N_16835,N_16841);
and U17022 (N_17022,N_16855,N_16933);
xnor U17023 (N_17023,N_16874,N_16870);
nand U17024 (N_17024,N_16807,N_16958);
xnor U17025 (N_17025,N_16839,N_16860);
or U17026 (N_17026,N_16892,N_16809);
nor U17027 (N_17027,N_16908,N_16818);
nor U17028 (N_17028,N_16854,N_16812);
xor U17029 (N_17029,N_16885,N_16941);
or U17030 (N_17030,N_16919,N_16876);
nor U17031 (N_17031,N_16935,N_16846);
nor U17032 (N_17032,N_16833,N_16954);
and U17033 (N_17033,N_16883,N_16845);
and U17034 (N_17034,N_16928,N_16862);
or U17035 (N_17035,N_16888,N_16867);
or U17036 (N_17036,N_16866,N_16934);
and U17037 (N_17037,N_16910,N_16849);
and U17038 (N_17038,N_16943,N_16930);
nor U17039 (N_17039,N_16929,N_16838);
nor U17040 (N_17040,N_16952,N_16829);
or U17041 (N_17041,N_16823,N_16867);
xor U17042 (N_17042,N_16807,N_16846);
and U17043 (N_17043,N_16805,N_16839);
nor U17044 (N_17044,N_16821,N_16959);
and U17045 (N_17045,N_16910,N_16840);
or U17046 (N_17046,N_16901,N_16805);
xor U17047 (N_17047,N_16860,N_16928);
xnor U17048 (N_17048,N_16929,N_16935);
and U17049 (N_17049,N_16814,N_16915);
and U17050 (N_17050,N_16868,N_16952);
nor U17051 (N_17051,N_16879,N_16917);
xnor U17052 (N_17052,N_16953,N_16853);
nor U17053 (N_17053,N_16842,N_16955);
xnor U17054 (N_17054,N_16895,N_16890);
and U17055 (N_17055,N_16923,N_16839);
xor U17056 (N_17056,N_16891,N_16873);
xor U17057 (N_17057,N_16879,N_16924);
or U17058 (N_17058,N_16851,N_16801);
or U17059 (N_17059,N_16954,N_16853);
nand U17060 (N_17060,N_16832,N_16887);
xor U17061 (N_17061,N_16896,N_16891);
nor U17062 (N_17062,N_16938,N_16931);
nor U17063 (N_17063,N_16921,N_16935);
or U17064 (N_17064,N_16856,N_16804);
and U17065 (N_17065,N_16818,N_16884);
nor U17066 (N_17066,N_16917,N_16814);
nor U17067 (N_17067,N_16929,N_16872);
or U17068 (N_17068,N_16836,N_16803);
xnor U17069 (N_17069,N_16905,N_16832);
nand U17070 (N_17070,N_16914,N_16844);
nand U17071 (N_17071,N_16937,N_16852);
nand U17072 (N_17072,N_16917,N_16855);
nor U17073 (N_17073,N_16928,N_16836);
or U17074 (N_17074,N_16820,N_16861);
xnor U17075 (N_17075,N_16937,N_16840);
xor U17076 (N_17076,N_16920,N_16863);
or U17077 (N_17077,N_16868,N_16918);
and U17078 (N_17078,N_16954,N_16863);
or U17079 (N_17079,N_16833,N_16803);
and U17080 (N_17080,N_16849,N_16946);
or U17081 (N_17081,N_16901,N_16949);
xor U17082 (N_17082,N_16868,N_16865);
or U17083 (N_17083,N_16878,N_16958);
and U17084 (N_17084,N_16933,N_16941);
nand U17085 (N_17085,N_16901,N_16856);
nand U17086 (N_17086,N_16955,N_16805);
nor U17087 (N_17087,N_16955,N_16838);
nand U17088 (N_17088,N_16943,N_16826);
xor U17089 (N_17089,N_16897,N_16853);
or U17090 (N_17090,N_16912,N_16957);
and U17091 (N_17091,N_16915,N_16810);
nor U17092 (N_17092,N_16859,N_16854);
nor U17093 (N_17093,N_16816,N_16819);
and U17094 (N_17094,N_16868,N_16812);
xor U17095 (N_17095,N_16941,N_16875);
nor U17096 (N_17096,N_16884,N_16954);
nand U17097 (N_17097,N_16940,N_16909);
and U17098 (N_17098,N_16936,N_16827);
nand U17099 (N_17099,N_16923,N_16862);
and U17100 (N_17100,N_16870,N_16894);
or U17101 (N_17101,N_16886,N_16837);
nor U17102 (N_17102,N_16819,N_16855);
nand U17103 (N_17103,N_16875,N_16856);
nand U17104 (N_17104,N_16863,N_16805);
xor U17105 (N_17105,N_16897,N_16836);
or U17106 (N_17106,N_16881,N_16932);
nand U17107 (N_17107,N_16941,N_16894);
nand U17108 (N_17108,N_16812,N_16927);
or U17109 (N_17109,N_16888,N_16865);
nor U17110 (N_17110,N_16958,N_16890);
nor U17111 (N_17111,N_16811,N_16802);
or U17112 (N_17112,N_16824,N_16925);
and U17113 (N_17113,N_16845,N_16939);
and U17114 (N_17114,N_16821,N_16901);
and U17115 (N_17115,N_16818,N_16903);
nand U17116 (N_17116,N_16883,N_16820);
or U17117 (N_17117,N_16906,N_16894);
and U17118 (N_17118,N_16858,N_16931);
nand U17119 (N_17119,N_16879,N_16858);
or U17120 (N_17120,N_16995,N_17055);
and U17121 (N_17121,N_17119,N_16999);
xnor U17122 (N_17122,N_17063,N_17032);
and U17123 (N_17123,N_17109,N_17016);
xor U17124 (N_17124,N_16984,N_16968);
nand U17125 (N_17125,N_17011,N_17027);
and U17126 (N_17126,N_17097,N_17064);
xor U17127 (N_17127,N_17001,N_16973);
and U17128 (N_17128,N_17031,N_17103);
nor U17129 (N_17129,N_16992,N_16972);
and U17130 (N_17130,N_17082,N_17081);
nand U17131 (N_17131,N_17009,N_17037);
xnor U17132 (N_17132,N_17076,N_16960);
or U17133 (N_17133,N_17091,N_17042);
nand U17134 (N_17134,N_17101,N_17023);
nand U17135 (N_17135,N_16988,N_17086);
and U17136 (N_17136,N_17043,N_16967);
and U17137 (N_17137,N_17072,N_17053);
xnor U17138 (N_17138,N_17030,N_16985);
and U17139 (N_17139,N_16990,N_17073);
nand U17140 (N_17140,N_17051,N_16969);
xor U17141 (N_17141,N_17071,N_17007);
nand U17142 (N_17142,N_17029,N_17116);
xnor U17143 (N_17143,N_17094,N_17098);
or U17144 (N_17144,N_17036,N_16966);
xor U17145 (N_17145,N_17033,N_17035);
nand U17146 (N_17146,N_17002,N_17087);
or U17147 (N_17147,N_17056,N_17021);
or U17148 (N_17148,N_17078,N_17117);
or U17149 (N_17149,N_16963,N_17118);
nor U17150 (N_17150,N_17099,N_17065);
xor U17151 (N_17151,N_17034,N_17059);
xnor U17152 (N_17152,N_17005,N_16970);
xor U17153 (N_17153,N_16974,N_16971);
xor U17154 (N_17154,N_17017,N_17084);
or U17155 (N_17155,N_16981,N_16989);
and U17156 (N_17156,N_17112,N_17083);
or U17157 (N_17157,N_17004,N_17093);
nand U17158 (N_17158,N_17077,N_17058);
nand U17159 (N_17159,N_17049,N_17050);
nand U17160 (N_17160,N_17019,N_17041);
and U17161 (N_17161,N_17113,N_17044);
or U17162 (N_17162,N_17038,N_16975);
xnor U17163 (N_17163,N_16983,N_16982);
or U17164 (N_17164,N_17025,N_17024);
xnor U17165 (N_17165,N_17045,N_16986);
nor U17166 (N_17166,N_17010,N_17114);
or U17167 (N_17167,N_17090,N_17079);
or U17168 (N_17168,N_17026,N_17046);
xor U17169 (N_17169,N_16977,N_17085);
nand U17170 (N_17170,N_17105,N_17100);
xnor U17171 (N_17171,N_16993,N_17092);
nor U17172 (N_17172,N_17062,N_17048);
nor U17173 (N_17173,N_16979,N_17052);
or U17174 (N_17174,N_17104,N_17088);
and U17175 (N_17175,N_17040,N_17068);
nor U17176 (N_17176,N_17047,N_16961);
nor U17177 (N_17177,N_17061,N_17080);
and U17178 (N_17178,N_16996,N_17106);
nand U17179 (N_17179,N_17008,N_17028);
nand U17180 (N_17180,N_16987,N_17102);
or U17181 (N_17181,N_17060,N_17012);
xnor U17182 (N_17182,N_17096,N_17015);
nand U17183 (N_17183,N_17089,N_17054);
nand U17184 (N_17184,N_17018,N_17014);
nand U17185 (N_17185,N_16976,N_17111);
xor U17186 (N_17186,N_16964,N_16998);
xnor U17187 (N_17187,N_16980,N_17067);
nand U17188 (N_17188,N_17039,N_17115);
nand U17189 (N_17189,N_17069,N_17057);
xor U17190 (N_17190,N_17107,N_17022);
and U17191 (N_17191,N_16997,N_17013);
and U17192 (N_17192,N_17110,N_17006);
nand U17193 (N_17193,N_16965,N_16962);
nand U17194 (N_17194,N_17095,N_16991);
and U17195 (N_17195,N_16994,N_17000);
or U17196 (N_17196,N_17075,N_17074);
xnor U17197 (N_17197,N_17066,N_17108);
nor U17198 (N_17198,N_17020,N_17003);
nand U17199 (N_17199,N_17070,N_16978);
xnor U17200 (N_17200,N_17052,N_17106);
and U17201 (N_17201,N_17098,N_17054);
nor U17202 (N_17202,N_16972,N_17095);
nand U17203 (N_17203,N_17102,N_16984);
nor U17204 (N_17204,N_16970,N_17036);
xnor U17205 (N_17205,N_17117,N_16975);
or U17206 (N_17206,N_16981,N_17053);
xnor U17207 (N_17207,N_17112,N_17056);
xnor U17208 (N_17208,N_17114,N_17053);
nand U17209 (N_17209,N_17036,N_16965);
and U17210 (N_17210,N_17064,N_17025);
xnor U17211 (N_17211,N_17111,N_17092);
and U17212 (N_17212,N_16990,N_17021);
xnor U17213 (N_17213,N_17061,N_16975);
nor U17214 (N_17214,N_16992,N_17083);
and U17215 (N_17215,N_17092,N_17001);
and U17216 (N_17216,N_17100,N_17059);
or U17217 (N_17217,N_17085,N_16971);
or U17218 (N_17218,N_17019,N_17076);
and U17219 (N_17219,N_17006,N_17080);
and U17220 (N_17220,N_17106,N_17024);
nand U17221 (N_17221,N_17052,N_16994);
nand U17222 (N_17222,N_16971,N_17052);
or U17223 (N_17223,N_16980,N_16974);
or U17224 (N_17224,N_17046,N_17118);
or U17225 (N_17225,N_16973,N_17093);
and U17226 (N_17226,N_16964,N_17082);
xor U17227 (N_17227,N_17061,N_17036);
nand U17228 (N_17228,N_17029,N_17111);
xor U17229 (N_17229,N_16963,N_17088);
xor U17230 (N_17230,N_17034,N_17029);
and U17231 (N_17231,N_17002,N_17068);
nand U17232 (N_17232,N_17057,N_17055);
xnor U17233 (N_17233,N_17106,N_16968);
or U17234 (N_17234,N_17056,N_17011);
or U17235 (N_17235,N_17031,N_17105);
xor U17236 (N_17236,N_17068,N_17099);
xnor U17237 (N_17237,N_17013,N_16987);
and U17238 (N_17238,N_17050,N_17014);
nand U17239 (N_17239,N_17004,N_17106);
and U17240 (N_17240,N_16962,N_17045);
nor U17241 (N_17241,N_17082,N_17005);
xnor U17242 (N_17242,N_17114,N_17031);
nor U17243 (N_17243,N_17118,N_16992);
xor U17244 (N_17244,N_17102,N_17111);
and U17245 (N_17245,N_17065,N_16980);
or U17246 (N_17246,N_17054,N_17052);
and U17247 (N_17247,N_17078,N_17093);
xor U17248 (N_17248,N_17027,N_16998);
or U17249 (N_17249,N_17050,N_17069);
nand U17250 (N_17250,N_16983,N_17094);
nand U17251 (N_17251,N_17003,N_17092);
or U17252 (N_17252,N_17047,N_16989);
xor U17253 (N_17253,N_17003,N_17055);
xnor U17254 (N_17254,N_16976,N_16980);
or U17255 (N_17255,N_16978,N_17056);
xor U17256 (N_17256,N_16961,N_16988);
nand U17257 (N_17257,N_17046,N_17070);
nor U17258 (N_17258,N_17024,N_16969);
nor U17259 (N_17259,N_16977,N_17114);
and U17260 (N_17260,N_17042,N_17037);
and U17261 (N_17261,N_17005,N_16985);
xor U17262 (N_17262,N_17092,N_17040);
nand U17263 (N_17263,N_16989,N_17091);
xor U17264 (N_17264,N_17020,N_17027);
nor U17265 (N_17265,N_17064,N_16976);
nand U17266 (N_17266,N_16998,N_17116);
xor U17267 (N_17267,N_17084,N_17093);
or U17268 (N_17268,N_17039,N_17068);
nand U17269 (N_17269,N_17047,N_17096);
or U17270 (N_17270,N_17063,N_17010);
and U17271 (N_17271,N_16967,N_17041);
or U17272 (N_17272,N_17069,N_17100);
xor U17273 (N_17273,N_17024,N_17107);
and U17274 (N_17274,N_17034,N_17077);
and U17275 (N_17275,N_17032,N_17099);
or U17276 (N_17276,N_17119,N_16993);
and U17277 (N_17277,N_17030,N_16980);
or U17278 (N_17278,N_17013,N_17069);
and U17279 (N_17279,N_16975,N_17086);
xnor U17280 (N_17280,N_17187,N_17202);
and U17281 (N_17281,N_17253,N_17146);
nor U17282 (N_17282,N_17227,N_17197);
nor U17283 (N_17283,N_17175,N_17120);
and U17284 (N_17284,N_17261,N_17248);
xnor U17285 (N_17285,N_17134,N_17161);
or U17286 (N_17286,N_17208,N_17219);
nor U17287 (N_17287,N_17266,N_17142);
xnor U17288 (N_17288,N_17238,N_17239);
nand U17289 (N_17289,N_17153,N_17190);
xnor U17290 (N_17290,N_17254,N_17184);
xor U17291 (N_17291,N_17240,N_17165);
nand U17292 (N_17292,N_17252,N_17233);
and U17293 (N_17293,N_17243,N_17232);
and U17294 (N_17294,N_17270,N_17207);
xor U17295 (N_17295,N_17216,N_17277);
xnor U17296 (N_17296,N_17228,N_17185);
xnor U17297 (N_17297,N_17265,N_17133);
and U17298 (N_17298,N_17150,N_17127);
and U17299 (N_17299,N_17180,N_17163);
or U17300 (N_17300,N_17145,N_17172);
xor U17301 (N_17301,N_17279,N_17214);
nand U17302 (N_17302,N_17132,N_17181);
nor U17303 (N_17303,N_17147,N_17173);
or U17304 (N_17304,N_17192,N_17205);
nor U17305 (N_17305,N_17151,N_17182);
or U17306 (N_17306,N_17176,N_17274);
nor U17307 (N_17307,N_17158,N_17201);
nand U17308 (N_17308,N_17138,N_17267);
or U17309 (N_17309,N_17244,N_17188);
xor U17310 (N_17310,N_17191,N_17149);
xnor U17311 (N_17311,N_17218,N_17234);
xor U17312 (N_17312,N_17256,N_17263);
nor U17313 (N_17313,N_17121,N_17196);
nand U17314 (N_17314,N_17213,N_17141);
nand U17315 (N_17315,N_17143,N_17194);
nand U17316 (N_17316,N_17221,N_17168);
nor U17317 (N_17317,N_17260,N_17209);
nand U17318 (N_17318,N_17223,N_17174);
xor U17319 (N_17319,N_17245,N_17135);
nand U17320 (N_17320,N_17264,N_17156);
xnor U17321 (N_17321,N_17272,N_17278);
xor U17322 (N_17322,N_17271,N_17262);
nand U17323 (N_17323,N_17250,N_17215);
and U17324 (N_17324,N_17235,N_17211);
nor U17325 (N_17325,N_17129,N_17128);
nand U17326 (N_17326,N_17178,N_17251);
nand U17327 (N_17327,N_17206,N_17183);
nor U17328 (N_17328,N_17164,N_17162);
nor U17329 (N_17329,N_17159,N_17130);
nand U17330 (N_17330,N_17249,N_17241);
nand U17331 (N_17331,N_17257,N_17231);
and U17332 (N_17332,N_17167,N_17255);
and U17333 (N_17333,N_17230,N_17179);
or U17334 (N_17334,N_17124,N_17247);
xnor U17335 (N_17335,N_17148,N_17144);
and U17336 (N_17336,N_17210,N_17195);
and U17337 (N_17337,N_17212,N_17204);
xor U17338 (N_17338,N_17269,N_17122);
xnor U17339 (N_17339,N_17131,N_17203);
xor U17340 (N_17340,N_17226,N_17140);
xnor U17341 (N_17341,N_17222,N_17225);
xnor U17342 (N_17342,N_17273,N_17276);
and U17343 (N_17343,N_17189,N_17199);
or U17344 (N_17344,N_17258,N_17160);
nor U17345 (N_17345,N_17123,N_17217);
or U17346 (N_17346,N_17154,N_17157);
and U17347 (N_17347,N_17242,N_17229);
or U17348 (N_17348,N_17236,N_17139);
xor U17349 (N_17349,N_17275,N_17136);
nor U17350 (N_17350,N_17198,N_17155);
xnor U17351 (N_17351,N_17237,N_17200);
nand U17352 (N_17352,N_17268,N_17125);
xor U17353 (N_17353,N_17259,N_17193);
nor U17354 (N_17354,N_17170,N_17169);
nand U17355 (N_17355,N_17166,N_17220);
nand U17356 (N_17356,N_17246,N_17224);
or U17357 (N_17357,N_17171,N_17126);
xnor U17358 (N_17358,N_17177,N_17137);
nand U17359 (N_17359,N_17152,N_17186);
or U17360 (N_17360,N_17139,N_17218);
and U17361 (N_17361,N_17156,N_17188);
and U17362 (N_17362,N_17169,N_17130);
nand U17363 (N_17363,N_17123,N_17169);
xnor U17364 (N_17364,N_17207,N_17224);
or U17365 (N_17365,N_17142,N_17221);
xnor U17366 (N_17366,N_17146,N_17205);
nor U17367 (N_17367,N_17195,N_17265);
and U17368 (N_17368,N_17276,N_17153);
nand U17369 (N_17369,N_17170,N_17141);
xor U17370 (N_17370,N_17182,N_17133);
xor U17371 (N_17371,N_17248,N_17204);
or U17372 (N_17372,N_17238,N_17194);
nand U17373 (N_17373,N_17143,N_17195);
nor U17374 (N_17374,N_17204,N_17142);
and U17375 (N_17375,N_17202,N_17145);
and U17376 (N_17376,N_17122,N_17208);
or U17377 (N_17377,N_17158,N_17178);
or U17378 (N_17378,N_17263,N_17274);
xor U17379 (N_17379,N_17179,N_17131);
nand U17380 (N_17380,N_17245,N_17267);
xor U17381 (N_17381,N_17261,N_17140);
nor U17382 (N_17382,N_17278,N_17195);
nand U17383 (N_17383,N_17137,N_17259);
or U17384 (N_17384,N_17197,N_17233);
or U17385 (N_17385,N_17200,N_17239);
xnor U17386 (N_17386,N_17252,N_17209);
xor U17387 (N_17387,N_17186,N_17187);
or U17388 (N_17388,N_17227,N_17232);
nand U17389 (N_17389,N_17213,N_17128);
or U17390 (N_17390,N_17274,N_17217);
and U17391 (N_17391,N_17232,N_17155);
nor U17392 (N_17392,N_17256,N_17208);
or U17393 (N_17393,N_17211,N_17241);
nand U17394 (N_17394,N_17193,N_17275);
and U17395 (N_17395,N_17227,N_17168);
nor U17396 (N_17396,N_17143,N_17190);
nand U17397 (N_17397,N_17162,N_17184);
nor U17398 (N_17398,N_17141,N_17279);
and U17399 (N_17399,N_17204,N_17193);
xnor U17400 (N_17400,N_17173,N_17217);
xnor U17401 (N_17401,N_17177,N_17131);
nor U17402 (N_17402,N_17213,N_17158);
or U17403 (N_17403,N_17216,N_17147);
nor U17404 (N_17404,N_17184,N_17153);
and U17405 (N_17405,N_17147,N_17124);
or U17406 (N_17406,N_17171,N_17204);
nand U17407 (N_17407,N_17253,N_17217);
or U17408 (N_17408,N_17226,N_17151);
xnor U17409 (N_17409,N_17160,N_17155);
or U17410 (N_17410,N_17225,N_17221);
nor U17411 (N_17411,N_17215,N_17161);
xor U17412 (N_17412,N_17155,N_17214);
xor U17413 (N_17413,N_17151,N_17215);
nor U17414 (N_17414,N_17187,N_17120);
nor U17415 (N_17415,N_17225,N_17226);
xnor U17416 (N_17416,N_17160,N_17173);
nand U17417 (N_17417,N_17212,N_17202);
nor U17418 (N_17418,N_17175,N_17174);
xnor U17419 (N_17419,N_17157,N_17165);
xnor U17420 (N_17420,N_17127,N_17174);
nand U17421 (N_17421,N_17174,N_17229);
nand U17422 (N_17422,N_17184,N_17178);
nor U17423 (N_17423,N_17222,N_17218);
and U17424 (N_17424,N_17217,N_17120);
nor U17425 (N_17425,N_17206,N_17136);
or U17426 (N_17426,N_17218,N_17251);
nor U17427 (N_17427,N_17177,N_17267);
nand U17428 (N_17428,N_17186,N_17270);
nand U17429 (N_17429,N_17132,N_17227);
xor U17430 (N_17430,N_17146,N_17208);
or U17431 (N_17431,N_17165,N_17253);
or U17432 (N_17432,N_17179,N_17146);
or U17433 (N_17433,N_17254,N_17268);
xnor U17434 (N_17434,N_17195,N_17125);
nand U17435 (N_17435,N_17241,N_17152);
and U17436 (N_17436,N_17270,N_17196);
nand U17437 (N_17437,N_17236,N_17232);
xor U17438 (N_17438,N_17143,N_17202);
nand U17439 (N_17439,N_17180,N_17204);
nand U17440 (N_17440,N_17332,N_17385);
and U17441 (N_17441,N_17362,N_17298);
nor U17442 (N_17442,N_17351,N_17397);
or U17443 (N_17443,N_17408,N_17372);
or U17444 (N_17444,N_17416,N_17296);
and U17445 (N_17445,N_17354,N_17302);
xnor U17446 (N_17446,N_17308,N_17359);
nand U17447 (N_17447,N_17411,N_17338);
and U17448 (N_17448,N_17369,N_17292);
nand U17449 (N_17449,N_17407,N_17391);
nand U17450 (N_17450,N_17341,N_17426);
nand U17451 (N_17451,N_17421,N_17393);
and U17452 (N_17452,N_17400,N_17427);
xnor U17453 (N_17453,N_17312,N_17422);
and U17454 (N_17454,N_17365,N_17290);
nor U17455 (N_17455,N_17431,N_17323);
and U17456 (N_17456,N_17363,N_17318);
nand U17457 (N_17457,N_17381,N_17295);
and U17458 (N_17458,N_17353,N_17281);
or U17459 (N_17459,N_17322,N_17378);
and U17460 (N_17460,N_17331,N_17280);
nor U17461 (N_17461,N_17300,N_17357);
and U17462 (N_17462,N_17291,N_17337);
and U17463 (N_17463,N_17383,N_17424);
or U17464 (N_17464,N_17382,N_17410);
nand U17465 (N_17465,N_17430,N_17425);
xor U17466 (N_17466,N_17414,N_17343);
xnor U17467 (N_17467,N_17373,N_17311);
or U17468 (N_17468,N_17345,N_17394);
and U17469 (N_17469,N_17380,N_17395);
nand U17470 (N_17470,N_17396,N_17384);
or U17471 (N_17471,N_17433,N_17439);
and U17472 (N_17472,N_17435,N_17375);
and U17473 (N_17473,N_17304,N_17321);
and U17474 (N_17474,N_17402,N_17428);
nand U17475 (N_17475,N_17314,N_17417);
nand U17476 (N_17476,N_17434,N_17437);
and U17477 (N_17477,N_17342,N_17293);
or U17478 (N_17478,N_17401,N_17317);
nand U17479 (N_17479,N_17324,N_17330);
or U17480 (N_17480,N_17307,N_17285);
or U17481 (N_17481,N_17301,N_17305);
nor U17482 (N_17482,N_17297,N_17392);
nor U17483 (N_17483,N_17355,N_17346);
or U17484 (N_17484,N_17299,N_17348);
or U17485 (N_17485,N_17289,N_17333);
or U17486 (N_17486,N_17339,N_17418);
or U17487 (N_17487,N_17374,N_17377);
and U17488 (N_17488,N_17356,N_17366);
or U17489 (N_17489,N_17406,N_17294);
or U17490 (N_17490,N_17315,N_17386);
and U17491 (N_17491,N_17286,N_17412);
or U17492 (N_17492,N_17361,N_17306);
xor U17493 (N_17493,N_17303,N_17328);
xor U17494 (N_17494,N_17282,N_17320);
nand U17495 (N_17495,N_17310,N_17404);
and U17496 (N_17496,N_17329,N_17344);
nor U17497 (N_17497,N_17429,N_17287);
and U17498 (N_17498,N_17379,N_17288);
xnor U17499 (N_17499,N_17368,N_17399);
xor U17500 (N_17500,N_17316,N_17347);
and U17501 (N_17501,N_17325,N_17376);
xnor U17502 (N_17502,N_17349,N_17283);
xor U17503 (N_17503,N_17423,N_17350);
xor U17504 (N_17504,N_17309,N_17398);
nand U17505 (N_17505,N_17313,N_17371);
nand U17506 (N_17506,N_17409,N_17327);
and U17507 (N_17507,N_17360,N_17420);
xor U17508 (N_17508,N_17319,N_17436);
and U17509 (N_17509,N_17352,N_17415);
nand U17510 (N_17510,N_17336,N_17284);
and U17511 (N_17511,N_17403,N_17364);
nand U17512 (N_17512,N_17387,N_17388);
xnor U17513 (N_17513,N_17389,N_17326);
xor U17514 (N_17514,N_17438,N_17390);
nand U17515 (N_17515,N_17358,N_17419);
xor U17516 (N_17516,N_17432,N_17340);
xor U17517 (N_17517,N_17334,N_17335);
nand U17518 (N_17518,N_17370,N_17367);
nor U17519 (N_17519,N_17413,N_17405);
and U17520 (N_17520,N_17347,N_17332);
and U17521 (N_17521,N_17380,N_17387);
and U17522 (N_17522,N_17328,N_17436);
xnor U17523 (N_17523,N_17379,N_17354);
xnor U17524 (N_17524,N_17428,N_17366);
and U17525 (N_17525,N_17423,N_17316);
nand U17526 (N_17526,N_17344,N_17418);
nand U17527 (N_17527,N_17319,N_17367);
nand U17528 (N_17528,N_17300,N_17304);
or U17529 (N_17529,N_17326,N_17359);
and U17530 (N_17530,N_17302,N_17413);
and U17531 (N_17531,N_17325,N_17360);
nand U17532 (N_17532,N_17377,N_17394);
and U17533 (N_17533,N_17407,N_17424);
xor U17534 (N_17534,N_17328,N_17309);
or U17535 (N_17535,N_17371,N_17376);
xor U17536 (N_17536,N_17434,N_17328);
nand U17537 (N_17537,N_17325,N_17302);
nand U17538 (N_17538,N_17374,N_17280);
and U17539 (N_17539,N_17324,N_17373);
nor U17540 (N_17540,N_17421,N_17281);
or U17541 (N_17541,N_17322,N_17421);
nor U17542 (N_17542,N_17386,N_17437);
and U17543 (N_17543,N_17362,N_17358);
nor U17544 (N_17544,N_17323,N_17303);
xnor U17545 (N_17545,N_17368,N_17377);
nor U17546 (N_17546,N_17282,N_17337);
and U17547 (N_17547,N_17338,N_17355);
and U17548 (N_17548,N_17314,N_17285);
nand U17549 (N_17549,N_17381,N_17284);
and U17550 (N_17550,N_17292,N_17431);
nand U17551 (N_17551,N_17384,N_17305);
nand U17552 (N_17552,N_17424,N_17340);
or U17553 (N_17553,N_17393,N_17350);
xnor U17554 (N_17554,N_17343,N_17346);
and U17555 (N_17555,N_17438,N_17297);
or U17556 (N_17556,N_17306,N_17400);
nor U17557 (N_17557,N_17362,N_17282);
nor U17558 (N_17558,N_17383,N_17321);
and U17559 (N_17559,N_17333,N_17382);
nor U17560 (N_17560,N_17430,N_17341);
or U17561 (N_17561,N_17393,N_17292);
and U17562 (N_17562,N_17387,N_17329);
xnor U17563 (N_17563,N_17439,N_17306);
or U17564 (N_17564,N_17422,N_17344);
and U17565 (N_17565,N_17362,N_17402);
nand U17566 (N_17566,N_17288,N_17377);
or U17567 (N_17567,N_17391,N_17397);
xor U17568 (N_17568,N_17311,N_17340);
xor U17569 (N_17569,N_17285,N_17351);
and U17570 (N_17570,N_17390,N_17316);
nand U17571 (N_17571,N_17433,N_17348);
xor U17572 (N_17572,N_17387,N_17339);
xnor U17573 (N_17573,N_17314,N_17387);
xor U17574 (N_17574,N_17310,N_17350);
xnor U17575 (N_17575,N_17431,N_17404);
or U17576 (N_17576,N_17301,N_17402);
and U17577 (N_17577,N_17362,N_17408);
nand U17578 (N_17578,N_17289,N_17334);
nor U17579 (N_17579,N_17295,N_17409);
or U17580 (N_17580,N_17319,N_17291);
nand U17581 (N_17581,N_17386,N_17318);
or U17582 (N_17582,N_17382,N_17291);
nand U17583 (N_17583,N_17353,N_17350);
nor U17584 (N_17584,N_17436,N_17326);
xor U17585 (N_17585,N_17425,N_17356);
nor U17586 (N_17586,N_17298,N_17317);
nor U17587 (N_17587,N_17284,N_17400);
xnor U17588 (N_17588,N_17435,N_17355);
nand U17589 (N_17589,N_17423,N_17331);
xnor U17590 (N_17590,N_17354,N_17322);
and U17591 (N_17591,N_17358,N_17434);
nor U17592 (N_17592,N_17318,N_17365);
xor U17593 (N_17593,N_17434,N_17298);
nand U17594 (N_17594,N_17305,N_17425);
nand U17595 (N_17595,N_17326,N_17413);
nor U17596 (N_17596,N_17437,N_17336);
nor U17597 (N_17597,N_17402,N_17325);
nor U17598 (N_17598,N_17284,N_17286);
or U17599 (N_17599,N_17332,N_17333);
nor U17600 (N_17600,N_17460,N_17539);
xnor U17601 (N_17601,N_17512,N_17454);
xor U17602 (N_17602,N_17508,N_17537);
nor U17603 (N_17603,N_17472,N_17585);
or U17604 (N_17604,N_17484,N_17485);
xor U17605 (N_17605,N_17463,N_17474);
or U17606 (N_17606,N_17448,N_17497);
and U17607 (N_17607,N_17501,N_17452);
nand U17608 (N_17608,N_17502,N_17503);
xnor U17609 (N_17609,N_17492,N_17581);
nand U17610 (N_17610,N_17552,N_17576);
or U17611 (N_17611,N_17531,N_17464);
and U17612 (N_17612,N_17498,N_17466);
or U17613 (N_17613,N_17596,N_17476);
or U17614 (N_17614,N_17483,N_17496);
and U17615 (N_17615,N_17459,N_17520);
nand U17616 (N_17616,N_17550,N_17443);
and U17617 (N_17617,N_17440,N_17444);
or U17618 (N_17618,N_17574,N_17468);
nor U17619 (N_17619,N_17481,N_17456);
nor U17620 (N_17620,N_17594,N_17457);
and U17621 (N_17621,N_17546,N_17458);
nand U17622 (N_17622,N_17568,N_17562);
and U17623 (N_17623,N_17528,N_17595);
nor U17624 (N_17624,N_17489,N_17553);
and U17625 (N_17625,N_17522,N_17572);
xor U17626 (N_17626,N_17511,N_17519);
or U17627 (N_17627,N_17455,N_17535);
nor U17628 (N_17628,N_17525,N_17534);
nand U17629 (N_17629,N_17447,N_17549);
or U17630 (N_17630,N_17565,N_17449);
and U17631 (N_17631,N_17577,N_17532);
nor U17632 (N_17632,N_17588,N_17545);
or U17633 (N_17633,N_17518,N_17465);
and U17634 (N_17634,N_17490,N_17516);
xnor U17635 (N_17635,N_17590,N_17541);
nand U17636 (N_17636,N_17530,N_17591);
xnor U17637 (N_17637,N_17471,N_17462);
or U17638 (N_17638,N_17487,N_17488);
xnor U17639 (N_17639,N_17555,N_17510);
nand U17640 (N_17640,N_17597,N_17495);
nand U17641 (N_17641,N_17566,N_17479);
nand U17642 (N_17642,N_17482,N_17446);
nand U17643 (N_17643,N_17505,N_17544);
xnor U17644 (N_17644,N_17451,N_17569);
nand U17645 (N_17645,N_17477,N_17579);
nand U17646 (N_17646,N_17515,N_17582);
nor U17647 (N_17647,N_17571,N_17564);
and U17648 (N_17648,N_17575,N_17523);
nor U17649 (N_17649,N_17567,N_17551);
xnor U17650 (N_17650,N_17538,N_17580);
nor U17651 (N_17651,N_17586,N_17587);
nand U17652 (N_17652,N_17441,N_17467);
nand U17653 (N_17653,N_17542,N_17494);
xor U17654 (N_17654,N_17517,N_17470);
nor U17655 (N_17655,N_17558,N_17469);
or U17656 (N_17656,N_17527,N_17493);
and U17657 (N_17657,N_17513,N_17486);
xor U17658 (N_17658,N_17599,N_17593);
nand U17659 (N_17659,N_17560,N_17557);
or U17660 (N_17660,N_17500,N_17526);
and U17661 (N_17661,N_17554,N_17540);
nor U17662 (N_17662,N_17453,N_17559);
or U17663 (N_17663,N_17556,N_17583);
nor U17664 (N_17664,N_17543,N_17442);
nand U17665 (N_17665,N_17478,N_17533);
or U17666 (N_17666,N_17473,N_17578);
nor U17667 (N_17667,N_17461,N_17529);
or U17668 (N_17668,N_17524,N_17598);
nand U17669 (N_17669,N_17570,N_17480);
xor U17670 (N_17670,N_17573,N_17584);
nand U17671 (N_17671,N_17491,N_17514);
xnor U17672 (N_17672,N_17521,N_17506);
xnor U17673 (N_17673,N_17561,N_17589);
nor U17674 (N_17674,N_17548,N_17547);
nand U17675 (N_17675,N_17504,N_17475);
xor U17676 (N_17676,N_17450,N_17499);
and U17677 (N_17677,N_17592,N_17536);
and U17678 (N_17678,N_17563,N_17445);
and U17679 (N_17679,N_17509,N_17507);
nand U17680 (N_17680,N_17529,N_17592);
or U17681 (N_17681,N_17553,N_17461);
xor U17682 (N_17682,N_17539,N_17532);
or U17683 (N_17683,N_17592,N_17493);
or U17684 (N_17684,N_17505,N_17477);
or U17685 (N_17685,N_17566,N_17560);
nand U17686 (N_17686,N_17489,N_17547);
or U17687 (N_17687,N_17485,N_17465);
and U17688 (N_17688,N_17585,N_17517);
and U17689 (N_17689,N_17482,N_17595);
or U17690 (N_17690,N_17578,N_17480);
and U17691 (N_17691,N_17545,N_17555);
nand U17692 (N_17692,N_17518,N_17499);
or U17693 (N_17693,N_17595,N_17474);
nand U17694 (N_17694,N_17577,N_17505);
nor U17695 (N_17695,N_17521,N_17575);
or U17696 (N_17696,N_17599,N_17448);
and U17697 (N_17697,N_17464,N_17462);
nand U17698 (N_17698,N_17464,N_17591);
nand U17699 (N_17699,N_17515,N_17552);
nand U17700 (N_17700,N_17598,N_17579);
and U17701 (N_17701,N_17544,N_17448);
and U17702 (N_17702,N_17530,N_17446);
nand U17703 (N_17703,N_17471,N_17570);
nand U17704 (N_17704,N_17466,N_17581);
xor U17705 (N_17705,N_17509,N_17544);
nor U17706 (N_17706,N_17530,N_17487);
xor U17707 (N_17707,N_17451,N_17573);
nor U17708 (N_17708,N_17548,N_17521);
nor U17709 (N_17709,N_17510,N_17558);
xor U17710 (N_17710,N_17469,N_17523);
nand U17711 (N_17711,N_17580,N_17462);
or U17712 (N_17712,N_17598,N_17482);
and U17713 (N_17713,N_17523,N_17588);
or U17714 (N_17714,N_17592,N_17511);
xor U17715 (N_17715,N_17563,N_17517);
nand U17716 (N_17716,N_17507,N_17475);
nand U17717 (N_17717,N_17468,N_17490);
xor U17718 (N_17718,N_17540,N_17541);
nor U17719 (N_17719,N_17592,N_17579);
xnor U17720 (N_17720,N_17476,N_17451);
and U17721 (N_17721,N_17467,N_17440);
nor U17722 (N_17722,N_17537,N_17560);
and U17723 (N_17723,N_17501,N_17467);
nand U17724 (N_17724,N_17457,N_17572);
and U17725 (N_17725,N_17594,N_17590);
or U17726 (N_17726,N_17597,N_17554);
nor U17727 (N_17727,N_17533,N_17509);
nand U17728 (N_17728,N_17564,N_17590);
xor U17729 (N_17729,N_17460,N_17546);
nand U17730 (N_17730,N_17593,N_17522);
nor U17731 (N_17731,N_17455,N_17544);
or U17732 (N_17732,N_17563,N_17510);
xor U17733 (N_17733,N_17547,N_17486);
nor U17734 (N_17734,N_17447,N_17557);
xnor U17735 (N_17735,N_17470,N_17490);
nand U17736 (N_17736,N_17595,N_17519);
and U17737 (N_17737,N_17566,N_17481);
or U17738 (N_17738,N_17495,N_17468);
xnor U17739 (N_17739,N_17586,N_17484);
or U17740 (N_17740,N_17563,N_17443);
nand U17741 (N_17741,N_17519,N_17454);
or U17742 (N_17742,N_17516,N_17479);
xor U17743 (N_17743,N_17456,N_17465);
xnor U17744 (N_17744,N_17459,N_17488);
nor U17745 (N_17745,N_17548,N_17450);
xnor U17746 (N_17746,N_17478,N_17474);
xor U17747 (N_17747,N_17541,N_17459);
and U17748 (N_17748,N_17548,N_17489);
nand U17749 (N_17749,N_17505,N_17459);
xnor U17750 (N_17750,N_17540,N_17471);
nor U17751 (N_17751,N_17582,N_17453);
and U17752 (N_17752,N_17502,N_17552);
xnor U17753 (N_17753,N_17534,N_17539);
or U17754 (N_17754,N_17444,N_17540);
xor U17755 (N_17755,N_17490,N_17442);
or U17756 (N_17756,N_17550,N_17471);
and U17757 (N_17757,N_17527,N_17598);
xnor U17758 (N_17758,N_17520,N_17550);
xor U17759 (N_17759,N_17582,N_17462);
xor U17760 (N_17760,N_17656,N_17739);
or U17761 (N_17761,N_17711,N_17715);
nand U17762 (N_17762,N_17707,N_17696);
nor U17763 (N_17763,N_17678,N_17757);
xor U17764 (N_17764,N_17694,N_17751);
or U17765 (N_17765,N_17759,N_17753);
xor U17766 (N_17766,N_17755,N_17705);
xor U17767 (N_17767,N_17667,N_17601);
and U17768 (N_17768,N_17687,N_17653);
xor U17769 (N_17769,N_17735,N_17756);
xnor U17770 (N_17770,N_17740,N_17673);
nand U17771 (N_17771,N_17713,N_17622);
or U17772 (N_17772,N_17642,N_17691);
nand U17773 (N_17773,N_17638,N_17657);
nor U17774 (N_17774,N_17731,N_17664);
nor U17775 (N_17775,N_17719,N_17637);
or U17776 (N_17776,N_17723,N_17744);
xor U17777 (N_17777,N_17745,N_17714);
nand U17778 (N_17778,N_17615,N_17602);
nor U17779 (N_17779,N_17698,N_17724);
and U17780 (N_17780,N_17647,N_17750);
nor U17781 (N_17781,N_17618,N_17612);
nor U17782 (N_17782,N_17743,N_17649);
or U17783 (N_17783,N_17654,N_17725);
nor U17784 (N_17784,N_17669,N_17600);
or U17785 (N_17785,N_17662,N_17749);
xnor U17786 (N_17786,N_17604,N_17677);
xnor U17787 (N_17787,N_17644,N_17701);
and U17788 (N_17788,N_17730,N_17699);
or U17789 (N_17789,N_17611,N_17681);
nor U17790 (N_17790,N_17721,N_17617);
or U17791 (N_17791,N_17646,N_17729);
nor U17792 (N_17792,N_17732,N_17634);
or U17793 (N_17793,N_17629,N_17668);
and U17794 (N_17794,N_17613,N_17675);
nor U17795 (N_17795,N_17736,N_17660);
xor U17796 (N_17796,N_17748,N_17693);
nor U17797 (N_17797,N_17628,N_17663);
or U17798 (N_17798,N_17607,N_17625);
or U17799 (N_17799,N_17703,N_17605);
and U17800 (N_17800,N_17710,N_17686);
nand U17801 (N_17801,N_17722,N_17709);
or U17802 (N_17802,N_17754,N_17620);
nor U17803 (N_17803,N_17623,N_17674);
nand U17804 (N_17804,N_17648,N_17737);
and U17805 (N_17805,N_17643,N_17685);
and U17806 (N_17806,N_17733,N_17672);
nand U17807 (N_17807,N_17692,N_17684);
or U17808 (N_17808,N_17700,N_17614);
xnor U17809 (N_17809,N_17632,N_17631);
or U17810 (N_17810,N_17704,N_17608);
nor U17811 (N_17811,N_17697,N_17688);
nor U17812 (N_17812,N_17616,N_17658);
xnor U17813 (N_17813,N_17746,N_17727);
or U17814 (N_17814,N_17726,N_17640);
and U17815 (N_17815,N_17633,N_17627);
xor U17816 (N_17816,N_17650,N_17621);
or U17817 (N_17817,N_17747,N_17734);
nand U17818 (N_17818,N_17758,N_17670);
nand U17819 (N_17819,N_17651,N_17652);
nor U17820 (N_17820,N_17741,N_17720);
or U17821 (N_17821,N_17636,N_17639);
nor U17822 (N_17822,N_17738,N_17645);
or U17823 (N_17823,N_17717,N_17671);
or U17824 (N_17824,N_17603,N_17716);
nand U17825 (N_17825,N_17641,N_17702);
or U17826 (N_17826,N_17680,N_17661);
nor U17827 (N_17827,N_17706,N_17666);
and U17828 (N_17828,N_17708,N_17624);
and U17829 (N_17829,N_17690,N_17619);
nor U17830 (N_17830,N_17682,N_17659);
or U17831 (N_17831,N_17610,N_17606);
nand U17832 (N_17832,N_17695,N_17676);
nor U17833 (N_17833,N_17626,N_17635);
and U17834 (N_17834,N_17712,N_17655);
xnor U17835 (N_17835,N_17752,N_17728);
or U17836 (N_17836,N_17679,N_17742);
xor U17837 (N_17837,N_17683,N_17665);
xor U17838 (N_17838,N_17609,N_17630);
xnor U17839 (N_17839,N_17718,N_17689);
or U17840 (N_17840,N_17630,N_17642);
xnor U17841 (N_17841,N_17700,N_17620);
nor U17842 (N_17842,N_17730,N_17720);
or U17843 (N_17843,N_17640,N_17660);
and U17844 (N_17844,N_17659,N_17632);
nand U17845 (N_17845,N_17649,N_17722);
nor U17846 (N_17846,N_17718,N_17622);
xnor U17847 (N_17847,N_17700,N_17634);
xnor U17848 (N_17848,N_17658,N_17602);
or U17849 (N_17849,N_17725,N_17653);
or U17850 (N_17850,N_17628,N_17643);
nand U17851 (N_17851,N_17740,N_17720);
nor U17852 (N_17852,N_17709,N_17614);
and U17853 (N_17853,N_17678,N_17632);
and U17854 (N_17854,N_17729,N_17631);
nor U17855 (N_17855,N_17637,N_17715);
nand U17856 (N_17856,N_17710,N_17727);
nor U17857 (N_17857,N_17759,N_17610);
or U17858 (N_17858,N_17718,N_17748);
xor U17859 (N_17859,N_17623,N_17622);
or U17860 (N_17860,N_17726,N_17677);
and U17861 (N_17861,N_17610,N_17703);
and U17862 (N_17862,N_17616,N_17702);
or U17863 (N_17863,N_17734,N_17742);
xor U17864 (N_17864,N_17644,N_17684);
nor U17865 (N_17865,N_17754,N_17689);
nor U17866 (N_17866,N_17631,N_17677);
and U17867 (N_17867,N_17657,N_17664);
nand U17868 (N_17868,N_17707,N_17612);
nand U17869 (N_17869,N_17734,N_17687);
or U17870 (N_17870,N_17686,N_17687);
and U17871 (N_17871,N_17613,N_17667);
and U17872 (N_17872,N_17714,N_17708);
nand U17873 (N_17873,N_17642,N_17659);
and U17874 (N_17874,N_17704,N_17708);
nor U17875 (N_17875,N_17728,N_17691);
nand U17876 (N_17876,N_17629,N_17667);
and U17877 (N_17877,N_17694,N_17635);
or U17878 (N_17878,N_17728,N_17646);
xor U17879 (N_17879,N_17754,N_17713);
xor U17880 (N_17880,N_17621,N_17730);
or U17881 (N_17881,N_17744,N_17613);
xor U17882 (N_17882,N_17647,N_17622);
xnor U17883 (N_17883,N_17652,N_17639);
or U17884 (N_17884,N_17609,N_17637);
or U17885 (N_17885,N_17682,N_17617);
or U17886 (N_17886,N_17688,N_17728);
and U17887 (N_17887,N_17614,N_17604);
nand U17888 (N_17888,N_17672,N_17614);
and U17889 (N_17889,N_17631,N_17687);
nor U17890 (N_17890,N_17695,N_17631);
nor U17891 (N_17891,N_17746,N_17693);
or U17892 (N_17892,N_17740,N_17612);
or U17893 (N_17893,N_17691,N_17651);
nand U17894 (N_17894,N_17729,N_17691);
nand U17895 (N_17895,N_17682,N_17725);
nand U17896 (N_17896,N_17733,N_17675);
nor U17897 (N_17897,N_17649,N_17718);
and U17898 (N_17898,N_17757,N_17699);
or U17899 (N_17899,N_17699,N_17660);
or U17900 (N_17900,N_17658,N_17618);
xor U17901 (N_17901,N_17701,N_17622);
nor U17902 (N_17902,N_17666,N_17617);
xor U17903 (N_17903,N_17620,N_17606);
and U17904 (N_17904,N_17720,N_17639);
nor U17905 (N_17905,N_17755,N_17758);
or U17906 (N_17906,N_17706,N_17670);
or U17907 (N_17907,N_17737,N_17606);
nand U17908 (N_17908,N_17640,N_17678);
and U17909 (N_17909,N_17632,N_17743);
or U17910 (N_17910,N_17614,N_17748);
xnor U17911 (N_17911,N_17727,N_17644);
nand U17912 (N_17912,N_17645,N_17712);
or U17913 (N_17913,N_17673,N_17606);
nand U17914 (N_17914,N_17660,N_17624);
and U17915 (N_17915,N_17637,N_17622);
and U17916 (N_17916,N_17664,N_17602);
or U17917 (N_17917,N_17646,N_17645);
or U17918 (N_17918,N_17716,N_17739);
xnor U17919 (N_17919,N_17680,N_17730);
and U17920 (N_17920,N_17839,N_17832);
xnor U17921 (N_17921,N_17845,N_17835);
nand U17922 (N_17922,N_17770,N_17858);
and U17923 (N_17923,N_17802,N_17906);
or U17924 (N_17924,N_17890,N_17883);
xor U17925 (N_17925,N_17813,N_17804);
nor U17926 (N_17926,N_17903,N_17869);
and U17927 (N_17927,N_17812,N_17917);
nor U17928 (N_17928,N_17901,N_17766);
or U17929 (N_17929,N_17829,N_17786);
or U17930 (N_17930,N_17795,N_17817);
nand U17931 (N_17931,N_17872,N_17768);
nor U17932 (N_17932,N_17761,N_17871);
nand U17933 (N_17933,N_17873,N_17898);
nor U17934 (N_17934,N_17852,N_17830);
nand U17935 (N_17935,N_17821,N_17851);
or U17936 (N_17936,N_17831,N_17911);
and U17937 (N_17937,N_17876,N_17914);
nor U17938 (N_17938,N_17815,N_17806);
or U17939 (N_17939,N_17865,N_17913);
nor U17940 (N_17940,N_17788,N_17767);
and U17941 (N_17941,N_17827,N_17916);
xor U17942 (N_17942,N_17868,N_17819);
nand U17943 (N_17943,N_17822,N_17790);
and U17944 (N_17944,N_17769,N_17863);
xor U17945 (N_17945,N_17820,N_17881);
xor U17946 (N_17946,N_17789,N_17902);
and U17947 (N_17947,N_17785,N_17884);
and U17948 (N_17948,N_17774,N_17895);
nand U17949 (N_17949,N_17919,N_17844);
nand U17950 (N_17950,N_17866,N_17824);
and U17951 (N_17951,N_17885,N_17826);
nand U17952 (N_17952,N_17892,N_17896);
or U17953 (N_17953,N_17814,N_17847);
or U17954 (N_17954,N_17860,N_17915);
and U17955 (N_17955,N_17909,N_17805);
nand U17956 (N_17956,N_17803,N_17772);
nand U17957 (N_17957,N_17838,N_17807);
and U17958 (N_17958,N_17801,N_17879);
nand U17959 (N_17959,N_17837,N_17793);
xnor U17960 (N_17960,N_17808,N_17777);
nand U17961 (N_17961,N_17787,N_17862);
nor U17962 (N_17962,N_17904,N_17800);
nand U17963 (N_17963,N_17842,N_17825);
and U17964 (N_17964,N_17854,N_17849);
and U17965 (N_17965,N_17810,N_17784);
and U17966 (N_17966,N_17828,N_17875);
and U17967 (N_17967,N_17908,N_17877);
or U17968 (N_17968,N_17763,N_17891);
nand U17969 (N_17969,N_17771,N_17781);
and U17970 (N_17970,N_17840,N_17765);
nand U17971 (N_17971,N_17846,N_17823);
or U17972 (N_17972,N_17912,N_17870);
or U17973 (N_17973,N_17809,N_17782);
xnor U17974 (N_17974,N_17880,N_17762);
nor U17975 (N_17975,N_17794,N_17843);
xnor U17976 (N_17976,N_17836,N_17773);
xor U17977 (N_17977,N_17893,N_17816);
or U17978 (N_17978,N_17867,N_17859);
nand U17979 (N_17979,N_17888,N_17811);
xor U17980 (N_17980,N_17897,N_17841);
or U17981 (N_17981,N_17900,N_17882);
xor U17982 (N_17982,N_17760,N_17894);
and U17983 (N_17983,N_17899,N_17797);
or U17984 (N_17984,N_17848,N_17855);
nor U17985 (N_17985,N_17799,N_17864);
or U17986 (N_17986,N_17779,N_17798);
or U17987 (N_17987,N_17764,N_17918);
nor U17988 (N_17988,N_17775,N_17791);
and U17989 (N_17989,N_17886,N_17850);
xnor U17990 (N_17990,N_17905,N_17874);
nor U17991 (N_17991,N_17833,N_17856);
and U17992 (N_17992,N_17792,N_17796);
xnor U17993 (N_17993,N_17889,N_17818);
xor U17994 (N_17994,N_17887,N_17780);
nor U17995 (N_17995,N_17857,N_17853);
nor U17996 (N_17996,N_17878,N_17776);
or U17997 (N_17997,N_17861,N_17778);
nor U17998 (N_17998,N_17907,N_17783);
xor U17999 (N_17999,N_17834,N_17910);
nor U18000 (N_18000,N_17774,N_17790);
xnor U18001 (N_18001,N_17877,N_17887);
or U18002 (N_18002,N_17785,N_17910);
or U18003 (N_18003,N_17783,N_17794);
nand U18004 (N_18004,N_17784,N_17857);
and U18005 (N_18005,N_17851,N_17767);
xor U18006 (N_18006,N_17918,N_17908);
xnor U18007 (N_18007,N_17892,N_17874);
and U18008 (N_18008,N_17833,N_17825);
xor U18009 (N_18009,N_17780,N_17797);
xor U18010 (N_18010,N_17903,N_17894);
xor U18011 (N_18011,N_17765,N_17834);
xor U18012 (N_18012,N_17915,N_17900);
or U18013 (N_18013,N_17769,N_17856);
xnor U18014 (N_18014,N_17872,N_17859);
and U18015 (N_18015,N_17788,N_17906);
and U18016 (N_18016,N_17824,N_17791);
nor U18017 (N_18017,N_17792,N_17910);
xnor U18018 (N_18018,N_17897,N_17833);
nor U18019 (N_18019,N_17876,N_17772);
nor U18020 (N_18020,N_17850,N_17863);
nor U18021 (N_18021,N_17763,N_17879);
xnor U18022 (N_18022,N_17817,N_17796);
xor U18023 (N_18023,N_17893,N_17899);
nor U18024 (N_18024,N_17865,N_17898);
and U18025 (N_18025,N_17778,N_17833);
and U18026 (N_18026,N_17776,N_17898);
nand U18027 (N_18027,N_17869,N_17817);
and U18028 (N_18028,N_17866,N_17788);
nor U18029 (N_18029,N_17785,N_17829);
and U18030 (N_18030,N_17779,N_17835);
xor U18031 (N_18031,N_17775,N_17833);
and U18032 (N_18032,N_17794,N_17910);
and U18033 (N_18033,N_17908,N_17792);
nand U18034 (N_18034,N_17803,N_17795);
xnor U18035 (N_18035,N_17810,N_17827);
nand U18036 (N_18036,N_17781,N_17835);
or U18037 (N_18037,N_17902,N_17808);
and U18038 (N_18038,N_17788,N_17869);
or U18039 (N_18039,N_17832,N_17878);
nor U18040 (N_18040,N_17805,N_17770);
nand U18041 (N_18041,N_17898,N_17822);
or U18042 (N_18042,N_17872,N_17871);
nand U18043 (N_18043,N_17845,N_17789);
nand U18044 (N_18044,N_17807,N_17859);
and U18045 (N_18045,N_17861,N_17849);
and U18046 (N_18046,N_17883,N_17814);
and U18047 (N_18047,N_17793,N_17869);
nor U18048 (N_18048,N_17898,N_17761);
nand U18049 (N_18049,N_17886,N_17849);
nand U18050 (N_18050,N_17804,N_17868);
or U18051 (N_18051,N_17881,N_17847);
xnor U18052 (N_18052,N_17828,N_17901);
nor U18053 (N_18053,N_17877,N_17899);
nor U18054 (N_18054,N_17774,N_17824);
and U18055 (N_18055,N_17839,N_17901);
or U18056 (N_18056,N_17809,N_17824);
xor U18057 (N_18057,N_17808,N_17812);
nor U18058 (N_18058,N_17804,N_17794);
or U18059 (N_18059,N_17804,N_17774);
xnor U18060 (N_18060,N_17894,N_17895);
nand U18061 (N_18061,N_17807,N_17900);
nor U18062 (N_18062,N_17863,N_17829);
nand U18063 (N_18063,N_17802,N_17907);
nand U18064 (N_18064,N_17780,N_17789);
nor U18065 (N_18065,N_17912,N_17841);
xor U18066 (N_18066,N_17768,N_17790);
nand U18067 (N_18067,N_17873,N_17882);
nand U18068 (N_18068,N_17802,N_17822);
or U18069 (N_18069,N_17821,N_17909);
or U18070 (N_18070,N_17787,N_17871);
nand U18071 (N_18071,N_17811,N_17789);
nand U18072 (N_18072,N_17897,N_17780);
xnor U18073 (N_18073,N_17859,N_17800);
nand U18074 (N_18074,N_17788,N_17822);
and U18075 (N_18075,N_17901,N_17836);
and U18076 (N_18076,N_17773,N_17762);
xnor U18077 (N_18077,N_17839,N_17898);
or U18078 (N_18078,N_17818,N_17822);
xnor U18079 (N_18079,N_17903,N_17863);
xnor U18080 (N_18080,N_17995,N_18014);
nor U18081 (N_18081,N_18048,N_17950);
nor U18082 (N_18082,N_18045,N_17926);
and U18083 (N_18083,N_18039,N_17967);
nand U18084 (N_18084,N_17984,N_18059);
xor U18085 (N_18085,N_18035,N_17954);
nor U18086 (N_18086,N_18078,N_18023);
nor U18087 (N_18087,N_17977,N_18053);
nor U18088 (N_18088,N_17932,N_17951);
and U18089 (N_18089,N_18060,N_18016);
or U18090 (N_18090,N_17979,N_18062);
nand U18091 (N_18091,N_18019,N_17968);
and U18092 (N_18092,N_18012,N_17961);
or U18093 (N_18093,N_17945,N_17982);
nand U18094 (N_18094,N_18033,N_18057);
and U18095 (N_18095,N_18043,N_17929);
xnor U18096 (N_18096,N_18038,N_17974);
or U18097 (N_18097,N_18052,N_18024);
nor U18098 (N_18098,N_18037,N_18027);
nand U18099 (N_18099,N_18074,N_17994);
and U18100 (N_18100,N_18065,N_18069);
or U18101 (N_18101,N_17920,N_18032);
nor U18102 (N_18102,N_17940,N_18070);
nor U18103 (N_18103,N_17997,N_18010);
nor U18104 (N_18104,N_18058,N_17937);
or U18105 (N_18105,N_17957,N_18034);
or U18106 (N_18106,N_18073,N_17980);
and U18107 (N_18107,N_17975,N_18063);
and U18108 (N_18108,N_17966,N_18046);
nor U18109 (N_18109,N_17987,N_18077);
nand U18110 (N_18110,N_17928,N_17962);
xor U18111 (N_18111,N_18008,N_17973);
or U18112 (N_18112,N_18018,N_18005);
xnor U18113 (N_18113,N_17934,N_17930);
and U18114 (N_18114,N_18009,N_17993);
nand U18115 (N_18115,N_17996,N_18000);
nand U18116 (N_18116,N_17921,N_18072);
nand U18117 (N_18117,N_17981,N_17960);
nand U18118 (N_18118,N_17925,N_18028);
xnor U18119 (N_18119,N_17956,N_17985);
xor U18120 (N_18120,N_17958,N_17941);
nor U18121 (N_18121,N_17988,N_17991);
xnor U18122 (N_18122,N_18029,N_17936);
nor U18123 (N_18123,N_17986,N_18050);
nor U18124 (N_18124,N_18064,N_18056);
and U18125 (N_18125,N_18079,N_17922);
and U18126 (N_18126,N_17969,N_18025);
xnor U18127 (N_18127,N_17992,N_17998);
nand U18128 (N_18128,N_18007,N_18020);
and U18129 (N_18129,N_18054,N_17933);
or U18130 (N_18130,N_18001,N_17959);
and U18131 (N_18131,N_17976,N_18026);
or U18132 (N_18132,N_18041,N_17949);
nand U18133 (N_18133,N_17965,N_17952);
xor U18134 (N_18134,N_18067,N_18068);
or U18135 (N_18135,N_18030,N_18051);
xnor U18136 (N_18136,N_18002,N_18011);
nand U18137 (N_18137,N_18055,N_17948);
and U18138 (N_18138,N_17990,N_17946);
and U18139 (N_18139,N_18044,N_18004);
and U18140 (N_18140,N_17970,N_17955);
nand U18141 (N_18141,N_17935,N_17938);
xor U18142 (N_18142,N_17944,N_18022);
or U18143 (N_18143,N_17924,N_18021);
nand U18144 (N_18144,N_17964,N_18049);
nand U18145 (N_18145,N_17989,N_18040);
or U18146 (N_18146,N_17983,N_18061);
or U18147 (N_18147,N_17923,N_17942);
xnor U18148 (N_18148,N_18015,N_18047);
or U18149 (N_18149,N_18006,N_17947);
nor U18150 (N_18150,N_17943,N_18003);
xor U18151 (N_18151,N_18066,N_18071);
and U18152 (N_18152,N_18036,N_17972);
nand U18153 (N_18153,N_17999,N_18017);
nand U18154 (N_18154,N_17953,N_18013);
xnor U18155 (N_18155,N_17971,N_18042);
xnor U18156 (N_18156,N_18076,N_17931);
xor U18157 (N_18157,N_17939,N_17963);
or U18158 (N_18158,N_18075,N_17927);
nor U18159 (N_18159,N_17978,N_18031);
nand U18160 (N_18160,N_18056,N_17935);
or U18161 (N_18161,N_17949,N_18020);
and U18162 (N_18162,N_18058,N_18013);
and U18163 (N_18163,N_17924,N_18017);
or U18164 (N_18164,N_18077,N_18073);
nor U18165 (N_18165,N_17978,N_17948);
or U18166 (N_18166,N_17945,N_18062);
nand U18167 (N_18167,N_18026,N_17920);
and U18168 (N_18168,N_18028,N_17953);
xor U18169 (N_18169,N_17957,N_17981);
nor U18170 (N_18170,N_18008,N_17966);
nor U18171 (N_18171,N_17928,N_18005);
nand U18172 (N_18172,N_17980,N_17921);
and U18173 (N_18173,N_17961,N_17942);
and U18174 (N_18174,N_17995,N_17969);
and U18175 (N_18175,N_18027,N_17980);
and U18176 (N_18176,N_18030,N_17926);
nand U18177 (N_18177,N_18071,N_17984);
nor U18178 (N_18178,N_17979,N_17981);
and U18179 (N_18179,N_17929,N_18008);
or U18180 (N_18180,N_18050,N_18053);
nand U18181 (N_18181,N_18040,N_18029);
nor U18182 (N_18182,N_17949,N_17957);
nand U18183 (N_18183,N_18066,N_18060);
or U18184 (N_18184,N_18051,N_18068);
nand U18185 (N_18185,N_18020,N_18038);
xor U18186 (N_18186,N_17988,N_18016);
nor U18187 (N_18187,N_17953,N_18042);
or U18188 (N_18188,N_18013,N_18075);
nand U18189 (N_18189,N_18014,N_18022);
or U18190 (N_18190,N_18042,N_17940);
and U18191 (N_18191,N_18039,N_17989);
nand U18192 (N_18192,N_18003,N_17925);
nand U18193 (N_18193,N_17927,N_18019);
nor U18194 (N_18194,N_17966,N_18060);
xnor U18195 (N_18195,N_17933,N_18073);
or U18196 (N_18196,N_18052,N_17958);
or U18197 (N_18197,N_17961,N_17980);
nor U18198 (N_18198,N_17988,N_18019);
or U18199 (N_18199,N_17923,N_17946);
nor U18200 (N_18200,N_17926,N_18007);
or U18201 (N_18201,N_18031,N_17935);
xnor U18202 (N_18202,N_18041,N_17928);
nand U18203 (N_18203,N_17923,N_18014);
xor U18204 (N_18204,N_18034,N_18036);
nand U18205 (N_18205,N_17987,N_17926);
and U18206 (N_18206,N_17998,N_18066);
and U18207 (N_18207,N_18048,N_18034);
and U18208 (N_18208,N_17992,N_17956);
nand U18209 (N_18209,N_18008,N_17964);
nor U18210 (N_18210,N_18001,N_18035);
nand U18211 (N_18211,N_18072,N_18029);
or U18212 (N_18212,N_18066,N_18013);
nand U18213 (N_18213,N_17949,N_17938);
nor U18214 (N_18214,N_18038,N_17995);
xor U18215 (N_18215,N_18039,N_18013);
and U18216 (N_18216,N_17984,N_17935);
nor U18217 (N_18217,N_18002,N_18059);
xnor U18218 (N_18218,N_17948,N_18030);
or U18219 (N_18219,N_18014,N_18075);
nand U18220 (N_18220,N_18036,N_17996);
and U18221 (N_18221,N_18059,N_18063);
nand U18222 (N_18222,N_17934,N_17998);
and U18223 (N_18223,N_18019,N_18075);
nand U18224 (N_18224,N_18028,N_18021);
nand U18225 (N_18225,N_18059,N_17999);
nand U18226 (N_18226,N_17929,N_18010);
xnor U18227 (N_18227,N_17961,N_18005);
or U18228 (N_18228,N_17971,N_18020);
xnor U18229 (N_18229,N_18057,N_17951);
xor U18230 (N_18230,N_17970,N_17933);
or U18231 (N_18231,N_17959,N_18068);
nor U18232 (N_18232,N_17922,N_18076);
or U18233 (N_18233,N_18022,N_18006);
xnor U18234 (N_18234,N_18025,N_17921);
xnor U18235 (N_18235,N_17941,N_17953);
and U18236 (N_18236,N_17948,N_17934);
or U18237 (N_18237,N_18042,N_18027);
nor U18238 (N_18238,N_18079,N_17991);
and U18239 (N_18239,N_18018,N_18073);
or U18240 (N_18240,N_18164,N_18237);
xor U18241 (N_18241,N_18147,N_18209);
and U18242 (N_18242,N_18190,N_18116);
and U18243 (N_18243,N_18191,N_18127);
and U18244 (N_18244,N_18124,N_18146);
nor U18245 (N_18245,N_18125,N_18167);
and U18246 (N_18246,N_18133,N_18180);
or U18247 (N_18247,N_18122,N_18213);
nor U18248 (N_18248,N_18169,N_18115);
nor U18249 (N_18249,N_18113,N_18210);
and U18250 (N_18250,N_18198,N_18212);
nand U18251 (N_18251,N_18231,N_18086);
and U18252 (N_18252,N_18188,N_18087);
xor U18253 (N_18253,N_18197,N_18138);
and U18254 (N_18254,N_18107,N_18189);
nor U18255 (N_18255,N_18217,N_18101);
nand U18256 (N_18256,N_18193,N_18238);
or U18257 (N_18257,N_18137,N_18083);
and U18258 (N_18258,N_18159,N_18131);
nor U18259 (N_18259,N_18218,N_18153);
or U18260 (N_18260,N_18096,N_18233);
nor U18261 (N_18261,N_18216,N_18226);
and U18262 (N_18262,N_18187,N_18205);
nor U18263 (N_18263,N_18104,N_18091);
xor U18264 (N_18264,N_18183,N_18105);
xor U18265 (N_18265,N_18128,N_18223);
xor U18266 (N_18266,N_18139,N_18150);
xor U18267 (N_18267,N_18160,N_18173);
nor U18268 (N_18268,N_18082,N_18102);
nor U18269 (N_18269,N_18080,N_18154);
xor U18270 (N_18270,N_18219,N_18103);
nor U18271 (N_18271,N_18228,N_18156);
and U18272 (N_18272,N_18192,N_18089);
and U18273 (N_18273,N_18204,N_18227);
xor U18274 (N_18274,N_18157,N_18222);
nor U18275 (N_18275,N_18140,N_18119);
nand U18276 (N_18276,N_18170,N_18081);
nor U18277 (N_18277,N_18232,N_18179);
nand U18278 (N_18278,N_18144,N_18126);
nor U18279 (N_18279,N_18224,N_18120);
or U18280 (N_18280,N_18200,N_18136);
and U18281 (N_18281,N_18098,N_18203);
nand U18282 (N_18282,N_18172,N_18130);
xnor U18283 (N_18283,N_18141,N_18099);
or U18284 (N_18284,N_18132,N_18129);
and U18285 (N_18285,N_18100,N_18201);
and U18286 (N_18286,N_18094,N_18143);
nor U18287 (N_18287,N_18109,N_18106);
and U18288 (N_18288,N_18110,N_18239);
nor U18289 (N_18289,N_18234,N_18084);
and U18290 (N_18290,N_18090,N_18134);
nor U18291 (N_18291,N_18162,N_18117);
nand U18292 (N_18292,N_18155,N_18148);
nor U18293 (N_18293,N_18114,N_18161);
xor U18294 (N_18294,N_18158,N_18166);
xnor U18295 (N_18295,N_18165,N_18206);
or U18296 (N_18296,N_18152,N_18085);
or U18297 (N_18297,N_18168,N_18185);
xnor U18298 (N_18298,N_18194,N_18184);
xnor U18299 (N_18299,N_18118,N_18108);
nor U18300 (N_18300,N_18178,N_18214);
and U18301 (N_18301,N_18182,N_18171);
nor U18302 (N_18302,N_18195,N_18221);
and U18303 (N_18303,N_18111,N_18145);
nand U18304 (N_18304,N_18215,N_18095);
nand U18305 (N_18305,N_18220,N_18225);
and U18306 (N_18306,N_18229,N_18175);
nor U18307 (N_18307,N_18207,N_18199);
nor U18308 (N_18308,N_18177,N_18202);
or U18309 (N_18309,N_18112,N_18211);
and U18310 (N_18310,N_18121,N_18230);
nand U18311 (N_18311,N_18088,N_18142);
and U18312 (N_18312,N_18208,N_18163);
xor U18313 (N_18313,N_18235,N_18174);
and U18314 (N_18314,N_18149,N_18123);
nor U18315 (N_18315,N_18135,N_18097);
xor U18316 (N_18316,N_18176,N_18092);
xnor U18317 (N_18317,N_18181,N_18093);
or U18318 (N_18318,N_18196,N_18186);
nand U18319 (N_18319,N_18236,N_18151);
or U18320 (N_18320,N_18135,N_18136);
and U18321 (N_18321,N_18139,N_18163);
xnor U18322 (N_18322,N_18186,N_18210);
and U18323 (N_18323,N_18188,N_18140);
or U18324 (N_18324,N_18138,N_18180);
and U18325 (N_18325,N_18208,N_18125);
and U18326 (N_18326,N_18109,N_18126);
nor U18327 (N_18327,N_18080,N_18100);
or U18328 (N_18328,N_18232,N_18205);
nand U18329 (N_18329,N_18173,N_18187);
or U18330 (N_18330,N_18198,N_18191);
or U18331 (N_18331,N_18099,N_18082);
xor U18332 (N_18332,N_18108,N_18119);
nor U18333 (N_18333,N_18237,N_18092);
nor U18334 (N_18334,N_18189,N_18182);
and U18335 (N_18335,N_18099,N_18140);
or U18336 (N_18336,N_18089,N_18216);
nor U18337 (N_18337,N_18168,N_18222);
nand U18338 (N_18338,N_18237,N_18219);
xnor U18339 (N_18339,N_18097,N_18237);
nand U18340 (N_18340,N_18144,N_18106);
nand U18341 (N_18341,N_18214,N_18209);
and U18342 (N_18342,N_18180,N_18179);
xnor U18343 (N_18343,N_18167,N_18215);
or U18344 (N_18344,N_18112,N_18214);
or U18345 (N_18345,N_18128,N_18135);
and U18346 (N_18346,N_18096,N_18148);
nand U18347 (N_18347,N_18234,N_18096);
nor U18348 (N_18348,N_18089,N_18146);
xor U18349 (N_18349,N_18226,N_18129);
or U18350 (N_18350,N_18222,N_18172);
nor U18351 (N_18351,N_18192,N_18129);
nor U18352 (N_18352,N_18148,N_18214);
and U18353 (N_18353,N_18177,N_18205);
xnor U18354 (N_18354,N_18216,N_18206);
nand U18355 (N_18355,N_18174,N_18148);
nand U18356 (N_18356,N_18145,N_18205);
and U18357 (N_18357,N_18210,N_18143);
nor U18358 (N_18358,N_18127,N_18154);
nor U18359 (N_18359,N_18138,N_18235);
xor U18360 (N_18360,N_18098,N_18082);
xor U18361 (N_18361,N_18190,N_18139);
nor U18362 (N_18362,N_18175,N_18125);
xor U18363 (N_18363,N_18145,N_18130);
nand U18364 (N_18364,N_18181,N_18205);
or U18365 (N_18365,N_18221,N_18178);
or U18366 (N_18366,N_18166,N_18184);
xnor U18367 (N_18367,N_18105,N_18186);
or U18368 (N_18368,N_18201,N_18187);
nor U18369 (N_18369,N_18201,N_18123);
xor U18370 (N_18370,N_18236,N_18226);
or U18371 (N_18371,N_18130,N_18229);
xnor U18372 (N_18372,N_18137,N_18219);
or U18373 (N_18373,N_18083,N_18116);
and U18374 (N_18374,N_18209,N_18213);
nand U18375 (N_18375,N_18107,N_18162);
nand U18376 (N_18376,N_18083,N_18128);
nor U18377 (N_18377,N_18144,N_18148);
nor U18378 (N_18378,N_18081,N_18235);
nor U18379 (N_18379,N_18176,N_18112);
and U18380 (N_18380,N_18123,N_18151);
or U18381 (N_18381,N_18167,N_18164);
xnor U18382 (N_18382,N_18131,N_18139);
and U18383 (N_18383,N_18082,N_18236);
and U18384 (N_18384,N_18236,N_18139);
nand U18385 (N_18385,N_18084,N_18198);
xor U18386 (N_18386,N_18203,N_18096);
and U18387 (N_18387,N_18236,N_18183);
and U18388 (N_18388,N_18187,N_18220);
nand U18389 (N_18389,N_18119,N_18123);
nor U18390 (N_18390,N_18172,N_18163);
xnor U18391 (N_18391,N_18159,N_18125);
nand U18392 (N_18392,N_18092,N_18230);
xnor U18393 (N_18393,N_18095,N_18114);
xnor U18394 (N_18394,N_18238,N_18143);
nor U18395 (N_18395,N_18181,N_18172);
xor U18396 (N_18396,N_18226,N_18091);
or U18397 (N_18397,N_18102,N_18127);
and U18398 (N_18398,N_18177,N_18146);
xor U18399 (N_18399,N_18190,N_18124);
nand U18400 (N_18400,N_18399,N_18374);
and U18401 (N_18401,N_18349,N_18253);
xnor U18402 (N_18402,N_18257,N_18284);
xor U18403 (N_18403,N_18323,N_18328);
and U18404 (N_18404,N_18268,N_18281);
nor U18405 (N_18405,N_18321,N_18370);
nand U18406 (N_18406,N_18359,N_18299);
or U18407 (N_18407,N_18337,N_18397);
or U18408 (N_18408,N_18251,N_18311);
nand U18409 (N_18409,N_18378,N_18394);
xor U18410 (N_18410,N_18391,N_18388);
xor U18411 (N_18411,N_18269,N_18316);
nand U18412 (N_18412,N_18304,N_18305);
xnor U18413 (N_18413,N_18243,N_18271);
nand U18414 (N_18414,N_18315,N_18261);
xnor U18415 (N_18415,N_18373,N_18355);
nor U18416 (N_18416,N_18371,N_18390);
xor U18417 (N_18417,N_18358,N_18283);
and U18418 (N_18418,N_18276,N_18332);
nor U18419 (N_18419,N_18350,N_18383);
nor U18420 (N_18420,N_18326,N_18293);
nor U18421 (N_18421,N_18295,N_18317);
xnor U18422 (N_18422,N_18312,N_18335);
xor U18423 (N_18423,N_18297,N_18354);
nand U18424 (N_18424,N_18396,N_18372);
nand U18425 (N_18425,N_18338,N_18368);
or U18426 (N_18426,N_18260,N_18292);
and U18427 (N_18427,N_18398,N_18365);
xnor U18428 (N_18428,N_18314,N_18362);
and U18429 (N_18429,N_18348,N_18262);
xor U18430 (N_18430,N_18353,N_18385);
or U18431 (N_18431,N_18301,N_18366);
nor U18432 (N_18432,N_18298,N_18361);
nand U18433 (N_18433,N_18287,N_18320);
xor U18434 (N_18434,N_18346,N_18329);
xor U18435 (N_18435,N_18351,N_18306);
nor U18436 (N_18436,N_18339,N_18267);
xor U18437 (N_18437,N_18270,N_18303);
and U18438 (N_18438,N_18285,N_18254);
and U18439 (N_18439,N_18322,N_18341);
or U18440 (N_18440,N_18245,N_18249);
nor U18441 (N_18441,N_18296,N_18376);
nor U18442 (N_18442,N_18282,N_18264);
and U18443 (N_18443,N_18291,N_18302);
and U18444 (N_18444,N_18381,N_18336);
nand U18445 (N_18445,N_18278,N_18308);
or U18446 (N_18446,N_18369,N_18246);
xor U18447 (N_18447,N_18356,N_18380);
or U18448 (N_18448,N_18265,N_18334);
xnor U18449 (N_18449,N_18343,N_18333);
nand U18450 (N_18450,N_18392,N_18247);
nor U18451 (N_18451,N_18273,N_18263);
or U18452 (N_18452,N_18331,N_18255);
and U18453 (N_18453,N_18286,N_18364);
nor U18454 (N_18454,N_18330,N_18300);
nor U18455 (N_18455,N_18244,N_18279);
nand U18456 (N_18456,N_18241,N_18250);
xnor U18457 (N_18457,N_18325,N_18363);
nor U18458 (N_18458,N_18290,N_18375);
and U18459 (N_18459,N_18387,N_18318);
nor U18460 (N_18460,N_18344,N_18389);
and U18461 (N_18461,N_18324,N_18340);
and U18462 (N_18462,N_18252,N_18377);
and U18463 (N_18463,N_18289,N_18395);
xor U18464 (N_18464,N_18347,N_18275);
xor U18465 (N_18465,N_18242,N_18310);
or U18466 (N_18466,N_18367,N_18357);
nand U18467 (N_18467,N_18342,N_18386);
and U18468 (N_18468,N_18319,N_18266);
nor U18469 (N_18469,N_18327,N_18379);
nand U18470 (N_18470,N_18384,N_18345);
nor U18471 (N_18471,N_18307,N_18258);
and U18472 (N_18472,N_18280,N_18309);
xnor U18473 (N_18473,N_18294,N_18288);
or U18474 (N_18474,N_18382,N_18393);
nand U18475 (N_18475,N_18352,N_18274);
and U18476 (N_18476,N_18277,N_18240);
nand U18477 (N_18477,N_18248,N_18360);
nand U18478 (N_18478,N_18256,N_18313);
xor U18479 (N_18479,N_18272,N_18259);
xor U18480 (N_18480,N_18352,N_18391);
nor U18481 (N_18481,N_18280,N_18356);
xnor U18482 (N_18482,N_18259,N_18319);
or U18483 (N_18483,N_18341,N_18244);
or U18484 (N_18484,N_18365,N_18374);
and U18485 (N_18485,N_18379,N_18325);
and U18486 (N_18486,N_18322,N_18291);
or U18487 (N_18487,N_18340,N_18259);
or U18488 (N_18488,N_18254,N_18396);
xor U18489 (N_18489,N_18341,N_18309);
nor U18490 (N_18490,N_18371,N_18255);
or U18491 (N_18491,N_18265,N_18343);
nand U18492 (N_18492,N_18244,N_18262);
nand U18493 (N_18493,N_18262,N_18391);
nand U18494 (N_18494,N_18345,N_18268);
and U18495 (N_18495,N_18263,N_18342);
and U18496 (N_18496,N_18375,N_18310);
nor U18497 (N_18497,N_18365,N_18294);
nor U18498 (N_18498,N_18275,N_18319);
nor U18499 (N_18499,N_18325,N_18241);
nor U18500 (N_18500,N_18289,N_18397);
nor U18501 (N_18501,N_18286,N_18387);
or U18502 (N_18502,N_18339,N_18280);
or U18503 (N_18503,N_18333,N_18320);
nand U18504 (N_18504,N_18272,N_18340);
nor U18505 (N_18505,N_18379,N_18340);
nor U18506 (N_18506,N_18356,N_18277);
nand U18507 (N_18507,N_18389,N_18241);
nor U18508 (N_18508,N_18373,N_18316);
nor U18509 (N_18509,N_18264,N_18363);
or U18510 (N_18510,N_18301,N_18281);
xnor U18511 (N_18511,N_18298,N_18329);
or U18512 (N_18512,N_18257,N_18396);
nand U18513 (N_18513,N_18261,N_18348);
nor U18514 (N_18514,N_18368,N_18394);
xor U18515 (N_18515,N_18314,N_18257);
nor U18516 (N_18516,N_18367,N_18398);
nor U18517 (N_18517,N_18380,N_18316);
nor U18518 (N_18518,N_18348,N_18347);
and U18519 (N_18519,N_18264,N_18280);
and U18520 (N_18520,N_18399,N_18335);
xnor U18521 (N_18521,N_18357,N_18259);
and U18522 (N_18522,N_18372,N_18367);
or U18523 (N_18523,N_18348,N_18353);
and U18524 (N_18524,N_18327,N_18370);
and U18525 (N_18525,N_18339,N_18316);
and U18526 (N_18526,N_18256,N_18356);
and U18527 (N_18527,N_18296,N_18291);
or U18528 (N_18528,N_18299,N_18327);
nor U18529 (N_18529,N_18351,N_18316);
nor U18530 (N_18530,N_18384,N_18286);
nand U18531 (N_18531,N_18305,N_18271);
and U18532 (N_18532,N_18318,N_18290);
xor U18533 (N_18533,N_18316,N_18383);
and U18534 (N_18534,N_18304,N_18269);
and U18535 (N_18535,N_18281,N_18305);
xnor U18536 (N_18536,N_18352,N_18286);
xor U18537 (N_18537,N_18329,N_18353);
nor U18538 (N_18538,N_18254,N_18325);
or U18539 (N_18539,N_18399,N_18362);
xnor U18540 (N_18540,N_18381,N_18296);
xor U18541 (N_18541,N_18310,N_18294);
nor U18542 (N_18542,N_18397,N_18315);
xor U18543 (N_18543,N_18246,N_18376);
or U18544 (N_18544,N_18249,N_18376);
nand U18545 (N_18545,N_18321,N_18388);
nor U18546 (N_18546,N_18344,N_18274);
nor U18547 (N_18547,N_18336,N_18341);
and U18548 (N_18548,N_18305,N_18292);
and U18549 (N_18549,N_18259,N_18254);
and U18550 (N_18550,N_18269,N_18252);
nor U18551 (N_18551,N_18367,N_18362);
nor U18552 (N_18552,N_18298,N_18393);
or U18553 (N_18553,N_18336,N_18338);
or U18554 (N_18554,N_18394,N_18345);
nor U18555 (N_18555,N_18325,N_18383);
xor U18556 (N_18556,N_18379,N_18269);
and U18557 (N_18557,N_18264,N_18291);
or U18558 (N_18558,N_18359,N_18381);
nor U18559 (N_18559,N_18277,N_18305);
xnor U18560 (N_18560,N_18443,N_18517);
xor U18561 (N_18561,N_18492,N_18467);
nand U18562 (N_18562,N_18462,N_18552);
nand U18563 (N_18563,N_18486,N_18428);
xnor U18564 (N_18564,N_18556,N_18466);
nor U18565 (N_18565,N_18518,N_18461);
nand U18566 (N_18566,N_18465,N_18439);
nor U18567 (N_18567,N_18407,N_18498);
nor U18568 (N_18568,N_18490,N_18472);
xor U18569 (N_18569,N_18422,N_18406);
xor U18570 (N_18570,N_18501,N_18513);
xor U18571 (N_18571,N_18503,N_18511);
nand U18572 (N_18572,N_18499,N_18433);
nand U18573 (N_18573,N_18489,N_18448);
and U18574 (N_18574,N_18452,N_18417);
nand U18575 (N_18575,N_18453,N_18480);
nand U18576 (N_18576,N_18478,N_18434);
nor U18577 (N_18577,N_18488,N_18557);
nor U18578 (N_18578,N_18539,N_18463);
nand U18579 (N_18579,N_18431,N_18401);
and U18580 (N_18580,N_18482,N_18532);
or U18581 (N_18581,N_18468,N_18505);
and U18582 (N_18582,N_18429,N_18496);
xor U18583 (N_18583,N_18476,N_18451);
xor U18584 (N_18584,N_18514,N_18544);
and U18585 (N_18585,N_18507,N_18542);
or U18586 (N_18586,N_18546,N_18446);
and U18587 (N_18587,N_18420,N_18533);
or U18588 (N_18588,N_18415,N_18403);
nor U18589 (N_18589,N_18430,N_18522);
nor U18590 (N_18590,N_18504,N_18421);
nand U18591 (N_18591,N_18512,N_18545);
nand U18592 (N_18592,N_18436,N_18456);
xnor U18593 (N_18593,N_18536,N_18502);
xor U18594 (N_18594,N_18409,N_18437);
or U18595 (N_18595,N_18454,N_18470);
xor U18596 (N_18596,N_18553,N_18543);
xor U18597 (N_18597,N_18487,N_18445);
xor U18598 (N_18598,N_18554,N_18460);
and U18599 (N_18599,N_18509,N_18419);
nand U18600 (N_18600,N_18550,N_18519);
nor U18601 (N_18601,N_18413,N_18508);
nand U18602 (N_18602,N_18551,N_18469);
nor U18603 (N_18603,N_18540,N_18515);
nand U18604 (N_18604,N_18495,N_18494);
nand U18605 (N_18605,N_18425,N_18491);
or U18606 (N_18606,N_18475,N_18405);
nand U18607 (N_18607,N_18441,N_18516);
nand U18608 (N_18608,N_18500,N_18555);
nor U18609 (N_18609,N_18541,N_18538);
nand U18610 (N_18610,N_18457,N_18458);
xnor U18611 (N_18611,N_18537,N_18427);
or U18612 (N_18612,N_18524,N_18464);
and U18613 (N_18613,N_18400,N_18444);
nand U18614 (N_18614,N_18423,N_18526);
nor U18615 (N_18615,N_18529,N_18479);
nor U18616 (N_18616,N_18474,N_18527);
nand U18617 (N_18617,N_18435,N_18424);
nor U18618 (N_18618,N_18497,N_18411);
xor U18619 (N_18619,N_18449,N_18459);
nand U18620 (N_18620,N_18530,N_18477);
or U18621 (N_18621,N_18520,N_18447);
and U18622 (N_18622,N_18481,N_18432);
and U18623 (N_18623,N_18455,N_18548);
and U18624 (N_18624,N_18408,N_18559);
or U18625 (N_18625,N_18410,N_18440);
or U18626 (N_18626,N_18506,N_18483);
nor U18627 (N_18627,N_18521,N_18484);
nor U18628 (N_18628,N_18402,N_18414);
xor U18629 (N_18629,N_18531,N_18528);
xnor U18630 (N_18630,N_18493,N_18485);
or U18631 (N_18631,N_18473,N_18471);
nor U18632 (N_18632,N_18549,N_18558);
nand U18633 (N_18633,N_18416,N_18450);
xnor U18634 (N_18634,N_18418,N_18404);
nor U18635 (N_18635,N_18442,N_18547);
and U18636 (N_18636,N_18525,N_18510);
and U18637 (N_18637,N_18535,N_18523);
and U18638 (N_18638,N_18438,N_18412);
nand U18639 (N_18639,N_18426,N_18534);
or U18640 (N_18640,N_18498,N_18422);
nor U18641 (N_18641,N_18559,N_18417);
xor U18642 (N_18642,N_18535,N_18553);
nand U18643 (N_18643,N_18465,N_18464);
xor U18644 (N_18644,N_18443,N_18543);
or U18645 (N_18645,N_18476,N_18481);
xnor U18646 (N_18646,N_18415,N_18478);
and U18647 (N_18647,N_18448,N_18431);
xnor U18648 (N_18648,N_18409,N_18517);
xor U18649 (N_18649,N_18400,N_18445);
nor U18650 (N_18650,N_18535,N_18456);
xnor U18651 (N_18651,N_18408,N_18475);
and U18652 (N_18652,N_18515,N_18472);
nand U18653 (N_18653,N_18419,N_18474);
nor U18654 (N_18654,N_18516,N_18412);
xnor U18655 (N_18655,N_18509,N_18492);
xor U18656 (N_18656,N_18557,N_18469);
or U18657 (N_18657,N_18431,N_18557);
and U18658 (N_18658,N_18425,N_18513);
and U18659 (N_18659,N_18533,N_18486);
nand U18660 (N_18660,N_18406,N_18508);
or U18661 (N_18661,N_18459,N_18413);
and U18662 (N_18662,N_18505,N_18425);
nor U18663 (N_18663,N_18431,N_18517);
and U18664 (N_18664,N_18450,N_18544);
or U18665 (N_18665,N_18404,N_18456);
xor U18666 (N_18666,N_18431,N_18450);
xor U18667 (N_18667,N_18416,N_18549);
xor U18668 (N_18668,N_18435,N_18404);
and U18669 (N_18669,N_18441,N_18415);
nand U18670 (N_18670,N_18492,N_18421);
nand U18671 (N_18671,N_18514,N_18482);
xor U18672 (N_18672,N_18527,N_18558);
nand U18673 (N_18673,N_18543,N_18514);
or U18674 (N_18674,N_18553,N_18465);
xnor U18675 (N_18675,N_18549,N_18556);
nand U18676 (N_18676,N_18492,N_18541);
xor U18677 (N_18677,N_18502,N_18493);
nor U18678 (N_18678,N_18438,N_18405);
nand U18679 (N_18679,N_18557,N_18429);
nor U18680 (N_18680,N_18437,N_18533);
xor U18681 (N_18681,N_18548,N_18421);
or U18682 (N_18682,N_18445,N_18523);
or U18683 (N_18683,N_18466,N_18486);
nand U18684 (N_18684,N_18499,N_18484);
nor U18685 (N_18685,N_18556,N_18435);
and U18686 (N_18686,N_18518,N_18524);
nor U18687 (N_18687,N_18501,N_18524);
nand U18688 (N_18688,N_18526,N_18457);
nand U18689 (N_18689,N_18483,N_18539);
xor U18690 (N_18690,N_18487,N_18524);
nand U18691 (N_18691,N_18427,N_18502);
nor U18692 (N_18692,N_18550,N_18410);
or U18693 (N_18693,N_18431,N_18501);
or U18694 (N_18694,N_18459,N_18539);
nand U18695 (N_18695,N_18507,N_18470);
and U18696 (N_18696,N_18457,N_18483);
xnor U18697 (N_18697,N_18427,N_18483);
or U18698 (N_18698,N_18500,N_18513);
nor U18699 (N_18699,N_18436,N_18476);
nand U18700 (N_18700,N_18424,N_18480);
nand U18701 (N_18701,N_18442,N_18519);
and U18702 (N_18702,N_18438,N_18511);
nor U18703 (N_18703,N_18508,N_18408);
or U18704 (N_18704,N_18518,N_18500);
nand U18705 (N_18705,N_18456,N_18472);
xor U18706 (N_18706,N_18439,N_18511);
xor U18707 (N_18707,N_18466,N_18498);
xnor U18708 (N_18708,N_18510,N_18437);
xor U18709 (N_18709,N_18524,N_18471);
nor U18710 (N_18710,N_18501,N_18454);
nor U18711 (N_18711,N_18525,N_18453);
or U18712 (N_18712,N_18531,N_18527);
or U18713 (N_18713,N_18463,N_18477);
nor U18714 (N_18714,N_18541,N_18544);
or U18715 (N_18715,N_18510,N_18419);
nor U18716 (N_18716,N_18515,N_18440);
nor U18717 (N_18717,N_18456,N_18444);
and U18718 (N_18718,N_18553,N_18459);
nor U18719 (N_18719,N_18445,N_18466);
nor U18720 (N_18720,N_18618,N_18583);
xor U18721 (N_18721,N_18581,N_18574);
and U18722 (N_18722,N_18703,N_18570);
nor U18723 (N_18723,N_18684,N_18693);
nor U18724 (N_18724,N_18612,N_18650);
nand U18725 (N_18725,N_18580,N_18655);
nand U18726 (N_18726,N_18672,N_18635);
nor U18727 (N_18727,N_18665,N_18718);
nand U18728 (N_18728,N_18615,N_18603);
or U18729 (N_18729,N_18670,N_18631);
and U18730 (N_18730,N_18594,N_18659);
and U18731 (N_18731,N_18634,N_18698);
and U18732 (N_18732,N_18563,N_18586);
and U18733 (N_18733,N_18644,N_18576);
xnor U18734 (N_18734,N_18628,N_18687);
nor U18735 (N_18735,N_18652,N_18696);
nor U18736 (N_18736,N_18619,N_18675);
xor U18737 (N_18737,N_18588,N_18716);
or U18738 (N_18738,N_18613,N_18700);
nor U18739 (N_18739,N_18719,N_18704);
nand U18740 (N_18740,N_18707,N_18682);
and U18741 (N_18741,N_18651,N_18609);
and U18742 (N_18742,N_18564,N_18676);
xor U18743 (N_18743,N_18691,N_18569);
or U18744 (N_18744,N_18604,N_18711);
and U18745 (N_18745,N_18712,N_18661);
nor U18746 (N_18746,N_18579,N_18677);
nand U18747 (N_18747,N_18606,N_18705);
xnor U18748 (N_18748,N_18647,N_18646);
nor U18749 (N_18749,N_18686,N_18610);
xnor U18750 (N_18750,N_18657,N_18597);
nand U18751 (N_18751,N_18598,N_18714);
nand U18752 (N_18752,N_18595,N_18648);
or U18753 (N_18753,N_18688,N_18640);
nand U18754 (N_18754,N_18664,N_18654);
or U18755 (N_18755,N_18689,N_18614);
nor U18756 (N_18756,N_18625,N_18577);
nand U18757 (N_18757,N_18596,N_18633);
xor U18758 (N_18758,N_18717,N_18575);
and U18759 (N_18759,N_18666,N_18573);
or U18760 (N_18760,N_18590,N_18641);
or U18761 (N_18761,N_18566,N_18599);
and U18762 (N_18762,N_18680,N_18568);
nand U18763 (N_18763,N_18674,N_18611);
xor U18764 (N_18764,N_18600,N_18645);
nor U18765 (N_18765,N_18715,N_18593);
or U18766 (N_18766,N_18649,N_18710);
nand U18767 (N_18767,N_18624,N_18582);
and U18768 (N_18768,N_18673,N_18626);
nand U18769 (N_18769,N_18621,N_18620);
or U18770 (N_18770,N_18629,N_18591);
and U18771 (N_18771,N_18605,N_18608);
nand U18772 (N_18772,N_18678,N_18685);
and U18773 (N_18773,N_18607,N_18571);
or U18774 (N_18774,N_18669,N_18632);
and U18775 (N_18775,N_18709,N_18587);
or U18776 (N_18776,N_18706,N_18630);
xnor U18777 (N_18777,N_18638,N_18660);
xnor U18778 (N_18778,N_18565,N_18681);
xnor U18779 (N_18779,N_18699,N_18589);
or U18780 (N_18780,N_18572,N_18601);
nand U18781 (N_18781,N_18617,N_18637);
and U18782 (N_18782,N_18622,N_18642);
xnor U18783 (N_18783,N_18697,N_18690);
and U18784 (N_18784,N_18695,N_18623);
xor U18785 (N_18785,N_18592,N_18643);
and U18786 (N_18786,N_18562,N_18692);
and U18787 (N_18787,N_18656,N_18663);
or U18788 (N_18788,N_18567,N_18683);
or U18789 (N_18789,N_18679,N_18639);
nor U18790 (N_18790,N_18668,N_18585);
nor U18791 (N_18791,N_18671,N_18662);
xor U18792 (N_18792,N_18708,N_18702);
nor U18793 (N_18793,N_18584,N_18701);
nor U18794 (N_18794,N_18667,N_18578);
nand U18795 (N_18795,N_18694,N_18627);
or U18796 (N_18796,N_18560,N_18713);
xnor U18797 (N_18797,N_18616,N_18602);
xor U18798 (N_18798,N_18636,N_18561);
xor U18799 (N_18799,N_18658,N_18653);
xnor U18800 (N_18800,N_18714,N_18676);
xnor U18801 (N_18801,N_18593,N_18698);
nand U18802 (N_18802,N_18699,N_18626);
or U18803 (N_18803,N_18625,N_18696);
and U18804 (N_18804,N_18560,N_18669);
nand U18805 (N_18805,N_18676,N_18634);
xor U18806 (N_18806,N_18598,N_18590);
nor U18807 (N_18807,N_18594,N_18614);
nor U18808 (N_18808,N_18707,N_18573);
or U18809 (N_18809,N_18652,N_18609);
nand U18810 (N_18810,N_18642,N_18581);
and U18811 (N_18811,N_18590,N_18575);
and U18812 (N_18812,N_18659,N_18670);
nand U18813 (N_18813,N_18613,N_18708);
and U18814 (N_18814,N_18712,N_18705);
nand U18815 (N_18815,N_18685,N_18701);
xor U18816 (N_18816,N_18605,N_18700);
or U18817 (N_18817,N_18618,N_18567);
nand U18818 (N_18818,N_18567,N_18561);
or U18819 (N_18819,N_18670,N_18624);
nor U18820 (N_18820,N_18681,N_18714);
nand U18821 (N_18821,N_18612,N_18639);
or U18822 (N_18822,N_18701,N_18686);
nor U18823 (N_18823,N_18655,N_18649);
and U18824 (N_18824,N_18591,N_18701);
nand U18825 (N_18825,N_18649,N_18719);
nor U18826 (N_18826,N_18620,N_18719);
nor U18827 (N_18827,N_18598,N_18668);
nor U18828 (N_18828,N_18593,N_18563);
and U18829 (N_18829,N_18608,N_18655);
xor U18830 (N_18830,N_18591,N_18562);
nand U18831 (N_18831,N_18702,N_18592);
or U18832 (N_18832,N_18610,N_18662);
nor U18833 (N_18833,N_18696,N_18690);
nand U18834 (N_18834,N_18606,N_18592);
nand U18835 (N_18835,N_18682,N_18706);
nor U18836 (N_18836,N_18650,N_18692);
nor U18837 (N_18837,N_18628,N_18636);
xor U18838 (N_18838,N_18693,N_18701);
nor U18839 (N_18839,N_18673,N_18566);
xor U18840 (N_18840,N_18692,N_18581);
and U18841 (N_18841,N_18572,N_18704);
nand U18842 (N_18842,N_18645,N_18607);
xor U18843 (N_18843,N_18617,N_18694);
or U18844 (N_18844,N_18641,N_18596);
or U18845 (N_18845,N_18702,N_18602);
nand U18846 (N_18846,N_18682,N_18636);
nor U18847 (N_18847,N_18606,N_18605);
nor U18848 (N_18848,N_18646,N_18717);
or U18849 (N_18849,N_18693,N_18709);
and U18850 (N_18850,N_18653,N_18563);
and U18851 (N_18851,N_18686,N_18605);
xnor U18852 (N_18852,N_18683,N_18628);
xnor U18853 (N_18853,N_18625,N_18633);
nor U18854 (N_18854,N_18595,N_18611);
and U18855 (N_18855,N_18657,N_18562);
or U18856 (N_18856,N_18702,N_18630);
nor U18857 (N_18857,N_18578,N_18708);
xnor U18858 (N_18858,N_18589,N_18579);
or U18859 (N_18859,N_18714,N_18596);
xor U18860 (N_18860,N_18608,N_18649);
nor U18861 (N_18861,N_18679,N_18690);
nand U18862 (N_18862,N_18696,N_18589);
nor U18863 (N_18863,N_18567,N_18674);
and U18864 (N_18864,N_18623,N_18588);
xnor U18865 (N_18865,N_18592,N_18607);
nor U18866 (N_18866,N_18666,N_18719);
nand U18867 (N_18867,N_18588,N_18698);
xor U18868 (N_18868,N_18629,N_18704);
xnor U18869 (N_18869,N_18664,N_18629);
nor U18870 (N_18870,N_18675,N_18560);
nor U18871 (N_18871,N_18658,N_18668);
or U18872 (N_18872,N_18632,N_18663);
nand U18873 (N_18873,N_18602,N_18701);
xnor U18874 (N_18874,N_18657,N_18645);
nand U18875 (N_18875,N_18593,N_18706);
nor U18876 (N_18876,N_18563,N_18651);
nand U18877 (N_18877,N_18641,N_18709);
nand U18878 (N_18878,N_18572,N_18599);
or U18879 (N_18879,N_18665,N_18636);
nor U18880 (N_18880,N_18857,N_18871);
or U18881 (N_18881,N_18746,N_18776);
nand U18882 (N_18882,N_18837,N_18773);
nand U18883 (N_18883,N_18793,N_18797);
xnor U18884 (N_18884,N_18838,N_18750);
xnor U18885 (N_18885,N_18825,N_18847);
nor U18886 (N_18886,N_18754,N_18788);
nand U18887 (N_18887,N_18804,N_18873);
xor U18888 (N_18888,N_18751,N_18849);
nand U18889 (N_18889,N_18785,N_18761);
and U18890 (N_18890,N_18824,N_18815);
or U18891 (N_18891,N_18778,N_18813);
or U18892 (N_18892,N_18802,N_18855);
xnor U18893 (N_18893,N_18859,N_18774);
nand U18894 (N_18894,N_18811,N_18744);
and U18895 (N_18895,N_18737,N_18800);
and U18896 (N_18896,N_18872,N_18787);
nor U18897 (N_18897,N_18875,N_18820);
nor U18898 (N_18898,N_18741,N_18752);
nand U18899 (N_18899,N_18852,N_18867);
and U18900 (N_18900,N_18817,N_18870);
nand U18901 (N_18901,N_18742,N_18836);
nand U18902 (N_18902,N_18879,N_18844);
and U18903 (N_18903,N_18869,N_18759);
or U18904 (N_18904,N_18828,N_18853);
xnor U18905 (N_18905,N_18768,N_18868);
xnor U18906 (N_18906,N_18856,N_18822);
nor U18907 (N_18907,N_18808,N_18803);
nand U18908 (N_18908,N_18767,N_18736);
or U18909 (N_18909,N_18770,N_18833);
nor U18910 (N_18910,N_18726,N_18848);
and U18911 (N_18911,N_18721,N_18720);
xor U18912 (N_18912,N_18860,N_18722);
or U18913 (N_18913,N_18733,N_18777);
or U18914 (N_18914,N_18863,N_18794);
nor U18915 (N_18915,N_18772,N_18858);
nor U18916 (N_18916,N_18753,N_18831);
and U18917 (N_18917,N_18723,N_18783);
nand U18918 (N_18918,N_18795,N_18729);
xnor U18919 (N_18919,N_18786,N_18732);
nor U18920 (N_18920,N_18758,N_18814);
nand U18921 (N_18921,N_18835,N_18841);
xor U18922 (N_18922,N_18830,N_18818);
xnor U18923 (N_18923,N_18784,N_18730);
or U18924 (N_18924,N_18791,N_18827);
xor U18925 (N_18925,N_18842,N_18780);
and U18926 (N_18926,N_18799,N_18725);
xnor U18927 (N_18927,N_18756,N_18747);
and U18928 (N_18928,N_18861,N_18739);
nor U18929 (N_18929,N_18864,N_18823);
xnor U18930 (N_18930,N_18738,N_18766);
nand U18931 (N_18931,N_18829,N_18832);
nor U18932 (N_18932,N_18789,N_18878);
xnor U18933 (N_18933,N_18865,N_18792);
nand U18934 (N_18934,N_18782,N_18735);
nor U18935 (N_18935,N_18796,N_18812);
nand U18936 (N_18936,N_18805,N_18816);
and U18937 (N_18937,N_18755,N_18771);
xor U18938 (N_18938,N_18760,N_18740);
or U18939 (N_18939,N_18840,N_18809);
or U18940 (N_18940,N_18762,N_18763);
or U18941 (N_18941,N_18810,N_18854);
xor U18942 (N_18942,N_18839,N_18775);
xor U18943 (N_18943,N_18845,N_18728);
nand U18944 (N_18944,N_18819,N_18731);
xor U18945 (N_18945,N_18790,N_18850);
nor U18946 (N_18946,N_18798,N_18748);
nand U18947 (N_18947,N_18821,N_18745);
nand U18948 (N_18948,N_18769,N_18806);
and U18949 (N_18949,N_18826,N_18764);
or U18950 (N_18950,N_18749,N_18866);
or U18951 (N_18951,N_18876,N_18779);
nand U18952 (N_18952,N_18724,N_18834);
nand U18953 (N_18953,N_18843,N_18846);
and U18954 (N_18954,N_18765,N_18727);
nor U18955 (N_18955,N_18734,N_18781);
nand U18956 (N_18956,N_18877,N_18851);
xor U18957 (N_18957,N_18801,N_18862);
nor U18958 (N_18958,N_18743,N_18757);
and U18959 (N_18959,N_18874,N_18807);
or U18960 (N_18960,N_18733,N_18871);
nor U18961 (N_18961,N_18762,N_18792);
nor U18962 (N_18962,N_18795,N_18827);
nand U18963 (N_18963,N_18732,N_18756);
nand U18964 (N_18964,N_18872,N_18747);
xnor U18965 (N_18965,N_18855,N_18869);
or U18966 (N_18966,N_18760,N_18872);
xor U18967 (N_18967,N_18740,N_18785);
nand U18968 (N_18968,N_18848,N_18813);
nand U18969 (N_18969,N_18858,N_18829);
nor U18970 (N_18970,N_18843,N_18852);
or U18971 (N_18971,N_18821,N_18781);
nor U18972 (N_18972,N_18779,N_18774);
or U18973 (N_18973,N_18723,N_18745);
nand U18974 (N_18974,N_18769,N_18851);
and U18975 (N_18975,N_18735,N_18758);
xor U18976 (N_18976,N_18737,N_18780);
nor U18977 (N_18977,N_18806,N_18741);
xor U18978 (N_18978,N_18786,N_18871);
nand U18979 (N_18979,N_18841,N_18758);
xor U18980 (N_18980,N_18868,N_18723);
and U18981 (N_18981,N_18854,N_18808);
nand U18982 (N_18982,N_18827,N_18757);
and U18983 (N_18983,N_18751,N_18761);
nor U18984 (N_18984,N_18771,N_18856);
nor U18985 (N_18985,N_18798,N_18803);
and U18986 (N_18986,N_18731,N_18736);
xor U18987 (N_18987,N_18724,N_18799);
or U18988 (N_18988,N_18804,N_18844);
nor U18989 (N_18989,N_18740,N_18808);
nand U18990 (N_18990,N_18744,N_18791);
nor U18991 (N_18991,N_18734,N_18793);
xor U18992 (N_18992,N_18816,N_18747);
xor U18993 (N_18993,N_18829,N_18799);
and U18994 (N_18994,N_18734,N_18817);
nand U18995 (N_18995,N_18730,N_18865);
nor U18996 (N_18996,N_18737,N_18746);
xnor U18997 (N_18997,N_18727,N_18733);
and U18998 (N_18998,N_18851,N_18760);
nor U18999 (N_18999,N_18851,N_18853);
nand U19000 (N_19000,N_18721,N_18754);
or U19001 (N_19001,N_18729,N_18852);
or U19002 (N_19002,N_18775,N_18749);
and U19003 (N_19003,N_18861,N_18850);
nand U19004 (N_19004,N_18823,N_18738);
or U19005 (N_19005,N_18819,N_18801);
nor U19006 (N_19006,N_18876,N_18767);
nand U19007 (N_19007,N_18758,N_18868);
nor U19008 (N_19008,N_18740,N_18758);
nor U19009 (N_19009,N_18827,N_18744);
xor U19010 (N_19010,N_18750,N_18738);
nor U19011 (N_19011,N_18809,N_18816);
xnor U19012 (N_19012,N_18801,N_18762);
nor U19013 (N_19013,N_18763,N_18743);
nor U19014 (N_19014,N_18843,N_18809);
or U19015 (N_19015,N_18875,N_18851);
or U19016 (N_19016,N_18787,N_18749);
nor U19017 (N_19017,N_18746,N_18828);
nor U19018 (N_19018,N_18794,N_18723);
and U19019 (N_19019,N_18805,N_18839);
nor U19020 (N_19020,N_18839,N_18798);
or U19021 (N_19021,N_18869,N_18852);
nand U19022 (N_19022,N_18833,N_18756);
and U19023 (N_19023,N_18837,N_18747);
nor U19024 (N_19024,N_18728,N_18808);
xnor U19025 (N_19025,N_18824,N_18830);
and U19026 (N_19026,N_18785,N_18860);
and U19027 (N_19027,N_18873,N_18740);
nand U19028 (N_19028,N_18731,N_18850);
nand U19029 (N_19029,N_18824,N_18776);
xor U19030 (N_19030,N_18806,N_18796);
nand U19031 (N_19031,N_18756,N_18837);
nand U19032 (N_19032,N_18876,N_18800);
nor U19033 (N_19033,N_18812,N_18737);
nor U19034 (N_19034,N_18772,N_18784);
and U19035 (N_19035,N_18814,N_18757);
nand U19036 (N_19036,N_18874,N_18823);
nor U19037 (N_19037,N_18864,N_18789);
and U19038 (N_19038,N_18796,N_18817);
and U19039 (N_19039,N_18828,N_18783);
xor U19040 (N_19040,N_18881,N_18930);
nor U19041 (N_19041,N_18988,N_19013);
nor U19042 (N_19042,N_18996,N_18925);
nand U19043 (N_19043,N_19000,N_18961);
or U19044 (N_19044,N_18926,N_18940);
nor U19045 (N_19045,N_19002,N_19006);
xnor U19046 (N_19046,N_18934,N_18973);
xnor U19047 (N_19047,N_18891,N_18979);
nor U19048 (N_19048,N_18883,N_18982);
nor U19049 (N_19049,N_18950,N_19014);
nor U19050 (N_19050,N_18956,N_18880);
xnor U19051 (N_19051,N_18966,N_18970);
xor U19052 (N_19052,N_18999,N_19027);
nor U19053 (N_19053,N_19015,N_18944);
xnor U19054 (N_19054,N_18887,N_18928);
nand U19055 (N_19055,N_18886,N_19026);
or U19056 (N_19056,N_18986,N_18943);
and U19057 (N_19057,N_18935,N_18993);
or U19058 (N_19058,N_18914,N_19005);
and U19059 (N_19059,N_18987,N_18909);
or U19060 (N_19060,N_18965,N_18985);
and U19061 (N_19061,N_18898,N_19028);
nor U19062 (N_19062,N_18964,N_18937);
nand U19063 (N_19063,N_18907,N_18908);
or U19064 (N_19064,N_18974,N_19020);
or U19065 (N_19065,N_18902,N_18906);
nor U19066 (N_19066,N_18962,N_18959);
or U19067 (N_19067,N_18945,N_18913);
nand U19068 (N_19068,N_18995,N_18983);
and U19069 (N_19069,N_19021,N_18894);
nand U19070 (N_19070,N_18960,N_18948);
nor U19071 (N_19071,N_18918,N_18884);
or U19072 (N_19072,N_18968,N_19019);
and U19073 (N_19073,N_18949,N_18941);
and U19074 (N_19074,N_19033,N_18912);
xnor U19075 (N_19075,N_18903,N_18922);
nor U19076 (N_19076,N_19038,N_18992);
nand U19077 (N_19077,N_18927,N_18981);
xnor U19078 (N_19078,N_18929,N_18910);
nor U19079 (N_19079,N_19004,N_18997);
nand U19080 (N_19080,N_19031,N_19009);
nand U19081 (N_19081,N_19017,N_18984);
xor U19082 (N_19082,N_18947,N_18897);
and U19083 (N_19083,N_18932,N_19035);
and U19084 (N_19084,N_18977,N_18899);
and U19085 (N_19085,N_18952,N_18980);
or U19086 (N_19086,N_18975,N_18917);
or U19087 (N_19087,N_18900,N_19032);
nor U19088 (N_19088,N_18969,N_18957);
xnor U19089 (N_19089,N_19001,N_19011);
and U19090 (N_19090,N_18905,N_18936);
nor U19091 (N_19091,N_18921,N_19024);
xnor U19092 (N_19092,N_18951,N_19039);
nand U19093 (N_19093,N_19029,N_19022);
nor U19094 (N_19094,N_19012,N_19003);
nor U19095 (N_19095,N_18978,N_18904);
nor U19096 (N_19096,N_18923,N_18890);
nand U19097 (N_19097,N_18990,N_18946);
xor U19098 (N_19098,N_18971,N_19036);
or U19099 (N_19099,N_18958,N_18933);
nor U19100 (N_19100,N_18991,N_18955);
nand U19101 (N_19101,N_18916,N_18931);
nand U19102 (N_19102,N_18888,N_19008);
and U19103 (N_19103,N_19037,N_18901);
or U19104 (N_19104,N_18989,N_18924);
nor U19105 (N_19105,N_19007,N_19018);
nand U19106 (N_19106,N_18882,N_18942);
nor U19107 (N_19107,N_18939,N_18976);
and U19108 (N_19108,N_19030,N_18919);
xor U19109 (N_19109,N_18963,N_18892);
or U19110 (N_19110,N_18885,N_19034);
nor U19111 (N_19111,N_18896,N_18967);
xor U19112 (N_19112,N_18953,N_18938);
and U19113 (N_19113,N_18972,N_18954);
and U19114 (N_19114,N_19023,N_18893);
and U19115 (N_19115,N_18911,N_19016);
xnor U19116 (N_19116,N_19010,N_19025);
or U19117 (N_19117,N_18915,N_18994);
nand U19118 (N_19118,N_18920,N_18895);
xor U19119 (N_19119,N_18998,N_18889);
nor U19120 (N_19120,N_18989,N_18887);
nor U19121 (N_19121,N_19008,N_18993);
xor U19122 (N_19122,N_19003,N_18935);
nor U19123 (N_19123,N_19000,N_19025);
nor U19124 (N_19124,N_18929,N_19029);
xnor U19125 (N_19125,N_18952,N_18999);
nand U19126 (N_19126,N_18993,N_18887);
xnor U19127 (N_19127,N_18972,N_18882);
xnor U19128 (N_19128,N_18907,N_18939);
nor U19129 (N_19129,N_18899,N_18987);
xnor U19130 (N_19130,N_18973,N_18919);
or U19131 (N_19131,N_18963,N_19006);
or U19132 (N_19132,N_19023,N_18987);
nor U19133 (N_19133,N_18929,N_18960);
or U19134 (N_19134,N_18933,N_19019);
xnor U19135 (N_19135,N_18881,N_18992);
nand U19136 (N_19136,N_18889,N_19028);
nor U19137 (N_19137,N_18984,N_19005);
nand U19138 (N_19138,N_18986,N_18951);
or U19139 (N_19139,N_18943,N_18922);
or U19140 (N_19140,N_19013,N_18979);
xnor U19141 (N_19141,N_18973,N_18930);
and U19142 (N_19142,N_18923,N_19013);
xor U19143 (N_19143,N_18880,N_19003);
and U19144 (N_19144,N_19005,N_19034);
nand U19145 (N_19145,N_19010,N_18993);
and U19146 (N_19146,N_18950,N_19018);
xor U19147 (N_19147,N_18977,N_18959);
and U19148 (N_19148,N_18909,N_18981);
nor U19149 (N_19149,N_18981,N_18941);
or U19150 (N_19150,N_18955,N_18917);
and U19151 (N_19151,N_18934,N_18974);
nor U19152 (N_19152,N_18903,N_18941);
nand U19153 (N_19153,N_19036,N_18958);
nor U19154 (N_19154,N_18933,N_18902);
and U19155 (N_19155,N_19024,N_18904);
and U19156 (N_19156,N_19011,N_18907);
and U19157 (N_19157,N_18982,N_18949);
nand U19158 (N_19158,N_18945,N_18927);
or U19159 (N_19159,N_18969,N_18882);
nor U19160 (N_19160,N_19016,N_18930);
xor U19161 (N_19161,N_18965,N_18952);
and U19162 (N_19162,N_18922,N_18949);
nand U19163 (N_19163,N_19004,N_18970);
or U19164 (N_19164,N_18935,N_19039);
nor U19165 (N_19165,N_18924,N_18910);
xor U19166 (N_19166,N_18935,N_19012);
nor U19167 (N_19167,N_18992,N_19001);
xnor U19168 (N_19168,N_18963,N_18943);
xor U19169 (N_19169,N_18948,N_19027);
xor U19170 (N_19170,N_18940,N_18966);
or U19171 (N_19171,N_18948,N_18925);
or U19172 (N_19172,N_19015,N_18945);
nor U19173 (N_19173,N_18921,N_18885);
xor U19174 (N_19174,N_18894,N_19028);
xor U19175 (N_19175,N_18958,N_19035);
or U19176 (N_19176,N_18994,N_18941);
or U19177 (N_19177,N_18969,N_19037);
or U19178 (N_19178,N_19028,N_18925);
nand U19179 (N_19179,N_18935,N_18917);
or U19180 (N_19180,N_18994,N_18887);
xor U19181 (N_19181,N_18906,N_19008);
and U19182 (N_19182,N_18922,N_19034);
or U19183 (N_19183,N_19013,N_18925);
xor U19184 (N_19184,N_18927,N_18982);
xnor U19185 (N_19185,N_18992,N_18985);
xor U19186 (N_19186,N_18896,N_18981);
nand U19187 (N_19187,N_19026,N_18992);
nand U19188 (N_19188,N_18939,N_18889);
xor U19189 (N_19189,N_18993,N_18968);
or U19190 (N_19190,N_18914,N_19009);
nand U19191 (N_19191,N_18936,N_18987);
xor U19192 (N_19192,N_19013,N_18958);
or U19193 (N_19193,N_18884,N_18982);
nor U19194 (N_19194,N_18959,N_18956);
nand U19195 (N_19195,N_19039,N_18944);
nand U19196 (N_19196,N_18943,N_18989);
nor U19197 (N_19197,N_18977,N_19037);
nor U19198 (N_19198,N_18923,N_18918);
nand U19199 (N_19199,N_18983,N_19027);
xnor U19200 (N_19200,N_19096,N_19045);
and U19201 (N_19201,N_19143,N_19119);
xor U19202 (N_19202,N_19122,N_19161);
nand U19203 (N_19203,N_19063,N_19171);
nor U19204 (N_19204,N_19107,N_19129);
nor U19205 (N_19205,N_19139,N_19044);
xnor U19206 (N_19206,N_19042,N_19155);
or U19207 (N_19207,N_19162,N_19173);
xor U19208 (N_19208,N_19126,N_19098);
nor U19209 (N_19209,N_19131,N_19087);
nand U19210 (N_19210,N_19144,N_19078);
and U19211 (N_19211,N_19170,N_19184);
and U19212 (N_19212,N_19051,N_19121);
and U19213 (N_19213,N_19114,N_19159);
xnor U19214 (N_19214,N_19056,N_19123);
and U19215 (N_19215,N_19169,N_19187);
or U19216 (N_19216,N_19108,N_19125);
nor U19217 (N_19217,N_19136,N_19174);
nand U19218 (N_19218,N_19116,N_19040);
nor U19219 (N_19219,N_19175,N_19158);
or U19220 (N_19220,N_19167,N_19093);
or U19221 (N_19221,N_19057,N_19165);
nand U19222 (N_19222,N_19166,N_19142);
or U19223 (N_19223,N_19196,N_19141);
nor U19224 (N_19224,N_19061,N_19132);
nor U19225 (N_19225,N_19047,N_19157);
xor U19226 (N_19226,N_19113,N_19095);
nand U19227 (N_19227,N_19140,N_19194);
xor U19228 (N_19228,N_19100,N_19146);
and U19229 (N_19229,N_19163,N_19052);
or U19230 (N_19230,N_19058,N_19124);
nand U19231 (N_19231,N_19150,N_19178);
xor U19232 (N_19232,N_19179,N_19074);
and U19233 (N_19233,N_19172,N_19177);
xnor U19234 (N_19234,N_19067,N_19079);
and U19235 (N_19235,N_19076,N_19064);
nor U19236 (N_19236,N_19153,N_19069);
xor U19237 (N_19237,N_19128,N_19183);
or U19238 (N_19238,N_19043,N_19197);
xor U19239 (N_19239,N_19070,N_19086);
nand U19240 (N_19240,N_19109,N_19138);
xnor U19241 (N_19241,N_19115,N_19059);
or U19242 (N_19242,N_19110,N_19101);
or U19243 (N_19243,N_19071,N_19112);
nand U19244 (N_19244,N_19160,N_19182);
nand U19245 (N_19245,N_19198,N_19077);
nor U19246 (N_19246,N_19083,N_19065);
nor U19247 (N_19247,N_19117,N_19148);
nor U19248 (N_19248,N_19081,N_19068);
nor U19249 (N_19249,N_19062,N_19049);
nand U19250 (N_19250,N_19080,N_19066);
nor U19251 (N_19251,N_19130,N_19099);
nand U19252 (N_19252,N_19156,N_19041);
nor U19253 (N_19253,N_19105,N_19106);
nand U19254 (N_19254,N_19164,N_19192);
or U19255 (N_19255,N_19089,N_19154);
xnor U19256 (N_19256,N_19090,N_19050);
nand U19257 (N_19257,N_19127,N_19046);
and U19258 (N_19258,N_19082,N_19091);
nand U19259 (N_19259,N_19060,N_19188);
nor U19260 (N_19260,N_19191,N_19135);
or U19261 (N_19261,N_19133,N_19152);
nand U19262 (N_19262,N_19085,N_19055);
xnor U19263 (N_19263,N_19084,N_19137);
and U19264 (N_19264,N_19088,N_19193);
and U19265 (N_19265,N_19151,N_19075);
nand U19266 (N_19266,N_19053,N_19168);
xnor U19267 (N_19267,N_19120,N_19054);
nand U19268 (N_19268,N_19048,N_19102);
nand U19269 (N_19269,N_19195,N_19199);
or U19270 (N_19270,N_19190,N_19104);
nand U19271 (N_19271,N_19103,N_19073);
and U19272 (N_19272,N_19072,N_19097);
nor U19273 (N_19273,N_19111,N_19118);
nor U19274 (N_19274,N_19186,N_19092);
xnor U19275 (N_19275,N_19181,N_19185);
nor U19276 (N_19276,N_19149,N_19147);
nand U19277 (N_19277,N_19176,N_19189);
nand U19278 (N_19278,N_19134,N_19145);
xnor U19279 (N_19279,N_19094,N_19180);
nand U19280 (N_19280,N_19182,N_19167);
nor U19281 (N_19281,N_19180,N_19118);
or U19282 (N_19282,N_19101,N_19129);
xor U19283 (N_19283,N_19193,N_19192);
or U19284 (N_19284,N_19051,N_19044);
and U19285 (N_19285,N_19139,N_19136);
xnor U19286 (N_19286,N_19060,N_19086);
and U19287 (N_19287,N_19170,N_19194);
nor U19288 (N_19288,N_19141,N_19162);
nand U19289 (N_19289,N_19187,N_19153);
xnor U19290 (N_19290,N_19057,N_19152);
nor U19291 (N_19291,N_19098,N_19151);
nor U19292 (N_19292,N_19123,N_19181);
nor U19293 (N_19293,N_19052,N_19197);
xnor U19294 (N_19294,N_19056,N_19114);
nor U19295 (N_19295,N_19146,N_19067);
nand U19296 (N_19296,N_19137,N_19162);
nand U19297 (N_19297,N_19142,N_19169);
and U19298 (N_19298,N_19160,N_19096);
or U19299 (N_19299,N_19132,N_19123);
or U19300 (N_19300,N_19068,N_19054);
nand U19301 (N_19301,N_19192,N_19169);
or U19302 (N_19302,N_19116,N_19104);
and U19303 (N_19303,N_19155,N_19182);
nand U19304 (N_19304,N_19085,N_19135);
xor U19305 (N_19305,N_19154,N_19193);
or U19306 (N_19306,N_19139,N_19182);
nand U19307 (N_19307,N_19150,N_19054);
xor U19308 (N_19308,N_19088,N_19174);
or U19309 (N_19309,N_19093,N_19182);
nor U19310 (N_19310,N_19196,N_19083);
and U19311 (N_19311,N_19172,N_19085);
or U19312 (N_19312,N_19095,N_19076);
or U19313 (N_19313,N_19146,N_19191);
or U19314 (N_19314,N_19178,N_19113);
and U19315 (N_19315,N_19163,N_19089);
and U19316 (N_19316,N_19179,N_19121);
and U19317 (N_19317,N_19162,N_19189);
and U19318 (N_19318,N_19099,N_19073);
nor U19319 (N_19319,N_19044,N_19105);
or U19320 (N_19320,N_19187,N_19102);
and U19321 (N_19321,N_19183,N_19050);
and U19322 (N_19322,N_19143,N_19152);
or U19323 (N_19323,N_19181,N_19061);
and U19324 (N_19324,N_19185,N_19093);
and U19325 (N_19325,N_19175,N_19079);
and U19326 (N_19326,N_19127,N_19097);
or U19327 (N_19327,N_19081,N_19098);
and U19328 (N_19328,N_19122,N_19172);
and U19329 (N_19329,N_19166,N_19065);
or U19330 (N_19330,N_19130,N_19171);
or U19331 (N_19331,N_19083,N_19047);
nor U19332 (N_19332,N_19157,N_19191);
xnor U19333 (N_19333,N_19170,N_19104);
xnor U19334 (N_19334,N_19150,N_19155);
nand U19335 (N_19335,N_19052,N_19111);
nor U19336 (N_19336,N_19106,N_19144);
nor U19337 (N_19337,N_19074,N_19085);
nand U19338 (N_19338,N_19163,N_19107);
and U19339 (N_19339,N_19044,N_19195);
or U19340 (N_19340,N_19154,N_19060);
nand U19341 (N_19341,N_19079,N_19153);
nand U19342 (N_19342,N_19111,N_19065);
or U19343 (N_19343,N_19145,N_19118);
and U19344 (N_19344,N_19136,N_19170);
or U19345 (N_19345,N_19158,N_19146);
nand U19346 (N_19346,N_19092,N_19101);
or U19347 (N_19347,N_19084,N_19054);
or U19348 (N_19348,N_19150,N_19176);
and U19349 (N_19349,N_19048,N_19145);
nor U19350 (N_19350,N_19174,N_19051);
or U19351 (N_19351,N_19117,N_19073);
and U19352 (N_19352,N_19094,N_19165);
xor U19353 (N_19353,N_19091,N_19095);
and U19354 (N_19354,N_19157,N_19081);
nand U19355 (N_19355,N_19105,N_19066);
nor U19356 (N_19356,N_19151,N_19163);
and U19357 (N_19357,N_19060,N_19082);
and U19358 (N_19358,N_19103,N_19134);
nor U19359 (N_19359,N_19119,N_19150);
or U19360 (N_19360,N_19247,N_19307);
nor U19361 (N_19361,N_19358,N_19254);
xor U19362 (N_19362,N_19280,N_19272);
and U19363 (N_19363,N_19268,N_19230);
or U19364 (N_19364,N_19265,N_19210);
xor U19365 (N_19365,N_19236,N_19337);
nand U19366 (N_19366,N_19352,N_19346);
nor U19367 (N_19367,N_19240,N_19305);
nor U19368 (N_19368,N_19279,N_19330);
xnor U19369 (N_19369,N_19244,N_19239);
or U19370 (N_19370,N_19238,N_19260);
xnor U19371 (N_19371,N_19294,N_19271);
and U19372 (N_19372,N_19324,N_19219);
nand U19373 (N_19373,N_19215,N_19251);
nor U19374 (N_19374,N_19201,N_19243);
or U19375 (N_19375,N_19204,N_19354);
and U19376 (N_19376,N_19297,N_19349);
nand U19377 (N_19377,N_19235,N_19220);
xor U19378 (N_19378,N_19314,N_19225);
xor U19379 (N_19379,N_19345,N_19291);
and U19380 (N_19380,N_19350,N_19233);
and U19381 (N_19381,N_19348,N_19332);
nand U19382 (N_19382,N_19224,N_19317);
nand U19383 (N_19383,N_19299,N_19290);
xnor U19384 (N_19384,N_19275,N_19285);
and U19385 (N_19385,N_19329,N_19355);
nor U19386 (N_19386,N_19340,N_19287);
or U19387 (N_19387,N_19266,N_19298);
nand U19388 (N_19388,N_19232,N_19216);
or U19389 (N_19389,N_19259,N_19269);
xor U19390 (N_19390,N_19208,N_19320);
nor U19391 (N_19391,N_19263,N_19283);
or U19392 (N_19392,N_19356,N_19327);
and U19393 (N_19393,N_19231,N_19200);
xnor U19394 (N_19394,N_19336,N_19343);
nor U19395 (N_19395,N_19300,N_19262);
or U19396 (N_19396,N_19341,N_19325);
nor U19397 (N_19397,N_19318,N_19289);
nand U19398 (N_19398,N_19255,N_19292);
nor U19399 (N_19399,N_19237,N_19357);
or U19400 (N_19400,N_19311,N_19347);
xor U19401 (N_19401,N_19214,N_19264);
nand U19402 (N_19402,N_19202,N_19316);
or U19403 (N_19403,N_19301,N_19277);
xor U19404 (N_19404,N_19303,N_19295);
and U19405 (N_19405,N_19226,N_19248);
or U19406 (N_19406,N_19221,N_19218);
nor U19407 (N_19407,N_19284,N_19322);
and U19408 (N_19408,N_19242,N_19227);
xnor U19409 (N_19409,N_19222,N_19326);
xor U19410 (N_19410,N_19209,N_19313);
nor U19411 (N_19411,N_19246,N_19267);
nand U19412 (N_19412,N_19217,N_19296);
or U19413 (N_19413,N_19308,N_19353);
xnor U19414 (N_19414,N_19312,N_19234);
xnor U19415 (N_19415,N_19212,N_19250);
or U19416 (N_19416,N_19228,N_19257);
nor U19417 (N_19417,N_19333,N_19278);
nor U19418 (N_19418,N_19321,N_19252);
nand U19419 (N_19419,N_19359,N_19223);
nand U19420 (N_19420,N_19229,N_19203);
nand U19421 (N_19421,N_19288,N_19319);
nand U19422 (N_19422,N_19351,N_19344);
and U19423 (N_19423,N_19213,N_19276);
nand U19424 (N_19424,N_19310,N_19245);
xor U19425 (N_19425,N_19323,N_19206);
or U19426 (N_19426,N_19335,N_19334);
or U19427 (N_19427,N_19241,N_19293);
nor U19428 (N_19428,N_19302,N_19282);
nor U19429 (N_19429,N_19304,N_19286);
nor U19430 (N_19430,N_19270,N_19261);
and U19431 (N_19431,N_19258,N_19328);
xnor U19432 (N_19432,N_19249,N_19331);
nor U19433 (N_19433,N_19339,N_19274);
or U19434 (N_19434,N_19306,N_19253);
and U19435 (N_19435,N_19273,N_19207);
nand U19436 (N_19436,N_19205,N_19309);
or U19437 (N_19437,N_19342,N_19211);
nand U19438 (N_19438,N_19281,N_19315);
nor U19439 (N_19439,N_19256,N_19338);
nand U19440 (N_19440,N_19204,N_19281);
and U19441 (N_19441,N_19326,N_19233);
or U19442 (N_19442,N_19202,N_19261);
and U19443 (N_19443,N_19312,N_19228);
xor U19444 (N_19444,N_19287,N_19220);
or U19445 (N_19445,N_19284,N_19297);
or U19446 (N_19446,N_19305,N_19220);
and U19447 (N_19447,N_19264,N_19317);
nand U19448 (N_19448,N_19314,N_19329);
nor U19449 (N_19449,N_19283,N_19244);
xor U19450 (N_19450,N_19335,N_19253);
and U19451 (N_19451,N_19240,N_19315);
and U19452 (N_19452,N_19233,N_19236);
or U19453 (N_19453,N_19308,N_19329);
nand U19454 (N_19454,N_19329,N_19260);
xor U19455 (N_19455,N_19316,N_19241);
nand U19456 (N_19456,N_19212,N_19236);
xnor U19457 (N_19457,N_19207,N_19309);
or U19458 (N_19458,N_19346,N_19285);
nor U19459 (N_19459,N_19265,N_19250);
nor U19460 (N_19460,N_19275,N_19337);
nand U19461 (N_19461,N_19318,N_19311);
and U19462 (N_19462,N_19328,N_19220);
xnor U19463 (N_19463,N_19203,N_19338);
nand U19464 (N_19464,N_19233,N_19273);
nand U19465 (N_19465,N_19331,N_19203);
and U19466 (N_19466,N_19287,N_19359);
xnor U19467 (N_19467,N_19254,N_19244);
nor U19468 (N_19468,N_19247,N_19212);
nor U19469 (N_19469,N_19324,N_19284);
or U19470 (N_19470,N_19286,N_19357);
or U19471 (N_19471,N_19293,N_19298);
or U19472 (N_19472,N_19286,N_19354);
xor U19473 (N_19473,N_19208,N_19203);
nor U19474 (N_19474,N_19205,N_19276);
xor U19475 (N_19475,N_19258,N_19269);
nand U19476 (N_19476,N_19260,N_19296);
nand U19477 (N_19477,N_19299,N_19324);
nor U19478 (N_19478,N_19243,N_19326);
xnor U19479 (N_19479,N_19218,N_19324);
nor U19480 (N_19480,N_19323,N_19261);
or U19481 (N_19481,N_19227,N_19222);
or U19482 (N_19482,N_19212,N_19307);
and U19483 (N_19483,N_19205,N_19240);
and U19484 (N_19484,N_19223,N_19336);
or U19485 (N_19485,N_19235,N_19236);
xor U19486 (N_19486,N_19295,N_19216);
or U19487 (N_19487,N_19239,N_19263);
and U19488 (N_19488,N_19240,N_19271);
or U19489 (N_19489,N_19317,N_19287);
and U19490 (N_19490,N_19342,N_19299);
nand U19491 (N_19491,N_19297,N_19350);
or U19492 (N_19492,N_19230,N_19263);
nor U19493 (N_19493,N_19274,N_19324);
nor U19494 (N_19494,N_19357,N_19289);
xnor U19495 (N_19495,N_19253,N_19318);
nand U19496 (N_19496,N_19275,N_19278);
and U19497 (N_19497,N_19208,N_19303);
or U19498 (N_19498,N_19347,N_19281);
nor U19499 (N_19499,N_19306,N_19211);
xor U19500 (N_19500,N_19215,N_19345);
xnor U19501 (N_19501,N_19260,N_19208);
nor U19502 (N_19502,N_19300,N_19277);
and U19503 (N_19503,N_19310,N_19206);
or U19504 (N_19504,N_19293,N_19254);
xnor U19505 (N_19505,N_19244,N_19285);
and U19506 (N_19506,N_19264,N_19217);
nand U19507 (N_19507,N_19304,N_19242);
and U19508 (N_19508,N_19239,N_19303);
nand U19509 (N_19509,N_19345,N_19280);
or U19510 (N_19510,N_19314,N_19303);
or U19511 (N_19511,N_19312,N_19233);
nor U19512 (N_19512,N_19238,N_19271);
or U19513 (N_19513,N_19276,N_19235);
nand U19514 (N_19514,N_19262,N_19241);
nor U19515 (N_19515,N_19249,N_19292);
and U19516 (N_19516,N_19320,N_19256);
xor U19517 (N_19517,N_19313,N_19237);
or U19518 (N_19518,N_19223,N_19207);
and U19519 (N_19519,N_19256,N_19236);
xor U19520 (N_19520,N_19446,N_19404);
xnor U19521 (N_19521,N_19459,N_19429);
xor U19522 (N_19522,N_19391,N_19440);
nand U19523 (N_19523,N_19431,N_19500);
nor U19524 (N_19524,N_19448,N_19490);
xor U19525 (N_19525,N_19464,N_19360);
xor U19526 (N_19526,N_19513,N_19465);
xnor U19527 (N_19527,N_19518,N_19410);
nand U19528 (N_19528,N_19373,N_19478);
nor U19529 (N_19529,N_19496,N_19408);
nor U19530 (N_19530,N_19378,N_19432);
or U19531 (N_19531,N_19427,N_19503);
nor U19532 (N_19532,N_19475,N_19425);
xnor U19533 (N_19533,N_19382,N_19415);
or U19534 (N_19534,N_19435,N_19483);
xnor U19535 (N_19535,N_19460,N_19441);
nor U19536 (N_19536,N_19477,N_19470);
nor U19537 (N_19537,N_19456,N_19388);
nor U19538 (N_19538,N_19514,N_19376);
xnor U19539 (N_19539,N_19380,N_19406);
and U19540 (N_19540,N_19368,N_19419);
xnor U19541 (N_19541,N_19467,N_19366);
nor U19542 (N_19542,N_19442,N_19507);
and U19543 (N_19543,N_19371,N_19369);
or U19544 (N_19544,N_19422,N_19519);
nor U19545 (N_19545,N_19384,N_19455);
xnor U19546 (N_19546,N_19430,N_19449);
and U19547 (N_19547,N_19486,N_19481);
or U19548 (N_19548,N_19372,N_19361);
and U19549 (N_19549,N_19454,N_19386);
and U19550 (N_19550,N_19396,N_19472);
and U19551 (N_19551,N_19511,N_19428);
and U19552 (N_19552,N_19392,N_19497);
nand U19553 (N_19553,N_19479,N_19484);
xor U19554 (N_19554,N_19461,N_19405);
and U19555 (N_19555,N_19482,N_19379);
or U19556 (N_19556,N_19385,N_19375);
nand U19557 (N_19557,N_19444,N_19466);
nand U19558 (N_19558,N_19416,N_19468);
or U19559 (N_19559,N_19504,N_19399);
nand U19560 (N_19560,N_19499,N_19510);
nand U19561 (N_19561,N_19393,N_19493);
xor U19562 (N_19562,N_19515,N_19364);
xnor U19563 (N_19563,N_19502,N_19395);
nand U19564 (N_19564,N_19426,N_19495);
or U19565 (N_19565,N_19506,N_19407);
nor U19566 (N_19566,N_19485,N_19409);
nand U19567 (N_19567,N_19443,N_19417);
and U19568 (N_19568,N_19452,N_19457);
nand U19569 (N_19569,N_19420,N_19474);
and U19570 (N_19570,N_19411,N_19492);
nor U19571 (N_19571,N_19505,N_19402);
nor U19572 (N_19572,N_19381,N_19400);
or U19573 (N_19573,N_19480,N_19494);
nand U19574 (N_19574,N_19383,N_19473);
nor U19575 (N_19575,N_19390,N_19398);
nand U19576 (N_19576,N_19451,N_19374);
or U19577 (N_19577,N_19471,N_19387);
and U19578 (N_19578,N_19362,N_19487);
xnor U19579 (N_19579,N_19516,N_19447);
xnor U19580 (N_19580,N_19450,N_19517);
nor U19581 (N_19581,N_19438,N_19401);
or U19582 (N_19582,N_19489,N_19434);
xnor U19583 (N_19583,N_19508,N_19445);
nand U19584 (N_19584,N_19509,N_19458);
nor U19585 (N_19585,N_19453,N_19365);
xnor U19586 (N_19586,N_19367,N_19476);
or U19587 (N_19587,N_19418,N_19370);
nor U19588 (N_19588,N_19436,N_19498);
xnor U19589 (N_19589,N_19363,N_19394);
nor U19590 (N_19590,N_19433,N_19421);
and U19591 (N_19591,N_19389,N_19512);
nor U19592 (N_19592,N_19491,N_19414);
xnor U19593 (N_19593,N_19423,N_19501);
and U19594 (N_19594,N_19437,N_19424);
nor U19595 (N_19595,N_19403,N_19377);
nor U19596 (N_19596,N_19397,N_19463);
and U19597 (N_19597,N_19413,N_19488);
xnor U19598 (N_19598,N_19462,N_19412);
nand U19599 (N_19599,N_19439,N_19469);
nor U19600 (N_19600,N_19470,N_19371);
xor U19601 (N_19601,N_19420,N_19518);
nand U19602 (N_19602,N_19512,N_19387);
and U19603 (N_19603,N_19460,N_19462);
nor U19604 (N_19604,N_19483,N_19404);
nor U19605 (N_19605,N_19395,N_19433);
xnor U19606 (N_19606,N_19504,N_19453);
nor U19607 (N_19607,N_19417,N_19362);
nor U19608 (N_19608,N_19387,N_19433);
and U19609 (N_19609,N_19459,N_19490);
or U19610 (N_19610,N_19388,N_19430);
and U19611 (N_19611,N_19381,N_19419);
nand U19612 (N_19612,N_19404,N_19376);
xor U19613 (N_19613,N_19365,N_19510);
nor U19614 (N_19614,N_19379,N_19425);
and U19615 (N_19615,N_19510,N_19405);
nor U19616 (N_19616,N_19461,N_19477);
or U19617 (N_19617,N_19392,N_19455);
nor U19618 (N_19618,N_19386,N_19515);
or U19619 (N_19619,N_19473,N_19409);
and U19620 (N_19620,N_19417,N_19391);
xor U19621 (N_19621,N_19470,N_19459);
xnor U19622 (N_19622,N_19471,N_19505);
nand U19623 (N_19623,N_19382,N_19507);
nand U19624 (N_19624,N_19477,N_19410);
nor U19625 (N_19625,N_19435,N_19412);
xnor U19626 (N_19626,N_19398,N_19478);
and U19627 (N_19627,N_19412,N_19468);
xor U19628 (N_19628,N_19423,N_19518);
xnor U19629 (N_19629,N_19442,N_19401);
nand U19630 (N_19630,N_19390,N_19439);
and U19631 (N_19631,N_19360,N_19408);
and U19632 (N_19632,N_19479,N_19451);
xnor U19633 (N_19633,N_19478,N_19472);
nand U19634 (N_19634,N_19471,N_19487);
nor U19635 (N_19635,N_19508,N_19484);
or U19636 (N_19636,N_19370,N_19383);
nor U19637 (N_19637,N_19379,N_19486);
nor U19638 (N_19638,N_19370,N_19368);
and U19639 (N_19639,N_19467,N_19510);
and U19640 (N_19640,N_19433,N_19462);
or U19641 (N_19641,N_19398,N_19497);
or U19642 (N_19642,N_19451,N_19420);
nand U19643 (N_19643,N_19507,N_19398);
nor U19644 (N_19644,N_19426,N_19513);
or U19645 (N_19645,N_19442,N_19371);
or U19646 (N_19646,N_19397,N_19425);
and U19647 (N_19647,N_19483,N_19516);
nand U19648 (N_19648,N_19392,N_19502);
nor U19649 (N_19649,N_19397,N_19458);
or U19650 (N_19650,N_19496,N_19460);
or U19651 (N_19651,N_19491,N_19366);
xor U19652 (N_19652,N_19452,N_19398);
xor U19653 (N_19653,N_19515,N_19471);
nor U19654 (N_19654,N_19412,N_19373);
nor U19655 (N_19655,N_19451,N_19405);
xor U19656 (N_19656,N_19441,N_19400);
xor U19657 (N_19657,N_19365,N_19487);
xnor U19658 (N_19658,N_19421,N_19436);
xnor U19659 (N_19659,N_19474,N_19490);
and U19660 (N_19660,N_19481,N_19420);
nor U19661 (N_19661,N_19461,N_19377);
nor U19662 (N_19662,N_19425,N_19484);
and U19663 (N_19663,N_19455,N_19510);
xor U19664 (N_19664,N_19474,N_19363);
or U19665 (N_19665,N_19400,N_19458);
xnor U19666 (N_19666,N_19500,N_19475);
xor U19667 (N_19667,N_19497,N_19461);
and U19668 (N_19668,N_19431,N_19511);
nand U19669 (N_19669,N_19469,N_19518);
or U19670 (N_19670,N_19480,N_19409);
or U19671 (N_19671,N_19362,N_19437);
nor U19672 (N_19672,N_19493,N_19446);
xor U19673 (N_19673,N_19378,N_19413);
nor U19674 (N_19674,N_19432,N_19430);
nor U19675 (N_19675,N_19407,N_19409);
xnor U19676 (N_19676,N_19426,N_19396);
or U19677 (N_19677,N_19509,N_19364);
and U19678 (N_19678,N_19400,N_19492);
xor U19679 (N_19679,N_19397,N_19486);
or U19680 (N_19680,N_19521,N_19665);
nand U19681 (N_19681,N_19547,N_19587);
and U19682 (N_19682,N_19673,N_19533);
nor U19683 (N_19683,N_19544,N_19607);
nor U19684 (N_19684,N_19550,N_19634);
xnor U19685 (N_19685,N_19568,N_19605);
or U19686 (N_19686,N_19576,N_19558);
xnor U19687 (N_19687,N_19623,N_19647);
nor U19688 (N_19688,N_19584,N_19604);
or U19689 (N_19689,N_19597,N_19659);
and U19690 (N_19690,N_19581,N_19552);
nor U19691 (N_19691,N_19598,N_19572);
nor U19692 (N_19692,N_19535,N_19556);
nor U19693 (N_19693,N_19608,N_19593);
or U19694 (N_19694,N_19588,N_19583);
xnor U19695 (N_19695,N_19624,N_19592);
nor U19696 (N_19696,N_19649,N_19632);
xor U19697 (N_19697,N_19655,N_19662);
and U19698 (N_19698,N_19609,N_19525);
nand U19699 (N_19699,N_19667,N_19548);
nor U19700 (N_19700,N_19668,N_19633);
nand U19701 (N_19701,N_19560,N_19612);
nand U19702 (N_19702,N_19606,N_19637);
or U19703 (N_19703,N_19651,N_19557);
or U19704 (N_19704,N_19575,N_19636);
nand U19705 (N_19705,N_19528,N_19677);
and U19706 (N_19706,N_19554,N_19627);
nor U19707 (N_19707,N_19582,N_19546);
xor U19708 (N_19708,N_19621,N_19644);
and U19709 (N_19709,N_19566,N_19561);
or U19710 (N_19710,N_19646,N_19524);
xnor U19711 (N_19711,N_19617,N_19589);
nor U19712 (N_19712,N_19594,N_19578);
nand U19713 (N_19713,N_19615,N_19553);
nor U19714 (N_19714,N_19601,N_19603);
nor U19715 (N_19715,N_19564,N_19643);
and U19716 (N_19716,N_19529,N_19551);
xor U19717 (N_19717,N_19642,N_19611);
and U19718 (N_19718,N_19658,N_19559);
or U19719 (N_19719,N_19574,N_19657);
and U19720 (N_19720,N_19674,N_19676);
nand U19721 (N_19721,N_19650,N_19540);
nor U19722 (N_19722,N_19549,N_19602);
nor U19723 (N_19723,N_19570,N_19579);
or U19724 (N_19724,N_19590,N_19675);
nand U19725 (N_19725,N_19563,N_19670);
and U19726 (N_19726,N_19613,N_19616);
nand U19727 (N_19727,N_19653,N_19671);
nand U19728 (N_19728,N_19573,N_19539);
nor U19729 (N_19729,N_19620,N_19577);
and U19730 (N_19730,N_19585,N_19625);
or U19731 (N_19731,N_19523,N_19619);
and U19732 (N_19732,N_19640,N_19654);
xnor U19733 (N_19733,N_19520,N_19538);
nand U19734 (N_19734,N_19660,N_19522);
and U19735 (N_19735,N_19536,N_19586);
nor U19736 (N_19736,N_19663,N_19638);
nor U19737 (N_19737,N_19618,N_19530);
or U19738 (N_19738,N_19543,N_19562);
nand U19739 (N_19739,N_19645,N_19567);
nand U19740 (N_19740,N_19648,N_19629);
nand U19741 (N_19741,N_19641,N_19595);
xnor U19742 (N_19742,N_19532,N_19537);
nand U19743 (N_19743,N_19542,N_19652);
nor U19744 (N_19744,N_19669,N_19639);
and U19745 (N_19745,N_19630,N_19596);
nor U19746 (N_19746,N_19678,N_19565);
nor U19747 (N_19747,N_19580,N_19679);
nor U19748 (N_19748,N_19614,N_19628);
or U19749 (N_19749,N_19610,N_19666);
xnor U19750 (N_19750,N_19545,N_19600);
or U19751 (N_19751,N_19569,N_19599);
and U19752 (N_19752,N_19672,N_19555);
nand U19753 (N_19753,N_19622,N_19571);
and U19754 (N_19754,N_19526,N_19661);
nor U19755 (N_19755,N_19664,N_19591);
nand U19756 (N_19756,N_19541,N_19635);
and U19757 (N_19757,N_19656,N_19527);
and U19758 (N_19758,N_19626,N_19534);
and U19759 (N_19759,N_19631,N_19531);
xnor U19760 (N_19760,N_19547,N_19528);
nor U19761 (N_19761,N_19610,N_19533);
or U19762 (N_19762,N_19646,N_19637);
xnor U19763 (N_19763,N_19545,N_19638);
nor U19764 (N_19764,N_19531,N_19521);
nor U19765 (N_19765,N_19627,N_19536);
nor U19766 (N_19766,N_19618,N_19632);
and U19767 (N_19767,N_19562,N_19566);
and U19768 (N_19768,N_19539,N_19659);
xnor U19769 (N_19769,N_19635,N_19561);
nor U19770 (N_19770,N_19525,N_19651);
xor U19771 (N_19771,N_19658,N_19670);
nor U19772 (N_19772,N_19542,N_19559);
xnor U19773 (N_19773,N_19631,N_19598);
nor U19774 (N_19774,N_19635,N_19628);
xor U19775 (N_19775,N_19572,N_19587);
or U19776 (N_19776,N_19677,N_19592);
or U19777 (N_19777,N_19598,N_19531);
nor U19778 (N_19778,N_19628,N_19578);
xnor U19779 (N_19779,N_19639,N_19663);
or U19780 (N_19780,N_19543,N_19560);
or U19781 (N_19781,N_19563,N_19654);
or U19782 (N_19782,N_19617,N_19522);
or U19783 (N_19783,N_19620,N_19613);
and U19784 (N_19784,N_19677,N_19652);
or U19785 (N_19785,N_19604,N_19663);
and U19786 (N_19786,N_19619,N_19590);
xnor U19787 (N_19787,N_19660,N_19600);
xor U19788 (N_19788,N_19606,N_19542);
nor U19789 (N_19789,N_19618,N_19575);
nand U19790 (N_19790,N_19672,N_19569);
nor U19791 (N_19791,N_19604,N_19628);
and U19792 (N_19792,N_19560,N_19634);
or U19793 (N_19793,N_19672,N_19563);
or U19794 (N_19794,N_19583,N_19672);
nor U19795 (N_19795,N_19542,N_19560);
nor U19796 (N_19796,N_19523,N_19584);
xnor U19797 (N_19797,N_19585,N_19609);
nand U19798 (N_19798,N_19639,N_19588);
xor U19799 (N_19799,N_19530,N_19521);
nor U19800 (N_19800,N_19545,N_19588);
nor U19801 (N_19801,N_19669,N_19577);
nand U19802 (N_19802,N_19634,N_19556);
xnor U19803 (N_19803,N_19549,N_19615);
nand U19804 (N_19804,N_19566,N_19528);
nand U19805 (N_19805,N_19597,N_19576);
nor U19806 (N_19806,N_19594,N_19662);
nor U19807 (N_19807,N_19678,N_19673);
and U19808 (N_19808,N_19529,N_19525);
nor U19809 (N_19809,N_19643,N_19585);
and U19810 (N_19810,N_19535,N_19673);
or U19811 (N_19811,N_19572,N_19535);
nand U19812 (N_19812,N_19630,N_19619);
and U19813 (N_19813,N_19561,N_19611);
and U19814 (N_19814,N_19658,N_19576);
xor U19815 (N_19815,N_19666,N_19552);
and U19816 (N_19816,N_19642,N_19637);
xor U19817 (N_19817,N_19585,N_19570);
or U19818 (N_19818,N_19663,N_19659);
nand U19819 (N_19819,N_19530,N_19676);
nor U19820 (N_19820,N_19588,N_19541);
nand U19821 (N_19821,N_19627,N_19679);
nand U19822 (N_19822,N_19564,N_19524);
or U19823 (N_19823,N_19666,N_19527);
nor U19824 (N_19824,N_19628,N_19665);
xor U19825 (N_19825,N_19668,N_19625);
or U19826 (N_19826,N_19612,N_19656);
xnor U19827 (N_19827,N_19613,N_19584);
or U19828 (N_19828,N_19548,N_19565);
and U19829 (N_19829,N_19560,N_19551);
and U19830 (N_19830,N_19598,N_19659);
or U19831 (N_19831,N_19630,N_19652);
nor U19832 (N_19832,N_19607,N_19589);
and U19833 (N_19833,N_19531,N_19544);
or U19834 (N_19834,N_19524,N_19614);
nor U19835 (N_19835,N_19649,N_19614);
xor U19836 (N_19836,N_19649,N_19607);
nand U19837 (N_19837,N_19630,N_19651);
nor U19838 (N_19838,N_19549,N_19556);
and U19839 (N_19839,N_19560,N_19533);
and U19840 (N_19840,N_19722,N_19830);
and U19841 (N_19841,N_19768,N_19711);
nor U19842 (N_19842,N_19764,N_19693);
and U19843 (N_19843,N_19833,N_19705);
and U19844 (N_19844,N_19834,N_19818);
nor U19845 (N_19845,N_19728,N_19813);
nor U19846 (N_19846,N_19797,N_19757);
and U19847 (N_19847,N_19788,N_19742);
nor U19848 (N_19848,N_19782,N_19785);
nand U19849 (N_19849,N_19831,N_19791);
xor U19850 (N_19850,N_19789,N_19832);
nand U19851 (N_19851,N_19766,N_19718);
xor U19852 (N_19852,N_19765,N_19695);
xnor U19853 (N_19853,N_19809,N_19773);
xor U19854 (N_19854,N_19721,N_19746);
nor U19855 (N_19855,N_19822,N_19755);
nor U19856 (N_19856,N_19786,N_19681);
or U19857 (N_19857,N_19752,N_19688);
or U19858 (N_19858,N_19686,N_19716);
or U19859 (N_19859,N_19698,N_19814);
nor U19860 (N_19860,N_19747,N_19826);
xnor U19861 (N_19861,N_19827,N_19729);
or U19862 (N_19862,N_19710,N_19808);
xor U19863 (N_19863,N_19720,N_19800);
and U19864 (N_19864,N_19704,N_19749);
nor U19865 (N_19865,N_19811,N_19709);
nor U19866 (N_19866,N_19776,N_19798);
or U19867 (N_19867,N_19683,N_19707);
and U19868 (N_19868,N_19815,N_19825);
and U19869 (N_19869,N_19682,N_19781);
or U19870 (N_19870,N_19696,N_19812);
nand U19871 (N_19871,N_19684,N_19802);
nand U19872 (N_19872,N_19769,N_19741);
or U19873 (N_19873,N_19738,N_19706);
xor U19874 (N_19874,N_19807,N_19767);
xnor U19875 (N_19875,N_19734,N_19803);
and U19876 (N_19876,N_19771,N_19794);
xor U19877 (N_19877,N_19816,N_19839);
or U19878 (N_19878,N_19689,N_19737);
or U19879 (N_19879,N_19837,N_19719);
or U19880 (N_19880,N_19730,N_19753);
and U19881 (N_19881,N_19743,N_19701);
or U19882 (N_19882,N_19784,N_19817);
xnor U19883 (N_19883,N_19732,N_19714);
and U19884 (N_19884,N_19787,N_19733);
nand U19885 (N_19885,N_19713,N_19799);
or U19886 (N_19886,N_19770,N_19692);
and U19887 (N_19887,N_19751,N_19823);
or U19888 (N_19888,N_19775,N_19685);
nor U19889 (N_19889,N_19762,N_19806);
xnor U19890 (N_19890,N_19715,N_19758);
xor U19891 (N_19891,N_19779,N_19820);
and U19892 (N_19892,N_19805,N_19736);
and U19893 (N_19893,N_19744,N_19703);
and U19894 (N_19894,N_19810,N_19801);
and U19895 (N_19895,N_19819,N_19778);
xor U19896 (N_19896,N_19793,N_19724);
or U19897 (N_19897,N_19694,N_19739);
or U19898 (N_19898,N_19700,N_19804);
nor U19899 (N_19899,N_19780,N_19726);
nand U19900 (N_19900,N_19763,N_19836);
or U19901 (N_19901,N_19756,N_19783);
and U19902 (N_19902,N_19690,N_19829);
and U19903 (N_19903,N_19761,N_19774);
nor U19904 (N_19904,N_19699,N_19754);
nor U19905 (N_19905,N_19759,N_19727);
or U19906 (N_19906,N_19697,N_19702);
and U19907 (N_19907,N_19687,N_19680);
nand U19908 (N_19908,N_19795,N_19835);
nor U19909 (N_19909,N_19838,N_19717);
nand U19910 (N_19910,N_19723,N_19828);
or U19911 (N_19911,N_19790,N_19725);
xnor U19912 (N_19912,N_19745,N_19708);
or U19913 (N_19913,N_19824,N_19796);
nor U19914 (N_19914,N_19731,N_19691);
or U19915 (N_19915,N_19777,N_19792);
nand U19916 (N_19916,N_19740,N_19712);
nor U19917 (N_19917,N_19760,N_19821);
and U19918 (N_19918,N_19750,N_19748);
or U19919 (N_19919,N_19772,N_19735);
nor U19920 (N_19920,N_19837,N_19783);
or U19921 (N_19921,N_19690,N_19729);
xor U19922 (N_19922,N_19808,N_19690);
or U19923 (N_19923,N_19693,N_19837);
xnor U19924 (N_19924,N_19800,N_19731);
nor U19925 (N_19925,N_19730,N_19809);
and U19926 (N_19926,N_19752,N_19797);
or U19927 (N_19927,N_19806,N_19750);
and U19928 (N_19928,N_19727,N_19735);
nand U19929 (N_19929,N_19832,N_19805);
nor U19930 (N_19930,N_19812,N_19735);
or U19931 (N_19931,N_19710,N_19688);
nand U19932 (N_19932,N_19738,N_19703);
or U19933 (N_19933,N_19712,N_19816);
nor U19934 (N_19934,N_19799,N_19839);
and U19935 (N_19935,N_19691,N_19680);
and U19936 (N_19936,N_19739,N_19683);
nand U19937 (N_19937,N_19822,N_19700);
nor U19938 (N_19938,N_19815,N_19716);
nand U19939 (N_19939,N_19696,N_19714);
and U19940 (N_19940,N_19826,N_19817);
nor U19941 (N_19941,N_19748,N_19797);
or U19942 (N_19942,N_19798,N_19801);
and U19943 (N_19943,N_19691,N_19764);
xnor U19944 (N_19944,N_19811,N_19737);
and U19945 (N_19945,N_19777,N_19754);
or U19946 (N_19946,N_19770,N_19767);
xor U19947 (N_19947,N_19758,N_19805);
or U19948 (N_19948,N_19721,N_19700);
xnor U19949 (N_19949,N_19708,N_19823);
nand U19950 (N_19950,N_19734,N_19818);
nand U19951 (N_19951,N_19689,N_19693);
nor U19952 (N_19952,N_19807,N_19697);
nor U19953 (N_19953,N_19723,N_19777);
or U19954 (N_19954,N_19697,N_19830);
xor U19955 (N_19955,N_19741,N_19703);
or U19956 (N_19956,N_19766,N_19801);
nor U19957 (N_19957,N_19801,N_19826);
and U19958 (N_19958,N_19757,N_19809);
or U19959 (N_19959,N_19696,N_19725);
nor U19960 (N_19960,N_19819,N_19817);
xor U19961 (N_19961,N_19744,N_19756);
and U19962 (N_19962,N_19819,N_19804);
nand U19963 (N_19963,N_19767,N_19813);
nand U19964 (N_19964,N_19825,N_19786);
and U19965 (N_19965,N_19794,N_19709);
nor U19966 (N_19966,N_19791,N_19688);
nor U19967 (N_19967,N_19795,N_19723);
nor U19968 (N_19968,N_19758,N_19706);
nand U19969 (N_19969,N_19695,N_19782);
and U19970 (N_19970,N_19745,N_19819);
or U19971 (N_19971,N_19732,N_19724);
xor U19972 (N_19972,N_19712,N_19810);
xnor U19973 (N_19973,N_19729,N_19715);
or U19974 (N_19974,N_19723,N_19715);
nand U19975 (N_19975,N_19697,N_19794);
and U19976 (N_19976,N_19702,N_19729);
nor U19977 (N_19977,N_19744,N_19773);
nor U19978 (N_19978,N_19705,N_19744);
nor U19979 (N_19979,N_19743,N_19720);
nand U19980 (N_19980,N_19834,N_19687);
nor U19981 (N_19981,N_19752,N_19798);
nor U19982 (N_19982,N_19820,N_19707);
nor U19983 (N_19983,N_19683,N_19823);
nor U19984 (N_19984,N_19701,N_19718);
nand U19985 (N_19985,N_19747,N_19794);
nor U19986 (N_19986,N_19785,N_19706);
nand U19987 (N_19987,N_19826,N_19824);
xnor U19988 (N_19988,N_19802,N_19771);
or U19989 (N_19989,N_19713,N_19787);
and U19990 (N_19990,N_19756,N_19812);
and U19991 (N_19991,N_19803,N_19802);
and U19992 (N_19992,N_19839,N_19819);
nand U19993 (N_19993,N_19798,N_19684);
nor U19994 (N_19994,N_19839,N_19762);
nor U19995 (N_19995,N_19680,N_19732);
nand U19996 (N_19996,N_19734,N_19777);
nor U19997 (N_19997,N_19699,N_19766);
nand U19998 (N_19998,N_19737,N_19807);
or U19999 (N_19999,N_19700,N_19719);
and UO_0 (O_0,N_19958,N_19949);
or UO_1 (O_1,N_19950,N_19966);
and UO_2 (O_2,N_19849,N_19888);
xnor UO_3 (O_3,N_19922,N_19940);
and UO_4 (O_4,N_19901,N_19970);
xor UO_5 (O_5,N_19868,N_19998);
and UO_6 (O_6,N_19963,N_19904);
nor UO_7 (O_7,N_19864,N_19858);
and UO_8 (O_8,N_19905,N_19895);
and UO_9 (O_9,N_19915,N_19969);
nand UO_10 (O_10,N_19981,N_19846);
xor UO_11 (O_11,N_19920,N_19861);
nor UO_12 (O_12,N_19926,N_19947);
nand UO_13 (O_13,N_19857,N_19840);
and UO_14 (O_14,N_19885,N_19870);
nor UO_15 (O_15,N_19860,N_19989);
xor UO_16 (O_16,N_19965,N_19909);
nand UO_17 (O_17,N_19929,N_19863);
and UO_18 (O_18,N_19900,N_19985);
or UO_19 (O_19,N_19884,N_19906);
and UO_20 (O_20,N_19976,N_19956);
nor UO_21 (O_21,N_19918,N_19961);
nor UO_22 (O_22,N_19960,N_19903);
or UO_23 (O_23,N_19973,N_19944);
xor UO_24 (O_24,N_19933,N_19982);
nand UO_25 (O_25,N_19879,N_19913);
nand UO_26 (O_26,N_19843,N_19853);
nand UO_27 (O_27,N_19942,N_19978);
or UO_28 (O_28,N_19893,N_19877);
nor UO_29 (O_29,N_19980,N_19996);
and UO_30 (O_30,N_19862,N_19934);
nor UO_31 (O_31,N_19971,N_19919);
nand UO_32 (O_32,N_19931,N_19859);
nor UO_33 (O_33,N_19995,N_19943);
or UO_34 (O_34,N_19937,N_19991);
or UO_35 (O_35,N_19867,N_19880);
nor UO_36 (O_36,N_19842,N_19964);
nand UO_37 (O_37,N_19923,N_19921);
or UO_38 (O_38,N_19911,N_19951);
xnor UO_39 (O_39,N_19898,N_19962);
and UO_40 (O_40,N_19854,N_19852);
xor UO_41 (O_41,N_19955,N_19959);
and UO_42 (O_42,N_19994,N_19939);
nand UO_43 (O_43,N_19850,N_19845);
xnor UO_44 (O_44,N_19882,N_19897);
xor UO_45 (O_45,N_19841,N_19914);
nand UO_46 (O_46,N_19986,N_19935);
nand UO_47 (O_47,N_19872,N_19992);
nor UO_48 (O_48,N_19881,N_19952);
nor UO_49 (O_49,N_19987,N_19948);
nand UO_50 (O_50,N_19945,N_19907);
and UO_51 (O_51,N_19924,N_19957);
or UO_52 (O_52,N_19856,N_19938);
and UO_53 (O_53,N_19878,N_19902);
xor UO_54 (O_54,N_19889,N_19848);
or UO_55 (O_55,N_19874,N_19925);
nand UO_56 (O_56,N_19855,N_19917);
xnor UO_57 (O_57,N_19984,N_19977);
and UO_58 (O_58,N_19967,N_19930);
nand UO_59 (O_59,N_19896,N_19869);
or UO_60 (O_60,N_19997,N_19993);
xnor UO_61 (O_61,N_19891,N_19871);
nand UO_62 (O_62,N_19953,N_19873);
nor UO_63 (O_63,N_19890,N_19908);
xor UO_64 (O_64,N_19975,N_19876);
or UO_65 (O_65,N_19968,N_19886);
nand UO_66 (O_66,N_19972,N_19892);
xnor UO_67 (O_67,N_19927,N_19999);
nand UO_68 (O_68,N_19910,N_19979);
nor UO_69 (O_69,N_19954,N_19988);
nor UO_70 (O_70,N_19916,N_19912);
and UO_71 (O_71,N_19936,N_19883);
nand UO_72 (O_72,N_19899,N_19932);
and UO_73 (O_73,N_19928,N_19847);
nor UO_74 (O_74,N_19894,N_19887);
nor UO_75 (O_75,N_19875,N_19974);
xnor UO_76 (O_76,N_19990,N_19851);
xor UO_77 (O_77,N_19865,N_19983);
and UO_78 (O_78,N_19866,N_19941);
or UO_79 (O_79,N_19844,N_19946);
or UO_80 (O_80,N_19877,N_19923);
or UO_81 (O_81,N_19852,N_19952);
and UO_82 (O_82,N_19891,N_19845);
nand UO_83 (O_83,N_19934,N_19848);
or UO_84 (O_84,N_19864,N_19887);
and UO_85 (O_85,N_19870,N_19929);
nor UO_86 (O_86,N_19918,N_19871);
and UO_87 (O_87,N_19937,N_19959);
and UO_88 (O_88,N_19866,N_19888);
nor UO_89 (O_89,N_19957,N_19976);
nand UO_90 (O_90,N_19965,N_19954);
xnor UO_91 (O_91,N_19888,N_19936);
nor UO_92 (O_92,N_19882,N_19970);
or UO_93 (O_93,N_19998,N_19968);
or UO_94 (O_94,N_19890,N_19863);
nor UO_95 (O_95,N_19943,N_19870);
xnor UO_96 (O_96,N_19956,N_19985);
or UO_97 (O_97,N_19955,N_19942);
nand UO_98 (O_98,N_19863,N_19970);
nor UO_99 (O_99,N_19921,N_19922);
xnor UO_100 (O_100,N_19913,N_19877);
nor UO_101 (O_101,N_19913,N_19937);
xor UO_102 (O_102,N_19997,N_19863);
and UO_103 (O_103,N_19989,N_19887);
nand UO_104 (O_104,N_19870,N_19867);
nand UO_105 (O_105,N_19873,N_19977);
and UO_106 (O_106,N_19863,N_19954);
or UO_107 (O_107,N_19914,N_19957);
nand UO_108 (O_108,N_19913,N_19956);
nor UO_109 (O_109,N_19947,N_19973);
nand UO_110 (O_110,N_19900,N_19853);
or UO_111 (O_111,N_19886,N_19908);
or UO_112 (O_112,N_19852,N_19891);
nor UO_113 (O_113,N_19859,N_19867);
nor UO_114 (O_114,N_19911,N_19964);
and UO_115 (O_115,N_19901,N_19951);
nand UO_116 (O_116,N_19904,N_19921);
xor UO_117 (O_117,N_19989,N_19899);
nand UO_118 (O_118,N_19944,N_19843);
xor UO_119 (O_119,N_19962,N_19849);
nand UO_120 (O_120,N_19936,N_19876);
nor UO_121 (O_121,N_19977,N_19948);
nand UO_122 (O_122,N_19847,N_19976);
or UO_123 (O_123,N_19956,N_19894);
and UO_124 (O_124,N_19912,N_19915);
xor UO_125 (O_125,N_19873,N_19914);
and UO_126 (O_126,N_19947,N_19879);
nand UO_127 (O_127,N_19842,N_19962);
nand UO_128 (O_128,N_19939,N_19976);
or UO_129 (O_129,N_19950,N_19861);
or UO_130 (O_130,N_19878,N_19946);
nor UO_131 (O_131,N_19863,N_19877);
and UO_132 (O_132,N_19983,N_19977);
nand UO_133 (O_133,N_19958,N_19993);
xor UO_134 (O_134,N_19907,N_19927);
nand UO_135 (O_135,N_19991,N_19974);
xor UO_136 (O_136,N_19972,N_19979);
and UO_137 (O_137,N_19997,N_19852);
or UO_138 (O_138,N_19874,N_19917);
nand UO_139 (O_139,N_19877,N_19849);
nor UO_140 (O_140,N_19862,N_19933);
and UO_141 (O_141,N_19933,N_19928);
nor UO_142 (O_142,N_19948,N_19929);
xnor UO_143 (O_143,N_19983,N_19940);
nor UO_144 (O_144,N_19894,N_19983);
and UO_145 (O_145,N_19959,N_19889);
nand UO_146 (O_146,N_19880,N_19983);
nand UO_147 (O_147,N_19981,N_19843);
nand UO_148 (O_148,N_19847,N_19905);
and UO_149 (O_149,N_19854,N_19898);
nor UO_150 (O_150,N_19928,N_19990);
xor UO_151 (O_151,N_19985,N_19952);
nand UO_152 (O_152,N_19986,N_19966);
nand UO_153 (O_153,N_19984,N_19942);
nor UO_154 (O_154,N_19952,N_19942);
and UO_155 (O_155,N_19886,N_19930);
xnor UO_156 (O_156,N_19900,N_19876);
xnor UO_157 (O_157,N_19984,N_19941);
and UO_158 (O_158,N_19911,N_19893);
nand UO_159 (O_159,N_19889,N_19986);
nor UO_160 (O_160,N_19911,N_19902);
xnor UO_161 (O_161,N_19914,N_19945);
nor UO_162 (O_162,N_19943,N_19852);
nor UO_163 (O_163,N_19880,N_19995);
or UO_164 (O_164,N_19907,N_19897);
nor UO_165 (O_165,N_19875,N_19925);
xnor UO_166 (O_166,N_19866,N_19966);
and UO_167 (O_167,N_19888,N_19963);
nor UO_168 (O_168,N_19883,N_19892);
nor UO_169 (O_169,N_19888,N_19857);
or UO_170 (O_170,N_19858,N_19922);
and UO_171 (O_171,N_19888,N_19952);
and UO_172 (O_172,N_19939,N_19986);
nor UO_173 (O_173,N_19910,N_19916);
nand UO_174 (O_174,N_19986,N_19944);
xnor UO_175 (O_175,N_19945,N_19853);
xnor UO_176 (O_176,N_19985,N_19923);
nand UO_177 (O_177,N_19890,N_19897);
nand UO_178 (O_178,N_19995,N_19969);
nand UO_179 (O_179,N_19871,N_19929);
xnor UO_180 (O_180,N_19930,N_19994);
nand UO_181 (O_181,N_19914,N_19906);
xnor UO_182 (O_182,N_19969,N_19949);
or UO_183 (O_183,N_19998,N_19947);
and UO_184 (O_184,N_19924,N_19888);
nand UO_185 (O_185,N_19909,N_19916);
or UO_186 (O_186,N_19877,N_19844);
or UO_187 (O_187,N_19905,N_19928);
and UO_188 (O_188,N_19923,N_19864);
nor UO_189 (O_189,N_19944,N_19977);
xor UO_190 (O_190,N_19886,N_19852);
or UO_191 (O_191,N_19962,N_19868);
xor UO_192 (O_192,N_19950,N_19903);
xor UO_193 (O_193,N_19973,N_19955);
xor UO_194 (O_194,N_19883,N_19938);
or UO_195 (O_195,N_19893,N_19931);
or UO_196 (O_196,N_19946,N_19898);
nor UO_197 (O_197,N_19840,N_19924);
nor UO_198 (O_198,N_19938,N_19879);
nand UO_199 (O_199,N_19889,N_19863);
and UO_200 (O_200,N_19923,N_19958);
nor UO_201 (O_201,N_19973,N_19856);
or UO_202 (O_202,N_19874,N_19850);
and UO_203 (O_203,N_19897,N_19887);
nor UO_204 (O_204,N_19944,N_19976);
nand UO_205 (O_205,N_19991,N_19865);
xnor UO_206 (O_206,N_19986,N_19982);
or UO_207 (O_207,N_19845,N_19902);
and UO_208 (O_208,N_19903,N_19852);
and UO_209 (O_209,N_19883,N_19954);
or UO_210 (O_210,N_19852,N_19843);
and UO_211 (O_211,N_19992,N_19905);
nor UO_212 (O_212,N_19865,N_19968);
xnor UO_213 (O_213,N_19962,N_19993);
and UO_214 (O_214,N_19860,N_19881);
and UO_215 (O_215,N_19937,N_19905);
and UO_216 (O_216,N_19852,N_19932);
nor UO_217 (O_217,N_19989,N_19959);
nand UO_218 (O_218,N_19909,N_19973);
and UO_219 (O_219,N_19859,N_19892);
and UO_220 (O_220,N_19991,N_19993);
and UO_221 (O_221,N_19899,N_19884);
or UO_222 (O_222,N_19844,N_19996);
nand UO_223 (O_223,N_19849,N_19868);
nand UO_224 (O_224,N_19973,N_19921);
nor UO_225 (O_225,N_19961,N_19996);
xnor UO_226 (O_226,N_19972,N_19995);
nor UO_227 (O_227,N_19899,N_19942);
xor UO_228 (O_228,N_19896,N_19860);
or UO_229 (O_229,N_19896,N_19906);
or UO_230 (O_230,N_19982,N_19984);
nand UO_231 (O_231,N_19842,N_19876);
nand UO_232 (O_232,N_19996,N_19898);
nor UO_233 (O_233,N_19922,N_19872);
or UO_234 (O_234,N_19927,N_19992);
xnor UO_235 (O_235,N_19854,N_19982);
xnor UO_236 (O_236,N_19936,N_19940);
nor UO_237 (O_237,N_19971,N_19892);
nor UO_238 (O_238,N_19963,N_19937);
nor UO_239 (O_239,N_19953,N_19950);
nor UO_240 (O_240,N_19944,N_19946);
nand UO_241 (O_241,N_19930,N_19841);
nand UO_242 (O_242,N_19934,N_19846);
or UO_243 (O_243,N_19885,N_19994);
or UO_244 (O_244,N_19991,N_19924);
and UO_245 (O_245,N_19933,N_19867);
nand UO_246 (O_246,N_19900,N_19856);
nand UO_247 (O_247,N_19932,N_19928);
xor UO_248 (O_248,N_19933,N_19865);
and UO_249 (O_249,N_19978,N_19857);
nor UO_250 (O_250,N_19977,N_19935);
or UO_251 (O_251,N_19845,N_19941);
or UO_252 (O_252,N_19983,N_19864);
xor UO_253 (O_253,N_19929,N_19894);
or UO_254 (O_254,N_19917,N_19896);
xor UO_255 (O_255,N_19998,N_19990);
and UO_256 (O_256,N_19853,N_19854);
nand UO_257 (O_257,N_19970,N_19919);
xnor UO_258 (O_258,N_19956,N_19899);
xnor UO_259 (O_259,N_19947,N_19984);
xor UO_260 (O_260,N_19840,N_19994);
or UO_261 (O_261,N_19847,N_19894);
xnor UO_262 (O_262,N_19987,N_19962);
nand UO_263 (O_263,N_19991,N_19873);
nand UO_264 (O_264,N_19934,N_19917);
xnor UO_265 (O_265,N_19989,N_19847);
xor UO_266 (O_266,N_19923,N_19970);
nand UO_267 (O_267,N_19846,N_19861);
nand UO_268 (O_268,N_19979,N_19970);
or UO_269 (O_269,N_19935,N_19951);
xor UO_270 (O_270,N_19996,N_19946);
xnor UO_271 (O_271,N_19856,N_19942);
xor UO_272 (O_272,N_19978,N_19926);
or UO_273 (O_273,N_19891,N_19941);
xor UO_274 (O_274,N_19984,N_19854);
nor UO_275 (O_275,N_19924,N_19963);
xnor UO_276 (O_276,N_19894,N_19842);
and UO_277 (O_277,N_19849,N_19911);
nor UO_278 (O_278,N_19998,N_19862);
nand UO_279 (O_279,N_19997,N_19864);
and UO_280 (O_280,N_19852,N_19951);
or UO_281 (O_281,N_19918,N_19948);
or UO_282 (O_282,N_19883,N_19989);
xor UO_283 (O_283,N_19872,N_19997);
nand UO_284 (O_284,N_19978,N_19936);
xor UO_285 (O_285,N_19943,N_19954);
or UO_286 (O_286,N_19901,N_19895);
nor UO_287 (O_287,N_19950,N_19924);
and UO_288 (O_288,N_19869,N_19991);
xor UO_289 (O_289,N_19896,N_19899);
nand UO_290 (O_290,N_19941,N_19893);
and UO_291 (O_291,N_19879,N_19994);
nand UO_292 (O_292,N_19979,N_19887);
nor UO_293 (O_293,N_19948,N_19934);
nand UO_294 (O_294,N_19998,N_19926);
nor UO_295 (O_295,N_19942,N_19865);
or UO_296 (O_296,N_19884,N_19938);
xor UO_297 (O_297,N_19937,N_19966);
or UO_298 (O_298,N_19946,N_19887);
or UO_299 (O_299,N_19974,N_19893);
xor UO_300 (O_300,N_19899,N_19856);
xor UO_301 (O_301,N_19959,N_19934);
or UO_302 (O_302,N_19953,N_19932);
nand UO_303 (O_303,N_19983,N_19918);
xnor UO_304 (O_304,N_19905,N_19943);
and UO_305 (O_305,N_19992,N_19984);
and UO_306 (O_306,N_19893,N_19847);
nand UO_307 (O_307,N_19914,N_19953);
or UO_308 (O_308,N_19840,N_19859);
nand UO_309 (O_309,N_19865,N_19893);
nor UO_310 (O_310,N_19845,N_19890);
nand UO_311 (O_311,N_19856,N_19928);
or UO_312 (O_312,N_19852,N_19957);
xnor UO_313 (O_313,N_19988,N_19875);
or UO_314 (O_314,N_19958,N_19924);
nor UO_315 (O_315,N_19959,N_19971);
or UO_316 (O_316,N_19995,N_19902);
and UO_317 (O_317,N_19929,N_19874);
xor UO_318 (O_318,N_19978,N_19973);
and UO_319 (O_319,N_19930,N_19950);
nor UO_320 (O_320,N_19860,N_19978);
or UO_321 (O_321,N_19898,N_19881);
and UO_322 (O_322,N_19848,N_19943);
or UO_323 (O_323,N_19948,N_19879);
or UO_324 (O_324,N_19939,N_19950);
nor UO_325 (O_325,N_19986,N_19922);
xnor UO_326 (O_326,N_19983,N_19948);
nor UO_327 (O_327,N_19993,N_19939);
or UO_328 (O_328,N_19910,N_19915);
and UO_329 (O_329,N_19846,N_19997);
xnor UO_330 (O_330,N_19872,N_19908);
xnor UO_331 (O_331,N_19957,N_19915);
or UO_332 (O_332,N_19857,N_19847);
nand UO_333 (O_333,N_19848,N_19982);
or UO_334 (O_334,N_19878,N_19845);
xnor UO_335 (O_335,N_19847,N_19938);
xor UO_336 (O_336,N_19965,N_19913);
xnor UO_337 (O_337,N_19844,N_19912);
nor UO_338 (O_338,N_19855,N_19992);
or UO_339 (O_339,N_19984,N_19926);
or UO_340 (O_340,N_19986,N_19902);
xnor UO_341 (O_341,N_19996,N_19849);
and UO_342 (O_342,N_19957,N_19904);
nand UO_343 (O_343,N_19948,N_19906);
xor UO_344 (O_344,N_19882,N_19976);
nor UO_345 (O_345,N_19852,N_19953);
nand UO_346 (O_346,N_19928,N_19987);
nor UO_347 (O_347,N_19861,N_19845);
nor UO_348 (O_348,N_19921,N_19942);
or UO_349 (O_349,N_19878,N_19840);
xor UO_350 (O_350,N_19987,N_19906);
nand UO_351 (O_351,N_19950,N_19887);
and UO_352 (O_352,N_19904,N_19864);
xnor UO_353 (O_353,N_19965,N_19993);
nor UO_354 (O_354,N_19901,N_19979);
xor UO_355 (O_355,N_19952,N_19976);
nor UO_356 (O_356,N_19912,N_19974);
nor UO_357 (O_357,N_19979,N_19914);
nand UO_358 (O_358,N_19993,N_19902);
and UO_359 (O_359,N_19957,N_19865);
xor UO_360 (O_360,N_19901,N_19953);
nand UO_361 (O_361,N_19848,N_19882);
or UO_362 (O_362,N_19889,N_19934);
and UO_363 (O_363,N_19894,N_19964);
nor UO_364 (O_364,N_19882,N_19867);
nand UO_365 (O_365,N_19926,N_19844);
or UO_366 (O_366,N_19860,N_19937);
nand UO_367 (O_367,N_19945,N_19927);
nor UO_368 (O_368,N_19851,N_19929);
xor UO_369 (O_369,N_19885,N_19891);
or UO_370 (O_370,N_19971,N_19905);
nand UO_371 (O_371,N_19895,N_19848);
xnor UO_372 (O_372,N_19905,N_19927);
and UO_373 (O_373,N_19942,N_19924);
nor UO_374 (O_374,N_19884,N_19973);
nand UO_375 (O_375,N_19840,N_19908);
and UO_376 (O_376,N_19855,N_19914);
and UO_377 (O_377,N_19883,N_19937);
xnor UO_378 (O_378,N_19854,N_19901);
xor UO_379 (O_379,N_19905,N_19871);
nor UO_380 (O_380,N_19928,N_19891);
nor UO_381 (O_381,N_19968,N_19933);
xor UO_382 (O_382,N_19936,N_19882);
nor UO_383 (O_383,N_19978,N_19844);
or UO_384 (O_384,N_19949,N_19964);
xnor UO_385 (O_385,N_19864,N_19841);
nor UO_386 (O_386,N_19844,N_19958);
xor UO_387 (O_387,N_19931,N_19975);
nor UO_388 (O_388,N_19994,N_19986);
nand UO_389 (O_389,N_19923,N_19898);
and UO_390 (O_390,N_19897,N_19867);
nand UO_391 (O_391,N_19890,N_19965);
nand UO_392 (O_392,N_19871,N_19951);
xor UO_393 (O_393,N_19873,N_19984);
nor UO_394 (O_394,N_19859,N_19988);
nand UO_395 (O_395,N_19902,N_19922);
and UO_396 (O_396,N_19935,N_19958);
xnor UO_397 (O_397,N_19964,N_19893);
nor UO_398 (O_398,N_19967,N_19881);
nor UO_399 (O_399,N_19937,N_19892);
nand UO_400 (O_400,N_19898,N_19897);
or UO_401 (O_401,N_19993,N_19915);
nand UO_402 (O_402,N_19963,N_19982);
and UO_403 (O_403,N_19974,N_19884);
or UO_404 (O_404,N_19895,N_19954);
nand UO_405 (O_405,N_19939,N_19853);
or UO_406 (O_406,N_19964,N_19854);
nor UO_407 (O_407,N_19942,N_19903);
nor UO_408 (O_408,N_19992,N_19949);
xnor UO_409 (O_409,N_19874,N_19888);
and UO_410 (O_410,N_19938,N_19924);
or UO_411 (O_411,N_19873,N_19971);
and UO_412 (O_412,N_19893,N_19988);
or UO_413 (O_413,N_19873,N_19871);
and UO_414 (O_414,N_19873,N_19932);
nor UO_415 (O_415,N_19971,N_19988);
and UO_416 (O_416,N_19864,N_19946);
or UO_417 (O_417,N_19955,N_19847);
and UO_418 (O_418,N_19986,N_19843);
or UO_419 (O_419,N_19950,N_19865);
or UO_420 (O_420,N_19988,N_19958);
nand UO_421 (O_421,N_19940,N_19927);
xnor UO_422 (O_422,N_19896,N_19987);
or UO_423 (O_423,N_19911,N_19973);
xor UO_424 (O_424,N_19950,N_19946);
xnor UO_425 (O_425,N_19910,N_19905);
or UO_426 (O_426,N_19932,N_19965);
xor UO_427 (O_427,N_19854,N_19886);
xnor UO_428 (O_428,N_19958,N_19976);
xnor UO_429 (O_429,N_19935,N_19909);
xor UO_430 (O_430,N_19959,N_19925);
nor UO_431 (O_431,N_19928,N_19898);
nor UO_432 (O_432,N_19892,N_19918);
or UO_433 (O_433,N_19897,N_19916);
or UO_434 (O_434,N_19894,N_19900);
xnor UO_435 (O_435,N_19942,N_19877);
or UO_436 (O_436,N_19849,N_19920);
xor UO_437 (O_437,N_19841,N_19999);
nand UO_438 (O_438,N_19979,N_19937);
and UO_439 (O_439,N_19885,N_19974);
xor UO_440 (O_440,N_19875,N_19976);
xor UO_441 (O_441,N_19994,N_19898);
and UO_442 (O_442,N_19845,N_19971);
and UO_443 (O_443,N_19924,N_19946);
xnor UO_444 (O_444,N_19885,N_19938);
xnor UO_445 (O_445,N_19889,N_19936);
nor UO_446 (O_446,N_19921,N_19972);
or UO_447 (O_447,N_19843,N_19883);
nor UO_448 (O_448,N_19894,N_19988);
and UO_449 (O_449,N_19919,N_19841);
and UO_450 (O_450,N_19896,N_19873);
or UO_451 (O_451,N_19947,N_19934);
xor UO_452 (O_452,N_19893,N_19975);
nor UO_453 (O_453,N_19938,N_19840);
nor UO_454 (O_454,N_19879,N_19844);
nand UO_455 (O_455,N_19857,N_19988);
or UO_456 (O_456,N_19978,N_19991);
and UO_457 (O_457,N_19977,N_19990);
xnor UO_458 (O_458,N_19916,N_19911);
nor UO_459 (O_459,N_19944,N_19888);
nand UO_460 (O_460,N_19850,N_19924);
nand UO_461 (O_461,N_19847,N_19956);
xnor UO_462 (O_462,N_19840,N_19934);
xnor UO_463 (O_463,N_19949,N_19895);
xor UO_464 (O_464,N_19864,N_19897);
nand UO_465 (O_465,N_19984,N_19907);
and UO_466 (O_466,N_19843,N_19860);
xnor UO_467 (O_467,N_19961,N_19903);
nor UO_468 (O_468,N_19847,N_19904);
nor UO_469 (O_469,N_19966,N_19863);
nor UO_470 (O_470,N_19843,N_19958);
nand UO_471 (O_471,N_19878,N_19997);
nor UO_472 (O_472,N_19974,N_19956);
or UO_473 (O_473,N_19852,N_19935);
and UO_474 (O_474,N_19892,N_19967);
xnor UO_475 (O_475,N_19903,N_19907);
nor UO_476 (O_476,N_19886,N_19933);
and UO_477 (O_477,N_19906,N_19868);
xor UO_478 (O_478,N_19845,N_19937);
and UO_479 (O_479,N_19966,N_19889);
or UO_480 (O_480,N_19968,N_19875);
xnor UO_481 (O_481,N_19916,N_19937);
xnor UO_482 (O_482,N_19920,N_19863);
or UO_483 (O_483,N_19903,N_19926);
nor UO_484 (O_484,N_19924,N_19906);
or UO_485 (O_485,N_19981,N_19880);
xor UO_486 (O_486,N_19904,N_19868);
nor UO_487 (O_487,N_19934,N_19926);
xnor UO_488 (O_488,N_19902,N_19996);
or UO_489 (O_489,N_19969,N_19916);
or UO_490 (O_490,N_19984,N_19985);
xor UO_491 (O_491,N_19874,N_19992);
xor UO_492 (O_492,N_19992,N_19991);
and UO_493 (O_493,N_19883,N_19896);
nand UO_494 (O_494,N_19853,N_19931);
nand UO_495 (O_495,N_19998,N_19871);
or UO_496 (O_496,N_19878,N_19964);
xnor UO_497 (O_497,N_19870,N_19962);
nor UO_498 (O_498,N_19882,N_19851);
xnor UO_499 (O_499,N_19889,N_19964);
nor UO_500 (O_500,N_19944,N_19870);
or UO_501 (O_501,N_19921,N_19893);
and UO_502 (O_502,N_19943,N_19949);
nand UO_503 (O_503,N_19921,N_19998);
xor UO_504 (O_504,N_19910,N_19997);
or UO_505 (O_505,N_19857,N_19933);
nand UO_506 (O_506,N_19995,N_19898);
xor UO_507 (O_507,N_19944,N_19993);
and UO_508 (O_508,N_19887,N_19914);
or UO_509 (O_509,N_19953,N_19903);
nor UO_510 (O_510,N_19936,N_19864);
xor UO_511 (O_511,N_19962,N_19991);
or UO_512 (O_512,N_19897,N_19990);
nor UO_513 (O_513,N_19980,N_19950);
nor UO_514 (O_514,N_19847,N_19931);
and UO_515 (O_515,N_19934,N_19965);
nor UO_516 (O_516,N_19960,N_19961);
xnor UO_517 (O_517,N_19854,N_19932);
xnor UO_518 (O_518,N_19997,N_19858);
nand UO_519 (O_519,N_19901,N_19863);
nand UO_520 (O_520,N_19947,N_19941);
or UO_521 (O_521,N_19848,N_19972);
and UO_522 (O_522,N_19898,N_19992);
xnor UO_523 (O_523,N_19948,N_19920);
and UO_524 (O_524,N_19944,N_19864);
nor UO_525 (O_525,N_19896,N_19966);
nor UO_526 (O_526,N_19996,N_19913);
and UO_527 (O_527,N_19957,N_19926);
or UO_528 (O_528,N_19905,N_19897);
nand UO_529 (O_529,N_19971,N_19860);
xnor UO_530 (O_530,N_19860,N_19921);
or UO_531 (O_531,N_19937,N_19889);
or UO_532 (O_532,N_19988,N_19909);
or UO_533 (O_533,N_19848,N_19997);
nor UO_534 (O_534,N_19875,N_19990);
and UO_535 (O_535,N_19929,N_19932);
nand UO_536 (O_536,N_19875,N_19878);
or UO_537 (O_537,N_19991,N_19860);
nand UO_538 (O_538,N_19912,N_19887);
or UO_539 (O_539,N_19931,N_19878);
and UO_540 (O_540,N_19924,N_19982);
nand UO_541 (O_541,N_19885,N_19964);
or UO_542 (O_542,N_19954,N_19945);
or UO_543 (O_543,N_19935,N_19934);
or UO_544 (O_544,N_19966,N_19929);
nor UO_545 (O_545,N_19845,N_19934);
xor UO_546 (O_546,N_19928,N_19915);
or UO_547 (O_547,N_19997,N_19962);
nand UO_548 (O_548,N_19840,N_19978);
and UO_549 (O_549,N_19840,N_19861);
and UO_550 (O_550,N_19900,N_19851);
nor UO_551 (O_551,N_19981,N_19857);
and UO_552 (O_552,N_19939,N_19859);
or UO_553 (O_553,N_19947,N_19977);
and UO_554 (O_554,N_19860,N_19919);
or UO_555 (O_555,N_19881,N_19903);
and UO_556 (O_556,N_19950,N_19855);
nor UO_557 (O_557,N_19879,N_19989);
xnor UO_558 (O_558,N_19938,N_19976);
and UO_559 (O_559,N_19908,N_19912);
or UO_560 (O_560,N_19964,N_19877);
and UO_561 (O_561,N_19916,N_19869);
and UO_562 (O_562,N_19952,N_19934);
xnor UO_563 (O_563,N_19980,N_19973);
or UO_564 (O_564,N_19866,N_19956);
and UO_565 (O_565,N_19872,N_19920);
xor UO_566 (O_566,N_19868,N_19897);
or UO_567 (O_567,N_19926,N_19875);
nor UO_568 (O_568,N_19950,N_19843);
and UO_569 (O_569,N_19911,N_19846);
nand UO_570 (O_570,N_19918,N_19910);
and UO_571 (O_571,N_19880,N_19936);
nand UO_572 (O_572,N_19941,N_19914);
and UO_573 (O_573,N_19897,N_19872);
or UO_574 (O_574,N_19909,N_19932);
nor UO_575 (O_575,N_19953,N_19862);
nor UO_576 (O_576,N_19906,N_19843);
nor UO_577 (O_577,N_19984,N_19978);
nor UO_578 (O_578,N_19974,N_19920);
nand UO_579 (O_579,N_19912,N_19978);
nand UO_580 (O_580,N_19917,N_19994);
xnor UO_581 (O_581,N_19935,N_19940);
nand UO_582 (O_582,N_19874,N_19919);
xor UO_583 (O_583,N_19906,N_19932);
and UO_584 (O_584,N_19851,N_19959);
xor UO_585 (O_585,N_19857,N_19940);
and UO_586 (O_586,N_19933,N_19891);
xnor UO_587 (O_587,N_19857,N_19944);
and UO_588 (O_588,N_19844,N_19932);
xnor UO_589 (O_589,N_19843,N_19866);
nand UO_590 (O_590,N_19974,N_19963);
xor UO_591 (O_591,N_19915,N_19983);
nor UO_592 (O_592,N_19954,N_19865);
and UO_593 (O_593,N_19968,N_19955);
and UO_594 (O_594,N_19877,N_19914);
xnor UO_595 (O_595,N_19928,N_19871);
nand UO_596 (O_596,N_19854,N_19961);
or UO_597 (O_597,N_19949,N_19952);
or UO_598 (O_598,N_19953,N_19990);
nand UO_599 (O_599,N_19994,N_19871);
and UO_600 (O_600,N_19992,N_19961);
and UO_601 (O_601,N_19966,N_19898);
or UO_602 (O_602,N_19971,N_19841);
nand UO_603 (O_603,N_19990,N_19929);
or UO_604 (O_604,N_19854,N_19874);
and UO_605 (O_605,N_19889,N_19982);
or UO_606 (O_606,N_19896,N_19916);
nand UO_607 (O_607,N_19869,N_19936);
xnor UO_608 (O_608,N_19923,N_19937);
nand UO_609 (O_609,N_19900,N_19857);
nand UO_610 (O_610,N_19925,N_19996);
and UO_611 (O_611,N_19845,N_19997);
nor UO_612 (O_612,N_19929,N_19970);
nor UO_613 (O_613,N_19888,N_19898);
xor UO_614 (O_614,N_19991,N_19999);
or UO_615 (O_615,N_19930,N_19924);
or UO_616 (O_616,N_19987,N_19881);
nor UO_617 (O_617,N_19909,N_19985);
nor UO_618 (O_618,N_19939,N_19979);
nor UO_619 (O_619,N_19912,N_19895);
xnor UO_620 (O_620,N_19858,N_19968);
xnor UO_621 (O_621,N_19987,N_19934);
xor UO_622 (O_622,N_19936,N_19992);
and UO_623 (O_623,N_19855,N_19995);
xnor UO_624 (O_624,N_19994,N_19958);
or UO_625 (O_625,N_19994,N_19865);
nor UO_626 (O_626,N_19853,N_19952);
and UO_627 (O_627,N_19841,N_19911);
nand UO_628 (O_628,N_19937,N_19994);
or UO_629 (O_629,N_19873,N_19872);
or UO_630 (O_630,N_19846,N_19979);
or UO_631 (O_631,N_19972,N_19868);
or UO_632 (O_632,N_19907,N_19941);
nand UO_633 (O_633,N_19961,N_19873);
and UO_634 (O_634,N_19936,N_19853);
or UO_635 (O_635,N_19852,N_19938);
xnor UO_636 (O_636,N_19978,N_19875);
and UO_637 (O_637,N_19972,N_19882);
nand UO_638 (O_638,N_19972,N_19944);
xor UO_639 (O_639,N_19988,N_19933);
or UO_640 (O_640,N_19933,N_19950);
and UO_641 (O_641,N_19841,N_19866);
nand UO_642 (O_642,N_19914,N_19901);
nor UO_643 (O_643,N_19916,N_19873);
and UO_644 (O_644,N_19989,N_19909);
xnor UO_645 (O_645,N_19990,N_19886);
nand UO_646 (O_646,N_19923,N_19933);
nor UO_647 (O_647,N_19841,N_19915);
or UO_648 (O_648,N_19879,N_19866);
or UO_649 (O_649,N_19936,N_19965);
and UO_650 (O_650,N_19880,N_19997);
nor UO_651 (O_651,N_19961,N_19968);
xnor UO_652 (O_652,N_19931,N_19901);
nand UO_653 (O_653,N_19869,N_19855);
nor UO_654 (O_654,N_19964,N_19991);
nand UO_655 (O_655,N_19959,N_19909);
nor UO_656 (O_656,N_19993,N_19847);
or UO_657 (O_657,N_19940,N_19965);
or UO_658 (O_658,N_19926,N_19996);
nor UO_659 (O_659,N_19862,N_19971);
or UO_660 (O_660,N_19918,N_19914);
xor UO_661 (O_661,N_19891,N_19926);
nand UO_662 (O_662,N_19892,N_19924);
or UO_663 (O_663,N_19986,N_19969);
nand UO_664 (O_664,N_19850,N_19967);
or UO_665 (O_665,N_19943,N_19879);
and UO_666 (O_666,N_19895,N_19976);
and UO_667 (O_667,N_19898,N_19926);
nand UO_668 (O_668,N_19860,N_19910);
or UO_669 (O_669,N_19896,N_19938);
and UO_670 (O_670,N_19988,N_19986);
nor UO_671 (O_671,N_19847,N_19949);
nor UO_672 (O_672,N_19892,N_19983);
xnor UO_673 (O_673,N_19956,N_19960);
and UO_674 (O_674,N_19979,N_19923);
or UO_675 (O_675,N_19989,N_19892);
nand UO_676 (O_676,N_19999,N_19858);
or UO_677 (O_677,N_19995,N_19954);
nand UO_678 (O_678,N_19880,N_19842);
or UO_679 (O_679,N_19953,N_19863);
nor UO_680 (O_680,N_19869,N_19982);
and UO_681 (O_681,N_19896,N_19852);
nor UO_682 (O_682,N_19868,N_19852);
xor UO_683 (O_683,N_19876,N_19917);
and UO_684 (O_684,N_19978,N_19910);
nor UO_685 (O_685,N_19848,N_19915);
nand UO_686 (O_686,N_19979,N_19981);
xnor UO_687 (O_687,N_19937,N_19906);
and UO_688 (O_688,N_19904,N_19886);
xor UO_689 (O_689,N_19939,N_19903);
or UO_690 (O_690,N_19883,N_19975);
nor UO_691 (O_691,N_19938,N_19981);
or UO_692 (O_692,N_19946,N_19863);
and UO_693 (O_693,N_19844,N_19921);
or UO_694 (O_694,N_19847,N_19846);
xnor UO_695 (O_695,N_19965,N_19967);
and UO_696 (O_696,N_19898,N_19905);
xor UO_697 (O_697,N_19852,N_19912);
nor UO_698 (O_698,N_19987,N_19936);
nand UO_699 (O_699,N_19970,N_19861);
and UO_700 (O_700,N_19940,N_19853);
xor UO_701 (O_701,N_19869,N_19915);
xnor UO_702 (O_702,N_19849,N_19986);
nand UO_703 (O_703,N_19904,N_19917);
nor UO_704 (O_704,N_19982,N_19942);
xnor UO_705 (O_705,N_19903,N_19944);
xnor UO_706 (O_706,N_19848,N_19971);
nor UO_707 (O_707,N_19907,N_19862);
nand UO_708 (O_708,N_19959,N_19901);
or UO_709 (O_709,N_19946,N_19843);
nor UO_710 (O_710,N_19859,N_19866);
nand UO_711 (O_711,N_19860,N_19862);
xor UO_712 (O_712,N_19904,N_19841);
xnor UO_713 (O_713,N_19904,N_19855);
and UO_714 (O_714,N_19978,N_19982);
and UO_715 (O_715,N_19980,N_19848);
nor UO_716 (O_716,N_19894,N_19882);
xor UO_717 (O_717,N_19958,N_19913);
or UO_718 (O_718,N_19859,N_19919);
nand UO_719 (O_719,N_19972,N_19915);
xor UO_720 (O_720,N_19861,N_19955);
nor UO_721 (O_721,N_19858,N_19993);
xnor UO_722 (O_722,N_19905,N_19913);
nor UO_723 (O_723,N_19933,N_19986);
nand UO_724 (O_724,N_19967,N_19885);
nor UO_725 (O_725,N_19923,N_19934);
or UO_726 (O_726,N_19913,N_19981);
xnor UO_727 (O_727,N_19892,N_19861);
nand UO_728 (O_728,N_19866,N_19910);
or UO_729 (O_729,N_19904,N_19908);
or UO_730 (O_730,N_19891,N_19929);
or UO_731 (O_731,N_19963,N_19927);
xor UO_732 (O_732,N_19924,N_19857);
or UO_733 (O_733,N_19845,N_19915);
xor UO_734 (O_734,N_19999,N_19910);
nand UO_735 (O_735,N_19938,N_19977);
xnor UO_736 (O_736,N_19970,N_19873);
or UO_737 (O_737,N_19854,N_19976);
nor UO_738 (O_738,N_19872,N_19887);
and UO_739 (O_739,N_19901,N_19938);
nor UO_740 (O_740,N_19855,N_19899);
or UO_741 (O_741,N_19923,N_19931);
and UO_742 (O_742,N_19855,N_19971);
nor UO_743 (O_743,N_19881,N_19840);
nor UO_744 (O_744,N_19979,N_19930);
nor UO_745 (O_745,N_19873,N_19879);
nand UO_746 (O_746,N_19871,N_19860);
xor UO_747 (O_747,N_19966,N_19994);
or UO_748 (O_748,N_19956,N_19995);
xor UO_749 (O_749,N_19901,N_19899);
nor UO_750 (O_750,N_19904,N_19903);
and UO_751 (O_751,N_19928,N_19902);
nor UO_752 (O_752,N_19916,N_19948);
or UO_753 (O_753,N_19878,N_19959);
and UO_754 (O_754,N_19929,N_19921);
and UO_755 (O_755,N_19937,N_19982);
nand UO_756 (O_756,N_19918,N_19955);
and UO_757 (O_757,N_19978,N_19886);
and UO_758 (O_758,N_19971,N_19890);
and UO_759 (O_759,N_19867,N_19952);
or UO_760 (O_760,N_19941,N_19896);
nand UO_761 (O_761,N_19878,N_19980);
nor UO_762 (O_762,N_19868,N_19861);
or UO_763 (O_763,N_19900,N_19989);
xor UO_764 (O_764,N_19930,N_19986);
and UO_765 (O_765,N_19903,N_19958);
or UO_766 (O_766,N_19870,N_19876);
xnor UO_767 (O_767,N_19977,N_19897);
and UO_768 (O_768,N_19902,N_19953);
or UO_769 (O_769,N_19924,N_19866);
nand UO_770 (O_770,N_19878,N_19892);
or UO_771 (O_771,N_19920,N_19955);
or UO_772 (O_772,N_19964,N_19904);
or UO_773 (O_773,N_19991,N_19939);
and UO_774 (O_774,N_19933,N_19900);
nor UO_775 (O_775,N_19858,N_19948);
xnor UO_776 (O_776,N_19934,N_19937);
and UO_777 (O_777,N_19893,N_19908);
or UO_778 (O_778,N_19969,N_19931);
nand UO_779 (O_779,N_19952,N_19873);
and UO_780 (O_780,N_19996,N_19968);
or UO_781 (O_781,N_19953,N_19872);
and UO_782 (O_782,N_19911,N_19985);
nand UO_783 (O_783,N_19907,N_19851);
nor UO_784 (O_784,N_19862,N_19973);
nand UO_785 (O_785,N_19920,N_19967);
xnor UO_786 (O_786,N_19962,N_19956);
xor UO_787 (O_787,N_19896,N_19876);
or UO_788 (O_788,N_19973,N_19982);
or UO_789 (O_789,N_19971,N_19923);
and UO_790 (O_790,N_19841,N_19863);
nand UO_791 (O_791,N_19907,N_19952);
and UO_792 (O_792,N_19854,N_19907);
nor UO_793 (O_793,N_19936,N_19907);
nor UO_794 (O_794,N_19877,N_19937);
xor UO_795 (O_795,N_19948,N_19952);
nand UO_796 (O_796,N_19894,N_19990);
xnor UO_797 (O_797,N_19985,N_19960);
nand UO_798 (O_798,N_19855,N_19976);
xor UO_799 (O_799,N_19939,N_19882);
nor UO_800 (O_800,N_19963,N_19966);
or UO_801 (O_801,N_19871,N_19926);
and UO_802 (O_802,N_19941,N_19869);
and UO_803 (O_803,N_19859,N_19983);
or UO_804 (O_804,N_19900,N_19974);
or UO_805 (O_805,N_19989,N_19846);
or UO_806 (O_806,N_19883,N_19887);
nand UO_807 (O_807,N_19866,N_19874);
or UO_808 (O_808,N_19916,N_19901);
or UO_809 (O_809,N_19848,N_19985);
nand UO_810 (O_810,N_19863,N_19941);
nand UO_811 (O_811,N_19897,N_19846);
and UO_812 (O_812,N_19932,N_19994);
nand UO_813 (O_813,N_19902,N_19903);
or UO_814 (O_814,N_19840,N_19986);
or UO_815 (O_815,N_19862,N_19868);
nand UO_816 (O_816,N_19974,N_19865);
xnor UO_817 (O_817,N_19979,N_19871);
nor UO_818 (O_818,N_19879,N_19865);
nand UO_819 (O_819,N_19971,N_19869);
and UO_820 (O_820,N_19851,N_19870);
nor UO_821 (O_821,N_19983,N_19935);
nand UO_822 (O_822,N_19917,N_19979);
or UO_823 (O_823,N_19877,N_19956);
or UO_824 (O_824,N_19905,N_19864);
or UO_825 (O_825,N_19930,N_19881);
and UO_826 (O_826,N_19920,N_19856);
nand UO_827 (O_827,N_19952,N_19871);
or UO_828 (O_828,N_19906,N_19875);
nor UO_829 (O_829,N_19945,N_19913);
or UO_830 (O_830,N_19878,N_19999);
nand UO_831 (O_831,N_19949,N_19888);
nand UO_832 (O_832,N_19963,N_19891);
or UO_833 (O_833,N_19842,N_19983);
and UO_834 (O_834,N_19994,N_19926);
and UO_835 (O_835,N_19872,N_19939);
nor UO_836 (O_836,N_19876,N_19851);
or UO_837 (O_837,N_19910,N_19872);
xnor UO_838 (O_838,N_19852,N_19981);
xnor UO_839 (O_839,N_19966,N_19916);
nand UO_840 (O_840,N_19940,N_19848);
nor UO_841 (O_841,N_19996,N_19933);
nor UO_842 (O_842,N_19978,N_19885);
nand UO_843 (O_843,N_19905,N_19872);
and UO_844 (O_844,N_19894,N_19867);
nand UO_845 (O_845,N_19909,N_19900);
nor UO_846 (O_846,N_19994,N_19891);
nand UO_847 (O_847,N_19893,N_19986);
or UO_848 (O_848,N_19970,N_19961);
nor UO_849 (O_849,N_19923,N_19845);
and UO_850 (O_850,N_19994,N_19856);
or UO_851 (O_851,N_19939,N_19905);
and UO_852 (O_852,N_19965,N_19949);
and UO_853 (O_853,N_19998,N_19914);
and UO_854 (O_854,N_19970,N_19854);
and UO_855 (O_855,N_19943,N_19986);
nand UO_856 (O_856,N_19953,N_19894);
nor UO_857 (O_857,N_19901,N_19902);
or UO_858 (O_858,N_19891,N_19951);
xnor UO_859 (O_859,N_19947,N_19901);
or UO_860 (O_860,N_19936,N_19997);
nor UO_861 (O_861,N_19922,N_19857);
nand UO_862 (O_862,N_19921,N_19951);
nand UO_863 (O_863,N_19884,N_19923);
or UO_864 (O_864,N_19977,N_19980);
nand UO_865 (O_865,N_19959,N_19928);
nor UO_866 (O_866,N_19964,N_19873);
xor UO_867 (O_867,N_19840,N_19850);
xor UO_868 (O_868,N_19888,N_19992);
nand UO_869 (O_869,N_19852,N_19857);
nand UO_870 (O_870,N_19984,N_19870);
xnor UO_871 (O_871,N_19935,N_19880);
or UO_872 (O_872,N_19882,N_19914);
or UO_873 (O_873,N_19895,N_19887);
nand UO_874 (O_874,N_19862,N_19952);
and UO_875 (O_875,N_19857,N_19956);
and UO_876 (O_876,N_19986,N_19955);
nand UO_877 (O_877,N_19915,N_19867);
xor UO_878 (O_878,N_19891,N_19910);
nor UO_879 (O_879,N_19866,N_19855);
nor UO_880 (O_880,N_19863,N_19977);
or UO_881 (O_881,N_19905,N_19964);
nand UO_882 (O_882,N_19868,N_19887);
xor UO_883 (O_883,N_19981,N_19976);
nor UO_884 (O_884,N_19846,N_19943);
or UO_885 (O_885,N_19951,N_19976);
and UO_886 (O_886,N_19957,N_19860);
xor UO_887 (O_887,N_19948,N_19861);
and UO_888 (O_888,N_19918,N_19874);
xnor UO_889 (O_889,N_19935,N_19872);
nand UO_890 (O_890,N_19861,N_19849);
and UO_891 (O_891,N_19972,N_19855);
and UO_892 (O_892,N_19931,N_19913);
nand UO_893 (O_893,N_19969,N_19856);
and UO_894 (O_894,N_19858,N_19988);
and UO_895 (O_895,N_19891,N_19842);
nor UO_896 (O_896,N_19970,N_19985);
nand UO_897 (O_897,N_19876,N_19901);
nand UO_898 (O_898,N_19851,N_19949);
and UO_899 (O_899,N_19892,N_19841);
nor UO_900 (O_900,N_19909,N_19995);
nand UO_901 (O_901,N_19956,N_19920);
or UO_902 (O_902,N_19969,N_19924);
nand UO_903 (O_903,N_19991,N_19923);
nor UO_904 (O_904,N_19890,N_19898);
or UO_905 (O_905,N_19978,N_19945);
nor UO_906 (O_906,N_19929,N_19947);
nand UO_907 (O_907,N_19860,N_19987);
nor UO_908 (O_908,N_19895,N_19888);
nor UO_909 (O_909,N_19871,N_19936);
nand UO_910 (O_910,N_19995,N_19866);
and UO_911 (O_911,N_19997,N_19892);
and UO_912 (O_912,N_19853,N_19967);
or UO_913 (O_913,N_19859,N_19855);
xor UO_914 (O_914,N_19955,N_19924);
nand UO_915 (O_915,N_19916,N_19883);
nor UO_916 (O_916,N_19977,N_19900);
nand UO_917 (O_917,N_19937,N_19903);
and UO_918 (O_918,N_19994,N_19852);
and UO_919 (O_919,N_19981,N_19876);
nand UO_920 (O_920,N_19940,N_19947);
or UO_921 (O_921,N_19996,N_19870);
nand UO_922 (O_922,N_19993,N_19866);
or UO_923 (O_923,N_19975,N_19973);
nand UO_924 (O_924,N_19887,N_19865);
and UO_925 (O_925,N_19921,N_19902);
or UO_926 (O_926,N_19973,N_19919);
and UO_927 (O_927,N_19914,N_19869);
nand UO_928 (O_928,N_19858,N_19962);
xor UO_929 (O_929,N_19954,N_19890);
nor UO_930 (O_930,N_19974,N_19931);
nand UO_931 (O_931,N_19891,N_19937);
or UO_932 (O_932,N_19900,N_19966);
nand UO_933 (O_933,N_19985,N_19854);
and UO_934 (O_934,N_19889,N_19987);
or UO_935 (O_935,N_19998,N_19895);
xnor UO_936 (O_936,N_19952,N_19979);
xor UO_937 (O_937,N_19976,N_19889);
nand UO_938 (O_938,N_19854,N_19916);
or UO_939 (O_939,N_19978,N_19918);
and UO_940 (O_940,N_19852,N_19889);
nand UO_941 (O_941,N_19878,N_19883);
xor UO_942 (O_942,N_19985,N_19995);
and UO_943 (O_943,N_19972,N_19986);
and UO_944 (O_944,N_19868,N_19937);
and UO_945 (O_945,N_19949,N_19885);
nor UO_946 (O_946,N_19942,N_19874);
nand UO_947 (O_947,N_19950,N_19929);
xnor UO_948 (O_948,N_19947,N_19905);
nor UO_949 (O_949,N_19929,N_19887);
nor UO_950 (O_950,N_19978,N_19879);
nor UO_951 (O_951,N_19950,N_19948);
nor UO_952 (O_952,N_19939,N_19924);
and UO_953 (O_953,N_19882,N_19902);
nand UO_954 (O_954,N_19980,N_19981);
nand UO_955 (O_955,N_19879,N_19969);
or UO_956 (O_956,N_19938,N_19886);
and UO_957 (O_957,N_19975,N_19902);
nor UO_958 (O_958,N_19872,N_19861);
nor UO_959 (O_959,N_19957,N_19952);
or UO_960 (O_960,N_19857,N_19883);
and UO_961 (O_961,N_19923,N_19847);
xnor UO_962 (O_962,N_19894,N_19934);
nor UO_963 (O_963,N_19944,N_19992);
xor UO_964 (O_964,N_19869,N_19984);
or UO_965 (O_965,N_19999,N_19905);
xnor UO_966 (O_966,N_19979,N_19992);
or UO_967 (O_967,N_19933,N_19935);
nand UO_968 (O_968,N_19926,N_19849);
nor UO_969 (O_969,N_19864,N_19932);
nor UO_970 (O_970,N_19946,N_19936);
and UO_971 (O_971,N_19911,N_19850);
or UO_972 (O_972,N_19861,N_19998);
nand UO_973 (O_973,N_19975,N_19997);
or UO_974 (O_974,N_19871,N_19993);
or UO_975 (O_975,N_19990,N_19865);
or UO_976 (O_976,N_19942,N_19885);
and UO_977 (O_977,N_19883,N_19842);
nor UO_978 (O_978,N_19885,N_19892);
nand UO_979 (O_979,N_19908,N_19868);
xor UO_980 (O_980,N_19966,N_19993);
or UO_981 (O_981,N_19892,N_19925);
or UO_982 (O_982,N_19939,N_19909);
nand UO_983 (O_983,N_19989,N_19886);
nor UO_984 (O_984,N_19965,N_19879);
or UO_985 (O_985,N_19934,N_19864);
nor UO_986 (O_986,N_19893,N_19899);
and UO_987 (O_987,N_19939,N_19945);
or UO_988 (O_988,N_19999,N_19930);
and UO_989 (O_989,N_19878,N_19918);
nand UO_990 (O_990,N_19867,N_19977);
nor UO_991 (O_991,N_19970,N_19848);
or UO_992 (O_992,N_19965,N_19866);
xor UO_993 (O_993,N_19957,N_19993);
nor UO_994 (O_994,N_19929,N_19849);
or UO_995 (O_995,N_19858,N_19882);
nand UO_996 (O_996,N_19886,N_19876);
and UO_997 (O_997,N_19856,N_19968);
or UO_998 (O_998,N_19905,N_19873);
and UO_999 (O_999,N_19997,N_19893);
nand UO_1000 (O_1000,N_19891,N_19912);
xnor UO_1001 (O_1001,N_19868,N_19885);
xor UO_1002 (O_1002,N_19893,N_19848);
and UO_1003 (O_1003,N_19870,N_19954);
xnor UO_1004 (O_1004,N_19909,N_19901);
and UO_1005 (O_1005,N_19916,N_19902);
xor UO_1006 (O_1006,N_19996,N_19975);
or UO_1007 (O_1007,N_19931,N_19861);
nand UO_1008 (O_1008,N_19933,N_19909);
and UO_1009 (O_1009,N_19904,N_19974);
or UO_1010 (O_1010,N_19870,N_19855);
nor UO_1011 (O_1011,N_19881,N_19907);
nor UO_1012 (O_1012,N_19950,N_19851);
or UO_1013 (O_1013,N_19875,N_19945);
nor UO_1014 (O_1014,N_19886,N_19961);
or UO_1015 (O_1015,N_19999,N_19854);
or UO_1016 (O_1016,N_19924,N_19880);
and UO_1017 (O_1017,N_19980,N_19976);
nor UO_1018 (O_1018,N_19956,N_19914);
nor UO_1019 (O_1019,N_19922,N_19851);
or UO_1020 (O_1020,N_19946,N_19854);
xor UO_1021 (O_1021,N_19953,N_19846);
and UO_1022 (O_1022,N_19924,N_19913);
and UO_1023 (O_1023,N_19886,N_19986);
nor UO_1024 (O_1024,N_19851,N_19858);
nand UO_1025 (O_1025,N_19921,N_19980);
xor UO_1026 (O_1026,N_19991,N_19870);
and UO_1027 (O_1027,N_19919,N_19959);
nand UO_1028 (O_1028,N_19947,N_19930);
or UO_1029 (O_1029,N_19859,N_19956);
nor UO_1030 (O_1030,N_19978,N_19899);
and UO_1031 (O_1031,N_19889,N_19962);
or UO_1032 (O_1032,N_19874,N_19894);
and UO_1033 (O_1033,N_19853,N_19848);
and UO_1034 (O_1034,N_19877,N_19981);
or UO_1035 (O_1035,N_19892,N_19898);
nand UO_1036 (O_1036,N_19890,N_19961);
or UO_1037 (O_1037,N_19952,N_19861);
nand UO_1038 (O_1038,N_19873,N_19857);
or UO_1039 (O_1039,N_19914,N_19852);
nand UO_1040 (O_1040,N_19999,N_19923);
nand UO_1041 (O_1041,N_19937,N_19962);
xnor UO_1042 (O_1042,N_19905,N_19863);
and UO_1043 (O_1043,N_19879,N_19853);
or UO_1044 (O_1044,N_19945,N_19973);
nand UO_1045 (O_1045,N_19946,N_19884);
and UO_1046 (O_1046,N_19876,N_19844);
and UO_1047 (O_1047,N_19964,N_19891);
nand UO_1048 (O_1048,N_19955,N_19886);
and UO_1049 (O_1049,N_19901,N_19850);
nor UO_1050 (O_1050,N_19902,N_19847);
and UO_1051 (O_1051,N_19995,N_19879);
nor UO_1052 (O_1052,N_19908,N_19919);
nand UO_1053 (O_1053,N_19938,N_19844);
or UO_1054 (O_1054,N_19900,N_19871);
nand UO_1055 (O_1055,N_19971,N_19916);
xnor UO_1056 (O_1056,N_19911,N_19887);
nand UO_1057 (O_1057,N_19895,N_19864);
and UO_1058 (O_1058,N_19998,N_19997);
and UO_1059 (O_1059,N_19841,N_19853);
xor UO_1060 (O_1060,N_19986,N_19940);
nand UO_1061 (O_1061,N_19848,N_19885);
xor UO_1062 (O_1062,N_19884,N_19921);
nor UO_1063 (O_1063,N_19848,N_19899);
nor UO_1064 (O_1064,N_19892,N_19958);
nor UO_1065 (O_1065,N_19844,N_19869);
and UO_1066 (O_1066,N_19886,N_19920);
nand UO_1067 (O_1067,N_19973,N_19940);
and UO_1068 (O_1068,N_19992,N_19934);
nor UO_1069 (O_1069,N_19915,N_19866);
or UO_1070 (O_1070,N_19921,N_19957);
or UO_1071 (O_1071,N_19963,N_19884);
xor UO_1072 (O_1072,N_19967,N_19978);
or UO_1073 (O_1073,N_19872,N_19926);
nand UO_1074 (O_1074,N_19869,N_19878);
nand UO_1075 (O_1075,N_19919,N_19974);
and UO_1076 (O_1076,N_19931,N_19989);
and UO_1077 (O_1077,N_19893,N_19857);
nand UO_1078 (O_1078,N_19881,N_19964);
or UO_1079 (O_1079,N_19961,N_19989);
xor UO_1080 (O_1080,N_19899,N_19936);
and UO_1081 (O_1081,N_19996,N_19949);
and UO_1082 (O_1082,N_19935,N_19861);
nand UO_1083 (O_1083,N_19938,N_19978);
nor UO_1084 (O_1084,N_19973,N_19918);
nand UO_1085 (O_1085,N_19943,N_19977);
xor UO_1086 (O_1086,N_19995,N_19932);
and UO_1087 (O_1087,N_19998,N_19894);
or UO_1088 (O_1088,N_19985,N_19938);
xnor UO_1089 (O_1089,N_19898,N_19919);
nor UO_1090 (O_1090,N_19919,N_19865);
nand UO_1091 (O_1091,N_19888,N_19923);
nor UO_1092 (O_1092,N_19927,N_19895);
or UO_1093 (O_1093,N_19990,N_19942);
nor UO_1094 (O_1094,N_19996,N_19944);
xnor UO_1095 (O_1095,N_19944,N_19882);
xor UO_1096 (O_1096,N_19880,N_19881);
nor UO_1097 (O_1097,N_19844,N_19950);
nand UO_1098 (O_1098,N_19909,N_19991);
nor UO_1099 (O_1099,N_19919,N_19927);
or UO_1100 (O_1100,N_19961,N_19889);
or UO_1101 (O_1101,N_19956,N_19852);
xnor UO_1102 (O_1102,N_19970,N_19943);
xnor UO_1103 (O_1103,N_19995,N_19857);
nor UO_1104 (O_1104,N_19912,N_19938);
and UO_1105 (O_1105,N_19942,N_19879);
nand UO_1106 (O_1106,N_19899,N_19849);
xnor UO_1107 (O_1107,N_19878,N_19936);
xnor UO_1108 (O_1108,N_19908,N_19953);
nor UO_1109 (O_1109,N_19875,N_19887);
xnor UO_1110 (O_1110,N_19954,N_19957);
xor UO_1111 (O_1111,N_19884,N_19976);
nand UO_1112 (O_1112,N_19957,N_19869);
and UO_1113 (O_1113,N_19946,N_19865);
and UO_1114 (O_1114,N_19977,N_19906);
or UO_1115 (O_1115,N_19867,N_19931);
and UO_1116 (O_1116,N_19844,N_19969);
nor UO_1117 (O_1117,N_19957,N_19917);
nand UO_1118 (O_1118,N_19984,N_19877);
nor UO_1119 (O_1119,N_19900,N_19868);
and UO_1120 (O_1120,N_19986,N_19916);
nor UO_1121 (O_1121,N_19909,N_19880);
or UO_1122 (O_1122,N_19880,N_19974);
xor UO_1123 (O_1123,N_19843,N_19938);
nand UO_1124 (O_1124,N_19966,N_19844);
nand UO_1125 (O_1125,N_19999,N_19860);
and UO_1126 (O_1126,N_19906,N_19869);
nand UO_1127 (O_1127,N_19886,N_19878);
nand UO_1128 (O_1128,N_19941,N_19968);
or UO_1129 (O_1129,N_19860,N_19998);
xnor UO_1130 (O_1130,N_19846,N_19976);
nand UO_1131 (O_1131,N_19956,N_19944);
nor UO_1132 (O_1132,N_19955,N_19987);
and UO_1133 (O_1133,N_19854,N_19934);
and UO_1134 (O_1134,N_19922,N_19947);
and UO_1135 (O_1135,N_19966,N_19957);
and UO_1136 (O_1136,N_19951,N_19863);
nand UO_1137 (O_1137,N_19969,N_19966);
or UO_1138 (O_1138,N_19850,N_19979);
nor UO_1139 (O_1139,N_19925,N_19909);
or UO_1140 (O_1140,N_19930,N_19905);
xor UO_1141 (O_1141,N_19865,N_19876);
nand UO_1142 (O_1142,N_19854,N_19879);
nor UO_1143 (O_1143,N_19941,N_19958);
nor UO_1144 (O_1144,N_19896,N_19853);
and UO_1145 (O_1145,N_19928,N_19988);
xor UO_1146 (O_1146,N_19884,N_19957);
and UO_1147 (O_1147,N_19956,N_19957);
and UO_1148 (O_1148,N_19872,N_19912);
nand UO_1149 (O_1149,N_19997,N_19850);
and UO_1150 (O_1150,N_19881,N_19957);
or UO_1151 (O_1151,N_19853,N_19987);
nor UO_1152 (O_1152,N_19844,N_19885);
or UO_1153 (O_1153,N_19908,N_19918);
nand UO_1154 (O_1154,N_19981,N_19999);
nand UO_1155 (O_1155,N_19845,N_19930);
nand UO_1156 (O_1156,N_19842,N_19989);
or UO_1157 (O_1157,N_19858,N_19916);
nand UO_1158 (O_1158,N_19895,N_19938);
xnor UO_1159 (O_1159,N_19992,N_19882);
and UO_1160 (O_1160,N_19999,N_19990);
xor UO_1161 (O_1161,N_19900,N_19928);
nor UO_1162 (O_1162,N_19973,N_19892);
nand UO_1163 (O_1163,N_19962,N_19857);
nor UO_1164 (O_1164,N_19906,N_19981);
and UO_1165 (O_1165,N_19918,N_19866);
and UO_1166 (O_1166,N_19959,N_19871);
and UO_1167 (O_1167,N_19916,N_19866);
xnor UO_1168 (O_1168,N_19951,N_19853);
nand UO_1169 (O_1169,N_19923,N_19897);
nand UO_1170 (O_1170,N_19990,N_19997);
or UO_1171 (O_1171,N_19903,N_19863);
or UO_1172 (O_1172,N_19949,N_19982);
nand UO_1173 (O_1173,N_19897,N_19955);
nand UO_1174 (O_1174,N_19966,N_19936);
xnor UO_1175 (O_1175,N_19966,N_19943);
or UO_1176 (O_1176,N_19842,N_19981);
and UO_1177 (O_1177,N_19968,N_19853);
xnor UO_1178 (O_1178,N_19867,N_19987);
nor UO_1179 (O_1179,N_19917,N_19898);
xor UO_1180 (O_1180,N_19995,N_19842);
nor UO_1181 (O_1181,N_19942,N_19935);
nand UO_1182 (O_1182,N_19917,N_19853);
xnor UO_1183 (O_1183,N_19989,N_19866);
or UO_1184 (O_1184,N_19860,N_19920);
nor UO_1185 (O_1185,N_19950,N_19965);
or UO_1186 (O_1186,N_19886,N_19879);
nor UO_1187 (O_1187,N_19878,N_19933);
nand UO_1188 (O_1188,N_19933,N_19901);
nand UO_1189 (O_1189,N_19927,N_19928);
or UO_1190 (O_1190,N_19891,N_19876);
nor UO_1191 (O_1191,N_19953,N_19934);
or UO_1192 (O_1192,N_19969,N_19984);
nor UO_1193 (O_1193,N_19854,N_19845);
nor UO_1194 (O_1194,N_19925,N_19908);
nand UO_1195 (O_1195,N_19985,N_19977);
and UO_1196 (O_1196,N_19890,N_19847);
nand UO_1197 (O_1197,N_19905,N_19862);
nor UO_1198 (O_1198,N_19875,N_19954);
xor UO_1199 (O_1199,N_19883,N_19935);
or UO_1200 (O_1200,N_19847,N_19980);
or UO_1201 (O_1201,N_19982,N_19927);
and UO_1202 (O_1202,N_19867,N_19988);
nor UO_1203 (O_1203,N_19937,N_19975);
nand UO_1204 (O_1204,N_19914,N_19910);
nand UO_1205 (O_1205,N_19848,N_19939);
nand UO_1206 (O_1206,N_19971,N_19978);
nand UO_1207 (O_1207,N_19972,N_19973);
or UO_1208 (O_1208,N_19873,N_19869);
or UO_1209 (O_1209,N_19981,N_19978);
xnor UO_1210 (O_1210,N_19969,N_19849);
nand UO_1211 (O_1211,N_19975,N_19867);
and UO_1212 (O_1212,N_19892,N_19916);
nor UO_1213 (O_1213,N_19869,N_19886);
nand UO_1214 (O_1214,N_19990,N_19884);
xnor UO_1215 (O_1215,N_19874,N_19957);
nor UO_1216 (O_1216,N_19906,N_19956);
xor UO_1217 (O_1217,N_19951,N_19876);
or UO_1218 (O_1218,N_19951,N_19884);
nand UO_1219 (O_1219,N_19952,N_19913);
nand UO_1220 (O_1220,N_19927,N_19972);
xnor UO_1221 (O_1221,N_19923,N_19875);
nor UO_1222 (O_1222,N_19921,N_19857);
nand UO_1223 (O_1223,N_19949,N_19925);
nor UO_1224 (O_1224,N_19968,N_19861);
nand UO_1225 (O_1225,N_19888,N_19906);
and UO_1226 (O_1226,N_19882,N_19979);
nor UO_1227 (O_1227,N_19951,N_19928);
xor UO_1228 (O_1228,N_19905,N_19904);
nand UO_1229 (O_1229,N_19889,N_19941);
and UO_1230 (O_1230,N_19940,N_19937);
or UO_1231 (O_1231,N_19851,N_19957);
nand UO_1232 (O_1232,N_19851,N_19988);
and UO_1233 (O_1233,N_19950,N_19959);
or UO_1234 (O_1234,N_19906,N_19908);
nand UO_1235 (O_1235,N_19985,N_19849);
nand UO_1236 (O_1236,N_19884,N_19941);
nor UO_1237 (O_1237,N_19949,N_19858);
nor UO_1238 (O_1238,N_19872,N_19899);
and UO_1239 (O_1239,N_19994,N_19920);
nor UO_1240 (O_1240,N_19841,N_19943);
xnor UO_1241 (O_1241,N_19887,N_19971);
and UO_1242 (O_1242,N_19880,N_19943);
and UO_1243 (O_1243,N_19864,N_19938);
xnor UO_1244 (O_1244,N_19911,N_19894);
nand UO_1245 (O_1245,N_19978,N_19862);
nand UO_1246 (O_1246,N_19942,N_19904);
xnor UO_1247 (O_1247,N_19893,N_19860);
nor UO_1248 (O_1248,N_19952,N_19991);
or UO_1249 (O_1249,N_19882,N_19853);
and UO_1250 (O_1250,N_19933,N_19930);
or UO_1251 (O_1251,N_19886,N_19891);
or UO_1252 (O_1252,N_19896,N_19884);
nand UO_1253 (O_1253,N_19921,N_19981);
xnor UO_1254 (O_1254,N_19943,N_19931);
nand UO_1255 (O_1255,N_19971,N_19969);
nand UO_1256 (O_1256,N_19961,N_19962);
xor UO_1257 (O_1257,N_19916,N_19842);
nand UO_1258 (O_1258,N_19932,N_19951);
or UO_1259 (O_1259,N_19936,N_19905);
and UO_1260 (O_1260,N_19861,N_19855);
nor UO_1261 (O_1261,N_19876,N_19947);
xnor UO_1262 (O_1262,N_19954,N_19948);
and UO_1263 (O_1263,N_19989,N_19928);
or UO_1264 (O_1264,N_19976,N_19924);
nor UO_1265 (O_1265,N_19933,N_19977);
and UO_1266 (O_1266,N_19900,N_19952);
xnor UO_1267 (O_1267,N_19948,N_19975);
and UO_1268 (O_1268,N_19958,N_19902);
and UO_1269 (O_1269,N_19869,N_19992);
nor UO_1270 (O_1270,N_19947,N_19893);
nand UO_1271 (O_1271,N_19871,N_19971);
nor UO_1272 (O_1272,N_19994,N_19881);
and UO_1273 (O_1273,N_19863,N_19895);
nand UO_1274 (O_1274,N_19998,N_19850);
nand UO_1275 (O_1275,N_19859,N_19886);
and UO_1276 (O_1276,N_19879,N_19914);
and UO_1277 (O_1277,N_19998,N_19909);
xnor UO_1278 (O_1278,N_19857,N_19905);
nor UO_1279 (O_1279,N_19965,N_19991);
nand UO_1280 (O_1280,N_19987,N_19933);
xor UO_1281 (O_1281,N_19981,N_19866);
and UO_1282 (O_1282,N_19958,N_19991);
and UO_1283 (O_1283,N_19955,N_19849);
nand UO_1284 (O_1284,N_19864,N_19892);
xor UO_1285 (O_1285,N_19851,N_19996);
and UO_1286 (O_1286,N_19877,N_19899);
or UO_1287 (O_1287,N_19968,N_19879);
nand UO_1288 (O_1288,N_19891,N_19985);
or UO_1289 (O_1289,N_19946,N_19866);
nand UO_1290 (O_1290,N_19883,N_19855);
and UO_1291 (O_1291,N_19863,N_19914);
nor UO_1292 (O_1292,N_19873,N_19954);
and UO_1293 (O_1293,N_19888,N_19854);
and UO_1294 (O_1294,N_19913,N_19929);
nand UO_1295 (O_1295,N_19935,N_19965);
or UO_1296 (O_1296,N_19920,N_19968);
xnor UO_1297 (O_1297,N_19890,N_19952);
or UO_1298 (O_1298,N_19986,N_19850);
nand UO_1299 (O_1299,N_19855,N_19993);
or UO_1300 (O_1300,N_19928,N_19890);
and UO_1301 (O_1301,N_19962,N_19875);
or UO_1302 (O_1302,N_19894,N_19863);
nand UO_1303 (O_1303,N_19855,N_19964);
nor UO_1304 (O_1304,N_19852,N_19955);
and UO_1305 (O_1305,N_19856,N_19979);
xnor UO_1306 (O_1306,N_19926,N_19847);
nand UO_1307 (O_1307,N_19868,N_19975);
and UO_1308 (O_1308,N_19922,N_19933);
nand UO_1309 (O_1309,N_19991,N_19850);
nor UO_1310 (O_1310,N_19964,N_19927);
nor UO_1311 (O_1311,N_19972,N_19857);
nand UO_1312 (O_1312,N_19853,N_19942);
nor UO_1313 (O_1313,N_19959,N_19864);
or UO_1314 (O_1314,N_19869,N_19998);
nor UO_1315 (O_1315,N_19860,N_19874);
and UO_1316 (O_1316,N_19874,N_19906);
nand UO_1317 (O_1317,N_19917,N_19871);
and UO_1318 (O_1318,N_19843,N_19975);
nor UO_1319 (O_1319,N_19848,N_19973);
or UO_1320 (O_1320,N_19978,N_19985);
nand UO_1321 (O_1321,N_19985,N_19926);
xnor UO_1322 (O_1322,N_19862,N_19940);
or UO_1323 (O_1323,N_19900,N_19984);
nand UO_1324 (O_1324,N_19990,N_19923);
and UO_1325 (O_1325,N_19902,N_19957);
and UO_1326 (O_1326,N_19857,N_19943);
and UO_1327 (O_1327,N_19923,N_19903);
or UO_1328 (O_1328,N_19926,N_19927);
and UO_1329 (O_1329,N_19862,N_19967);
and UO_1330 (O_1330,N_19967,N_19985);
and UO_1331 (O_1331,N_19934,N_19925);
or UO_1332 (O_1332,N_19984,N_19840);
and UO_1333 (O_1333,N_19924,N_19935);
nor UO_1334 (O_1334,N_19851,N_19971);
xor UO_1335 (O_1335,N_19972,N_19841);
xnor UO_1336 (O_1336,N_19905,N_19888);
nand UO_1337 (O_1337,N_19977,N_19845);
or UO_1338 (O_1338,N_19944,N_19961);
nor UO_1339 (O_1339,N_19863,N_19867);
and UO_1340 (O_1340,N_19890,N_19874);
nor UO_1341 (O_1341,N_19981,N_19888);
nor UO_1342 (O_1342,N_19892,N_19858);
xnor UO_1343 (O_1343,N_19877,N_19953);
and UO_1344 (O_1344,N_19915,N_19994);
nand UO_1345 (O_1345,N_19948,N_19907);
and UO_1346 (O_1346,N_19898,N_19879);
xnor UO_1347 (O_1347,N_19948,N_19943);
or UO_1348 (O_1348,N_19916,N_19985);
nor UO_1349 (O_1349,N_19869,N_19922);
xnor UO_1350 (O_1350,N_19958,N_19980);
xor UO_1351 (O_1351,N_19901,N_19921);
or UO_1352 (O_1352,N_19954,N_19984);
nor UO_1353 (O_1353,N_19973,N_19985);
nand UO_1354 (O_1354,N_19893,N_19969);
or UO_1355 (O_1355,N_19898,N_19884);
and UO_1356 (O_1356,N_19856,N_19887);
nor UO_1357 (O_1357,N_19926,N_19932);
and UO_1358 (O_1358,N_19933,N_19874);
and UO_1359 (O_1359,N_19884,N_19968);
or UO_1360 (O_1360,N_19928,N_19938);
nor UO_1361 (O_1361,N_19941,N_19925);
nor UO_1362 (O_1362,N_19883,N_19931);
and UO_1363 (O_1363,N_19927,N_19952);
nor UO_1364 (O_1364,N_19998,N_19991);
xnor UO_1365 (O_1365,N_19922,N_19878);
and UO_1366 (O_1366,N_19955,N_19999);
nor UO_1367 (O_1367,N_19969,N_19859);
or UO_1368 (O_1368,N_19912,N_19894);
xor UO_1369 (O_1369,N_19869,N_19852);
nor UO_1370 (O_1370,N_19848,N_19930);
nor UO_1371 (O_1371,N_19979,N_19934);
nand UO_1372 (O_1372,N_19948,N_19909);
xnor UO_1373 (O_1373,N_19954,N_19923);
nand UO_1374 (O_1374,N_19916,N_19996);
nor UO_1375 (O_1375,N_19889,N_19935);
nand UO_1376 (O_1376,N_19957,N_19987);
and UO_1377 (O_1377,N_19870,N_19921);
and UO_1378 (O_1378,N_19990,N_19958);
nor UO_1379 (O_1379,N_19987,N_19858);
or UO_1380 (O_1380,N_19914,N_19974);
or UO_1381 (O_1381,N_19862,N_19968);
and UO_1382 (O_1382,N_19921,N_19984);
nand UO_1383 (O_1383,N_19911,N_19984);
xnor UO_1384 (O_1384,N_19964,N_19962);
and UO_1385 (O_1385,N_19862,N_19980);
xor UO_1386 (O_1386,N_19852,N_19998);
or UO_1387 (O_1387,N_19888,N_19865);
nand UO_1388 (O_1388,N_19889,N_19888);
nand UO_1389 (O_1389,N_19933,N_19939);
nor UO_1390 (O_1390,N_19938,N_19947);
nor UO_1391 (O_1391,N_19913,N_19899);
nor UO_1392 (O_1392,N_19998,N_19949);
nand UO_1393 (O_1393,N_19883,N_19945);
xnor UO_1394 (O_1394,N_19842,N_19857);
or UO_1395 (O_1395,N_19845,N_19956);
nand UO_1396 (O_1396,N_19876,N_19983);
nand UO_1397 (O_1397,N_19977,N_19949);
nor UO_1398 (O_1398,N_19891,N_19889);
nor UO_1399 (O_1399,N_19990,N_19840);
nand UO_1400 (O_1400,N_19995,N_19895);
xnor UO_1401 (O_1401,N_19922,N_19944);
nor UO_1402 (O_1402,N_19874,N_19904);
nand UO_1403 (O_1403,N_19933,N_19897);
and UO_1404 (O_1404,N_19962,N_19994);
nor UO_1405 (O_1405,N_19933,N_19842);
and UO_1406 (O_1406,N_19914,N_19925);
and UO_1407 (O_1407,N_19975,N_19966);
xor UO_1408 (O_1408,N_19884,N_19900);
xnor UO_1409 (O_1409,N_19873,N_19980);
and UO_1410 (O_1410,N_19844,N_19979);
nor UO_1411 (O_1411,N_19859,N_19914);
or UO_1412 (O_1412,N_19848,N_19917);
nand UO_1413 (O_1413,N_19855,N_19926);
nor UO_1414 (O_1414,N_19943,N_19874);
and UO_1415 (O_1415,N_19843,N_19851);
or UO_1416 (O_1416,N_19921,N_19974);
nor UO_1417 (O_1417,N_19852,N_19918);
and UO_1418 (O_1418,N_19874,N_19934);
nor UO_1419 (O_1419,N_19885,N_19904);
and UO_1420 (O_1420,N_19961,N_19950);
or UO_1421 (O_1421,N_19848,N_19901);
nor UO_1422 (O_1422,N_19921,N_19862);
xnor UO_1423 (O_1423,N_19964,N_19942);
and UO_1424 (O_1424,N_19920,N_19951);
or UO_1425 (O_1425,N_19858,N_19915);
and UO_1426 (O_1426,N_19982,N_19969);
nor UO_1427 (O_1427,N_19863,N_19949);
nand UO_1428 (O_1428,N_19853,N_19944);
and UO_1429 (O_1429,N_19936,N_19916);
and UO_1430 (O_1430,N_19877,N_19992);
or UO_1431 (O_1431,N_19868,N_19981);
and UO_1432 (O_1432,N_19984,N_19889);
or UO_1433 (O_1433,N_19913,N_19840);
nand UO_1434 (O_1434,N_19842,N_19941);
and UO_1435 (O_1435,N_19891,N_19981);
and UO_1436 (O_1436,N_19964,N_19995);
xnor UO_1437 (O_1437,N_19866,N_19987);
nand UO_1438 (O_1438,N_19962,N_19894);
xnor UO_1439 (O_1439,N_19907,N_19868);
nor UO_1440 (O_1440,N_19974,N_19925);
nor UO_1441 (O_1441,N_19844,N_19849);
or UO_1442 (O_1442,N_19859,N_19902);
or UO_1443 (O_1443,N_19927,N_19900);
or UO_1444 (O_1444,N_19985,N_19942);
and UO_1445 (O_1445,N_19919,N_19885);
xnor UO_1446 (O_1446,N_19882,N_19973);
nand UO_1447 (O_1447,N_19965,N_19923);
nand UO_1448 (O_1448,N_19892,N_19845);
and UO_1449 (O_1449,N_19982,N_19917);
nor UO_1450 (O_1450,N_19945,N_19935);
nand UO_1451 (O_1451,N_19968,N_19848);
xnor UO_1452 (O_1452,N_19893,N_19927);
and UO_1453 (O_1453,N_19862,N_19932);
or UO_1454 (O_1454,N_19880,N_19843);
or UO_1455 (O_1455,N_19869,N_19847);
and UO_1456 (O_1456,N_19855,N_19961);
nand UO_1457 (O_1457,N_19996,N_19845);
nor UO_1458 (O_1458,N_19939,N_19908);
nor UO_1459 (O_1459,N_19978,N_19947);
xnor UO_1460 (O_1460,N_19916,N_19930);
nand UO_1461 (O_1461,N_19998,N_19859);
xor UO_1462 (O_1462,N_19877,N_19870);
or UO_1463 (O_1463,N_19954,N_19952);
or UO_1464 (O_1464,N_19976,N_19945);
and UO_1465 (O_1465,N_19871,N_19958);
nor UO_1466 (O_1466,N_19855,N_19909);
and UO_1467 (O_1467,N_19992,N_19954);
nand UO_1468 (O_1468,N_19986,N_19975);
xnor UO_1469 (O_1469,N_19996,N_19876);
nand UO_1470 (O_1470,N_19910,N_19930);
xor UO_1471 (O_1471,N_19943,N_19856);
nand UO_1472 (O_1472,N_19969,N_19970);
or UO_1473 (O_1473,N_19964,N_19946);
and UO_1474 (O_1474,N_19880,N_19960);
and UO_1475 (O_1475,N_19987,N_19916);
nand UO_1476 (O_1476,N_19902,N_19915);
nor UO_1477 (O_1477,N_19954,N_19858);
nand UO_1478 (O_1478,N_19989,N_19962);
nor UO_1479 (O_1479,N_19960,N_19953);
and UO_1480 (O_1480,N_19913,N_19890);
and UO_1481 (O_1481,N_19901,N_19935);
nand UO_1482 (O_1482,N_19879,N_19919);
nand UO_1483 (O_1483,N_19858,N_19875);
xnor UO_1484 (O_1484,N_19960,N_19899);
and UO_1485 (O_1485,N_19903,N_19887);
xor UO_1486 (O_1486,N_19985,N_19930);
nand UO_1487 (O_1487,N_19972,N_19953);
and UO_1488 (O_1488,N_19875,N_19983);
or UO_1489 (O_1489,N_19954,N_19910);
and UO_1490 (O_1490,N_19859,N_19864);
nand UO_1491 (O_1491,N_19885,N_19862);
nor UO_1492 (O_1492,N_19865,N_19907);
nor UO_1493 (O_1493,N_19892,N_19953);
nor UO_1494 (O_1494,N_19870,N_19896);
or UO_1495 (O_1495,N_19959,N_19888);
xor UO_1496 (O_1496,N_19851,N_19968);
nand UO_1497 (O_1497,N_19912,N_19956);
nand UO_1498 (O_1498,N_19898,N_19867);
nand UO_1499 (O_1499,N_19910,N_19904);
nand UO_1500 (O_1500,N_19896,N_19991);
nand UO_1501 (O_1501,N_19869,N_19985);
nand UO_1502 (O_1502,N_19975,N_19915);
nor UO_1503 (O_1503,N_19955,N_19906);
xor UO_1504 (O_1504,N_19907,N_19995);
xnor UO_1505 (O_1505,N_19918,N_19885);
and UO_1506 (O_1506,N_19958,N_19877);
xnor UO_1507 (O_1507,N_19843,N_19934);
or UO_1508 (O_1508,N_19896,N_19856);
nor UO_1509 (O_1509,N_19844,N_19862);
xnor UO_1510 (O_1510,N_19965,N_19843);
or UO_1511 (O_1511,N_19907,N_19848);
nand UO_1512 (O_1512,N_19955,N_19887);
nand UO_1513 (O_1513,N_19947,N_19887);
and UO_1514 (O_1514,N_19920,N_19896);
nand UO_1515 (O_1515,N_19891,N_19908);
nand UO_1516 (O_1516,N_19860,N_19939);
and UO_1517 (O_1517,N_19906,N_19912);
xnor UO_1518 (O_1518,N_19973,N_19961);
xor UO_1519 (O_1519,N_19856,N_19883);
and UO_1520 (O_1520,N_19995,N_19976);
xor UO_1521 (O_1521,N_19935,N_19971);
nor UO_1522 (O_1522,N_19968,N_19866);
xor UO_1523 (O_1523,N_19967,N_19953);
nor UO_1524 (O_1524,N_19964,N_19924);
and UO_1525 (O_1525,N_19892,N_19931);
nand UO_1526 (O_1526,N_19931,N_19955);
or UO_1527 (O_1527,N_19840,N_19989);
and UO_1528 (O_1528,N_19996,N_19862);
and UO_1529 (O_1529,N_19958,N_19964);
xnor UO_1530 (O_1530,N_19855,N_19968);
and UO_1531 (O_1531,N_19865,N_19872);
xnor UO_1532 (O_1532,N_19909,N_19904);
and UO_1533 (O_1533,N_19935,N_19893);
and UO_1534 (O_1534,N_19930,N_19891);
or UO_1535 (O_1535,N_19939,N_19948);
or UO_1536 (O_1536,N_19890,N_19991);
nand UO_1537 (O_1537,N_19973,N_19957);
nand UO_1538 (O_1538,N_19955,N_19916);
nor UO_1539 (O_1539,N_19901,N_19972);
and UO_1540 (O_1540,N_19859,N_19982);
or UO_1541 (O_1541,N_19862,N_19895);
and UO_1542 (O_1542,N_19907,N_19943);
and UO_1543 (O_1543,N_19932,N_19956);
nor UO_1544 (O_1544,N_19864,N_19956);
and UO_1545 (O_1545,N_19996,N_19969);
nand UO_1546 (O_1546,N_19914,N_19870);
nor UO_1547 (O_1547,N_19924,N_19928);
xnor UO_1548 (O_1548,N_19891,N_19879);
or UO_1549 (O_1549,N_19929,N_19935);
or UO_1550 (O_1550,N_19900,N_19875);
or UO_1551 (O_1551,N_19899,N_19967);
xnor UO_1552 (O_1552,N_19986,N_19848);
or UO_1553 (O_1553,N_19907,N_19914);
xnor UO_1554 (O_1554,N_19859,N_19992);
xor UO_1555 (O_1555,N_19964,N_19935);
nor UO_1556 (O_1556,N_19963,N_19900);
xnor UO_1557 (O_1557,N_19886,N_19850);
or UO_1558 (O_1558,N_19851,N_19903);
and UO_1559 (O_1559,N_19951,N_19981);
nor UO_1560 (O_1560,N_19936,N_19986);
nor UO_1561 (O_1561,N_19874,N_19995);
or UO_1562 (O_1562,N_19881,N_19884);
or UO_1563 (O_1563,N_19928,N_19912);
or UO_1564 (O_1564,N_19979,N_19889);
xnor UO_1565 (O_1565,N_19909,N_19852);
nand UO_1566 (O_1566,N_19982,N_19858);
or UO_1567 (O_1567,N_19891,N_19939);
and UO_1568 (O_1568,N_19914,N_19917);
and UO_1569 (O_1569,N_19883,N_19925);
nand UO_1570 (O_1570,N_19967,N_19936);
nor UO_1571 (O_1571,N_19855,N_19875);
xnor UO_1572 (O_1572,N_19975,N_19858);
nand UO_1573 (O_1573,N_19981,N_19967);
or UO_1574 (O_1574,N_19961,N_19913);
xnor UO_1575 (O_1575,N_19861,N_19938);
nand UO_1576 (O_1576,N_19985,N_19906);
xor UO_1577 (O_1577,N_19909,N_19937);
xnor UO_1578 (O_1578,N_19954,N_19991);
or UO_1579 (O_1579,N_19926,N_19878);
or UO_1580 (O_1580,N_19854,N_19862);
nor UO_1581 (O_1581,N_19937,N_19989);
nand UO_1582 (O_1582,N_19906,N_19889);
nand UO_1583 (O_1583,N_19988,N_19882);
or UO_1584 (O_1584,N_19923,N_19900);
or UO_1585 (O_1585,N_19877,N_19882);
and UO_1586 (O_1586,N_19902,N_19981);
nand UO_1587 (O_1587,N_19998,N_19960);
and UO_1588 (O_1588,N_19888,N_19931);
or UO_1589 (O_1589,N_19901,N_19898);
nand UO_1590 (O_1590,N_19972,N_19866);
xnor UO_1591 (O_1591,N_19900,N_19981);
xnor UO_1592 (O_1592,N_19950,N_19979);
and UO_1593 (O_1593,N_19979,N_19866);
or UO_1594 (O_1594,N_19977,N_19957);
nor UO_1595 (O_1595,N_19970,N_19975);
or UO_1596 (O_1596,N_19878,N_19976);
xor UO_1597 (O_1597,N_19910,N_19927);
nor UO_1598 (O_1598,N_19906,N_19957);
nor UO_1599 (O_1599,N_19876,N_19922);
xnor UO_1600 (O_1600,N_19959,N_19915);
nand UO_1601 (O_1601,N_19993,N_19842);
or UO_1602 (O_1602,N_19948,N_19963);
or UO_1603 (O_1603,N_19862,N_19866);
xnor UO_1604 (O_1604,N_19993,N_19865);
and UO_1605 (O_1605,N_19906,N_19946);
nor UO_1606 (O_1606,N_19949,N_19912);
nand UO_1607 (O_1607,N_19845,N_19910);
nand UO_1608 (O_1608,N_19893,N_19898);
and UO_1609 (O_1609,N_19959,N_19922);
and UO_1610 (O_1610,N_19927,N_19868);
nand UO_1611 (O_1611,N_19882,N_19978);
nand UO_1612 (O_1612,N_19902,N_19938);
nor UO_1613 (O_1613,N_19927,N_19863);
xor UO_1614 (O_1614,N_19924,N_19945);
or UO_1615 (O_1615,N_19906,N_19923);
and UO_1616 (O_1616,N_19924,N_19968);
xnor UO_1617 (O_1617,N_19890,N_19974);
nand UO_1618 (O_1618,N_19915,N_19998);
xnor UO_1619 (O_1619,N_19933,N_19859);
and UO_1620 (O_1620,N_19909,N_19928);
or UO_1621 (O_1621,N_19996,N_19935);
xor UO_1622 (O_1622,N_19871,N_19887);
nor UO_1623 (O_1623,N_19870,N_19905);
nor UO_1624 (O_1624,N_19964,N_19968);
or UO_1625 (O_1625,N_19954,N_19955);
or UO_1626 (O_1626,N_19868,N_19873);
nand UO_1627 (O_1627,N_19997,N_19979);
nand UO_1628 (O_1628,N_19877,N_19855);
nand UO_1629 (O_1629,N_19859,N_19958);
nor UO_1630 (O_1630,N_19953,N_19959);
nor UO_1631 (O_1631,N_19897,N_19840);
and UO_1632 (O_1632,N_19863,N_19902);
nand UO_1633 (O_1633,N_19932,N_19866);
nor UO_1634 (O_1634,N_19964,N_19853);
or UO_1635 (O_1635,N_19877,N_19852);
xor UO_1636 (O_1636,N_19929,N_19885);
and UO_1637 (O_1637,N_19848,N_19880);
xor UO_1638 (O_1638,N_19987,N_19990);
nor UO_1639 (O_1639,N_19926,N_19869);
nor UO_1640 (O_1640,N_19988,N_19972);
or UO_1641 (O_1641,N_19991,N_19875);
nand UO_1642 (O_1642,N_19845,N_19840);
nor UO_1643 (O_1643,N_19939,N_19867);
nand UO_1644 (O_1644,N_19966,N_19861);
xnor UO_1645 (O_1645,N_19990,N_19878);
or UO_1646 (O_1646,N_19966,N_19922);
xnor UO_1647 (O_1647,N_19964,N_19990);
and UO_1648 (O_1648,N_19960,N_19851);
nor UO_1649 (O_1649,N_19921,N_19932);
and UO_1650 (O_1650,N_19965,N_19930);
and UO_1651 (O_1651,N_19988,N_19981);
or UO_1652 (O_1652,N_19999,N_19851);
xnor UO_1653 (O_1653,N_19910,N_19874);
nand UO_1654 (O_1654,N_19896,N_19862);
nand UO_1655 (O_1655,N_19978,N_19915);
and UO_1656 (O_1656,N_19891,N_19932);
xor UO_1657 (O_1657,N_19976,N_19864);
xnor UO_1658 (O_1658,N_19926,N_19858);
or UO_1659 (O_1659,N_19867,N_19907);
or UO_1660 (O_1660,N_19948,N_19971);
nor UO_1661 (O_1661,N_19881,N_19869);
nor UO_1662 (O_1662,N_19939,N_19968);
nand UO_1663 (O_1663,N_19867,N_19843);
or UO_1664 (O_1664,N_19980,N_19991);
and UO_1665 (O_1665,N_19908,N_19883);
nor UO_1666 (O_1666,N_19974,N_19873);
or UO_1667 (O_1667,N_19941,N_19847);
nor UO_1668 (O_1668,N_19936,N_19910);
nand UO_1669 (O_1669,N_19900,N_19916);
and UO_1670 (O_1670,N_19843,N_19968);
or UO_1671 (O_1671,N_19990,N_19922);
and UO_1672 (O_1672,N_19933,N_19913);
nand UO_1673 (O_1673,N_19840,N_19982);
or UO_1674 (O_1674,N_19989,N_19995);
xnor UO_1675 (O_1675,N_19952,N_19945);
nand UO_1676 (O_1676,N_19915,N_19849);
and UO_1677 (O_1677,N_19934,N_19908);
and UO_1678 (O_1678,N_19998,N_19961);
or UO_1679 (O_1679,N_19872,N_19848);
or UO_1680 (O_1680,N_19930,N_19995);
xor UO_1681 (O_1681,N_19857,N_19915);
xor UO_1682 (O_1682,N_19915,N_19850);
xnor UO_1683 (O_1683,N_19888,N_19869);
or UO_1684 (O_1684,N_19847,N_19903);
xnor UO_1685 (O_1685,N_19862,N_19977);
nand UO_1686 (O_1686,N_19846,N_19899);
nand UO_1687 (O_1687,N_19872,N_19993);
nand UO_1688 (O_1688,N_19921,N_19842);
nand UO_1689 (O_1689,N_19851,N_19958);
and UO_1690 (O_1690,N_19926,N_19874);
and UO_1691 (O_1691,N_19852,N_19881);
nand UO_1692 (O_1692,N_19881,N_19857);
xor UO_1693 (O_1693,N_19857,N_19977);
and UO_1694 (O_1694,N_19855,N_19933);
and UO_1695 (O_1695,N_19903,N_19996);
nand UO_1696 (O_1696,N_19949,N_19907);
and UO_1697 (O_1697,N_19870,N_19920);
or UO_1698 (O_1698,N_19898,N_19965);
nor UO_1699 (O_1699,N_19939,N_19899);
or UO_1700 (O_1700,N_19992,N_19941);
xnor UO_1701 (O_1701,N_19941,N_19982);
xor UO_1702 (O_1702,N_19973,N_19851);
xor UO_1703 (O_1703,N_19954,N_19934);
and UO_1704 (O_1704,N_19915,N_19970);
nor UO_1705 (O_1705,N_19878,N_19996);
or UO_1706 (O_1706,N_19857,N_19910);
or UO_1707 (O_1707,N_19978,N_19897);
or UO_1708 (O_1708,N_19841,N_19865);
nor UO_1709 (O_1709,N_19924,N_19918);
and UO_1710 (O_1710,N_19926,N_19921);
nand UO_1711 (O_1711,N_19847,N_19901);
and UO_1712 (O_1712,N_19980,N_19989);
nand UO_1713 (O_1713,N_19852,N_19983);
nor UO_1714 (O_1714,N_19843,N_19953);
and UO_1715 (O_1715,N_19987,N_19983);
nand UO_1716 (O_1716,N_19854,N_19868);
and UO_1717 (O_1717,N_19880,N_19970);
nor UO_1718 (O_1718,N_19891,N_19942);
or UO_1719 (O_1719,N_19872,N_19961);
nor UO_1720 (O_1720,N_19846,N_19910);
xor UO_1721 (O_1721,N_19919,N_19977);
xnor UO_1722 (O_1722,N_19938,N_19880);
or UO_1723 (O_1723,N_19950,N_19993);
nor UO_1724 (O_1724,N_19860,N_19976);
nand UO_1725 (O_1725,N_19942,N_19897);
xor UO_1726 (O_1726,N_19932,N_19969);
nand UO_1727 (O_1727,N_19924,N_19841);
nor UO_1728 (O_1728,N_19901,N_19883);
or UO_1729 (O_1729,N_19867,N_19850);
and UO_1730 (O_1730,N_19884,N_19929);
xor UO_1731 (O_1731,N_19912,N_19934);
nand UO_1732 (O_1732,N_19917,N_19985);
nand UO_1733 (O_1733,N_19986,N_19957);
and UO_1734 (O_1734,N_19877,N_19940);
nand UO_1735 (O_1735,N_19862,N_19908);
or UO_1736 (O_1736,N_19858,N_19971);
xor UO_1737 (O_1737,N_19967,N_19946);
or UO_1738 (O_1738,N_19921,N_19876);
xnor UO_1739 (O_1739,N_19878,N_19916);
or UO_1740 (O_1740,N_19938,N_19922);
nand UO_1741 (O_1741,N_19869,N_19866);
nor UO_1742 (O_1742,N_19883,N_19940);
xnor UO_1743 (O_1743,N_19893,N_19840);
nor UO_1744 (O_1744,N_19882,N_19878);
or UO_1745 (O_1745,N_19914,N_19943);
nor UO_1746 (O_1746,N_19935,N_19926);
and UO_1747 (O_1747,N_19884,N_19902);
or UO_1748 (O_1748,N_19980,N_19859);
and UO_1749 (O_1749,N_19931,N_19920);
and UO_1750 (O_1750,N_19944,N_19912);
and UO_1751 (O_1751,N_19912,N_19851);
nor UO_1752 (O_1752,N_19927,N_19957);
nor UO_1753 (O_1753,N_19926,N_19917);
and UO_1754 (O_1754,N_19955,N_19889);
nor UO_1755 (O_1755,N_19885,N_19954);
xor UO_1756 (O_1756,N_19984,N_19955);
and UO_1757 (O_1757,N_19970,N_19842);
nand UO_1758 (O_1758,N_19914,N_19898);
xnor UO_1759 (O_1759,N_19970,N_19987);
xor UO_1760 (O_1760,N_19955,N_19882);
xor UO_1761 (O_1761,N_19921,N_19956);
or UO_1762 (O_1762,N_19914,N_19904);
or UO_1763 (O_1763,N_19956,N_19891);
and UO_1764 (O_1764,N_19911,N_19891);
or UO_1765 (O_1765,N_19951,N_19994);
or UO_1766 (O_1766,N_19851,N_19875);
nor UO_1767 (O_1767,N_19928,N_19884);
and UO_1768 (O_1768,N_19991,N_19967);
xor UO_1769 (O_1769,N_19900,N_19976);
nor UO_1770 (O_1770,N_19960,N_19858);
and UO_1771 (O_1771,N_19951,N_19970);
xor UO_1772 (O_1772,N_19885,N_19916);
or UO_1773 (O_1773,N_19866,N_19970);
and UO_1774 (O_1774,N_19888,N_19995);
xnor UO_1775 (O_1775,N_19893,N_19904);
xor UO_1776 (O_1776,N_19840,N_19980);
and UO_1777 (O_1777,N_19856,N_19937);
and UO_1778 (O_1778,N_19860,N_19903);
nand UO_1779 (O_1779,N_19992,N_19899);
or UO_1780 (O_1780,N_19977,N_19920);
nor UO_1781 (O_1781,N_19844,N_19860);
or UO_1782 (O_1782,N_19867,N_19924);
and UO_1783 (O_1783,N_19841,N_19997);
nor UO_1784 (O_1784,N_19989,N_19977);
nor UO_1785 (O_1785,N_19898,N_19921);
nand UO_1786 (O_1786,N_19875,N_19898);
and UO_1787 (O_1787,N_19934,N_19884);
or UO_1788 (O_1788,N_19915,N_19934);
nor UO_1789 (O_1789,N_19935,N_19845);
nor UO_1790 (O_1790,N_19979,N_19964);
nor UO_1791 (O_1791,N_19960,N_19846);
xor UO_1792 (O_1792,N_19881,N_19950);
nor UO_1793 (O_1793,N_19945,N_19977);
or UO_1794 (O_1794,N_19871,N_19841);
xor UO_1795 (O_1795,N_19877,N_19938);
nor UO_1796 (O_1796,N_19926,N_19971);
nor UO_1797 (O_1797,N_19970,N_19849);
or UO_1798 (O_1798,N_19875,N_19970);
or UO_1799 (O_1799,N_19934,N_19961);
or UO_1800 (O_1800,N_19943,N_19941);
or UO_1801 (O_1801,N_19968,N_19917);
and UO_1802 (O_1802,N_19882,N_19987);
and UO_1803 (O_1803,N_19894,N_19881);
or UO_1804 (O_1804,N_19911,N_19982);
nor UO_1805 (O_1805,N_19986,N_19861);
and UO_1806 (O_1806,N_19994,N_19866);
xnor UO_1807 (O_1807,N_19868,N_19892);
or UO_1808 (O_1808,N_19861,N_19900);
and UO_1809 (O_1809,N_19944,N_19950);
and UO_1810 (O_1810,N_19909,N_19895);
nor UO_1811 (O_1811,N_19978,N_19904);
nor UO_1812 (O_1812,N_19846,N_19856);
and UO_1813 (O_1813,N_19931,N_19899);
nor UO_1814 (O_1814,N_19855,N_19996);
nand UO_1815 (O_1815,N_19890,N_19951);
and UO_1816 (O_1816,N_19848,N_19854);
nand UO_1817 (O_1817,N_19921,N_19875);
xnor UO_1818 (O_1818,N_19914,N_19840);
or UO_1819 (O_1819,N_19968,N_19883);
and UO_1820 (O_1820,N_19857,N_19923);
xor UO_1821 (O_1821,N_19930,N_19889);
nand UO_1822 (O_1822,N_19972,N_19963);
xnor UO_1823 (O_1823,N_19927,N_19885);
nor UO_1824 (O_1824,N_19876,N_19909);
nor UO_1825 (O_1825,N_19958,N_19906);
nand UO_1826 (O_1826,N_19955,N_19862);
nor UO_1827 (O_1827,N_19887,N_19896);
nor UO_1828 (O_1828,N_19851,N_19915);
and UO_1829 (O_1829,N_19964,N_19883);
or UO_1830 (O_1830,N_19917,N_19971);
xor UO_1831 (O_1831,N_19981,N_19889);
nand UO_1832 (O_1832,N_19893,N_19970);
or UO_1833 (O_1833,N_19983,N_19976);
nor UO_1834 (O_1834,N_19980,N_19992);
nand UO_1835 (O_1835,N_19863,N_19897);
and UO_1836 (O_1836,N_19979,N_19888);
xnor UO_1837 (O_1837,N_19938,N_19956);
xnor UO_1838 (O_1838,N_19981,N_19844);
nand UO_1839 (O_1839,N_19993,N_19840);
or UO_1840 (O_1840,N_19948,N_19981);
and UO_1841 (O_1841,N_19892,N_19986);
xor UO_1842 (O_1842,N_19994,N_19854);
nand UO_1843 (O_1843,N_19868,N_19997);
nor UO_1844 (O_1844,N_19860,N_19840);
xnor UO_1845 (O_1845,N_19940,N_19907);
nand UO_1846 (O_1846,N_19912,N_19929);
or UO_1847 (O_1847,N_19873,N_19921);
or UO_1848 (O_1848,N_19996,N_19983);
nand UO_1849 (O_1849,N_19859,N_19986);
or UO_1850 (O_1850,N_19913,N_19857);
xnor UO_1851 (O_1851,N_19974,N_19930);
nand UO_1852 (O_1852,N_19968,N_19901);
xor UO_1853 (O_1853,N_19883,N_19900);
nand UO_1854 (O_1854,N_19856,N_19932);
and UO_1855 (O_1855,N_19984,N_19883);
nand UO_1856 (O_1856,N_19967,N_19871);
xnor UO_1857 (O_1857,N_19931,N_19972);
nor UO_1858 (O_1858,N_19843,N_19930);
xor UO_1859 (O_1859,N_19854,N_19894);
nor UO_1860 (O_1860,N_19894,N_19884);
and UO_1861 (O_1861,N_19959,N_19911);
or UO_1862 (O_1862,N_19843,N_19856);
nor UO_1863 (O_1863,N_19990,N_19970);
nand UO_1864 (O_1864,N_19862,N_19974);
and UO_1865 (O_1865,N_19956,N_19911);
xnor UO_1866 (O_1866,N_19995,N_19980);
and UO_1867 (O_1867,N_19966,N_19874);
xor UO_1868 (O_1868,N_19982,N_19910);
or UO_1869 (O_1869,N_19896,N_19993);
nor UO_1870 (O_1870,N_19992,N_19863);
nand UO_1871 (O_1871,N_19941,N_19868);
and UO_1872 (O_1872,N_19963,N_19960);
and UO_1873 (O_1873,N_19901,N_19910);
or UO_1874 (O_1874,N_19879,N_19959);
xor UO_1875 (O_1875,N_19907,N_19947);
nand UO_1876 (O_1876,N_19945,N_19862);
or UO_1877 (O_1877,N_19971,N_19947);
nor UO_1878 (O_1878,N_19856,N_19996);
nor UO_1879 (O_1879,N_19863,N_19888);
xor UO_1880 (O_1880,N_19840,N_19950);
or UO_1881 (O_1881,N_19855,N_19911);
or UO_1882 (O_1882,N_19990,N_19911);
nand UO_1883 (O_1883,N_19920,N_19875);
and UO_1884 (O_1884,N_19982,N_19998);
nor UO_1885 (O_1885,N_19987,N_19892);
nor UO_1886 (O_1886,N_19981,N_19919);
xor UO_1887 (O_1887,N_19940,N_19971);
and UO_1888 (O_1888,N_19877,N_19840);
xor UO_1889 (O_1889,N_19961,N_19858);
nand UO_1890 (O_1890,N_19915,N_19987);
xnor UO_1891 (O_1891,N_19907,N_19929);
and UO_1892 (O_1892,N_19840,N_19851);
nor UO_1893 (O_1893,N_19916,N_19970);
and UO_1894 (O_1894,N_19947,N_19900);
and UO_1895 (O_1895,N_19969,N_19933);
or UO_1896 (O_1896,N_19908,N_19958);
xor UO_1897 (O_1897,N_19893,N_19892);
and UO_1898 (O_1898,N_19945,N_19889);
xor UO_1899 (O_1899,N_19920,N_19973);
or UO_1900 (O_1900,N_19842,N_19874);
and UO_1901 (O_1901,N_19994,N_19997);
xor UO_1902 (O_1902,N_19951,N_19965);
xnor UO_1903 (O_1903,N_19941,N_19897);
nor UO_1904 (O_1904,N_19882,N_19903);
and UO_1905 (O_1905,N_19861,N_19973);
and UO_1906 (O_1906,N_19906,N_19962);
nand UO_1907 (O_1907,N_19970,N_19883);
xor UO_1908 (O_1908,N_19991,N_19942);
and UO_1909 (O_1909,N_19892,N_19877);
or UO_1910 (O_1910,N_19885,N_19960);
nor UO_1911 (O_1911,N_19858,N_19847);
nand UO_1912 (O_1912,N_19844,N_19925);
xor UO_1913 (O_1913,N_19913,N_19950);
and UO_1914 (O_1914,N_19899,N_19976);
and UO_1915 (O_1915,N_19909,N_19875);
and UO_1916 (O_1916,N_19917,N_19951);
xnor UO_1917 (O_1917,N_19926,N_19936);
and UO_1918 (O_1918,N_19848,N_19995);
xor UO_1919 (O_1919,N_19956,N_19924);
nor UO_1920 (O_1920,N_19923,N_19997);
and UO_1921 (O_1921,N_19859,N_19928);
or UO_1922 (O_1922,N_19920,N_19858);
nor UO_1923 (O_1923,N_19967,N_19875);
or UO_1924 (O_1924,N_19898,N_19935);
and UO_1925 (O_1925,N_19882,N_19859);
or UO_1926 (O_1926,N_19877,N_19856);
xnor UO_1927 (O_1927,N_19964,N_19989);
nand UO_1928 (O_1928,N_19915,N_19923);
nand UO_1929 (O_1929,N_19960,N_19968);
or UO_1930 (O_1930,N_19943,N_19866);
xor UO_1931 (O_1931,N_19972,N_19846);
or UO_1932 (O_1932,N_19882,N_19845);
nand UO_1933 (O_1933,N_19867,N_19919);
xnor UO_1934 (O_1934,N_19917,N_19928);
and UO_1935 (O_1935,N_19868,N_19947);
nand UO_1936 (O_1936,N_19972,N_19900);
nor UO_1937 (O_1937,N_19856,N_19951);
xor UO_1938 (O_1938,N_19915,N_19889);
xor UO_1939 (O_1939,N_19864,N_19933);
and UO_1940 (O_1940,N_19917,N_19952);
or UO_1941 (O_1941,N_19874,N_19864);
nor UO_1942 (O_1942,N_19993,N_19856);
and UO_1943 (O_1943,N_19989,N_19996);
xor UO_1944 (O_1944,N_19915,N_19881);
nor UO_1945 (O_1945,N_19897,N_19998);
nand UO_1946 (O_1946,N_19840,N_19842);
xor UO_1947 (O_1947,N_19855,N_19979);
or UO_1948 (O_1948,N_19952,N_19851);
nor UO_1949 (O_1949,N_19945,N_19972);
nor UO_1950 (O_1950,N_19917,N_19861);
nor UO_1951 (O_1951,N_19890,N_19980);
or UO_1952 (O_1952,N_19858,N_19903);
and UO_1953 (O_1953,N_19931,N_19930);
nor UO_1954 (O_1954,N_19897,N_19946);
nor UO_1955 (O_1955,N_19975,N_19953);
and UO_1956 (O_1956,N_19856,N_19998);
and UO_1957 (O_1957,N_19875,N_19903);
nand UO_1958 (O_1958,N_19973,N_19878);
nand UO_1959 (O_1959,N_19998,N_19893);
nor UO_1960 (O_1960,N_19897,N_19976);
xnor UO_1961 (O_1961,N_19881,N_19978);
nand UO_1962 (O_1962,N_19948,N_19979);
nor UO_1963 (O_1963,N_19880,N_19903);
and UO_1964 (O_1964,N_19927,N_19950);
or UO_1965 (O_1965,N_19927,N_19946);
and UO_1966 (O_1966,N_19905,N_19994);
or UO_1967 (O_1967,N_19906,N_19856);
or UO_1968 (O_1968,N_19918,N_19952);
xor UO_1969 (O_1969,N_19974,N_19984);
nor UO_1970 (O_1970,N_19968,N_19971);
xnor UO_1971 (O_1971,N_19896,N_19948);
xnor UO_1972 (O_1972,N_19888,N_19989);
nor UO_1973 (O_1973,N_19900,N_19979);
or UO_1974 (O_1974,N_19872,N_19970);
nand UO_1975 (O_1975,N_19938,N_19954);
and UO_1976 (O_1976,N_19928,N_19955);
or UO_1977 (O_1977,N_19875,N_19931);
nor UO_1978 (O_1978,N_19888,N_19843);
nand UO_1979 (O_1979,N_19986,N_19971);
nand UO_1980 (O_1980,N_19879,N_19970);
and UO_1981 (O_1981,N_19868,N_19939);
nand UO_1982 (O_1982,N_19892,N_19860);
nor UO_1983 (O_1983,N_19969,N_19922);
xor UO_1984 (O_1984,N_19994,N_19888);
or UO_1985 (O_1985,N_19881,N_19962);
and UO_1986 (O_1986,N_19853,N_19922);
xor UO_1987 (O_1987,N_19950,N_19925);
nand UO_1988 (O_1988,N_19882,N_19990);
and UO_1989 (O_1989,N_19997,N_19941);
xor UO_1990 (O_1990,N_19895,N_19936);
and UO_1991 (O_1991,N_19983,N_19937);
nand UO_1992 (O_1992,N_19899,N_19952);
or UO_1993 (O_1993,N_19852,N_19944);
nand UO_1994 (O_1994,N_19972,N_19930);
nor UO_1995 (O_1995,N_19952,N_19956);
xnor UO_1996 (O_1996,N_19969,N_19886);
nor UO_1997 (O_1997,N_19918,N_19868);
or UO_1998 (O_1998,N_19965,N_19984);
nor UO_1999 (O_1999,N_19897,N_19969);
xnor UO_2000 (O_2000,N_19969,N_19860);
or UO_2001 (O_2001,N_19934,N_19940);
nor UO_2002 (O_2002,N_19885,N_19859);
nand UO_2003 (O_2003,N_19898,N_19843);
and UO_2004 (O_2004,N_19858,N_19955);
xnor UO_2005 (O_2005,N_19852,N_19939);
and UO_2006 (O_2006,N_19971,N_19878);
or UO_2007 (O_2007,N_19983,N_19990);
xnor UO_2008 (O_2008,N_19937,N_19988);
or UO_2009 (O_2009,N_19971,N_19850);
and UO_2010 (O_2010,N_19948,N_19857);
and UO_2011 (O_2011,N_19870,N_19965);
nand UO_2012 (O_2012,N_19901,N_19983);
and UO_2013 (O_2013,N_19897,N_19889);
or UO_2014 (O_2014,N_19927,N_19998);
nand UO_2015 (O_2015,N_19980,N_19851);
xor UO_2016 (O_2016,N_19847,N_19958);
and UO_2017 (O_2017,N_19879,N_19902);
and UO_2018 (O_2018,N_19977,N_19841);
nor UO_2019 (O_2019,N_19856,N_19987);
nand UO_2020 (O_2020,N_19929,N_19865);
nand UO_2021 (O_2021,N_19925,N_19937);
xor UO_2022 (O_2022,N_19904,N_19982);
xnor UO_2023 (O_2023,N_19968,N_19977);
and UO_2024 (O_2024,N_19870,N_19889);
nand UO_2025 (O_2025,N_19991,N_19861);
and UO_2026 (O_2026,N_19885,N_19921);
or UO_2027 (O_2027,N_19875,N_19860);
nand UO_2028 (O_2028,N_19935,N_19844);
and UO_2029 (O_2029,N_19991,N_19932);
xnor UO_2030 (O_2030,N_19949,N_19939);
nand UO_2031 (O_2031,N_19886,N_19947);
xor UO_2032 (O_2032,N_19905,N_19969);
nand UO_2033 (O_2033,N_19928,N_19985);
nor UO_2034 (O_2034,N_19989,N_19949);
and UO_2035 (O_2035,N_19940,N_19987);
or UO_2036 (O_2036,N_19990,N_19934);
or UO_2037 (O_2037,N_19991,N_19948);
nor UO_2038 (O_2038,N_19846,N_19936);
or UO_2039 (O_2039,N_19931,N_19956);
nor UO_2040 (O_2040,N_19978,N_19902);
nand UO_2041 (O_2041,N_19993,N_19889);
nand UO_2042 (O_2042,N_19892,N_19903);
xor UO_2043 (O_2043,N_19902,N_19840);
nand UO_2044 (O_2044,N_19914,N_19895);
nand UO_2045 (O_2045,N_19969,N_19881);
and UO_2046 (O_2046,N_19971,N_19911);
xor UO_2047 (O_2047,N_19841,N_19907);
nand UO_2048 (O_2048,N_19906,N_19951);
xnor UO_2049 (O_2049,N_19981,N_19923);
or UO_2050 (O_2050,N_19925,N_19841);
or UO_2051 (O_2051,N_19869,N_19946);
nand UO_2052 (O_2052,N_19983,N_19885);
nor UO_2053 (O_2053,N_19875,N_19940);
and UO_2054 (O_2054,N_19931,N_19954);
xnor UO_2055 (O_2055,N_19991,N_19904);
xor UO_2056 (O_2056,N_19925,N_19879);
nor UO_2057 (O_2057,N_19925,N_19869);
xnor UO_2058 (O_2058,N_19950,N_19868);
xor UO_2059 (O_2059,N_19988,N_19910);
nand UO_2060 (O_2060,N_19842,N_19918);
xor UO_2061 (O_2061,N_19853,N_19888);
nand UO_2062 (O_2062,N_19872,N_19916);
nand UO_2063 (O_2063,N_19926,N_19900);
and UO_2064 (O_2064,N_19913,N_19986);
or UO_2065 (O_2065,N_19984,N_19960);
nor UO_2066 (O_2066,N_19865,N_19840);
nor UO_2067 (O_2067,N_19944,N_19895);
xnor UO_2068 (O_2068,N_19917,N_19910);
nand UO_2069 (O_2069,N_19953,N_19919);
or UO_2070 (O_2070,N_19894,N_19926);
or UO_2071 (O_2071,N_19901,N_19866);
and UO_2072 (O_2072,N_19859,N_19851);
and UO_2073 (O_2073,N_19879,N_19916);
nand UO_2074 (O_2074,N_19996,N_19924);
or UO_2075 (O_2075,N_19883,N_19891);
nand UO_2076 (O_2076,N_19883,N_19874);
or UO_2077 (O_2077,N_19970,N_19931);
nand UO_2078 (O_2078,N_19843,N_19882);
nand UO_2079 (O_2079,N_19922,N_19957);
or UO_2080 (O_2080,N_19984,N_19936);
and UO_2081 (O_2081,N_19917,N_19977);
nand UO_2082 (O_2082,N_19865,N_19981);
nor UO_2083 (O_2083,N_19954,N_19976);
nand UO_2084 (O_2084,N_19845,N_19852);
and UO_2085 (O_2085,N_19848,N_19888);
nand UO_2086 (O_2086,N_19878,N_19890);
or UO_2087 (O_2087,N_19907,N_19895);
xnor UO_2088 (O_2088,N_19846,N_19887);
or UO_2089 (O_2089,N_19881,N_19858);
xnor UO_2090 (O_2090,N_19901,N_19857);
xor UO_2091 (O_2091,N_19996,N_19971);
xnor UO_2092 (O_2092,N_19890,N_19929);
nand UO_2093 (O_2093,N_19946,N_19881);
nand UO_2094 (O_2094,N_19874,N_19935);
or UO_2095 (O_2095,N_19958,N_19864);
nor UO_2096 (O_2096,N_19873,N_19942);
nor UO_2097 (O_2097,N_19971,N_19984);
nand UO_2098 (O_2098,N_19849,N_19931);
and UO_2099 (O_2099,N_19928,N_19952);
nand UO_2100 (O_2100,N_19859,N_19852);
or UO_2101 (O_2101,N_19944,N_19941);
nand UO_2102 (O_2102,N_19962,N_19998);
and UO_2103 (O_2103,N_19909,N_19871);
nor UO_2104 (O_2104,N_19858,N_19956);
nor UO_2105 (O_2105,N_19852,N_19888);
nand UO_2106 (O_2106,N_19854,N_19864);
and UO_2107 (O_2107,N_19927,N_19876);
or UO_2108 (O_2108,N_19938,N_19898);
and UO_2109 (O_2109,N_19936,N_19866);
nor UO_2110 (O_2110,N_19969,N_19983);
and UO_2111 (O_2111,N_19960,N_19959);
or UO_2112 (O_2112,N_19936,N_19852);
and UO_2113 (O_2113,N_19893,N_19907);
or UO_2114 (O_2114,N_19981,N_19983);
nor UO_2115 (O_2115,N_19945,N_19997);
or UO_2116 (O_2116,N_19912,N_19847);
nor UO_2117 (O_2117,N_19890,N_19979);
and UO_2118 (O_2118,N_19872,N_19880);
nor UO_2119 (O_2119,N_19936,N_19964);
nand UO_2120 (O_2120,N_19899,N_19843);
and UO_2121 (O_2121,N_19883,N_19966);
and UO_2122 (O_2122,N_19930,N_19884);
nor UO_2123 (O_2123,N_19996,N_19970);
nor UO_2124 (O_2124,N_19873,N_19865);
xnor UO_2125 (O_2125,N_19871,N_19924);
and UO_2126 (O_2126,N_19960,N_19977);
xnor UO_2127 (O_2127,N_19841,N_19859);
nor UO_2128 (O_2128,N_19865,N_19903);
nor UO_2129 (O_2129,N_19962,N_19860);
nand UO_2130 (O_2130,N_19931,N_19894);
or UO_2131 (O_2131,N_19877,N_19970);
or UO_2132 (O_2132,N_19840,N_19999);
and UO_2133 (O_2133,N_19992,N_19982);
or UO_2134 (O_2134,N_19897,N_19971);
or UO_2135 (O_2135,N_19989,N_19952);
and UO_2136 (O_2136,N_19962,N_19981);
nand UO_2137 (O_2137,N_19860,N_19856);
nor UO_2138 (O_2138,N_19889,N_19884);
or UO_2139 (O_2139,N_19846,N_19941);
nor UO_2140 (O_2140,N_19994,N_19842);
and UO_2141 (O_2141,N_19871,N_19989);
and UO_2142 (O_2142,N_19874,N_19969);
or UO_2143 (O_2143,N_19982,N_19852);
xor UO_2144 (O_2144,N_19967,N_19916);
nor UO_2145 (O_2145,N_19997,N_19877);
and UO_2146 (O_2146,N_19876,N_19970);
and UO_2147 (O_2147,N_19912,N_19855);
or UO_2148 (O_2148,N_19970,N_19930);
xor UO_2149 (O_2149,N_19889,N_19949);
xor UO_2150 (O_2150,N_19996,N_19901);
nor UO_2151 (O_2151,N_19913,N_19858);
or UO_2152 (O_2152,N_19912,N_19945);
nor UO_2153 (O_2153,N_19924,N_19847);
nor UO_2154 (O_2154,N_19913,N_19898);
nor UO_2155 (O_2155,N_19875,N_19971);
nor UO_2156 (O_2156,N_19850,N_19904);
xor UO_2157 (O_2157,N_19917,N_19854);
nand UO_2158 (O_2158,N_19866,N_19975);
or UO_2159 (O_2159,N_19903,N_19891);
or UO_2160 (O_2160,N_19885,N_19936);
or UO_2161 (O_2161,N_19974,N_19864);
and UO_2162 (O_2162,N_19905,N_19987);
nor UO_2163 (O_2163,N_19914,N_19883);
xor UO_2164 (O_2164,N_19889,N_19860);
and UO_2165 (O_2165,N_19933,N_19853);
nand UO_2166 (O_2166,N_19877,N_19851);
and UO_2167 (O_2167,N_19857,N_19912);
xor UO_2168 (O_2168,N_19963,N_19868);
xor UO_2169 (O_2169,N_19951,N_19988);
or UO_2170 (O_2170,N_19962,N_19846);
xor UO_2171 (O_2171,N_19963,N_19947);
xor UO_2172 (O_2172,N_19977,N_19965);
xnor UO_2173 (O_2173,N_19958,N_19971);
and UO_2174 (O_2174,N_19931,N_19857);
nor UO_2175 (O_2175,N_19842,N_19913);
nor UO_2176 (O_2176,N_19948,N_19922);
or UO_2177 (O_2177,N_19907,N_19920);
nor UO_2178 (O_2178,N_19847,N_19946);
and UO_2179 (O_2179,N_19953,N_19883);
and UO_2180 (O_2180,N_19873,N_19862);
or UO_2181 (O_2181,N_19984,N_19993);
nand UO_2182 (O_2182,N_19891,N_19983);
nand UO_2183 (O_2183,N_19947,N_19920);
and UO_2184 (O_2184,N_19912,N_19897);
and UO_2185 (O_2185,N_19972,N_19987);
nor UO_2186 (O_2186,N_19990,N_19951);
nor UO_2187 (O_2187,N_19970,N_19924);
xnor UO_2188 (O_2188,N_19885,N_19989);
or UO_2189 (O_2189,N_19885,N_19897);
xor UO_2190 (O_2190,N_19999,N_19861);
nand UO_2191 (O_2191,N_19978,N_19937);
nor UO_2192 (O_2192,N_19892,N_19867);
and UO_2193 (O_2193,N_19944,N_19930);
nand UO_2194 (O_2194,N_19870,N_19864);
nor UO_2195 (O_2195,N_19879,N_19847);
nor UO_2196 (O_2196,N_19874,N_19967);
nor UO_2197 (O_2197,N_19889,N_19896);
nor UO_2198 (O_2198,N_19899,N_19879);
xnor UO_2199 (O_2199,N_19940,N_19921);
or UO_2200 (O_2200,N_19914,N_19987);
or UO_2201 (O_2201,N_19940,N_19882);
nor UO_2202 (O_2202,N_19840,N_19889);
or UO_2203 (O_2203,N_19930,N_19885);
xor UO_2204 (O_2204,N_19929,N_19855);
nor UO_2205 (O_2205,N_19978,N_19979);
or UO_2206 (O_2206,N_19985,N_19907);
nand UO_2207 (O_2207,N_19957,N_19912);
or UO_2208 (O_2208,N_19871,N_19881);
nand UO_2209 (O_2209,N_19892,N_19873);
nand UO_2210 (O_2210,N_19880,N_19851);
nor UO_2211 (O_2211,N_19854,N_19904);
nor UO_2212 (O_2212,N_19863,N_19962);
nand UO_2213 (O_2213,N_19881,N_19888);
nand UO_2214 (O_2214,N_19853,N_19995);
xnor UO_2215 (O_2215,N_19876,N_19879);
or UO_2216 (O_2216,N_19889,N_19948);
nor UO_2217 (O_2217,N_19987,N_19965);
nor UO_2218 (O_2218,N_19956,N_19871);
or UO_2219 (O_2219,N_19978,N_19900);
nor UO_2220 (O_2220,N_19860,N_19887);
or UO_2221 (O_2221,N_19916,N_19848);
or UO_2222 (O_2222,N_19984,N_19879);
xnor UO_2223 (O_2223,N_19945,N_19852);
xor UO_2224 (O_2224,N_19988,N_19977);
or UO_2225 (O_2225,N_19861,N_19899);
and UO_2226 (O_2226,N_19871,N_19992);
nand UO_2227 (O_2227,N_19881,N_19927);
xor UO_2228 (O_2228,N_19911,N_19944);
nor UO_2229 (O_2229,N_19947,N_19927);
nand UO_2230 (O_2230,N_19876,N_19882);
xor UO_2231 (O_2231,N_19902,N_19900);
xnor UO_2232 (O_2232,N_19937,N_19858);
xor UO_2233 (O_2233,N_19846,N_19871);
xnor UO_2234 (O_2234,N_19901,N_19884);
xnor UO_2235 (O_2235,N_19999,N_19961);
nor UO_2236 (O_2236,N_19924,N_19869);
nand UO_2237 (O_2237,N_19875,N_19868);
and UO_2238 (O_2238,N_19943,N_19891);
or UO_2239 (O_2239,N_19981,N_19987);
or UO_2240 (O_2240,N_19989,N_19976);
or UO_2241 (O_2241,N_19868,N_19948);
and UO_2242 (O_2242,N_19872,N_19857);
and UO_2243 (O_2243,N_19908,N_19900);
nand UO_2244 (O_2244,N_19913,N_19897);
nand UO_2245 (O_2245,N_19876,N_19858);
and UO_2246 (O_2246,N_19984,N_19991);
xnor UO_2247 (O_2247,N_19913,N_19940);
nor UO_2248 (O_2248,N_19937,N_19973);
xnor UO_2249 (O_2249,N_19932,N_19871);
and UO_2250 (O_2250,N_19926,N_19850);
xnor UO_2251 (O_2251,N_19939,N_19846);
xor UO_2252 (O_2252,N_19938,N_19866);
xor UO_2253 (O_2253,N_19930,N_19849);
xor UO_2254 (O_2254,N_19877,N_19894);
nand UO_2255 (O_2255,N_19936,N_19903);
and UO_2256 (O_2256,N_19879,N_19950);
and UO_2257 (O_2257,N_19927,N_19922);
nor UO_2258 (O_2258,N_19872,N_19982);
xnor UO_2259 (O_2259,N_19990,N_19955);
and UO_2260 (O_2260,N_19988,N_19957);
or UO_2261 (O_2261,N_19841,N_19867);
nor UO_2262 (O_2262,N_19897,N_19875);
and UO_2263 (O_2263,N_19918,N_19921);
nand UO_2264 (O_2264,N_19962,N_19939);
xor UO_2265 (O_2265,N_19863,N_19986);
or UO_2266 (O_2266,N_19859,N_19947);
xnor UO_2267 (O_2267,N_19990,N_19867);
or UO_2268 (O_2268,N_19903,N_19866);
xnor UO_2269 (O_2269,N_19879,N_19867);
or UO_2270 (O_2270,N_19949,N_19932);
nand UO_2271 (O_2271,N_19904,N_19880);
nor UO_2272 (O_2272,N_19901,N_19922);
or UO_2273 (O_2273,N_19983,N_19980);
nor UO_2274 (O_2274,N_19904,N_19872);
xor UO_2275 (O_2275,N_19910,N_19896);
or UO_2276 (O_2276,N_19882,N_19953);
nor UO_2277 (O_2277,N_19935,N_19972);
xor UO_2278 (O_2278,N_19955,N_19964);
and UO_2279 (O_2279,N_19962,N_19874);
and UO_2280 (O_2280,N_19849,N_19864);
xor UO_2281 (O_2281,N_19880,N_19992);
and UO_2282 (O_2282,N_19989,N_19875);
nand UO_2283 (O_2283,N_19934,N_19943);
or UO_2284 (O_2284,N_19979,N_19861);
nor UO_2285 (O_2285,N_19997,N_19879);
xor UO_2286 (O_2286,N_19995,N_19999);
nor UO_2287 (O_2287,N_19903,N_19871);
nor UO_2288 (O_2288,N_19937,N_19946);
or UO_2289 (O_2289,N_19996,N_19908);
or UO_2290 (O_2290,N_19893,N_19949);
nor UO_2291 (O_2291,N_19880,N_19917);
nand UO_2292 (O_2292,N_19898,N_19925);
and UO_2293 (O_2293,N_19908,N_19898);
nor UO_2294 (O_2294,N_19953,N_19887);
and UO_2295 (O_2295,N_19983,N_19958);
or UO_2296 (O_2296,N_19971,N_19924);
and UO_2297 (O_2297,N_19887,N_19972);
xor UO_2298 (O_2298,N_19866,N_19935);
nand UO_2299 (O_2299,N_19970,N_19928);
or UO_2300 (O_2300,N_19861,N_19930);
xnor UO_2301 (O_2301,N_19972,N_19954);
xor UO_2302 (O_2302,N_19880,N_19976);
and UO_2303 (O_2303,N_19880,N_19949);
or UO_2304 (O_2304,N_19876,N_19875);
or UO_2305 (O_2305,N_19991,N_19975);
or UO_2306 (O_2306,N_19922,N_19996);
nand UO_2307 (O_2307,N_19952,N_19950);
xnor UO_2308 (O_2308,N_19851,N_19865);
xnor UO_2309 (O_2309,N_19980,N_19893);
xnor UO_2310 (O_2310,N_19961,N_19902);
or UO_2311 (O_2311,N_19899,N_19842);
nor UO_2312 (O_2312,N_19847,N_19867);
nor UO_2313 (O_2313,N_19958,N_19920);
nand UO_2314 (O_2314,N_19955,N_19865);
nor UO_2315 (O_2315,N_19932,N_19865);
or UO_2316 (O_2316,N_19978,N_19977);
nor UO_2317 (O_2317,N_19918,N_19851);
xnor UO_2318 (O_2318,N_19948,N_19872);
nor UO_2319 (O_2319,N_19973,N_19938);
and UO_2320 (O_2320,N_19972,N_19957);
or UO_2321 (O_2321,N_19902,N_19862);
xor UO_2322 (O_2322,N_19906,N_19933);
nand UO_2323 (O_2323,N_19966,N_19991);
and UO_2324 (O_2324,N_19936,N_19847);
and UO_2325 (O_2325,N_19992,N_19957);
nand UO_2326 (O_2326,N_19854,N_19972);
nand UO_2327 (O_2327,N_19994,N_19876);
nor UO_2328 (O_2328,N_19850,N_19953);
xor UO_2329 (O_2329,N_19891,N_19860);
nand UO_2330 (O_2330,N_19920,N_19902);
or UO_2331 (O_2331,N_19999,N_19949);
and UO_2332 (O_2332,N_19881,N_19985);
and UO_2333 (O_2333,N_19851,N_19846);
nand UO_2334 (O_2334,N_19866,N_19894);
and UO_2335 (O_2335,N_19934,N_19977);
or UO_2336 (O_2336,N_19881,N_19849);
nor UO_2337 (O_2337,N_19916,N_19844);
and UO_2338 (O_2338,N_19963,N_19968);
nand UO_2339 (O_2339,N_19960,N_19894);
nand UO_2340 (O_2340,N_19948,N_19957);
or UO_2341 (O_2341,N_19996,N_19857);
xnor UO_2342 (O_2342,N_19916,N_19846);
and UO_2343 (O_2343,N_19890,N_19941);
nand UO_2344 (O_2344,N_19969,N_19892);
xnor UO_2345 (O_2345,N_19986,N_19867);
xor UO_2346 (O_2346,N_19977,N_19893);
nand UO_2347 (O_2347,N_19991,N_19852);
nor UO_2348 (O_2348,N_19914,N_19862);
or UO_2349 (O_2349,N_19997,N_19887);
xor UO_2350 (O_2350,N_19991,N_19892);
nor UO_2351 (O_2351,N_19848,N_19932);
nand UO_2352 (O_2352,N_19931,N_19968);
nand UO_2353 (O_2353,N_19895,N_19929);
nand UO_2354 (O_2354,N_19995,N_19852);
xor UO_2355 (O_2355,N_19917,N_19894);
xnor UO_2356 (O_2356,N_19955,N_19992);
xor UO_2357 (O_2357,N_19888,N_19937);
xnor UO_2358 (O_2358,N_19878,N_19861);
xor UO_2359 (O_2359,N_19954,N_19891);
nand UO_2360 (O_2360,N_19988,N_19923);
or UO_2361 (O_2361,N_19923,N_19896);
nor UO_2362 (O_2362,N_19905,N_19878);
and UO_2363 (O_2363,N_19891,N_19856);
nor UO_2364 (O_2364,N_19847,N_19845);
xor UO_2365 (O_2365,N_19938,N_19997);
or UO_2366 (O_2366,N_19860,N_19904);
or UO_2367 (O_2367,N_19883,N_19849);
nor UO_2368 (O_2368,N_19851,N_19942);
or UO_2369 (O_2369,N_19918,N_19849);
and UO_2370 (O_2370,N_19867,N_19934);
and UO_2371 (O_2371,N_19977,N_19910);
xnor UO_2372 (O_2372,N_19948,N_19917);
or UO_2373 (O_2373,N_19867,N_19974);
nand UO_2374 (O_2374,N_19959,N_19872);
nand UO_2375 (O_2375,N_19870,N_19840);
nor UO_2376 (O_2376,N_19841,N_19927);
or UO_2377 (O_2377,N_19937,N_19911);
nor UO_2378 (O_2378,N_19864,N_19844);
and UO_2379 (O_2379,N_19994,N_19867);
nor UO_2380 (O_2380,N_19886,N_19957);
or UO_2381 (O_2381,N_19915,N_19976);
nor UO_2382 (O_2382,N_19890,N_19983);
nor UO_2383 (O_2383,N_19989,N_19939);
or UO_2384 (O_2384,N_19888,N_19955);
nand UO_2385 (O_2385,N_19913,N_19927);
nand UO_2386 (O_2386,N_19908,N_19850);
xor UO_2387 (O_2387,N_19961,N_19948);
or UO_2388 (O_2388,N_19987,N_19995);
xor UO_2389 (O_2389,N_19902,N_19942);
or UO_2390 (O_2390,N_19932,N_19857);
and UO_2391 (O_2391,N_19977,N_19950);
or UO_2392 (O_2392,N_19909,N_19869);
and UO_2393 (O_2393,N_19934,N_19857);
xnor UO_2394 (O_2394,N_19855,N_19940);
xnor UO_2395 (O_2395,N_19873,N_19955);
and UO_2396 (O_2396,N_19864,N_19882);
and UO_2397 (O_2397,N_19903,N_19911);
or UO_2398 (O_2398,N_19959,N_19995);
or UO_2399 (O_2399,N_19968,N_19934);
nor UO_2400 (O_2400,N_19942,N_19892);
nor UO_2401 (O_2401,N_19980,N_19857);
and UO_2402 (O_2402,N_19880,N_19963);
or UO_2403 (O_2403,N_19952,N_19843);
nor UO_2404 (O_2404,N_19963,N_19877);
nand UO_2405 (O_2405,N_19844,N_19988);
or UO_2406 (O_2406,N_19982,N_19890);
and UO_2407 (O_2407,N_19886,N_19880);
xnor UO_2408 (O_2408,N_19976,N_19965);
xnor UO_2409 (O_2409,N_19951,N_19929);
and UO_2410 (O_2410,N_19987,N_19885);
and UO_2411 (O_2411,N_19888,N_19948);
xnor UO_2412 (O_2412,N_19880,N_19998);
nor UO_2413 (O_2413,N_19899,N_19998);
nor UO_2414 (O_2414,N_19951,N_19992);
xnor UO_2415 (O_2415,N_19849,N_19950);
nand UO_2416 (O_2416,N_19914,N_19975);
xnor UO_2417 (O_2417,N_19992,N_19910);
nand UO_2418 (O_2418,N_19946,N_19990);
nor UO_2419 (O_2419,N_19941,N_19851);
and UO_2420 (O_2420,N_19849,N_19867);
or UO_2421 (O_2421,N_19960,N_19924);
nor UO_2422 (O_2422,N_19895,N_19854);
nand UO_2423 (O_2423,N_19869,N_19892);
nand UO_2424 (O_2424,N_19991,N_19914);
and UO_2425 (O_2425,N_19860,N_19938);
xnor UO_2426 (O_2426,N_19902,N_19944);
and UO_2427 (O_2427,N_19843,N_19877);
nand UO_2428 (O_2428,N_19873,N_19891);
and UO_2429 (O_2429,N_19860,N_19945);
nor UO_2430 (O_2430,N_19857,N_19925);
xnor UO_2431 (O_2431,N_19872,N_19900);
xnor UO_2432 (O_2432,N_19962,N_19976);
and UO_2433 (O_2433,N_19979,N_19847);
and UO_2434 (O_2434,N_19882,N_19937);
nor UO_2435 (O_2435,N_19918,N_19936);
or UO_2436 (O_2436,N_19974,N_19995);
nor UO_2437 (O_2437,N_19928,N_19969);
xnor UO_2438 (O_2438,N_19968,N_19918);
nor UO_2439 (O_2439,N_19922,N_19923);
or UO_2440 (O_2440,N_19965,N_19887);
or UO_2441 (O_2441,N_19941,N_19931);
or UO_2442 (O_2442,N_19857,N_19871);
nor UO_2443 (O_2443,N_19853,N_19851);
and UO_2444 (O_2444,N_19974,N_19915);
xor UO_2445 (O_2445,N_19953,N_19936);
and UO_2446 (O_2446,N_19918,N_19926);
nand UO_2447 (O_2447,N_19994,N_19931);
or UO_2448 (O_2448,N_19903,N_19933);
nor UO_2449 (O_2449,N_19938,N_19862);
or UO_2450 (O_2450,N_19979,N_19956);
xnor UO_2451 (O_2451,N_19976,N_19927);
or UO_2452 (O_2452,N_19916,N_19882);
nand UO_2453 (O_2453,N_19865,N_19928);
and UO_2454 (O_2454,N_19886,N_19925);
and UO_2455 (O_2455,N_19967,N_19868);
or UO_2456 (O_2456,N_19976,N_19926);
nand UO_2457 (O_2457,N_19955,N_19907);
and UO_2458 (O_2458,N_19952,N_19870);
nand UO_2459 (O_2459,N_19935,N_19976);
or UO_2460 (O_2460,N_19940,N_19845);
and UO_2461 (O_2461,N_19938,N_19994);
nand UO_2462 (O_2462,N_19960,N_19925);
nand UO_2463 (O_2463,N_19887,N_19938);
or UO_2464 (O_2464,N_19946,N_19840);
nor UO_2465 (O_2465,N_19971,N_19952);
nand UO_2466 (O_2466,N_19924,N_19972);
or UO_2467 (O_2467,N_19994,N_19855);
nor UO_2468 (O_2468,N_19970,N_19965);
nand UO_2469 (O_2469,N_19998,N_19938);
nor UO_2470 (O_2470,N_19875,N_19938);
xor UO_2471 (O_2471,N_19857,N_19955);
and UO_2472 (O_2472,N_19847,N_19868);
xor UO_2473 (O_2473,N_19866,N_19973);
nor UO_2474 (O_2474,N_19852,N_19907);
xnor UO_2475 (O_2475,N_19987,N_19930);
nand UO_2476 (O_2476,N_19902,N_19924);
and UO_2477 (O_2477,N_19982,N_19918);
nand UO_2478 (O_2478,N_19850,N_19905);
xor UO_2479 (O_2479,N_19974,N_19866);
xor UO_2480 (O_2480,N_19941,N_19910);
xnor UO_2481 (O_2481,N_19910,N_19911);
or UO_2482 (O_2482,N_19998,N_19878);
nor UO_2483 (O_2483,N_19870,N_19979);
or UO_2484 (O_2484,N_19878,N_19867);
xnor UO_2485 (O_2485,N_19924,N_19905);
and UO_2486 (O_2486,N_19994,N_19900);
nor UO_2487 (O_2487,N_19911,N_19987);
nand UO_2488 (O_2488,N_19855,N_19842);
nand UO_2489 (O_2489,N_19917,N_19949);
nand UO_2490 (O_2490,N_19901,N_19907);
nand UO_2491 (O_2491,N_19870,N_19995);
and UO_2492 (O_2492,N_19982,N_19950);
nor UO_2493 (O_2493,N_19866,N_19913);
xnor UO_2494 (O_2494,N_19945,N_19917);
nor UO_2495 (O_2495,N_19885,N_19985);
and UO_2496 (O_2496,N_19840,N_19922);
xor UO_2497 (O_2497,N_19984,N_19913);
and UO_2498 (O_2498,N_19969,N_19840);
and UO_2499 (O_2499,N_19992,N_19935);
endmodule