module basic_500_3000_500_6_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_371,In_403);
and U1 (N_1,In_219,In_389);
xor U2 (N_2,In_245,In_373);
or U3 (N_3,In_137,In_125);
or U4 (N_4,In_187,In_301);
and U5 (N_5,In_40,In_101);
or U6 (N_6,In_434,In_383);
and U7 (N_7,In_406,In_188);
nand U8 (N_8,In_430,In_499);
nor U9 (N_9,In_378,In_443);
nand U10 (N_10,In_248,In_449);
nor U11 (N_11,In_362,In_484);
or U12 (N_12,In_237,In_220);
nor U13 (N_13,In_165,In_151);
nand U14 (N_14,In_10,In_441);
or U15 (N_15,In_316,In_61);
xor U16 (N_16,In_428,In_25);
nor U17 (N_17,In_281,In_416);
or U18 (N_18,In_217,In_154);
nand U19 (N_19,In_257,In_177);
and U20 (N_20,In_70,In_111);
and U21 (N_21,In_410,In_213);
or U22 (N_22,In_110,In_183);
or U23 (N_23,In_493,In_247);
nor U24 (N_24,In_469,In_81);
nor U25 (N_25,In_307,In_8);
or U26 (N_26,In_22,In_481);
and U27 (N_27,In_216,In_421);
or U28 (N_28,In_381,In_181);
and U29 (N_29,In_2,In_471);
nand U30 (N_30,In_205,In_162);
or U31 (N_31,In_84,In_190);
or U32 (N_32,In_118,In_488);
and U33 (N_33,In_38,In_114);
nor U34 (N_34,In_132,In_21);
nor U35 (N_35,In_436,In_20);
nor U36 (N_36,In_201,In_223);
and U37 (N_37,In_34,In_360);
nor U38 (N_38,In_108,In_292);
or U39 (N_39,In_282,In_455);
nor U40 (N_40,In_66,In_355);
or U41 (N_41,In_6,In_277);
nor U42 (N_42,In_429,In_51);
nand U43 (N_43,In_147,In_310);
nor U44 (N_44,In_446,In_106);
and U45 (N_45,In_340,In_149);
and U46 (N_46,In_184,In_57);
nor U47 (N_47,In_475,In_172);
nand U48 (N_48,In_329,In_414);
xor U49 (N_49,In_143,In_322);
xor U50 (N_50,In_180,In_45);
and U51 (N_51,In_327,In_46);
xor U52 (N_52,In_18,In_209);
nand U53 (N_53,In_269,In_227);
nor U54 (N_54,In_144,In_130);
nand U55 (N_55,In_454,In_466);
or U56 (N_56,In_325,In_343);
and U57 (N_57,In_226,In_13);
or U58 (N_58,In_192,In_287);
or U59 (N_59,In_126,In_391);
or U60 (N_60,In_11,In_313);
nor U61 (N_61,In_356,In_109);
nor U62 (N_62,In_342,In_120);
and U63 (N_63,In_480,In_367);
nand U64 (N_64,In_402,In_439);
nor U65 (N_65,In_370,In_385);
nor U66 (N_66,In_59,In_175);
nand U67 (N_67,In_255,In_453);
nand U68 (N_68,In_167,In_233);
and U69 (N_69,In_314,In_401);
nand U70 (N_70,In_423,In_275);
xnor U71 (N_71,In_358,In_462);
or U72 (N_72,In_200,In_95);
or U73 (N_73,In_107,In_256);
or U74 (N_74,In_212,In_295);
nor U75 (N_75,In_250,In_56);
or U76 (N_76,In_341,In_43);
and U77 (N_77,In_468,In_335);
nand U78 (N_78,In_16,In_196);
and U79 (N_79,In_451,In_85);
nand U80 (N_80,In_230,In_78);
nor U81 (N_81,In_288,In_131);
nand U82 (N_82,In_231,In_452);
and U83 (N_83,In_148,In_496);
and U84 (N_84,In_267,In_67);
nand U85 (N_85,In_89,In_311);
nor U86 (N_86,In_419,In_376);
nand U87 (N_87,In_17,In_160);
nor U88 (N_88,In_29,In_404);
or U89 (N_89,In_459,In_235);
or U90 (N_90,In_321,In_435);
and U91 (N_91,In_203,In_208);
nor U92 (N_92,In_418,In_1);
xnor U93 (N_93,In_15,In_444);
nand U94 (N_94,In_409,In_79);
xnor U95 (N_95,In_482,In_413);
or U96 (N_96,In_478,In_306);
or U97 (N_97,In_420,In_479);
or U98 (N_98,In_238,In_398);
nor U99 (N_99,In_41,In_39);
or U100 (N_100,In_344,In_476);
and U101 (N_101,In_19,In_268);
and U102 (N_102,In_374,In_372);
nor U103 (N_103,In_347,In_54);
or U104 (N_104,In_179,In_457);
nand U105 (N_105,In_387,In_133);
nor U106 (N_106,In_204,In_477);
nand U107 (N_107,In_442,In_396);
xor U108 (N_108,In_100,In_461);
nand U109 (N_109,In_332,In_166);
nand U110 (N_110,In_136,In_395);
or U111 (N_111,In_379,In_221);
nor U112 (N_112,In_12,In_49);
or U113 (N_113,In_470,In_198);
nand U114 (N_114,In_112,In_243);
nor U115 (N_115,In_252,In_440);
and U116 (N_116,In_189,In_486);
nor U117 (N_117,In_432,In_337);
and U118 (N_118,In_463,In_97);
nand U119 (N_119,In_393,In_353);
nor U120 (N_120,In_318,In_135);
xor U121 (N_121,In_73,In_244);
nand U122 (N_122,In_339,In_119);
and U123 (N_123,In_44,In_76);
nand U124 (N_124,In_465,In_173);
or U125 (N_125,In_142,In_88);
nand U126 (N_126,In_156,In_246);
nor U127 (N_127,In_124,In_102);
and U128 (N_128,In_346,In_7);
and U129 (N_129,In_87,In_309);
nor U130 (N_130,In_324,In_489);
nor U131 (N_131,In_146,In_152);
nor U132 (N_132,In_384,In_283);
nand U133 (N_133,In_30,In_53);
xnor U134 (N_134,In_261,In_333);
xnor U135 (N_135,In_141,In_169);
nand U136 (N_136,In_308,In_123);
and U137 (N_137,In_116,In_299);
nor U138 (N_138,In_357,In_456);
nand U139 (N_139,In_433,In_225);
or U140 (N_140,In_417,In_364);
nand U141 (N_141,In_350,In_359);
nor U142 (N_142,In_305,In_186);
nor U143 (N_143,In_161,In_315);
nor U144 (N_144,In_498,In_265);
and U145 (N_145,In_474,In_422);
and U146 (N_146,In_0,In_278);
nand U147 (N_147,In_331,In_338);
nor U148 (N_148,In_42,In_351);
and U149 (N_149,In_249,In_199);
and U150 (N_150,In_182,In_460);
xnor U151 (N_151,In_258,In_276);
or U152 (N_152,In_211,In_127);
or U153 (N_153,In_37,In_157);
and U154 (N_154,In_241,In_155);
nand U155 (N_155,In_363,In_103);
or U156 (N_156,In_392,In_289);
or U157 (N_157,In_5,In_28);
or U158 (N_158,In_382,In_60);
and U159 (N_159,In_407,In_467);
nor U160 (N_160,In_77,In_80);
nor U161 (N_161,In_485,In_214);
xnor U162 (N_162,In_266,In_386);
and U163 (N_163,In_83,In_352);
and U164 (N_164,In_96,In_72);
or U165 (N_165,In_236,In_336);
nand U166 (N_166,In_450,In_345);
or U167 (N_167,In_494,In_272);
nor U168 (N_168,In_368,In_239);
and U169 (N_169,In_113,In_458);
nand U170 (N_170,In_328,In_424);
nand U171 (N_171,In_411,In_264);
and U172 (N_172,In_437,In_464);
or U173 (N_173,In_399,In_296);
nor U174 (N_174,In_279,In_293);
nor U175 (N_175,In_490,In_23);
nor U176 (N_176,In_425,In_202);
nor U177 (N_177,In_242,In_27);
nand U178 (N_178,In_326,In_491);
nand U179 (N_179,In_117,In_286);
nor U180 (N_180,In_291,In_145);
or U181 (N_181,In_64,In_317);
nor U182 (N_182,In_426,In_365);
and U183 (N_183,In_104,In_193);
nand U184 (N_184,In_487,In_153);
and U185 (N_185,In_388,In_302);
and U186 (N_186,In_207,In_290);
and U187 (N_187,In_191,In_138);
nand U188 (N_188,In_380,In_115);
nand U189 (N_189,In_140,In_298);
or U190 (N_190,In_24,In_473);
nor U191 (N_191,In_32,In_3);
nor U192 (N_192,In_285,In_90);
and U193 (N_193,In_284,In_98);
or U194 (N_194,In_312,In_63);
nand U195 (N_195,In_320,In_222);
nand U196 (N_196,In_369,In_129);
and U197 (N_197,In_259,In_4);
xnor U198 (N_198,In_262,In_210);
or U199 (N_199,In_472,In_497);
and U200 (N_200,In_68,In_50);
or U201 (N_201,In_297,In_178);
and U202 (N_202,In_349,In_122);
or U203 (N_203,In_150,In_170);
nor U204 (N_204,In_224,In_300);
and U205 (N_205,In_323,In_93);
nor U206 (N_206,In_412,In_215);
and U207 (N_207,In_397,In_58);
or U208 (N_208,In_400,In_159);
and U209 (N_209,In_240,In_31);
or U210 (N_210,In_168,In_228);
and U211 (N_211,In_74,In_82);
nor U212 (N_212,In_394,In_495);
or U213 (N_213,In_94,In_354);
nand U214 (N_214,In_253,In_330);
nor U215 (N_215,In_105,In_377);
nor U216 (N_216,In_36,In_438);
and U217 (N_217,In_415,In_251);
or U218 (N_218,In_304,In_448);
or U219 (N_219,In_405,In_280);
nand U220 (N_220,In_195,In_128);
or U221 (N_221,In_75,In_62);
nor U222 (N_222,In_92,In_134);
and U223 (N_223,In_445,In_270);
and U224 (N_224,In_91,In_319);
nor U225 (N_225,In_232,In_206);
and U226 (N_226,In_273,In_303);
nand U227 (N_227,In_158,In_274);
or U228 (N_228,In_163,In_99);
or U229 (N_229,In_234,In_174);
and U230 (N_230,In_9,In_48);
nand U231 (N_231,In_35,In_194);
nor U232 (N_232,In_431,In_176);
nor U233 (N_233,In_47,In_348);
nand U234 (N_234,In_33,In_14);
nor U235 (N_235,In_171,In_254);
nor U236 (N_236,In_483,In_334);
or U237 (N_237,In_69,In_447);
nor U238 (N_238,In_52,In_26);
or U239 (N_239,In_65,In_390);
and U240 (N_240,In_361,In_294);
nand U241 (N_241,In_366,In_263);
nor U242 (N_242,In_427,In_164);
and U243 (N_243,In_218,In_260);
and U244 (N_244,In_121,In_375);
nand U245 (N_245,In_197,In_55);
nand U246 (N_246,In_229,In_492);
nand U247 (N_247,In_86,In_408);
and U248 (N_248,In_271,In_71);
and U249 (N_249,In_139,In_185);
nand U250 (N_250,In_82,In_37);
nand U251 (N_251,In_148,In_58);
xnor U252 (N_252,In_421,In_387);
nand U253 (N_253,In_95,In_348);
nand U254 (N_254,In_79,In_387);
and U255 (N_255,In_288,In_493);
and U256 (N_256,In_85,In_336);
nand U257 (N_257,In_119,In_231);
nor U258 (N_258,In_45,In_194);
nor U259 (N_259,In_15,In_225);
nand U260 (N_260,In_63,In_396);
nand U261 (N_261,In_449,In_120);
nor U262 (N_262,In_458,In_103);
nor U263 (N_263,In_282,In_201);
nor U264 (N_264,In_95,In_181);
and U265 (N_265,In_15,In_354);
nand U266 (N_266,In_358,In_250);
and U267 (N_267,In_320,In_181);
nor U268 (N_268,In_465,In_471);
nand U269 (N_269,In_299,In_312);
nand U270 (N_270,In_319,In_432);
nor U271 (N_271,In_376,In_109);
nand U272 (N_272,In_499,In_285);
nand U273 (N_273,In_433,In_47);
nor U274 (N_274,In_339,In_229);
nor U275 (N_275,In_341,In_165);
nand U276 (N_276,In_440,In_25);
or U277 (N_277,In_135,In_2);
and U278 (N_278,In_485,In_314);
and U279 (N_279,In_323,In_412);
nand U280 (N_280,In_70,In_434);
nor U281 (N_281,In_485,In_370);
nor U282 (N_282,In_122,In_138);
nor U283 (N_283,In_32,In_59);
nor U284 (N_284,In_67,In_397);
nor U285 (N_285,In_479,In_394);
and U286 (N_286,In_107,In_110);
nand U287 (N_287,In_35,In_5);
or U288 (N_288,In_122,In_401);
nand U289 (N_289,In_68,In_391);
nor U290 (N_290,In_82,In_212);
or U291 (N_291,In_97,In_200);
nand U292 (N_292,In_438,In_184);
or U293 (N_293,In_265,In_475);
nor U294 (N_294,In_208,In_405);
or U295 (N_295,In_122,In_205);
or U296 (N_296,In_59,In_229);
nand U297 (N_297,In_419,In_490);
nand U298 (N_298,In_36,In_245);
nor U299 (N_299,In_98,In_335);
nand U300 (N_300,In_337,In_52);
nor U301 (N_301,In_198,In_261);
nand U302 (N_302,In_43,In_395);
and U303 (N_303,In_151,In_195);
nand U304 (N_304,In_450,In_93);
and U305 (N_305,In_33,In_107);
and U306 (N_306,In_301,In_357);
nor U307 (N_307,In_326,In_302);
nor U308 (N_308,In_63,In_479);
and U309 (N_309,In_315,In_336);
nor U310 (N_310,In_372,In_496);
nand U311 (N_311,In_88,In_141);
nor U312 (N_312,In_255,In_239);
or U313 (N_313,In_377,In_250);
or U314 (N_314,In_278,In_471);
nand U315 (N_315,In_453,In_383);
and U316 (N_316,In_15,In_138);
and U317 (N_317,In_453,In_231);
nor U318 (N_318,In_62,In_100);
or U319 (N_319,In_297,In_305);
or U320 (N_320,In_260,In_450);
or U321 (N_321,In_311,In_384);
nand U322 (N_322,In_197,In_396);
nand U323 (N_323,In_449,In_466);
or U324 (N_324,In_294,In_175);
and U325 (N_325,In_27,In_195);
nand U326 (N_326,In_365,In_275);
or U327 (N_327,In_62,In_199);
nor U328 (N_328,In_360,In_201);
and U329 (N_329,In_381,In_38);
and U330 (N_330,In_55,In_133);
nand U331 (N_331,In_29,In_85);
nand U332 (N_332,In_19,In_393);
or U333 (N_333,In_196,In_341);
nand U334 (N_334,In_321,In_394);
and U335 (N_335,In_93,In_176);
nand U336 (N_336,In_179,In_255);
nand U337 (N_337,In_210,In_292);
or U338 (N_338,In_450,In_296);
nand U339 (N_339,In_313,In_244);
or U340 (N_340,In_84,In_267);
nand U341 (N_341,In_265,In_39);
or U342 (N_342,In_357,In_398);
or U343 (N_343,In_475,In_72);
or U344 (N_344,In_320,In_377);
xnor U345 (N_345,In_199,In_293);
nand U346 (N_346,In_403,In_163);
or U347 (N_347,In_102,In_290);
and U348 (N_348,In_15,In_410);
and U349 (N_349,In_334,In_104);
nor U350 (N_350,In_239,In_55);
or U351 (N_351,In_14,In_470);
xor U352 (N_352,In_298,In_356);
nand U353 (N_353,In_55,In_311);
xor U354 (N_354,In_9,In_95);
and U355 (N_355,In_371,In_192);
and U356 (N_356,In_85,In_171);
nor U357 (N_357,In_168,In_42);
nand U358 (N_358,In_328,In_195);
or U359 (N_359,In_340,In_239);
nor U360 (N_360,In_157,In_195);
nor U361 (N_361,In_401,In_319);
and U362 (N_362,In_386,In_186);
and U363 (N_363,In_76,In_116);
nor U364 (N_364,In_376,In_224);
nor U365 (N_365,In_345,In_298);
xnor U366 (N_366,In_121,In_236);
or U367 (N_367,In_244,In_326);
and U368 (N_368,In_259,In_63);
or U369 (N_369,In_91,In_259);
or U370 (N_370,In_0,In_461);
or U371 (N_371,In_286,In_470);
or U372 (N_372,In_302,In_403);
or U373 (N_373,In_203,In_481);
or U374 (N_374,In_404,In_347);
nand U375 (N_375,In_23,In_447);
or U376 (N_376,In_290,In_259);
or U377 (N_377,In_289,In_212);
nor U378 (N_378,In_113,In_89);
nand U379 (N_379,In_239,In_96);
nand U380 (N_380,In_38,In_174);
and U381 (N_381,In_233,In_467);
nor U382 (N_382,In_480,In_365);
or U383 (N_383,In_9,In_197);
or U384 (N_384,In_7,In_41);
nand U385 (N_385,In_159,In_299);
nand U386 (N_386,In_356,In_402);
or U387 (N_387,In_203,In_277);
and U388 (N_388,In_426,In_177);
or U389 (N_389,In_207,In_428);
nor U390 (N_390,In_49,In_68);
or U391 (N_391,In_341,In_290);
nor U392 (N_392,In_278,In_179);
and U393 (N_393,In_91,In_295);
nand U394 (N_394,In_135,In_485);
and U395 (N_395,In_122,In_209);
and U396 (N_396,In_44,In_465);
nand U397 (N_397,In_445,In_114);
xor U398 (N_398,In_387,In_32);
nand U399 (N_399,In_133,In_94);
nand U400 (N_400,In_372,In_215);
and U401 (N_401,In_288,In_225);
or U402 (N_402,In_166,In_211);
and U403 (N_403,In_122,In_100);
nor U404 (N_404,In_185,In_406);
and U405 (N_405,In_203,In_272);
or U406 (N_406,In_363,In_72);
or U407 (N_407,In_426,In_87);
nor U408 (N_408,In_334,In_70);
and U409 (N_409,In_401,In_47);
nand U410 (N_410,In_281,In_90);
nand U411 (N_411,In_152,In_341);
and U412 (N_412,In_298,In_324);
or U413 (N_413,In_387,In_86);
nor U414 (N_414,In_274,In_152);
and U415 (N_415,In_25,In_23);
nand U416 (N_416,In_277,In_213);
and U417 (N_417,In_417,In_34);
nor U418 (N_418,In_356,In_451);
nor U419 (N_419,In_202,In_349);
nand U420 (N_420,In_105,In_129);
nand U421 (N_421,In_66,In_202);
and U422 (N_422,In_365,In_273);
and U423 (N_423,In_440,In_476);
or U424 (N_424,In_282,In_253);
nand U425 (N_425,In_291,In_101);
and U426 (N_426,In_266,In_23);
or U427 (N_427,In_239,In_359);
and U428 (N_428,In_344,In_349);
or U429 (N_429,In_234,In_462);
nor U430 (N_430,In_89,In_185);
nor U431 (N_431,In_311,In_215);
and U432 (N_432,In_208,In_25);
nand U433 (N_433,In_127,In_224);
or U434 (N_434,In_79,In_21);
nand U435 (N_435,In_491,In_8);
or U436 (N_436,In_145,In_209);
nor U437 (N_437,In_260,In_163);
and U438 (N_438,In_275,In_394);
nand U439 (N_439,In_417,In_24);
nand U440 (N_440,In_12,In_336);
or U441 (N_441,In_54,In_384);
nand U442 (N_442,In_241,In_461);
and U443 (N_443,In_84,In_154);
nand U444 (N_444,In_215,In_345);
nand U445 (N_445,In_459,In_430);
nand U446 (N_446,In_384,In_133);
nand U447 (N_447,In_450,In_283);
nor U448 (N_448,In_210,In_128);
nand U449 (N_449,In_338,In_280);
or U450 (N_450,In_434,In_337);
or U451 (N_451,In_341,In_101);
and U452 (N_452,In_366,In_42);
nand U453 (N_453,In_164,In_97);
and U454 (N_454,In_261,In_484);
nor U455 (N_455,In_443,In_391);
nand U456 (N_456,In_258,In_480);
nor U457 (N_457,In_371,In_43);
and U458 (N_458,In_27,In_189);
nor U459 (N_459,In_97,In_499);
or U460 (N_460,In_292,In_134);
or U461 (N_461,In_422,In_417);
nor U462 (N_462,In_140,In_481);
or U463 (N_463,In_246,In_41);
xnor U464 (N_464,In_472,In_254);
nand U465 (N_465,In_170,In_428);
and U466 (N_466,In_124,In_32);
nor U467 (N_467,In_420,In_228);
nor U468 (N_468,In_159,In_36);
or U469 (N_469,In_432,In_265);
nand U470 (N_470,In_312,In_467);
nor U471 (N_471,In_230,In_324);
nand U472 (N_472,In_10,In_204);
nor U473 (N_473,In_134,In_206);
nor U474 (N_474,In_371,In_427);
or U475 (N_475,In_401,In_298);
nand U476 (N_476,In_238,In_201);
nand U477 (N_477,In_83,In_314);
nand U478 (N_478,In_471,In_192);
and U479 (N_479,In_311,In_457);
and U480 (N_480,In_301,In_245);
or U481 (N_481,In_213,In_446);
nand U482 (N_482,In_95,In_205);
nand U483 (N_483,In_174,In_269);
or U484 (N_484,In_13,In_406);
nor U485 (N_485,In_101,In_196);
nand U486 (N_486,In_210,In_434);
nand U487 (N_487,In_32,In_42);
or U488 (N_488,In_480,In_301);
nor U489 (N_489,In_88,In_41);
and U490 (N_490,In_84,In_431);
or U491 (N_491,In_239,In_323);
and U492 (N_492,In_409,In_201);
or U493 (N_493,In_383,In_318);
and U494 (N_494,In_340,In_475);
or U495 (N_495,In_15,In_184);
or U496 (N_496,In_304,In_317);
nand U497 (N_497,In_197,In_147);
and U498 (N_498,In_36,In_281);
and U499 (N_499,In_467,In_397);
and U500 (N_500,N_102,N_201);
and U501 (N_501,N_84,N_222);
nand U502 (N_502,N_412,N_147);
and U503 (N_503,N_492,N_255);
and U504 (N_504,N_337,N_256);
nor U505 (N_505,N_118,N_469);
nor U506 (N_506,N_314,N_493);
nor U507 (N_507,N_326,N_254);
nor U508 (N_508,N_413,N_290);
nor U509 (N_509,N_357,N_180);
nand U510 (N_510,N_460,N_345);
nand U511 (N_511,N_434,N_331);
and U512 (N_512,N_417,N_410);
or U513 (N_513,N_477,N_217);
and U514 (N_514,N_224,N_497);
and U515 (N_515,N_447,N_443);
xor U516 (N_516,N_258,N_248);
nor U517 (N_517,N_430,N_366);
and U518 (N_518,N_245,N_278);
and U519 (N_519,N_116,N_461);
nor U520 (N_520,N_372,N_313);
or U521 (N_521,N_327,N_394);
nor U522 (N_522,N_101,N_414);
nor U523 (N_523,N_252,N_106);
or U524 (N_524,N_479,N_296);
and U525 (N_525,N_288,N_480);
nor U526 (N_526,N_275,N_468);
nor U527 (N_527,N_453,N_73);
and U528 (N_528,N_317,N_368);
nand U529 (N_529,N_274,N_378);
nand U530 (N_530,N_161,N_298);
or U531 (N_531,N_243,N_232);
nor U532 (N_532,N_395,N_52);
and U533 (N_533,N_379,N_79);
nor U534 (N_534,N_125,N_42);
nor U535 (N_535,N_50,N_211);
xor U536 (N_536,N_303,N_316);
nand U537 (N_537,N_27,N_320);
and U538 (N_538,N_190,N_57);
and U539 (N_539,N_85,N_32);
and U540 (N_540,N_114,N_30);
and U541 (N_541,N_31,N_336);
nand U542 (N_542,N_38,N_415);
and U543 (N_543,N_115,N_310);
and U544 (N_544,N_53,N_104);
and U545 (N_545,N_127,N_486);
and U546 (N_546,N_140,N_433);
nor U547 (N_547,N_319,N_373);
or U548 (N_548,N_380,N_142);
nor U549 (N_549,N_33,N_163);
nand U550 (N_550,N_34,N_132);
nand U551 (N_551,N_156,N_152);
or U552 (N_552,N_407,N_382);
or U553 (N_553,N_426,N_351);
nor U554 (N_554,N_219,N_235);
nor U555 (N_555,N_482,N_11);
and U556 (N_556,N_498,N_44);
nand U557 (N_557,N_339,N_392);
or U558 (N_558,N_386,N_207);
or U559 (N_559,N_131,N_291);
nor U560 (N_560,N_247,N_409);
and U561 (N_561,N_158,N_164);
nor U562 (N_562,N_122,N_37);
and U563 (N_563,N_230,N_3);
or U564 (N_564,N_111,N_21);
nor U565 (N_565,N_133,N_26);
nor U566 (N_566,N_91,N_400);
nand U567 (N_567,N_408,N_401);
or U568 (N_568,N_173,N_175);
and U569 (N_569,N_178,N_39);
xnor U570 (N_570,N_450,N_444);
nand U571 (N_571,N_441,N_390);
nor U572 (N_572,N_82,N_198);
nor U573 (N_573,N_213,N_499);
or U574 (N_574,N_349,N_488);
and U575 (N_575,N_98,N_367);
and U576 (N_576,N_344,N_270);
or U577 (N_577,N_117,N_334);
or U578 (N_578,N_66,N_22);
nand U579 (N_579,N_148,N_437);
nand U580 (N_580,N_451,N_297);
and U581 (N_581,N_187,N_419);
and U582 (N_582,N_146,N_212);
or U583 (N_583,N_199,N_466);
nor U584 (N_584,N_472,N_280);
nor U585 (N_585,N_191,N_302);
nor U586 (N_586,N_424,N_216);
or U587 (N_587,N_177,N_110);
and U588 (N_588,N_277,N_257);
xor U589 (N_589,N_233,N_71);
nand U590 (N_590,N_397,N_90);
nor U591 (N_591,N_96,N_45);
or U592 (N_592,N_170,N_120);
nand U593 (N_593,N_353,N_86);
nand U594 (N_594,N_266,N_176);
nor U595 (N_595,N_13,N_128);
or U596 (N_596,N_143,N_234);
or U597 (N_597,N_287,N_202);
nand U598 (N_598,N_182,N_360);
nand U599 (N_599,N_321,N_0);
nor U600 (N_600,N_342,N_227);
or U601 (N_601,N_381,N_457);
nor U602 (N_602,N_483,N_136);
nand U603 (N_603,N_429,N_335);
and U604 (N_604,N_183,N_385);
and U605 (N_605,N_439,N_309);
and U606 (N_606,N_352,N_129);
or U607 (N_607,N_396,N_276);
or U608 (N_608,N_209,N_200);
nand U609 (N_609,N_325,N_49);
and U610 (N_610,N_259,N_387);
and U611 (N_611,N_369,N_484);
nor U612 (N_612,N_108,N_228);
and U613 (N_613,N_403,N_223);
nor U614 (N_614,N_43,N_289);
or U615 (N_615,N_56,N_193);
nand U616 (N_616,N_16,N_172);
xor U617 (N_617,N_364,N_312);
nand U618 (N_618,N_328,N_449);
or U619 (N_619,N_422,N_229);
xor U620 (N_620,N_99,N_206);
and U621 (N_621,N_29,N_197);
xnor U622 (N_622,N_463,N_446);
or U623 (N_623,N_55,N_20);
nand U624 (N_624,N_121,N_494);
nand U625 (N_625,N_10,N_225);
or U626 (N_626,N_307,N_487);
and U627 (N_627,N_62,N_241);
nand U628 (N_628,N_462,N_371);
or U629 (N_629,N_473,N_221);
or U630 (N_630,N_103,N_304);
nor U631 (N_631,N_398,N_188);
and U632 (N_632,N_124,N_467);
or U633 (N_633,N_428,N_340);
and U634 (N_634,N_240,N_195);
and U635 (N_635,N_14,N_406);
and U636 (N_636,N_231,N_470);
nand U637 (N_637,N_194,N_332);
or U638 (N_638,N_384,N_80);
nand U639 (N_639,N_294,N_456);
nor U640 (N_640,N_306,N_318);
or U641 (N_641,N_74,N_157);
and U642 (N_642,N_476,N_322);
and U643 (N_643,N_186,N_208);
or U644 (N_644,N_346,N_261);
and U645 (N_645,N_112,N_154);
nor U646 (N_646,N_279,N_347);
or U647 (N_647,N_226,N_391);
xor U648 (N_648,N_485,N_237);
and U649 (N_649,N_67,N_28);
nand U650 (N_650,N_354,N_474);
and U651 (N_651,N_475,N_455);
nor U652 (N_652,N_458,N_153);
and U653 (N_653,N_361,N_399);
and U654 (N_654,N_383,N_138);
and U655 (N_655,N_65,N_239);
and U656 (N_656,N_432,N_242);
nor U657 (N_657,N_192,N_249);
nand U658 (N_658,N_77,N_262);
nor U659 (N_659,N_36,N_160);
nor U660 (N_660,N_9,N_295);
nand U661 (N_661,N_141,N_47);
xnor U662 (N_662,N_496,N_4);
nor U663 (N_663,N_244,N_286);
nor U664 (N_664,N_139,N_251);
nor U665 (N_665,N_58,N_46);
nand U666 (N_666,N_5,N_78);
or U667 (N_667,N_362,N_445);
nand U668 (N_668,N_218,N_2);
nand U669 (N_669,N_436,N_459);
or U670 (N_670,N_388,N_405);
nor U671 (N_671,N_1,N_203);
nor U672 (N_672,N_283,N_169);
and U673 (N_673,N_418,N_358);
nand U674 (N_674,N_350,N_210);
nand U675 (N_675,N_92,N_238);
and U676 (N_676,N_393,N_60);
and U677 (N_677,N_19,N_25);
or U678 (N_678,N_365,N_355);
nand U679 (N_679,N_40,N_284);
nor U680 (N_680,N_72,N_12);
nor U681 (N_681,N_167,N_246);
and U682 (N_682,N_495,N_416);
nand U683 (N_683,N_389,N_423);
or U684 (N_684,N_442,N_48);
xor U685 (N_685,N_301,N_88);
nand U686 (N_686,N_435,N_171);
xnor U687 (N_687,N_324,N_490);
nor U688 (N_688,N_134,N_119);
nand U689 (N_689,N_151,N_8);
or U690 (N_690,N_293,N_265);
nand U691 (N_691,N_377,N_236);
nor U692 (N_692,N_24,N_64);
nor U693 (N_693,N_196,N_333);
or U694 (N_694,N_149,N_465);
and U695 (N_695,N_452,N_166);
nor U696 (N_696,N_63,N_93);
nand U697 (N_697,N_359,N_107);
nand U698 (N_698,N_144,N_97);
nand U699 (N_699,N_311,N_263);
or U700 (N_700,N_135,N_215);
or U701 (N_701,N_305,N_375);
nor U702 (N_702,N_330,N_425);
nand U703 (N_703,N_18,N_250);
and U704 (N_704,N_481,N_341);
and U705 (N_705,N_323,N_162);
nor U706 (N_706,N_68,N_329);
nand U707 (N_707,N_81,N_292);
nor U708 (N_708,N_271,N_150);
or U709 (N_709,N_431,N_126);
nand U710 (N_710,N_370,N_184);
and U711 (N_711,N_260,N_471);
xor U712 (N_712,N_165,N_179);
nor U713 (N_713,N_155,N_282);
and U714 (N_714,N_54,N_264);
xnor U715 (N_715,N_220,N_348);
nand U716 (N_716,N_105,N_109);
nand U717 (N_717,N_145,N_376);
nand U718 (N_718,N_402,N_427);
nand U719 (N_719,N_87,N_269);
and U720 (N_720,N_181,N_281);
or U721 (N_721,N_356,N_189);
nor U722 (N_722,N_338,N_41);
or U723 (N_723,N_69,N_100);
or U724 (N_724,N_137,N_6);
nor U725 (N_725,N_75,N_159);
nor U726 (N_726,N_421,N_94);
nor U727 (N_727,N_363,N_214);
nand U728 (N_728,N_464,N_285);
or U729 (N_729,N_17,N_130);
or U730 (N_730,N_272,N_35);
or U731 (N_731,N_440,N_7);
or U732 (N_732,N_315,N_59);
nor U733 (N_733,N_273,N_95);
and U734 (N_734,N_489,N_70);
nor U735 (N_735,N_89,N_204);
nand U736 (N_736,N_411,N_76);
nor U737 (N_737,N_51,N_123);
and U738 (N_738,N_83,N_491);
or U739 (N_739,N_454,N_268);
nand U740 (N_740,N_168,N_343);
nand U741 (N_741,N_448,N_299);
nor U742 (N_742,N_185,N_61);
and U743 (N_743,N_308,N_478);
and U744 (N_744,N_374,N_174);
or U745 (N_745,N_205,N_253);
and U746 (N_746,N_420,N_15);
or U747 (N_747,N_23,N_404);
and U748 (N_748,N_267,N_113);
or U749 (N_749,N_300,N_438);
or U750 (N_750,N_278,N_215);
or U751 (N_751,N_240,N_231);
and U752 (N_752,N_210,N_211);
or U753 (N_753,N_34,N_189);
nor U754 (N_754,N_198,N_147);
nor U755 (N_755,N_189,N_454);
or U756 (N_756,N_142,N_41);
nor U757 (N_757,N_52,N_281);
nor U758 (N_758,N_254,N_316);
nand U759 (N_759,N_208,N_274);
and U760 (N_760,N_368,N_220);
nand U761 (N_761,N_81,N_191);
or U762 (N_762,N_180,N_241);
xor U763 (N_763,N_260,N_307);
or U764 (N_764,N_343,N_425);
and U765 (N_765,N_409,N_257);
or U766 (N_766,N_177,N_391);
or U767 (N_767,N_306,N_435);
nand U768 (N_768,N_325,N_339);
nor U769 (N_769,N_153,N_454);
nand U770 (N_770,N_373,N_453);
and U771 (N_771,N_55,N_441);
or U772 (N_772,N_363,N_73);
and U773 (N_773,N_187,N_472);
and U774 (N_774,N_430,N_396);
and U775 (N_775,N_100,N_395);
nand U776 (N_776,N_343,N_330);
and U777 (N_777,N_75,N_198);
nand U778 (N_778,N_410,N_16);
nor U779 (N_779,N_137,N_17);
and U780 (N_780,N_313,N_424);
nor U781 (N_781,N_15,N_68);
nor U782 (N_782,N_485,N_303);
nor U783 (N_783,N_146,N_430);
xor U784 (N_784,N_180,N_95);
or U785 (N_785,N_183,N_18);
or U786 (N_786,N_226,N_67);
nand U787 (N_787,N_312,N_137);
and U788 (N_788,N_123,N_25);
and U789 (N_789,N_471,N_363);
or U790 (N_790,N_246,N_302);
nor U791 (N_791,N_186,N_457);
nor U792 (N_792,N_400,N_53);
or U793 (N_793,N_105,N_161);
or U794 (N_794,N_376,N_443);
nand U795 (N_795,N_238,N_267);
nor U796 (N_796,N_303,N_471);
and U797 (N_797,N_61,N_10);
and U798 (N_798,N_249,N_418);
nand U799 (N_799,N_154,N_102);
nand U800 (N_800,N_465,N_23);
and U801 (N_801,N_87,N_410);
and U802 (N_802,N_306,N_206);
nand U803 (N_803,N_334,N_149);
xnor U804 (N_804,N_407,N_327);
and U805 (N_805,N_175,N_353);
nand U806 (N_806,N_284,N_259);
nand U807 (N_807,N_320,N_91);
xnor U808 (N_808,N_24,N_255);
nor U809 (N_809,N_463,N_164);
nor U810 (N_810,N_273,N_221);
and U811 (N_811,N_163,N_383);
or U812 (N_812,N_354,N_210);
or U813 (N_813,N_109,N_400);
and U814 (N_814,N_334,N_183);
and U815 (N_815,N_136,N_390);
nor U816 (N_816,N_197,N_5);
nand U817 (N_817,N_4,N_374);
nor U818 (N_818,N_314,N_6);
and U819 (N_819,N_251,N_381);
or U820 (N_820,N_173,N_281);
and U821 (N_821,N_236,N_65);
nor U822 (N_822,N_351,N_373);
nand U823 (N_823,N_376,N_246);
or U824 (N_824,N_410,N_239);
or U825 (N_825,N_177,N_85);
nor U826 (N_826,N_366,N_219);
nor U827 (N_827,N_194,N_308);
or U828 (N_828,N_337,N_217);
or U829 (N_829,N_493,N_465);
or U830 (N_830,N_139,N_190);
and U831 (N_831,N_122,N_334);
nor U832 (N_832,N_379,N_154);
and U833 (N_833,N_8,N_343);
and U834 (N_834,N_69,N_96);
and U835 (N_835,N_53,N_12);
nor U836 (N_836,N_389,N_323);
nand U837 (N_837,N_319,N_262);
and U838 (N_838,N_352,N_233);
or U839 (N_839,N_17,N_426);
nor U840 (N_840,N_401,N_382);
or U841 (N_841,N_379,N_404);
and U842 (N_842,N_489,N_255);
and U843 (N_843,N_25,N_107);
or U844 (N_844,N_326,N_139);
and U845 (N_845,N_487,N_344);
nand U846 (N_846,N_215,N_228);
or U847 (N_847,N_367,N_62);
and U848 (N_848,N_9,N_43);
or U849 (N_849,N_231,N_298);
nand U850 (N_850,N_262,N_78);
nand U851 (N_851,N_376,N_83);
and U852 (N_852,N_234,N_308);
and U853 (N_853,N_449,N_17);
and U854 (N_854,N_156,N_183);
or U855 (N_855,N_431,N_301);
or U856 (N_856,N_414,N_245);
nand U857 (N_857,N_430,N_220);
or U858 (N_858,N_89,N_186);
and U859 (N_859,N_13,N_125);
and U860 (N_860,N_94,N_382);
and U861 (N_861,N_17,N_169);
and U862 (N_862,N_461,N_149);
and U863 (N_863,N_238,N_220);
and U864 (N_864,N_99,N_337);
or U865 (N_865,N_462,N_376);
nor U866 (N_866,N_402,N_404);
nand U867 (N_867,N_256,N_141);
nor U868 (N_868,N_375,N_2);
nor U869 (N_869,N_316,N_84);
nand U870 (N_870,N_270,N_430);
or U871 (N_871,N_136,N_156);
nor U872 (N_872,N_175,N_407);
and U873 (N_873,N_497,N_173);
xor U874 (N_874,N_433,N_336);
nand U875 (N_875,N_49,N_119);
xor U876 (N_876,N_169,N_400);
and U877 (N_877,N_200,N_126);
nor U878 (N_878,N_144,N_106);
nor U879 (N_879,N_285,N_445);
nor U880 (N_880,N_189,N_398);
nand U881 (N_881,N_493,N_136);
nor U882 (N_882,N_67,N_126);
or U883 (N_883,N_117,N_118);
xor U884 (N_884,N_392,N_317);
or U885 (N_885,N_139,N_45);
nor U886 (N_886,N_84,N_9);
nor U887 (N_887,N_223,N_407);
nor U888 (N_888,N_196,N_154);
or U889 (N_889,N_451,N_62);
or U890 (N_890,N_11,N_221);
or U891 (N_891,N_180,N_415);
and U892 (N_892,N_301,N_484);
and U893 (N_893,N_341,N_92);
and U894 (N_894,N_190,N_361);
xor U895 (N_895,N_249,N_344);
nand U896 (N_896,N_301,N_494);
and U897 (N_897,N_55,N_255);
or U898 (N_898,N_139,N_189);
nor U899 (N_899,N_210,N_103);
nor U900 (N_900,N_114,N_179);
nor U901 (N_901,N_402,N_348);
nand U902 (N_902,N_276,N_197);
nor U903 (N_903,N_98,N_464);
nor U904 (N_904,N_63,N_307);
nor U905 (N_905,N_127,N_52);
nor U906 (N_906,N_376,N_404);
or U907 (N_907,N_429,N_240);
and U908 (N_908,N_193,N_142);
nor U909 (N_909,N_425,N_295);
nand U910 (N_910,N_197,N_496);
or U911 (N_911,N_277,N_397);
and U912 (N_912,N_351,N_81);
nand U913 (N_913,N_269,N_418);
and U914 (N_914,N_125,N_457);
xnor U915 (N_915,N_38,N_44);
or U916 (N_916,N_201,N_336);
nor U917 (N_917,N_317,N_101);
nor U918 (N_918,N_375,N_128);
nor U919 (N_919,N_387,N_149);
or U920 (N_920,N_57,N_411);
or U921 (N_921,N_267,N_224);
or U922 (N_922,N_141,N_163);
nand U923 (N_923,N_382,N_332);
and U924 (N_924,N_420,N_169);
nand U925 (N_925,N_442,N_138);
nand U926 (N_926,N_161,N_182);
or U927 (N_927,N_225,N_38);
or U928 (N_928,N_232,N_183);
or U929 (N_929,N_369,N_106);
or U930 (N_930,N_267,N_378);
and U931 (N_931,N_279,N_439);
and U932 (N_932,N_324,N_328);
nor U933 (N_933,N_294,N_31);
or U934 (N_934,N_322,N_233);
nand U935 (N_935,N_271,N_311);
nor U936 (N_936,N_97,N_478);
and U937 (N_937,N_110,N_355);
or U938 (N_938,N_372,N_477);
nand U939 (N_939,N_111,N_5);
nor U940 (N_940,N_460,N_263);
or U941 (N_941,N_369,N_226);
xnor U942 (N_942,N_117,N_58);
nand U943 (N_943,N_215,N_249);
nand U944 (N_944,N_68,N_150);
nand U945 (N_945,N_205,N_370);
or U946 (N_946,N_268,N_70);
and U947 (N_947,N_65,N_219);
or U948 (N_948,N_388,N_155);
nand U949 (N_949,N_297,N_120);
nand U950 (N_950,N_350,N_433);
nor U951 (N_951,N_273,N_277);
nand U952 (N_952,N_146,N_300);
nor U953 (N_953,N_404,N_213);
nor U954 (N_954,N_302,N_419);
xnor U955 (N_955,N_380,N_202);
and U956 (N_956,N_225,N_449);
or U957 (N_957,N_146,N_466);
and U958 (N_958,N_439,N_466);
nand U959 (N_959,N_293,N_343);
and U960 (N_960,N_121,N_163);
nor U961 (N_961,N_481,N_127);
and U962 (N_962,N_170,N_140);
or U963 (N_963,N_170,N_383);
nor U964 (N_964,N_180,N_127);
and U965 (N_965,N_343,N_318);
nand U966 (N_966,N_214,N_38);
or U967 (N_967,N_24,N_65);
nand U968 (N_968,N_316,N_448);
and U969 (N_969,N_325,N_86);
and U970 (N_970,N_496,N_23);
nor U971 (N_971,N_215,N_25);
or U972 (N_972,N_166,N_155);
nand U973 (N_973,N_297,N_397);
xor U974 (N_974,N_25,N_369);
and U975 (N_975,N_74,N_238);
nor U976 (N_976,N_39,N_452);
nor U977 (N_977,N_230,N_224);
nor U978 (N_978,N_136,N_421);
or U979 (N_979,N_135,N_2);
nor U980 (N_980,N_368,N_383);
and U981 (N_981,N_437,N_480);
or U982 (N_982,N_141,N_456);
nand U983 (N_983,N_376,N_394);
nor U984 (N_984,N_81,N_115);
and U985 (N_985,N_159,N_348);
and U986 (N_986,N_42,N_116);
and U987 (N_987,N_185,N_390);
nor U988 (N_988,N_43,N_10);
nand U989 (N_989,N_443,N_308);
or U990 (N_990,N_400,N_210);
nor U991 (N_991,N_115,N_294);
or U992 (N_992,N_411,N_484);
and U993 (N_993,N_142,N_298);
nand U994 (N_994,N_249,N_161);
and U995 (N_995,N_283,N_229);
or U996 (N_996,N_98,N_484);
nor U997 (N_997,N_121,N_475);
and U998 (N_998,N_279,N_379);
nand U999 (N_999,N_202,N_247);
and U1000 (N_1000,N_907,N_789);
or U1001 (N_1001,N_602,N_849);
nand U1002 (N_1002,N_969,N_677);
nor U1003 (N_1003,N_857,N_589);
nand U1004 (N_1004,N_740,N_716);
and U1005 (N_1005,N_706,N_581);
or U1006 (N_1006,N_557,N_785);
and U1007 (N_1007,N_807,N_669);
and U1008 (N_1008,N_842,N_970);
or U1009 (N_1009,N_872,N_679);
xnor U1010 (N_1010,N_744,N_615);
nor U1011 (N_1011,N_814,N_665);
or U1012 (N_1012,N_966,N_548);
nand U1013 (N_1013,N_523,N_976);
nand U1014 (N_1014,N_537,N_648);
nand U1015 (N_1015,N_886,N_845);
and U1016 (N_1016,N_501,N_852);
and U1017 (N_1017,N_509,N_569);
nor U1018 (N_1018,N_882,N_865);
xnor U1019 (N_1019,N_894,N_580);
or U1020 (N_1020,N_993,N_978);
and U1021 (N_1021,N_796,N_588);
or U1022 (N_1022,N_968,N_577);
nand U1023 (N_1023,N_631,N_977);
xnor U1024 (N_1024,N_651,N_830);
or U1025 (N_1025,N_837,N_681);
nor U1026 (N_1026,N_660,N_753);
or U1027 (N_1027,N_554,N_728);
or U1028 (N_1028,N_749,N_988);
nand U1029 (N_1029,N_973,N_598);
and U1030 (N_1030,N_769,N_719);
nor U1031 (N_1031,N_795,N_752);
or U1032 (N_1032,N_914,N_793);
or U1033 (N_1033,N_871,N_559);
or U1034 (N_1034,N_819,N_955);
or U1035 (N_1035,N_779,N_881);
or U1036 (N_1036,N_790,N_685);
nor U1037 (N_1037,N_937,N_691);
nand U1038 (N_1038,N_764,N_880);
or U1039 (N_1039,N_739,N_659);
or U1040 (N_1040,N_906,N_941);
and U1041 (N_1041,N_763,N_626);
and U1042 (N_1042,N_515,N_636);
nand U1043 (N_1043,N_946,N_998);
nand U1044 (N_1044,N_956,N_902);
nor U1045 (N_1045,N_513,N_535);
nor U1046 (N_1046,N_713,N_990);
nor U1047 (N_1047,N_534,N_766);
and U1048 (N_1048,N_560,N_634);
nand U1049 (N_1049,N_806,N_999);
nor U1050 (N_1050,N_503,N_721);
nand U1051 (N_1051,N_673,N_675);
nand U1052 (N_1052,N_638,N_574);
or U1053 (N_1053,N_778,N_897);
nand U1054 (N_1054,N_575,N_889);
nor U1055 (N_1055,N_887,N_551);
nand U1056 (N_1056,N_985,N_612);
or U1057 (N_1057,N_817,N_715);
nand U1058 (N_1058,N_953,N_630);
or U1059 (N_1059,N_510,N_931);
nor U1060 (N_1060,N_952,N_687);
xnor U1061 (N_1061,N_986,N_875);
or U1062 (N_1062,N_570,N_682);
nand U1063 (N_1063,N_816,N_870);
nor U1064 (N_1064,N_755,N_811);
or U1065 (N_1065,N_947,N_639);
nor U1066 (N_1066,N_741,N_933);
and U1067 (N_1067,N_693,N_573);
nor U1068 (N_1068,N_661,N_583);
nor U1069 (N_1069,N_609,N_801);
or U1070 (N_1070,N_996,N_696);
nor U1071 (N_1071,N_858,N_737);
or U1072 (N_1072,N_767,N_962);
nand U1073 (N_1073,N_776,N_920);
and U1074 (N_1074,N_723,N_835);
nor U1075 (N_1075,N_909,N_502);
or U1076 (N_1076,N_777,N_797);
or U1077 (N_1077,N_949,N_618);
nand U1078 (N_1078,N_821,N_828);
nand U1079 (N_1079,N_957,N_622);
and U1080 (N_1080,N_771,N_926);
or U1081 (N_1081,N_561,N_683);
nor U1082 (N_1082,N_525,N_572);
or U1083 (N_1083,N_935,N_948);
nor U1084 (N_1084,N_809,N_844);
nand U1085 (N_1085,N_787,N_586);
nand U1086 (N_1086,N_649,N_900);
nor U1087 (N_1087,N_910,N_916);
or U1088 (N_1088,N_884,N_709);
nor U1089 (N_1089,N_748,N_975);
or U1090 (N_1090,N_918,N_788);
and U1091 (N_1091,N_928,N_831);
or U1092 (N_1092,N_507,N_550);
and U1093 (N_1093,N_624,N_934);
nand U1094 (N_1094,N_873,N_565);
or U1095 (N_1095,N_943,N_747);
nor U1096 (N_1096,N_840,N_803);
and U1097 (N_1097,N_915,N_862);
nand U1098 (N_1098,N_644,N_567);
or U1099 (N_1099,N_773,N_576);
nor U1100 (N_1100,N_734,N_658);
or U1101 (N_1101,N_584,N_695);
nand U1102 (N_1102,N_564,N_692);
nor U1103 (N_1103,N_994,N_710);
or U1104 (N_1104,N_768,N_594);
nand U1105 (N_1105,N_802,N_834);
nand U1106 (N_1106,N_655,N_836);
or U1107 (N_1107,N_984,N_827);
or U1108 (N_1108,N_867,N_629);
xnor U1109 (N_1109,N_725,N_979);
nand U1110 (N_1110,N_505,N_616);
or U1111 (N_1111,N_637,N_905);
or U1112 (N_1112,N_668,N_820);
or U1113 (N_1113,N_818,N_671);
nand U1114 (N_1114,N_783,N_841);
or U1115 (N_1115,N_772,N_971);
nand U1116 (N_1116,N_932,N_810);
and U1117 (N_1117,N_504,N_972);
nand U1118 (N_1118,N_982,N_846);
nand U1119 (N_1119,N_640,N_912);
nand U1120 (N_1120,N_959,N_874);
and U1121 (N_1121,N_829,N_758);
and U1122 (N_1122,N_607,N_899);
or U1123 (N_1123,N_605,N_582);
and U1124 (N_1124,N_712,N_813);
and U1125 (N_1125,N_542,N_526);
or U1126 (N_1126,N_717,N_743);
nand U1127 (N_1127,N_950,N_623);
or U1128 (N_1128,N_967,N_600);
nor U1129 (N_1129,N_954,N_539);
or U1130 (N_1130,N_686,N_617);
nor U1131 (N_1131,N_591,N_604);
nand U1132 (N_1132,N_908,N_621);
and U1133 (N_1133,N_891,N_705);
nand U1134 (N_1134,N_784,N_601);
or U1135 (N_1135,N_815,N_980);
nor U1136 (N_1136,N_863,N_930);
and U1137 (N_1137,N_500,N_558);
and U1138 (N_1138,N_650,N_786);
nor U1139 (N_1139,N_646,N_508);
nor U1140 (N_1140,N_724,N_878);
nand U1141 (N_1141,N_883,N_647);
nand U1142 (N_1142,N_632,N_593);
or U1143 (N_1143,N_869,N_775);
or U1144 (N_1144,N_855,N_531);
nand U1145 (N_1145,N_652,N_800);
and U1146 (N_1146,N_927,N_684);
nor U1147 (N_1147,N_825,N_854);
and U1148 (N_1148,N_642,N_832);
xor U1149 (N_1149,N_606,N_850);
or U1150 (N_1150,N_517,N_965);
and U1151 (N_1151,N_765,N_876);
nand U1152 (N_1152,N_822,N_613);
nor U1153 (N_1153,N_746,N_614);
nand U1154 (N_1154,N_942,N_553);
or U1155 (N_1155,N_656,N_864);
and U1156 (N_1156,N_545,N_851);
nor U1157 (N_1157,N_799,N_689);
nor U1158 (N_1158,N_524,N_536);
nand U1159 (N_1159,N_732,N_774);
or U1160 (N_1160,N_562,N_754);
nand U1161 (N_1161,N_913,N_805);
nor U1162 (N_1162,N_945,N_700);
nor U1163 (N_1163,N_987,N_662);
xnor U1164 (N_1164,N_518,N_512);
or U1165 (N_1165,N_745,N_963);
and U1166 (N_1166,N_633,N_533);
and U1167 (N_1167,N_722,N_530);
nand U1168 (N_1168,N_782,N_522);
or U1169 (N_1169,N_919,N_853);
nand U1170 (N_1170,N_547,N_736);
nand U1171 (N_1171,N_951,N_628);
nand U1172 (N_1172,N_995,N_917);
and U1173 (N_1173,N_888,N_911);
nor U1174 (N_1174,N_856,N_925);
and U1175 (N_1175,N_672,N_532);
or U1176 (N_1176,N_936,N_901);
or U1177 (N_1177,N_944,N_718);
or U1178 (N_1178,N_903,N_735);
nand U1179 (N_1179,N_895,N_833);
nor U1180 (N_1180,N_620,N_595);
and U1181 (N_1181,N_824,N_694);
and U1182 (N_1182,N_929,N_997);
nand U1183 (N_1183,N_610,N_592);
nor U1184 (N_1184,N_549,N_733);
or U1185 (N_1185,N_670,N_868);
xnor U1186 (N_1186,N_742,N_635);
or U1187 (N_1187,N_654,N_898);
and U1188 (N_1188,N_541,N_556);
or U1189 (N_1189,N_538,N_568);
and U1190 (N_1190,N_808,N_698);
nor U1191 (N_1191,N_627,N_688);
or U1192 (N_1192,N_860,N_540);
nor U1193 (N_1193,N_826,N_529);
nor U1194 (N_1194,N_579,N_751);
nand U1195 (N_1195,N_506,N_983);
nor U1196 (N_1196,N_603,N_519);
nor U1197 (N_1197,N_699,N_645);
nor U1198 (N_1198,N_893,N_738);
or U1199 (N_1199,N_958,N_521);
nand U1200 (N_1200,N_879,N_704);
nand U1201 (N_1201,N_770,N_608);
nand U1202 (N_1202,N_750,N_678);
nand U1203 (N_1203,N_896,N_759);
nand U1204 (N_1204,N_885,N_780);
nand U1205 (N_1205,N_964,N_701);
or U1206 (N_1206,N_904,N_804);
nor U1207 (N_1207,N_702,N_590);
nand U1208 (N_1208,N_877,N_555);
nand U1209 (N_1209,N_680,N_974);
nor U1210 (N_1210,N_697,N_791);
and U1211 (N_1211,N_757,N_991);
nand U1212 (N_1212,N_989,N_762);
xnor U1213 (N_1213,N_546,N_653);
xor U1214 (N_1214,N_848,N_619);
nor U1215 (N_1215,N_798,N_666);
or U1216 (N_1216,N_838,N_663);
and U1217 (N_1217,N_566,N_756);
nor U1218 (N_1218,N_667,N_664);
or U1219 (N_1219,N_921,N_707);
nand U1220 (N_1220,N_960,N_938);
xor U1221 (N_1221,N_597,N_520);
or U1222 (N_1222,N_528,N_794);
nand U1223 (N_1223,N_514,N_940);
nor U1224 (N_1224,N_961,N_516);
nor U1225 (N_1225,N_892,N_823);
or U1226 (N_1226,N_727,N_861);
nand U1227 (N_1227,N_676,N_711);
nand U1228 (N_1228,N_760,N_720);
and U1229 (N_1229,N_599,N_726);
nor U1230 (N_1230,N_839,N_596);
nand U1231 (N_1231,N_511,N_544);
nand U1232 (N_1232,N_563,N_761);
nor U1233 (N_1233,N_657,N_847);
nor U1234 (N_1234,N_641,N_674);
nor U1235 (N_1235,N_729,N_981);
xor U1236 (N_1236,N_792,N_923);
nor U1237 (N_1237,N_781,N_866);
and U1238 (N_1238,N_543,N_703);
nor U1239 (N_1239,N_611,N_812);
nor U1240 (N_1240,N_939,N_625);
nor U1241 (N_1241,N_585,N_578);
and U1242 (N_1242,N_714,N_527);
nand U1243 (N_1243,N_924,N_843);
or U1244 (N_1244,N_643,N_731);
nand U1245 (N_1245,N_859,N_552);
nand U1246 (N_1246,N_922,N_708);
nand U1247 (N_1247,N_992,N_730);
nor U1248 (N_1248,N_890,N_690);
or U1249 (N_1249,N_571,N_587);
nand U1250 (N_1250,N_597,N_532);
nor U1251 (N_1251,N_933,N_617);
nand U1252 (N_1252,N_550,N_823);
or U1253 (N_1253,N_503,N_528);
and U1254 (N_1254,N_683,N_730);
nand U1255 (N_1255,N_527,N_625);
and U1256 (N_1256,N_929,N_862);
nand U1257 (N_1257,N_801,N_885);
nor U1258 (N_1258,N_581,N_576);
or U1259 (N_1259,N_586,N_627);
nor U1260 (N_1260,N_828,N_924);
nor U1261 (N_1261,N_917,N_600);
or U1262 (N_1262,N_682,N_699);
nor U1263 (N_1263,N_994,N_983);
nor U1264 (N_1264,N_926,N_662);
or U1265 (N_1265,N_789,N_933);
nor U1266 (N_1266,N_596,N_805);
nand U1267 (N_1267,N_651,N_586);
xnor U1268 (N_1268,N_814,N_657);
nor U1269 (N_1269,N_553,N_668);
and U1270 (N_1270,N_597,N_807);
nor U1271 (N_1271,N_516,N_541);
nand U1272 (N_1272,N_652,N_798);
and U1273 (N_1273,N_768,N_521);
and U1274 (N_1274,N_759,N_792);
nand U1275 (N_1275,N_720,N_857);
and U1276 (N_1276,N_879,N_563);
nand U1277 (N_1277,N_515,N_587);
nor U1278 (N_1278,N_747,N_885);
xnor U1279 (N_1279,N_797,N_736);
xnor U1280 (N_1280,N_645,N_957);
nand U1281 (N_1281,N_658,N_840);
nor U1282 (N_1282,N_541,N_668);
and U1283 (N_1283,N_668,N_620);
nor U1284 (N_1284,N_903,N_650);
or U1285 (N_1285,N_833,N_958);
nor U1286 (N_1286,N_749,N_782);
nor U1287 (N_1287,N_622,N_962);
or U1288 (N_1288,N_835,N_760);
or U1289 (N_1289,N_859,N_923);
nor U1290 (N_1290,N_745,N_934);
and U1291 (N_1291,N_616,N_786);
and U1292 (N_1292,N_888,N_554);
or U1293 (N_1293,N_927,N_622);
nand U1294 (N_1294,N_718,N_873);
nand U1295 (N_1295,N_685,N_724);
xor U1296 (N_1296,N_518,N_971);
nor U1297 (N_1297,N_603,N_830);
nand U1298 (N_1298,N_507,N_882);
or U1299 (N_1299,N_859,N_935);
xnor U1300 (N_1300,N_822,N_798);
and U1301 (N_1301,N_967,N_972);
xor U1302 (N_1302,N_515,N_807);
or U1303 (N_1303,N_547,N_770);
or U1304 (N_1304,N_506,N_972);
xnor U1305 (N_1305,N_779,N_725);
nor U1306 (N_1306,N_783,N_844);
nor U1307 (N_1307,N_773,N_504);
or U1308 (N_1308,N_596,N_644);
nand U1309 (N_1309,N_527,N_561);
or U1310 (N_1310,N_726,N_603);
nand U1311 (N_1311,N_938,N_625);
or U1312 (N_1312,N_868,N_548);
and U1313 (N_1313,N_963,N_826);
nor U1314 (N_1314,N_749,N_973);
nor U1315 (N_1315,N_989,N_931);
nand U1316 (N_1316,N_959,N_801);
or U1317 (N_1317,N_964,N_766);
or U1318 (N_1318,N_850,N_648);
nor U1319 (N_1319,N_525,N_575);
nor U1320 (N_1320,N_769,N_550);
nor U1321 (N_1321,N_947,N_683);
nand U1322 (N_1322,N_867,N_667);
xnor U1323 (N_1323,N_752,N_566);
nand U1324 (N_1324,N_904,N_724);
nand U1325 (N_1325,N_597,N_810);
nor U1326 (N_1326,N_746,N_848);
nor U1327 (N_1327,N_933,N_783);
nand U1328 (N_1328,N_961,N_634);
and U1329 (N_1329,N_990,N_998);
nand U1330 (N_1330,N_803,N_805);
nor U1331 (N_1331,N_993,N_666);
and U1332 (N_1332,N_897,N_953);
or U1333 (N_1333,N_551,N_932);
nand U1334 (N_1334,N_883,N_746);
or U1335 (N_1335,N_895,N_884);
or U1336 (N_1336,N_688,N_559);
and U1337 (N_1337,N_840,N_829);
or U1338 (N_1338,N_554,N_569);
nand U1339 (N_1339,N_960,N_853);
nor U1340 (N_1340,N_679,N_596);
or U1341 (N_1341,N_847,N_661);
nor U1342 (N_1342,N_815,N_832);
and U1343 (N_1343,N_719,N_643);
nor U1344 (N_1344,N_679,N_717);
nand U1345 (N_1345,N_561,N_566);
and U1346 (N_1346,N_517,N_893);
or U1347 (N_1347,N_779,N_988);
nor U1348 (N_1348,N_747,N_964);
and U1349 (N_1349,N_599,N_750);
and U1350 (N_1350,N_684,N_803);
nand U1351 (N_1351,N_536,N_547);
xnor U1352 (N_1352,N_918,N_538);
nor U1353 (N_1353,N_575,N_858);
nand U1354 (N_1354,N_684,N_896);
nor U1355 (N_1355,N_897,N_524);
nand U1356 (N_1356,N_596,N_675);
nand U1357 (N_1357,N_865,N_660);
xor U1358 (N_1358,N_690,N_914);
or U1359 (N_1359,N_600,N_525);
and U1360 (N_1360,N_692,N_517);
and U1361 (N_1361,N_625,N_965);
nand U1362 (N_1362,N_578,N_572);
or U1363 (N_1363,N_570,N_565);
xor U1364 (N_1364,N_782,N_802);
or U1365 (N_1365,N_570,N_962);
and U1366 (N_1366,N_908,N_675);
or U1367 (N_1367,N_636,N_567);
or U1368 (N_1368,N_552,N_553);
and U1369 (N_1369,N_698,N_683);
and U1370 (N_1370,N_808,N_655);
and U1371 (N_1371,N_809,N_934);
or U1372 (N_1372,N_658,N_810);
and U1373 (N_1373,N_684,N_897);
or U1374 (N_1374,N_845,N_614);
and U1375 (N_1375,N_923,N_718);
nor U1376 (N_1376,N_603,N_920);
or U1377 (N_1377,N_757,N_633);
or U1378 (N_1378,N_641,N_782);
nor U1379 (N_1379,N_641,N_922);
and U1380 (N_1380,N_784,N_726);
and U1381 (N_1381,N_587,N_765);
and U1382 (N_1382,N_979,N_865);
and U1383 (N_1383,N_818,N_641);
nand U1384 (N_1384,N_551,N_507);
nand U1385 (N_1385,N_793,N_958);
or U1386 (N_1386,N_503,N_577);
and U1387 (N_1387,N_507,N_797);
or U1388 (N_1388,N_734,N_915);
nor U1389 (N_1389,N_636,N_660);
or U1390 (N_1390,N_965,N_819);
or U1391 (N_1391,N_710,N_927);
and U1392 (N_1392,N_846,N_870);
or U1393 (N_1393,N_662,N_529);
and U1394 (N_1394,N_644,N_704);
nand U1395 (N_1395,N_579,N_557);
nand U1396 (N_1396,N_614,N_769);
nand U1397 (N_1397,N_609,N_820);
and U1398 (N_1398,N_939,N_602);
nor U1399 (N_1399,N_537,N_643);
nand U1400 (N_1400,N_770,N_784);
or U1401 (N_1401,N_524,N_652);
and U1402 (N_1402,N_628,N_733);
nand U1403 (N_1403,N_663,N_815);
nor U1404 (N_1404,N_614,N_849);
nand U1405 (N_1405,N_523,N_615);
nand U1406 (N_1406,N_815,N_614);
nand U1407 (N_1407,N_662,N_951);
and U1408 (N_1408,N_711,N_567);
and U1409 (N_1409,N_913,N_638);
nor U1410 (N_1410,N_866,N_704);
nand U1411 (N_1411,N_749,N_620);
nand U1412 (N_1412,N_956,N_874);
or U1413 (N_1413,N_902,N_623);
and U1414 (N_1414,N_776,N_999);
nor U1415 (N_1415,N_504,N_531);
xnor U1416 (N_1416,N_957,N_610);
or U1417 (N_1417,N_548,N_692);
nor U1418 (N_1418,N_519,N_857);
nor U1419 (N_1419,N_513,N_724);
nor U1420 (N_1420,N_500,N_709);
xnor U1421 (N_1421,N_938,N_690);
nor U1422 (N_1422,N_991,N_521);
nand U1423 (N_1423,N_714,N_763);
or U1424 (N_1424,N_710,N_656);
nor U1425 (N_1425,N_669,N_934);
nor U1426 (N_1426,N_877,N_768);
nand U1427 (N_1427,N_718,N_641);
nor U1428 (N_1428,N_995,N_628);
or U1429 (N_1429,N_868,N_865);
nand U1430 (N_1430,N_634,N_842);
or U1431 (N_1431,N_880,N_569);
xor U1432 (N_1432,N_906,N_871);
nor U1433 (N_1433,N_509,N_795);
or U1434 (N_1434,N_542,N_587);
and U1435 (N_1435,N_582,N_938);
nor U1436 (N_1436,N_567,N_779);
and U1437 (N_1437,N_994,N_695);
nand U1438 (N_1438,N_577,N_627);
or U1439 (N_1439,N_999,N_861);
nand U1440 (N_1440,N_902,N_745);
or U1441 (N_1441,N_999,N_830);
nand U1442 (N_1442,N_582,N_734);
or U1443 (N_1443,N_557,N_506);
or U1444 (N_1444,N_981,N_697);
nor U1445 (N_1445,N_575,N_868);
nand U1446 (N_1446,N_531,N_768);
and U1447 (N_1447,N_681,N_848);
nand U1448 (N_1448,N_919,N_735);
nand U1449 (N_1449,N_912,N_748);
and U1450 (N_1450,N_764,N_561);
or U1451 (N_1451,N_966,N_615);
or U1452 (N_1452,N_680,N_832);
nor U1453 (N_1453,N_926,N_634);
nor U1454 (N_1454,N_509,N_904);
nand U1455 (N_1455,N_962,N_741);
or U1456 (N_1456,N_888,N_836);
and U1457 (N_1457,N_557,N_790);
and U1458 (N_1458,N_629,N_908);
or U1459 (N_1459,N_681,N_941);
or U1460 (N_1460,N_748,N_572);
xor U1461 (N_1461,N_657,N_696);
nand U1462 (N_1462,N_629,N_964);
or U1463 (N_1463,N_890,N_995);
and U1464 (N_1464,N_897,N_830);
nand U1465 (N_1465,N_853,N_586);
nor U1466 (N_1466,N_623,N_871);
and U1467 (N_1467,N_542,N_780);
and U1468 (N_1468,N_779,N_723);
and U1469 (N_1469,N_800,N_960);
or U1470 (N_1470,N_842,N_883);
nand U1471 (N_1471,N_801,N_795);
and U1472 (N_1472,N_847,N_809);
or U1473 (N_1473,N_662,N_831);
and U1474 (N_1474,N_702,N_863);
nor U1475 (N_1475,N_902,N_796);
nand U1476 (N_1476,N_863,N_777);
or U1477 (N_1477,N_630,N_904);
nor U1478 (N_1478,N_985,N_719);
and U1479 (N_1479,N_742,N_824);
or U1480 (N_1480,N_670,N_858);
nor U1481 (N_1481,N_896,N_735);
or U1482 (N_1482,N_826,N_691);
nand U1483 (N_1483,N_992,N_811);
and U1484 (N_1484,N_918,N_605);
and U1485 (N_1485,N_527,N_707);
and U1486 (N_1486,N_981,N_696);
nor U1487 (N_1487,N_522,N_752);
and U1488 (N_1488,N_776,N_678);
nor U1489 (N_1489,N_969,N_686);
or U1490 (N_1490,N_879,N_718);
nor U1491 (N_1491,N_969,N_641);
or U1492 (N_1492,N_524,N_563);
and U1493 (N_1493,N_844,N_608);
and U1494 (N_1494,N_886,N_644);
or U1495 (N_1495,N_875,N_896);
xnor U1496 (N_1496,N_605,N_725);
or U1497 (N_1497,N_876,N_642);
nor U1498 (N_1498,N_635,N_702);
nor U1499 (N_1499,N_966,N_580);
or U1500 (N_1500,N_1367,N_1410);
and U1501 (N_1501,N_1213,N_1087);
and U1502 (N_1502,N_1329,N_1337);
or U1503 (N_1503,N_1278,N_1413);
and U1504 (N_1504,N_1078,N_1046);
nor U1505 (N_1505,N_1149,N_1082);
and U1506 (N_1506,N_1028,N_1480);
nor U1507 (N_1507,N_1436,N_1336);
or U1508 (N_1508,N_1369,N_1225);
and U1509 (N_1509,N_1301,N_1447);
nand U1510 (N_1510,N_1492,N_1467);
and U1511 (N_1511,N_1152,N_1251);
or U1512 (N_1512,N_1014,N_1038);
or U1513 (N_1513,N_1274,N_1284);
and U1514 (N_1514,N_1496,N_1255);
nor U1515 (N_1515,N_1477,N_1323);
nor U1516 (N_1516,N_1299,N_1027);
and U1517 (N_1517,N_1338,N_1034);
nor U1518 (N_1518,N_1267,N_1229);
nor U1519 (N_1519,N_1228,N_1292);
nor U1520 (N_1520,N_1493,N_1384);
nor U1521 (N_1521,N_1201,N_1442);
and U1522 (N_1522,N_1309,N_1211);
or U1523 (N_1523,N_1463,N_1330);
nand U1524 (N_1524,N_1326,N_1308);
nand U1525 (N_1525,N_1091,N_1420);
nand U1526 (N_1526,N_1095,N_1187);
or U1527 (N_1527,N_1368,N_1482);
or U1528 (N_1528,N_1304,N_1281);
nor U1529 (N_1529,N_1069,N_1083);
nor U1530 (N_1530,N_1192,N_1464);
nor U1531 (N_1531,N_1489,N_1048);
nor U1532 (N_1532,N_1125,N_1448);
or U1533 (N_1533,N_1223,N_1216);
or U1534 (N_1534,N_1011,N_1212);
nand U1535 (N_1535,N_1004,N_1277);
or U1536 (N_1536,N_1075,N_1023);
or U1537 (N_1537,N_1037,N_1354);
nand U1538 (N_1538,N_1035,N_1250);
and U1539 (N_1539,N_1084,N_1065);
or U1540 (N_1540,N_1315,N_1360);
nor U1541 (N_1541,N_1389,N_1282);
nor U1542 (N_1542,N_1424,N_1425);
or U1543 (N_1543,N_1170,N_1194);
or U1544 (N_1544,N_1355,N_1172);
nand U1545 (N_1545,N_1182,N_1052);
nor U1546 (N_1546,N_1270,N_1099);
nand U1547 (N_1547,N_1268,N_1136);
nor U1548 (N_1548,N_1145,N_1141);
nor U1549 (N_1549,N_1311,N_1266);
and U1550 (N_1550,N_1321,N_1230);
xor U1551 (N_1551,N_1295,N_1407);
or U1552 (N_1552,N_1093,N_1039);
or U1553 (N_1553,N_1335,N_1332);
nand U1554 (N_1554,N_1352,N_1280);
or U1555 (N_1555,N_1422,N_1219);
nor U1556 (N_1556,N_1408,N_1426);
nor U1557 (N_1557,N_1462,N_1423);
and U1558 (N_1558,N_1207,N_1325);
nand U1559 (N_1559,N_1349,N_1409);
and U1560 (N_1560,N_1156,N_1148);
and U1561 (N_1561,N_1241,N_1001);
nor U1562 (N_1562,N_1124,N_1176);
nand U1563 (N_1563,N_1290,N_1167);
nand U1564 (N_1564,N_1179,N_1279);
and U1565 (N_1565,N_1236,N_1044);
and U1566 (N_1566,N_1071,N_1242);
nor U1567 (N_1567,N_1479,N_1066);
or U1568 (N_1568,N_1293,N_1380);
or U1569 (N_1569,N_1057,N_1262);
or U1570 (N_1570,N_1235,N_1215);
and U1571 (N_1571,N_1397,N_1399);
nand U1572 (N_1572,N_1047,N_1252);
or U1573 (N_1573,N_1025,N_1263);
xor U1574 (N_1574,N_1359,N_1395);
or U1575 (N_1575,N_1418,N_1351);
or U1576 (N_1576,N_1486,N_1246);
or U1577 (N_1577,N_1118,N_1029);
and U1578 (N_1578,N_1106,N_1112);
nand U1579 (N_1579,N_1288,N_1342);
nand U1580 (N_1580,N_1275,N_1077);
nor U1581 (N_1581,N_1319,N_1417);
or U1582 (N_1582,N_1166,N_1313);
nand U1583 (N_1583,N_1138,N_1400);
and U1584 (N_1584,N_1344,N_1440);
nor U1585 (N_1585,N_1098,N_1300);
and U1586 (N_1586,N_1457,N_1199);
and U1587 (N_1587,N_1053,N_1010);
nor U1588 (N_1588,N_1331,N_1232);
and U1589 (N_1589,N_1488,N_1161);
and U1590 (N_1590,N_1372,N_1312);
nor U1591 (N_1591,N_1238,N_1006);
or U1592 (N_1592,N_1226,N_1474);
and U1593 (N_1593,N_1155,N_1249);
xor U1594 (N_1594,N_1273,N_1364);
nor U1595 (N_1595,N_1411,N_1079);
and U1596 (N_1596,N_1348,N_1209);
nor U1597 (N_1597,N_1233,N_1195);
nand U1598 (N_1598,N_1080,N_1117);
nor U1599 (N_1599,N_1428,N_1391);
nor U1600 (N_1600,N_1345,N_1401);
nand U1601 (N_1601,N_1007,N_1473);
and U1602 (N_1602,N_1483,N_1461);
nand U1603 (N_1603,N_1013,N_1456);
nor U1604 (N_1604,N_1088,N_1198);
nor U1605 (N_1605,N_1421,N_1222);
nor U1606 (N_1606,N_1386,N_1142);
nand U1607 (N_1607,N_1185,N_1495);
and U1608 (N_1608,N_1043,N_1110);
xor U1609 (N_1609,N_1305,N_1478);
nor U1610 (N_1610,N_1020,N_1030);
nand U1611 (N_1611,N_1398,N_1476);
or U1612 (N_1612,N_1131,N_1339);
nand U1613 (N_1613,N_1024,N_1452);
nor U1614 (N_1614,N_1032,N_1294);
nand U1615 (N_1615,N_1171,N_1200);
nor U1616 (N_1616,N_1285,N_1116);
nor U1617 (N_1617,N_1427,N_1103);
or U1618 (N_1618,N_1127,N_1186);
nand U1619 (N_1619,N_1015,N_1322);
and U1620 (N_1620,N_1458,N_1143);
or U1621 (N_1621,N_1371,N_1206);
and U1622 (N_1622,N_1455,N_1049);
nand U1623 (N_1623,N_1202,N_1100);
nand U1624 (N_1624,N_1431,N_1220);
nor U1625 (N_1625,N_1434,N_1107);
or U1626 (N_1626,N_1439,N_1257);
and U1627 (N_1627,N_1302,N_1021);
nor U1628 (N_1628,N_1412,N_1113);
nand U1629 (N_1629,N_1433,N_1459);
or U1630 (N_1630,N_1494,N_1333);
nor U1631 (N_1631,N_1437,N_1260);
and U1632 (N_1632,N_1177,N_1385);
nand U1633 (N_1633,N_1314,N_1468);
nand U1634 (N_1634,N_1086,N_1383);
nand U1635 (N_1635,N_1115,N_1163);
or U1636 (N_1636,N_1231,N_1122);
and U1637 (N_1637,N_1214,N_1317);
or U1638 (N_1638,N_1221,N_1026);
or U1639 (N_1639,N_1271,N_1090);
and U1640 (N_1640,N_1050,N_1289);
nand U1641 (N_1641,N_1254,N_1296);
nand U1642 (N_1642,N_1074,N_1022);
nand U1643 (N_1643,N_1126,N_1366);
and U1644 (N_1644,N_1435,N_1162);
nor U1645 (N_1645,N_1016,N_1227);
nor U1646 (N_1646,N_1256,N_1460);
or U1647 (N_1647,N_1485,N_1160);
and U1648 (N_1648,N_1297,N_1303);
or U1649 (N_1649,N_1441,N_1390);
nor U1650 (N_1650,N_1076,N_1341);
or U1651 (N_1651,N_1188,N_1060);
nor U1652 (N_1652,N_1217,N_1358);
and U1653 (N_1653,N_1475,N_1340);
nor U1654 (N_1654,N_1361,N_1183);
nor U1655 (N_1655,N_1490,N_1153);
nand U1656 (N_1656,N_1133,N_1324);
and U1657 (N_1657,N_1234,N_1184);
and U1658 (N_1658,N_1276,N_1101);
or U1659 (N_1659,N_1469,N_1119);
and U1660 (N_1660,N_1283,N_1328);
or U1661 (N_1661,N_1144,N_1287);
nand U1662 (N_1662,N_1405,N_1121);
nand U1663 (N_1663,N_1362,N_1002);
and U1664 (N_1664,N_1062,N_1193);
nor U1665 (N_1665,N_1291,N_1416);
nor U1666 (N_1666,N_1393,N_1406);
nor U1667 (N_1667,N_1253,N_1269);
nor U1668 (N_1668,N_1146,N_1097);
or U1669 (N_1669,N_1379,N_1239);
nand U1670 (N_1670,N_1140,N_1123);
or U1671 (N_1671,N_1111,N_1104);
nor U1672 (N_1672,N_1147,N_1438);
nor U1673 (N_1673,N_1208,N_1357);
or U1674 (N_1674,N_1003,N_1108);
and U1675 (N_1675,N_1120,N_1033);
nor U1676 (N_1676,N_1472,N_1174);
nor U1677 (N_1677,N_1055,N_1382);
nor U1678 (N_1678,N_1307,N_1353);
nand U1679 (N_1679,N_1081,N_1102);
and U1680 (N_1680,N_1205,N_1135);
nand U1681 (N_1681,N_1471,N_1210);
nand U1682 (N_1682,N_1134,N_1224);
nand U1683 (N_1683,N_1310,N_1491);
nand U1684 (N_1684,N_1012,N_1068);
nand U1685 (N_1685,N_1388,N_1036);
or U1686 (N_1686,N_1403,N_1168);
or U1687 (N_1687,N_1430,N_1072);
or U1688 (N_1688,N_1204,N_1350);
nor U1689 (N_1689,N_1085,N_1445);
or U1690 (N_1690,N_1306,N_1094);
and U1691 (N_1691,N_1443,N_1203);
nor U1692 (N_1692,N_1320,N_1031);
nand U1693 (N_1693,N_1392,N_1181);
or U1694 (N_1694,N_1114,N_1197);
and U1695 (N_1695,N_1157,N_1404);
nor U1696 (N_1696,N_1040,N_1466);
or U1697 (N_1697,N_1298,N_1096);
and U1698 (N_1698,N_1465,N_1247);
or U1699 (N_1699,N_1377,N_1394);
xnor U1700 (N_1700,N_1240,N_1154);
nor U1701 (N_1701,N_1061,N_1381);
nand U1702 (N_1702,N_1419,N_1180);
nand U1703 (N_1703,N_1451,N_1376);
and U1704 (N_1704,N_1244,N_1196);
nor U1705 (N_1705,N_1158,N_1334);
or U1706 (N_1706,N_1051,N_1058);
and U1707 (N_1707,N_1432,N_1487);
or U1708 (N_1708,N_1092,N_1045);
and U1709 (N_1709,N_1370,N_1054);
nand U1710 (N_1710,N_1005,N_1259);
nor U1711 (N_1711,N_1318,N_1137);
nand U1712 (N_1712,N_1316,N_1173);
and U1713 (N_1713,N_1258,N_1446);
and U1714 (N_1714,N_1150,N_1165);
and U1715 (N_1715,N_1499,N_1063);
nand U1716 (N_1716,N_1415,N_1450);
nor U1717 (N_1717,N_1059,N_1132);
nand U1718 (N_1718,N_1151,N_1265);
or U1719 (N_1719,N_1105,N_1129);
and U1720 (N_1720,N_1041,N_1008);
nor U1721 (N_1721,N_1286,N_1089);
nor U1722 (N_1722,N_1414,N_1237);
nor U1723 (N_1723,N_1378,N_1128);
or U1724 (N_1724,N_1272,N_1190);
xor U1725 (N_1725,N_1363,N_1017);
nor U1726 (N_1726,N_1139,N_1327);
and U1727 (N_1727,N_1009,N_1454);
and U1728 (N_1728,N_1449,N_1164);
nand U1729 (N_1729,N_1073,N_1064);
or U1730 (N_1730,N_1264,N_1056);
nor U1731 (N_1731,N_1453,N_1484);
nor U1732 (N_1732,N_1243,N_1396);
nor U1733 (N_1733,N_1387,N_1191);
nand U1734 (N_1734,N_1042,N_1429);
or U1735 (N_1735,N_1248,N_1019);
xnor U1736 (N_1736,N_1373,N_1159);
or U1737 (N_1737,N_1130,N_1444);
and U1738 (N_1738,N_1343,N_1497);
xor U1739 (N_1739,N_1189,N_1374);
nand U1740 (N_1740,N_1169,N_1018);
nand U1741 (N_1741,N_1356,N_1375);
nand U1742 (N_1742,N_1175,N_1067);
nand U1743 (N_1743,N_1365,N_1470);
nor U1744 (N_1744,N_1402,N_1245);
and U1745 (N_1745,N_1070,N_1346);
nand U1746 (N_1746,N_1109,N_1347);
or U1747 (N_1747,N_1000,N_1498);
xnor U1748 (N_1748,N_1218,N_1481);
and U1749 (N_1749,N_1178,N_1261);
or U1750 (N_1750,N_1075,N_1318);
or U1751 (N_1751,N_1245,N_1098);
xnor U1752 (N_1752,N_1451,N_1084);
nor U1753 (N_1753,N_1362,N_1158);
nor U1754 (N_1754,N_1431,N_1459);
or U1755 (N_1755,N_1017,N_1090);
nor U1756 (N_1756,N_1170,N_1398);
and U1757 (N_1757,N_1023,N_1004);
and U1758 (N_1758,N_1252,N_1449);
nand U1759 (N_1759,N_1097,N_1413);
or U1760 (N_1760,N_1304,N_1289);
and U1761 (N_1761,N_1191,N_1235);
nor U1762 (N_1762,N_1251,N_1208);
and U1763 (N_1763,N_1032,N_1239);
nand U1764 (N_1764,N_1412,N_1489);
and U1765 (N_1765,N_1250,N_1351);
nand U1766 (N_1766,N_1051,N_1409);
or U1767 (N_1767,N_1494,N_1284);
nor U1768 (N_1768,N_1295,N_1204);
or U1769 (N_1769,N_1276,N_1372);
or U1770 (N_1770,N_1095,N_1214);
and U1771 (N_1771,N_1476,N_1487);
nand U1772 (N_1772,N_1117,N_1057);
nor U1773 (N_1773,N_1049,N_1460);
nor U1774 (N_1774,N_1287,N_1498);
nor U1775 (N_1775,N_1357,N_1138);
nand U1776 (N_1776,N_1273,N_1496);
nor U1777 (N_1777,N_1306,N_1402);
nand U1778 (N_1778,N_1096,N_1320);
or U1779 (N_1779,N_1272,N_1386);
nand U1780 (N_1780,N_1341,N_1132);
and U1781 (N_1781,N_1080,N_1199);
nor U1782 (N_1782,N_1467,N_1051);
nor U1783 (N_1783,N_1015,N_1440);
xnor U1784 (N_1784,N_1318,N_1367);
or U1785 (N_1785,N_1059,N_1269);
nor U1786 (N_1786,N_1223,N_1157);
nand U1787 (N_1787,N_1253,N_1319);
nor U1788 (N_1788,N_1158,N_1343);
and U1789 (N_1789,N_1482,N_1410);
and U1790 (N_1790,N_1208,N_1478);
nor U1791 (N_1791,N_1046,N_1329);
and U1792 (N_1792,N_1129,N_1360);
and U1793 (N_1793,N_1278,N_1449);
nand U1794 (N_1794,N_1458,N_1146);
or U1795 (N_1795,N_1152,N_1144);
nor U1796 (N_1796,N_1151,N_1307);
nand U1797 (N_1797,N_1261,N_1128);
nor U1798 (N_1798,N_1133,N_1127);
nand U1799 (N_1799,N_1118,N_1085);
nor U1800 (N_1800,N_1001,N_1004);
or U1801 (N_1801,N_1144,N_1161);
nand U1802 (N_1802,N_1135,N_1071);
or U1803 (N_1803,N_1442,N_1095);
nor U1804 (N_1804,N_1156,N_1036);
and U1805 (N_1805,N_1305,N_1411);
and U1806 (N_1806,N_1105,N_1416);
and U1807 (N_1807,N_1141,N_1370);
and U1808 (N_1808,N_1301,N_1422);
nand U1809 (N_1809,N_1189,N_1036);
and U1810 (N_1810,N_1250,N_1254);
and U1811 (N_1811,N_1347,N_1230);
and U1812 (N_1812,N_1343,N_1325);
and U1813 (N_1813,N_1058,N_1309);
and U1814 (N_1814,N_1134,N_1146);
nor U1815 (N_1815,N_1272,N_1047);
and U1816 (N_1816,N_1100,N_1057);
and U1817 (N_1817,N_1086,N_1405);
and U1818 (N_1818,N_1064,N_1323);
nand U1819 (N_1819,N_1080,N_1234);
nand U1820 (N_1820,N_1247,N_1306);
or U1821 (N_1821,N_1289,N_1023);
or U1822 (N_1822,N_1220,N_1134);
and U1823 (N_1823,N_1435,N_1118);
or U1824 (N_1824,N_1018,N_1383);
nor U1825 (N_1825,N_1063,N_1247);
or U1826 (N_1826,N_1314,N_1198);
or U1827 (N_1827,N_1304,N_1247);
or U1828 (N_1828,N_1248,N_1405);
nor U1829 (N_1829,N_1086,N_1477);
and U1830 (N_1830,N_1374,N_1265);
or U1831 (N_1831,N_1370,N_1358);
nand U1832 (N_1832,N_1053,N_1001);
and U1833 (N_1833,N_1454,N_1133);
nor U1834 (N_1834,N_1451,N_1127);
nor U1835 (N_1835,N_1160,N_1278);
and U1836 (N_1836,N_1411,N_1180);
nor U1837 (N_1837,N_1092,N_1196);
nor U1838 (N_1838,N_1161,N_1481);
or U1839 (N_1839,N_1316,N_1283);
or U1840 (N_1840,N_1020,N_1270);
or U1841 (N_1841,N_1041,N_1487);
nand U1842 (N_1842,N_1393,N_1416);
or U1843 (N_1843,N_1350,N_1213);
xnor U1844 (N_1844,N_1194,N_1237);
nand U1845 (N_1845,N_1407,N_1294);
or U1846 (N_1846,N_1239,N_1232);
nand U1847 (N_1847,N_1284,N_1381);
or U1848 (N_1848,N_1209,N_1489);
or U1849 (N_1849,N_1285,N_1083);
nor U1850 (N_1850,N_1098,N_1379);
nor U1851 (N_1851,N_1186,N_1082);
nand U1852 (N_1852,N_1087,N_1090);
or U1853 (N_1853,N_1074,N_1020);
and U1854 (N_1854,N_1260,N_1193);
nor U1855 (N_1855,N_1081,N_1120);
or U1856 (N_1856,N_1174,N_1382);
and U1857 (N_1857,N_1369,N_1107);
xnor U1858 (N_1858,N_1189,N_1468);
or U1859 (N_1859,N_1158,N_1374);
or U1860 (N_1860,N_1178,N_1427);
or U1861 (N_1861,N_1180,N_1152);
or U1862 (N_1862,N_1309,N_1272);
nand U1863 (N_1863,N_1478,N_1420);
or U1864 (N_1864,N_1087,N_1448);
nand U1865 (N_1865,N_1177,N_1336);
and U1866 (N_1866,N_1486,N_1204);
and U1867 (N_1867,N_1498,N_1311);
or U1868 (N_1868,N_1005,N_1175);
nand U1869 (N_1869,N_1016,N_1106);
nand U1870 (N_1870,N_1116,N_1000);
or U1871 (N_1871,N_1381,N_1252);
or U1872 (N_1872,N_1296,N_1208);
or U1873 (N_1873,N_1434,N_1058);
nor U1874 (N_1874,N_1452,N_1014);
or U1875 (N_1875,N_1129,N_1003);
nand U1876 (N_1876,N_1435,N_1261);
and U1877 (N_1877,N_1109,N_1034);
nand U1878 (N_1878,N_1287,N_1142);
nor U1879 (N_1879,N_1332,N_1499);
and U1880 (N_1880,N_1361,N_1248);
or U1881 (N_1881,N_1207,N_1343);
nor U1882 (N_1882,N_1193,N_1285);
nor U1883 (N_1883,N_1162,N_1429);
nand U1884 (N_1884,N_1065,N_1301);
nor U1885 (N_1885,N_1122,N_1461);
nor U1886 (N_1886,N_1328,N_1336);
nor U1887 (N_1887,N_1068,N_1452);
nand U1888 (N_1888,N_1007,N_1213);
and U1889 (N_1889,N_1257,N_1168);
or U1890 (N_1890,N_1078,N_1408);
and U1891 (N_1891,N_1034,N_1207);
xor U1892 (N_1892,N_1262,N_1042);
xor U1893 (N_1893,N_1021,N_1230);
nand U1894 (N_1894,N_1011,N_1098);
nor U1895 (N_1895,N_1222,N_1224);
or U1896 (N_1896,N_1029,N_1363);
and U1897 (N_1897,N_1444,N_1143);
or U1898 (N_1898,N_1411,N_1333);
nor U1899 (N_1899,N_1362,N_1393);
nor U1900 (N_1900,N_1174,N_1365);
nand U1901 (N_1901,N_1161,N_1316);
or U1902 (N_1902,N_1052,N_1141);
or U1903 (N_1903,N_1334,N_1474);
nor U1904 (N_1904,N_1149,N_1193);
nor U1905 (N_1905,N_1149,N_1225);
and U1906 (N_1906,N_1124,N_1471);
nor U1907 (N_1907,N_1367,N_1415);
xor U1908 (N_1908,N_1017,N_1071);
nand U1909 (N_1909,N_1366,N_1277);
nor U1910 (N_1910,N_1076,N_1166);
nand U1911 (N_1911,N_1344,N_1492);
nand U1912 (N_1912,N_1373,N_1417);
xnor U1913 (N_1913,N_1487,N_1468);
and U1914 (N_1914,N_1156,N_1479);
nor U1915 (N_1915,N_1409,N_1294);
or U1916 (N_1916,N_1292,N_1192);
nor U1917 (N_1917,N_1213,N_1084);
or U1918 (N_1918,N_1158,N_1076);
nor U1919 (N_1919,N_1494,N_1488);
or U1920 (N_1920,N_1021,N_1332);
nand U1921 (N_1921,N_1267,N_1442);
and U1922 (N_1922,N_1393,N_1117);
and U1923 (N_1923,N_1467,N_1347);
and U1924 (N_1924,N_1370,N_1479);
or U1925 (N_1925,N_1402,N_1261);
nand U1926 (N_1926,N_1453,N_1074);
or U1927 (N_1927,N_1256,N_1322);
xor U1928 (N_1928,N_1464,N_1491);
or U1929 (N_1929,N_1132,N_1447);
nor U1930 (N_1930,N_1193,N_1390);
nand U1931 (N_1931,N_1322,N_1198);
or U1932 (N_1932,N_1358,N_1211);
nand U1933 (N_1933,N_1067,N_1141);
nand U1934 (N_1934,N_1309,N_1333);
nor U1935 (N_1935,N_1157,N_1435);
and U1936 (N_1936,N_1287,N_1472);
nand U1937 (N_1937,N_1335,N_1484);
or U1938 (N_1938,N_1205,N_1401);
and U1939 (N_1939,N_1461,N_1238);
nor U1940 (N_1940,N_1389,N_1377);
and U1941 (N_1941,N_1442,N_1106);
nand U1942 (N_1942,N_1276,N_1474);
and U1943 (N_1943,N_1257,N_1419);
nor U1944 (N_1944,N_1095,N_1217);
and U1945 (N_1945,N_1265,N_1252);
or U1946 (N_1946,N_1209,N_1393);
and U1947 (N_1947,N_1170,N_1157);
nand U1948 (N_1948,N_1282,N_1274);
nor U1949 (N_1949,N_1457,N_1315);
nand U1950 (N_1950,N_1404,N_1291);
nor U1951 (N_1951,N_1447,N_1006);
nor U1952 (N_1952,N_1117,N_1455);
nand U1953 (N_1953,N_1187,N_1228);
and U1954 (N_1954,N_1210,N_1158);
nand U1955 (N_1955,N_1360,N_1479);
and U1956 (N_1956,N_1240,N_1270);
or U1957 (N_1957,N_1477,N_1094);
and U1958 (N_1958,N_1352,N_1219);
nand U1959 (N_1959,N_1334,N_1145);
and U1960 (N_1960,N_1474,N_1358);
nor U1961 (N_1961,N_1424,N_1168);
nor U1962 (N_1962,N_1483,N_1255);
nand U1963 (N_1963,N_1151,N_1204);
and U1964 (N_1964,N_1064,N_1362);
and U1965 (N_1965,N_1311,N_1263);
and U1966 (N_1966,N_1393,N_1137);
nor U1967 (N_1967,N_1103,N_1328);
nor U1968 (N_1968,N_1018,N_1206);
or U1969 (N_1969,N_1486,N_1050);
nand U1970 (N_1970,N_1057,N_1234);
or U1971 (N_1971,N_1398,N_1238);
or U1972 (N_1972,N_1427,N_1411);
nand U1973 (N_1973,N_1462,N_1155);
and U1974 (N_1974,N_1184,N_1395);
and U1975 (N_1975,N_1159,N_1193);
and U1976 (N_1976,N_1424,N_1056);
or U1977 (N_1977,N_1070,N_1215);
nor U1978 (N_1978,N_1100,N_1262);
and U1979 (N_1979,N_1493,N_1449);
and U1980 (N_1980,N_1048,N_1105);
nand U1981 (N_1981,N_1180,N_1257);
or U1982 (N_1982,N_1173,N_1407);
and U1983 (N_1983,N_1038,N_1463);
nor U1984 (N_1984,N_1070,N_1365);
or U1985 (N_1985,N_1007,N_1055);
or U1986 (N_1986,N_1462,N_1010);
nand U1987 (N_1987,N_1474,N_1043);
or U1988 (N_1988,N_1475,N_1031);
and U1989 (N_1989,N_1364,N_1402);
or U1990 (N_1990,N_1321,N_1168);
and U1991 (N_1991,N_1497,N_1107);
nor U1992 (N_1992,N_1459,N_1158);
or U1993 (N_1993,N_1014,N_1001);
nor U1994 (N_1994,N_1431,N_1332);
nor U1995 (N_1995,N_1288,N_1198);
xnor U1996 (N_1996,N_1312,N_1455);
nor U1997 (N_1997,N_1319,N_1284);
or U1998 (N_1998,N_1362,N_1045);
or U1999 (N_1999,N_1210,N_1382);
and U2000 (N_2000,N_1808,N_1908);
nand U2001 (N_2001,N_1547,N_1559);
nor U2002 (N_2002,N_1819,N_1974);
xnor U2003 (N_2003,N_1615,N_1922);
nor U2004 (N_2004,N_1971,N_1569);
nor U2005 (N_2005,N_1895,N_1620);
nand U2006 (N_2006,N_1767,N_1768);
nand U2007 (N_2007,N_1683,N_1590);
and U2008 (N_2008,N_1600,N_1891);
and U2009 (N_2009,N_1554,N_1715);
or U2010 (N_2010,N_1713,N_1961);
or U2011 (N_2011,N_1560,N_1950);
and U2012 (N_2012,N_1953,N_1704);
or U2013 (N_2013,N_1501,N_1697);
nor U2014 (N_2014,N_1770,N_1913);
and U2015 (N_2015,N_1845,N_1956);
nor U2016 (N_2016,N_1938,N_1840);
and U2017 (N_2017,N_1849,N_1670);
nor U2018 (N_2018,N_1608,N_1835);
nand U2019 (N_2019,N_1698,N_1717);
nand U2020 (N_2020,N_1732,N_1576);
nand U2021 (N_2021,N_1542,N_1662);
nand U2022 (N_2022,N_1567,N_1869);
nor U2023 (N_2023,N_1563,N_1759);
nand U2024 (N_2024,N_1667,N_1730);
or U2025 (N_2025,N_1774,N_1657);
nand U2026 (N_2026,N_1788,N_1694);
nand U2027 (N_2027,N_1613,N_1976);
nor U2028 (N_2028,N_1955,N_1844);
nor U2029 (N_2029,N_1733,N_1902);
nand U2030 (N_2030,N_1512,N_1872);
nand U2031 (N_2031,N_1566,N_1828);
nand U2032 (N_2032,N_1957,N_1843);
and U2033 (N_2033,N_1644,N_1522);
nand U2034 (N_2034,N_1777,N_1500);
nand U2035 (N_2035,N_1734,N_1538);
nand U2036 (N_2036,N_1751,N_1896);
nand U2037 (N_2037,N_1959,N_1886);
and U2038 (N_2038,N_1791,N_1612);
nor U2039 (N_2039,N_1518,N_1665);
and U2040 (N_2040,N_1664,N_1766);
and U2041 (N_2041,N_1632,N_1607);
or U2042 (N_2042,N_1631,N_1626);
nand U2043 (N_2043,N_1932,N_1969);
nand U2044 (N_2044,N_1963,N_1858);
and U2045 (N_2045,N_1830,N_1943);
nand U2046 (N_2046,N_1634,N_1760);
nor U2047 (N_2047,N_1682,N_1823);
nand U2048 (N_2048,N_1594,N_1587);
nor U2049 (N_2049,N_1786,N_1985);
nand U2050 (N_2050,N_1841,N_1801);
nand U2051 (N_2051,N_1978,N_1562);
and U2052 (N_2052,N_1710,N_1649);
or U2053 (N_2053,N_1919,N_1750);
or U2054 (N_2054,N_1848,N_1584);
xor U2055 (N_2055,N_1601,N_1537);
and U2056 (N_2056,N_1866,N_1528);
nor U2057 (N_2057,N_1889,N_1701);
and U2058 (N_2058,N_1689,N_1784);
nor U2059 (N_2059,N_1894,N_1806);
or U2060 (N_2060,N_1812,N_1571);
nor U2061 (N_2061,N_1755,N_1602);
and U2062 (N_2062,N_1946,N_1930);
nand U2063 (N_2063,N_1671,N_1720);
nor U2064 (N_2064,N_1798,N_1761);
and U2065 (N_2065,N_1785,N_1965);
nand U2066 (N_2066,N_1882,N_1708);
xnor U2067 (N_2067,N_1673,N_1624);
or U2068 (N_2068,N_1857,N_1826);
or U2069 (N_2069,N_1931,N_1979);
or U2070 (N_2070,N_1980,N_1599);
nor U2071 (N_2071,N_1617,N_1749);
and U2072 (N_2072,N_1853,N_1964);
nand U2073 (N_2073,N_1593,N_1691);
nand U2074 (N_2074,N_1640,N_1807);
nand U2075 (N_2075,N_1941,N_1577);
and U2076 (N_2076,N_1570,N_1778);
and U2077 (N_2077,N_1877,N_1868);
and U2078 (N_2078,N_1609,N_1970);
and U2079 (N_2079,N_1502,N_1592);
nand U2080 (N_2080,N_1532,N_1842);
or U2081 (N_2081,N_1580,N_1833);
or U2082 (N_2082,N_1586,N_1516);
or U2083 (N_2083,N_1897,N_1523);
nor U2084 (N_2084,N_1944,N_1513);
nor U2085 (N_2085,N_1771,N_1925);
or U2086 (N_2086,N_1503,N_1918);
nor U2087 (N_2087,N_1635,N_1529);
or U2088 (N_2088,N_1796,N_1727);
or U2089 (N_2089,N_1954,N_1616);
nor U2090 (N_2090,N_1747,N_1817);
nor U2091 (N_2091,N_1890,N_1618);
nor U2092 (N_2092,N_1669,N_1805);
and U2093 (N_2093,N_1934,N_1765);
nand U2094 (N_2094,N_1831,N_1726);
nand U2095 (N_2095,N_1855,N_1706);
nor U2096 (N_2096,N_1596,N_1851);
nand U2097 (N_2097,N_1573,N_1905);
nor U2098 (N_2098,N_1914,N_1824);
and U2099 (N_2099,N_1993,N_1642);
or U2100 (N_2100,N_1827,N_1603);
nor U2101 (N_2101,N_1816,N_1790);
or U2102 (N_2102,N_1783,N_1832);
or U2103 (N_2103,N_1546,N_1743);
and U2104 (N_2104,N_1935,N_1893);
nand U2105 (N_2105,N_1703,N_1535);
nor U2106 (N_2106,N_1622,N_1575);
or U2107 (N_2107,N_1994,N_1507);
and U2108 (N_2108,N_1531,N_1850);
and U2109 (N_2109,N_1558,N_1709);
and U2110 (N_2110,N_1654,N_1929);
nor U2111 (N_2111,N_1621,N_1863);
nor U2112 (N_2112,N_1779,N_1822);
nor U2113 (N_2113,N_1782,N_1677);
nor U2114 (N_2114,N_1773,N_1888);
and U2115 (N_2115,N_1564,N_1880);
nor U2116 (N_2116,N_1619,N_1871);
and U2117 (N_2117,N_1721,N_1948);
or U2118 (N_2118,N_1638,N_1656);
nand U2119 (N_2119,N_1561,N_1643);
nand U2120 (N_2120,N_1763,N_1998);
and U2121 (N_2121,N_1658,N_1627);
nor U2122 (N_2122,N_1937,N_1539);
and U2123 (N_2123,N_1676,N_1983);
and U2124 (N_2124,N_1879,N_1942);
and U2125 (N_2125,N_1549,N_1860);
nor U2126 (N_2126,N_1764,N_1614);
and U2127 (N_2127,N_1520,N_1544);
nand U2128 (N_2128,N_1996,N_1829);
or U2129 (N_2129,N_1949,N_1591);
and U2130 (N_2130,N_1920,N_1967);
or U2131 (N_2131,N_1675,N_1525);
and U2132 (N_2132,N_1540,N_1655);
nor U2133 (N_2133,N_1981,N_1916);
nand U2134 (N_2134,N_1506,N_1728);
or U2135 (N_2135,N_1997,N_1668);
and U2136 (N_2136,N_1660,N_1659);
or U2137 (N_2137,N_1991,N_1637);
and U2138 (N_2138,N_1821,N_1725);
or U2139 (N_2139,N_1722,N_1737);
nor U2140 (N_2140,N_1688,N_1907);
nand U2141 (N_2141,N_1530,N_1510);
or U2142 (N_2142,N_1511,N_1636);
or U2143 (N_2143,N_1903,N_1555);
nor U2144 (N_2144,N_1702,N_1952);
xnor U2145 (N_2145,N_1611,N_1864);
nand U2146 (N_2146,N_1958,N_1986);
nor U2147 (N_2147,N_1776,N_1738);
nand U2148 (N_2148,N_1606,N_1742);
nand U2149 (N_2149,N_1692,N_1900);
or U2150 (N_2150,N_1973,N_1653);
or U2151 (N_2151,N_1666,N_1705);
nor U2152 (N_2152,N_1582,N_1686);
nand U2153 (N_2153,N_1909,N_1651);
or U2154 (N_2154,N_1984,N_1881);
nand U2155 (N_2155,N_1536,N_1945);
and U2156 (N_2156,N_1574,N_1815);
nand U2157 (N_2157,N_1533,N_1859);
nor U2158 (N_2158,N_1792,N_1543);
or U2159 (N_2159,N_1534,N_1975);
and U2160 (N_2160,N_1820,N_1565);
nand U2161 (N_2161,N_1678,N_1700);
nor U2162 (N_2162,N_1699,N_1794);
or U2163 (N_2163,N_1995,N_1521);
nand U2164 (N_2164,N_1524,N_1878);
or U2165 (N_2165,N_1847,N_1772);
nand U2166 (N_2166,N_1723,N_1797);
nand U2167 (N_2167,N_1505,N_1923);
nor U2168 (N_2168,N_1745,N_1757);
nand U2169 (N_2169,N_1517,N_1679);
or U2170 (N_2170,N_1579,N_1589);
nand U2171 (N_2171,N_1799,N_1646);
nand U2172 (N_2172,N_1989,N_1527);
nor U2173 (N_2173,N_1610,N_1597);
and U2174 (N_2174,N_1652,N_1548);
nand U2175 (N_2175,N_1865,N_1924);
or U2176 (N_2176,N_1813,N_1837);
and U2177 (N_2177,N_1598,N_1883);
and U2178 (N_2178,N_1718,N_1867);
nand U2179 (N_2179,N_1650,N_1901);
nand U2180 (N_2180,N_1625,N_1982);
or U2181 (N_2181,N_1514,N_1758);
or U2182 (N_2182,N_1556,N_1545);
or U2183 (N_2183,N_1623,N_1836);
and U2184 (N_2184,N_1707,N_1787);
and U2185 (N_2185,N_1680,N_1695);
nand U2186 (N_2186,N_1581,N_1892);
or U2187 (N_2187,N_1648,N_1585);
or U2188 (N_2188,N_1915,N_1551);
nand U2189 (N_2189,N_1809,N_1550);
nand U2190 (N_2190,N_1862,N_1939);
nand U2191 (N_2191,N_1917,N_1714);
and U2192 (N_2192,N_1693,N_1712);
nand U2193 (N_2193,N_1553,N_1663);
nor U2194 (N_2194,N_1960,N_1735);
nor U2195 (N_2195,N_1804,N_1504);
nor U2196 (N_2196,N_1748,N_1988);
nand U2197 (N_2197,N_1795,N_1852);
and U2198 (N_2198,N_1854,N_1936);
and U2199 (N_2199,N_1887,N_1927);
nand U2200 (N_2200,N_1789,N_1933);
or U2201 (N_2201,N_1838,N_1793);
or U2202 (N_2202,N_1912,N_1834);
nand U2203 (N_2203,N_1861,N_1741);
or U2204 (N_2204,N_1595,N_1899);
nand U2205 (N_2205,N_1874,N_1508);
nor U2206 (N_2206,N_1810,N_1729);
nand U2207 (N_2207,N_1940,N_1769);
nor U2208 (N_2208,N_1583,N_1754);
and U2209 (N_2209,N_1696,N_1711);
nor U2210 (N_2210,N_1885,N_1674);
and U2211 (N_2211,N_1818,N_1968);
and U2212 (N_2212,N_1541,N_1781);
nor U2213 (N_2213,N_1762,N_1746);
nor U2214 (N_2214,N_1628,N_1588);
nand U2215 (N_2215,N_1681,N_1552);
or U2216 (N_2216,N_1629,N_1684);
nor U2217 (N_2217,N_1604,N_1811);
nor U2218 (N_2218,N_1724,N_1557);
or U2219 (N_2219,N_1992,N_1921);
or U2220 (N_2220,N_1962,N_1647);
nor U2221 (N_2221,N_1873,N_1633);
and U2222 (N_2222,N_1731,N_1977);
and U2223 (N_2223,N_1803,N_1875);
and U2224 (N_2224,N_1509,N_1987);
nand U2225 (N_2225,N_1578,N_1884);
or U2226 (N_2226,N_1870,N_1526);
nand U2227 (N_2227,N_1966,N_1972);
or U2228 (N_2228,N_1739,N_1572);
nor U2229 (N_2229,N_1775,N_1672);
and U2230 (N_2230,N_1802,N_1736);
or U2231 (N_2231,N_1999,N_1515);
and U2232 (N_2232,N_1814,N_1947);
or U2233 (N_2233,N_1605,N_1898);
nor U2234 (N_2234,N_1876,N_1800);
and U2235 (N_2235,N_1661,N_1690);
nand U2236 (N_2236,N_1752,N_1639);
or U2237 (N_2237,N_1856,N_1645);
nand U2238 (N_2238,N_1630,N_1568);
or U2239 (N_2239,N_1519,N_1904);
nor U2240 (N_2240,N_1716,N_1911);
and U2241 (N_2241,N_1780,N_1641);
or U2242 (N_2242,N_1740,N_1910);
nor U2243 (N_2243,N_1926,N_1951);
nand U2244 (N_2244,N_1756,N_1687);
or U2245 (N_2245,N_1753,N_1744);
or U2246 (N_2246,N_1906,N_1839);
and U2247 (N_2247,N_1928,N_1685);
and U2248 (N_2248,N_1825,N_1846);
nor U2249 (N_2249,N_1990,N_1719);
nand U2250 (N_2250,N_1737,N_1940);
or U2251 (N_2251,N_1736,N_1951);
and U2252 (N_2252,N_1691,N_1690);
xor U2253 (N_2253,N_1956,N_1967);
or U2254 (N_2254,N_1960,N_1714);
and U2255 (N_2255,N_1546,N_1505);
or U2256 (N_2256,N_1993,N_1572);
and U2257 (N_2257,N_1787,N_1853);
and U2258 (N_2258,N_1741,N_1752);
and U2259 (N_2259,N_1868,N_1817);
or U2260 (N_2260,N_1844,N_1619);
and U2261 (N_2261,N_1550,N_1953);
nor U2262 (N_2262,N_1956,N_1762);
nand U2263 (N_2263,N_1642,N_1979);
or U2264 (N_2264,N_1900,N_1864);
and U2265 (N_2265,N_1613,N_1919);
and U2266 (N_2266,N_1714,N_1616);
nand U2267 (N_2267,N_1875,N_1605);
and U2268 (N_2268,N_1884,N_1611);
or U2269 (N_2269,N_1554,N_1917);
nand U2270 (N_2270,N_1878,N_1547);
and U2271 (N_2271,N_1519,N_1603);
nor U2272 (N_2272,N_1998,N_1824);
nor U2273 (N_2273,N_1794,N_1774);
and U2274 (N_2274,N_1635,N_1815);
nor U2275 (N_2275,N_1553,N_1898);
nand U2276 (N_2276,N_1523,N_1511);
nor U2277 (N_2277,N_1910,N_1728);
xor U2278 (N_2278,N_1687,N_1535);
or U2279 (N_2279,N_1514,N_1581);
nand U2280 (N_2280,N_1707,N_1510);
and U2281 (N_2281,N_1605,N_1563);
nor U2282 (N_2282,N_1592,N_1936);
and U2283 (N_2283,N_1722,N_1876);
nor U2284 (N_2284,N_1996,N_1573);
and U2285 (N_2285,N_1734,N_1839);
or U2286 (N_2286,N_1726,N_1581);
xor U2287 (N_2287,N_1584,N_1956);
nor U2288 (N_2288,N_1764,N_1785);
nor U2289 (N_2289,N_1934,N_1559);
nand U2290 (N_2290,N_1953,N_1863);
and U2291 (N_2291,N_1984,N_1800);
or U2292 (N_2292,N_1698,N_1859);
or U2293 (N_2293,N_1583,N_1773);
xor U2294 (N_2294,N_1996,N_1697);
or U2295 (N_2295,N_1851,N_1545);
nand U2296 (N_2296,N_1930,N_1972);
nand U2297 (N_2297,N_1596,N_1928);
nor U2298 (N_2298,N_1955,N_1791);
or U2299 (N_2299,N_1732,N_1610);
nor U2300 (N_2300,N_1655,N_1976);
nor U2301 (N_2301,N_1592,N_1998);
or U2302 (N_2302,N_1692,N_1834);
or U2303 (N_2303,N_1651,N_1892);
xor U2304 (N_2304,N_1766,N_1558);
nand U2305 (N_2305,N_1872,N_1963);
or U2306 (N_2306,N_1990,N_1961);
nand U2307 (N_2307,N_1788,N_1818);
nand U2308 (N_2308,N_1625,N_1700);
or U2309 (N_2309,N_1871,N_1754);
or U2310 (N_2310,N_1545,N_1793);
nand U2311 (N_2311,N_1749,N_1951);
and U2312 (N_2312,N_1907,N_1797);
and U2313 (N_2313,N_1618,N_1944);
and U2314 (N_2314,N_1771,N_1510);
and U2315 (N_2315,N_1785,N_1657);
or U2316 (N_2316,N_1945,N_1841);
nand U2317 (N_2317,N_1792,N_1914);
and U2318 (N_2318,N_1950,N_1781);
nand U2319 (N_2319,N_1775,N_1508);
xnor U2320 (N_2320,N_1713,N_1695);
nor U2321 (N_2321,N_1698,N_1608);
and U2322 (N_2322,N_1653,N_1770);
xor U2323 (N_2323,N_1868,N_1600);
nand U2324 (N_2324,N_1844,N_1974);
nor U2325 (N_2325,N_1709,N_1633);
or U2326 (N_2326,N_1823,N_1972);
nand U2327 (N_2327,N_1798,N_1926);
and U2328 (N_2328,N_1620,N_1941);
and U2329 (N_2329,N_1509,N_1530);
and U2330 (N_2330,N_1719,N_1870);
nand U2331 (N_2331,N_1876,N_1719);
or U2332 (N_2332,N_1877,N_1724);
or U2333 (N_2333,N_1745,N_1808);
nor U2334 (N_2334,N_1945,N_1858);
xnor U2335 (N_2335,N_1717,N_1538);
and U2336 (N_2336,N_1545,N_1846);
and U2337 (N_2337,N_1785,N_1814);
and U2338 (N_2338,N_1983,N_1989);
or U2339 (N_2339,N_1767,N_1639);
and U2340 (N_2340,N_1739,N_1778);
nand U2341 (N_2341,N_1843,N_1548);
and U2342 (N_2342,N_1723,N_1520);
or U2343 (N_2343,N_1796,N_1765);
and U2344 (N_2344,N_1910,N_1523);
nor U2345 (N_2345,N_1994,N_1968);
nand U2346 (N_2346,N_1798,N_1715);
nand U2347 (N_2347,N_1934,N_1545);
or U2348 (N_2348,N_1924,N_1847);
nand U2349 (N_2349,N_1745,N_1568);
and U2350 (N_2350,N_1780,N_1712);
or U2351 (N_2351,N_1581,N_1530);
and U2352 (N_2352,N_1811,N_1572);
or U2353 (N_2353,N_1597,N_1954);
or U2354 (N_2354,N_1738,N_1549);
or U2355 (N_2355,N_1858,N_1710);
or U2356 (N_2356,N_1686,N_1744);
or U2357 (N_2357,N_1577,N_1657);
and U2358 (N_2358,N_1575,N_1682);
nor U2359 (N_2359,N_1954,N_1693);
nand U2360 (N_2360,N_1501,N_1746);
or U2361 (N_2361,N_1684,N_1879);
nor U2362 (N_2362,N_1802,N_1978);
and U2363 (N_2363,N_1991,N_1654);
nor U2364 (N_2364,N_1943,N_1532);
or U2365 (N_2365,N_1656,N_1571);
nand U2366 (N_2366,N_1609,N_1561);
and U2367 (N_2367,N_1863,N_1519);
or U2368 (N_2368,N_1677,N_1913);
and U2369 (N_2369,N_1755,N_1582);
or U2370 (N_2370,N_1520,N_1800);
and U2371 (N_2371,N_1689,N_1918);
and U2372 (N_2372,N_1811,N_1743);
and U2373 (N_2373,N_1831,N_1681);
or U2374 (N_2374,N_1654,N_1848);
or U2375 (N_2375,N_1665,N_1641);
nand U2376 (N_2376,N_1797,N_1765);
or U2377 (N_2377,N_1868,N_1671);
xor U2378 (N_2378,N_1862,N_1601);
or U2379 (N_2379,N_1682,N_1767);
nor U2380 (N_2380,N_1533,N_1861);
or U2381 (N_2381,N_1776,N_1825);
or U2382 (N_2382,N_1864,N_1672);
nor U2383 (N_2383,N_1724,N_1860);
xor U2384 (N_2384,N_1834,N_1840);
or U2385 (N_2385,N_1634,N_1799);
and U2386 (N_2386,N_1861,N_1556);
and U2387 (N_2387,N_1987,N_1947);
xor U2388 (N_2388,N_1618,N_1973);
and U2389 (N_2389,N_1916,N_1772);
nand U2390 (N_2390,N_1562,N_1969);
or U2391 (N_2391,N_1659,N_1668);
and U2392 (N_2392,N_1874,N_1517);
nor U2393 (N_2393,N_1993,N_1504);
and U2394 (N_2394,N_1747,N_1878);
nor U2395 (N_2395,N_1629,N_1706);
or U2396 (N_2396,N_1669,N_1624);
or U2397 (N_2397,N_1505,N_1806);
nor U2398 (N_2398,N_1818,N_1603);
or U2399 (N_2399,N_1715,N_1646);
and U2400 (N_2400,N_1529,N_1542);
nand U2401 (N_2401,N_1709,N_1551);
and U2402 (N_2402,N_1778,N_1742);
and U2403 (N_2403,N_1543,N_1784);
or U2404 (N_2404,N_1652,N_1651);
nand U2405 (N_2405,N_1928,N_1934);
nand U2406 (N_2406,N_1890,N_1889);
or U2407 (N_2407,N_1644,N_1607);
or U2408 (N_2408,N_1574,N_1725);
and U2409 (N_2409,N_1607,N_1795);
and U2410 (N_2410,N_1890,N_1514);
nor U2411 (N_2411,N_1613,N_1924);
or U2412 (N_2412,N_1978,N_1528);
or U2413 (N_2413,N_1989,N_1580);
or U2414 (N_2414,N_1713,N_1529);
nor U2415 (N_2415,N_1870,N_1955);
xor U2416 (N_2416,N_1505,N_1811);
nor U2417 (N_2417,N_1558,N_1955);
xnor U2418 (N_2418,N_1746,N_1527);
and U2419 (N_2419,N_1644,N_1659);
nor U2420 (N_2420,N_1604,N_1697);
nand U2421 (N_2421,N_1702,N_1967);
and U2422 (N_2422,N_1882,N_1812);
nand U2423 (N_2423,N_1691,N_1791);
nand U2424 (N_2424,N_1807,N_1888);
nor U2425 (N_2425,N_1848,N_1599);
nor U2426 (N_2426,N_1966,N_1582);
and U2427 (N_2427,N_1500,N_1875);
or U2428 (N_2428,N_1964,N_1657);
nor U2429 (N_2429,N_1982,N_1589);
or U2430 (N_2430,N_1841,N_1548);
nand U2431 (N_2431,N_1832,N_1667);
nand U2432 (N_2432,N_1813,N_1525);
nor U2433 (N_2433,N_1703,N_1649);
and U2434 (N_2434,N_1711,N_1599);
or U2435 (N_2435,N_1895,N_1801);
and U2436 (N_2436,N_1755,N_1617);
nand U2437 (N_2437,N_1864,N_1702);
nand U2438 (N_2438,N_1506,N_1752);
nand U2439 (N_2439,N_1813,N_1805);
or U2440 (N_2440,N_1836,N_1536);
nor U2441 (N_2441,N_1602,N_1921);
nor U2442 (N_2442,N_1631,N_1861);
or U2443 (N_2443,N_1667,N_1907);
and U2444 (N_2444,N_1807,N_1882);
and U2445 (N_2445,N_1607,N_1787);
or U2446 (N_2446,N_1875,N_1537);
and U2447 (N_2447,N_1878,N_1970);
or U2448 (N_2448,N_1906,N_1727);
nand U2449 (N_2449,N_1714,N_1973);
nor U2450 (N_2450,N_1930,N_1827);
xor U2451 (N_2451,N_1524,N_1639);
nor U2452 (N_2452,N_1529,N_1836);
or U2453 (N_2453,N_1613,N_1889);
nor U2454 (N_2454,N_1700,N_1765);
nor U2455 (N_2455,N_1502,N_1689);
and U2456 (N_2456,N_1868,N_1700);
nand U2457 (N_2457,N_1640,N_1923);
nor U2458 (N_2458,N_1663,N_1996);
nor U2459 (N_2459,N_1944,N_1802);
or U2460 (N_2460,N_1770,N_1717);
nor U2461 (N_2461,N_1870,N_1904);
xnor U2462 (N_2462,N_1796,N_1541);
nand U2463 (N_2463,N_1670,N_1900);
nor U2464 (N_2464,N_1867,N_1786);
or U2465 (N_2465,N_1968,N_1773);
nor U2466 (N_2466,N_1645,N_1907);
nor U2467 (N_2467,N_1644,N_1695);
nand U2468 (N_2468,N_1508,N_1644);
nand U2469 (N_2469,N_1563,N_1515);
and U2470 (N_2470,N_1743,N_1924);
nor U2471 (N_2471,N_1859,N_1834);
and U2472 (N_2472,N_1954,N_1878);
nand U2473 (N_2473,N_1832,N_1816);
or U2474 (N_2474,N_1891,N_1833);
and U2475 (N_2475,N_1923,N_1633);
or U2476 (N_2476,N_1945,N_1939);
nor U2477 (N_2477,N_1700,N_1703);
nor U2478 (N_2478,N_1963,N_1771);
or U2479 (N_2479,N_1524,N_1763);
and U2480 (N_2480,N_1532,N_1875);
or U2481 (N_2481,N_1531,N_1977);
or U2482 (N_2482,N_1736,N_1737);
nand U2483 (N_2483,N_1955,N_1853);
nor U2484 (N_2484,N_1556,N_1849);
nand U2485 (N_2485,N_1652,N_1760);
or U2486 (N_2486,N_1933,N_1778);
and U2487 (N_2487,N_1863,N_1820);
nor U2488 (N_2488,N_1614,N_1524);
xor U2489 (N_2489,N_1551,N_1985);
xor U2490 (N_2490,N_1672,N_1877);
nor U2491 (N_2491,N_1591,N_1587);
nand U2492 (N_2492,N_1865,N_1986);
and U2493 (N_2493,N_1627,N_1739);
or U2494 (N_2494,N_1977,N_1556);
or U2495 (N_2495,N_1747,N_1916);
nor U2496 (N_2496,N_1700,N_1752);
nor U2497 (N_2497,N_1884,N_1711);
and U2498 (N_2498,N_1923,N_1879);
nand U2499 (N_2499,N_1724,N_1727);
nor U2500 (N_2500,N_2389,N_2444);
and U2501 (N_2501,N_2057,N_2062);
nand U2502 (N_2502,N_2467,N_2055);
nor U2503 (N_2503,N_2319,N_2225);
nand U2504 (N_2504,N_2499,N_2068);
or U2505 (N_2505,N_2460,N_2231);
nand U2506 (N_2506,N_2164,N_2427);
nand U2507 (N_2507,N_2298,N_2259);
nor U2508 (N_2508,N_2161,N_2292);
xor U2509 (N_2509,N_2413,N_2490);
or U2510 (N_2510,N_2080,N_2311);
or U2511 (N_2511,N_2398,N_2375);
and U2512 (N_2512,N_2334,N_2027);
and U2513 (N_2513,N_2411,N_2173);
nand U2514 (N_2514,N_2123,N_2112);
nand U2515 (N_2515,N_2437,N_2064);
nand U2516 (N_2516,N_2299,N_2370);
and U2517 (N_2517,N_2442,N_2213);
nand U2518 (N_2518,N_2113,N_2354);
and U2519 (N_2519,N_2207,N_2449);
or U2520 (N_2520,N_2250,N_2122);
and U2521 (N_2521,N_2217,N_2177);
nand U2522 (N_2522,N_2220,N_2457);
or U2523 (N_2523,N_2234,N_2233);
nor U2524 (N_2524,N_2284,N_2328);
xnor U2525 (N_2525,N_2162,N_2070);
and U2526 (N_2526,N_2043,N_2422);
nand U2527 (N_2527,N_2235,N_2372);
xnor U2528 (N_2528,N_2265,N_2127);
and U2529 (N_2529,N_2324,N_2426);
nor U2530 (N_2530,N_2433,N_2380);
or U2531 (N_2531,N_2015,N_2353);
xor U2532 (N_2532,N_2039,N_2296);
or U2533 (N_2533,N_2211,N_2092);
nand U2534 (N_2534,N_2011,N_2331);
and U2535 (N_2535,N_2172,N_2240);
nor U2536 (N_2536,N_2119,N_2356);
nor U2537 (N_2537,N_2028,N_2425);
and U2538 (N_2538,N_2414,N_2218);
or U2539 (N_2539,N_2432,N_2263);
xor U2540 (N_2540,N_2362,N_2110);
nor U2541 (N_2541,N_2044,N_2190);
or U2542 (N_2542,N_2131,N_2048);
and U2543 (N_2543,N_2051,N_2232);
nor U2544 (N_2544,N_2184,N_2206);
nor U2545 (N_2545,N_2272,N_2209);
nand U2546 (N_2546,N_2087,N_2280);
xnor U2547 (N_2547,N_2321,N_2484);
and U2548 (N_2548,N_2409,N_2219);
nand U2549 (N_2549,N_2003,N_2019);
nor U2550 (N_2550,N_2496,N_2060);
nand U2551 (N_2551,N_2399,N_2182);
and U2552 (N_2552,N_2320,N_2175);
and U2553 (N_2553,N_2083,N_2135);
or U2554 (N_2554,N_2315,N_2492);
nand U2555 (N_2555,N_2293,N_2483);
nand U2556 (N_2556,N_2267,N_2448);
nand U2557 (N_2557,N_2488,N_2474);
and U2558 (N_2558,N_2104,N_2487);
nor U2559 (N_2559,N_2130,N_2063);
and U2560 (N_2560,N_2037,N_2408);
or U2561 (N_2561,N_2149,N_2035);
nor U2562 (N_2562,N_2086,N_2363);
xnor U2563 (N_2563,N_2046,N_2153);
nor U2564 (N_2564,N_2374,N_2199);
nor U2565 (N_2565,N_2243,N_2029);
and U2566 (N_2566,N_2458,N_2001);
nand U2567 (N_2567,N_2106,N_2108);
nand U2568 (N_2568,N_2396,N_2438);
or U2569 (N_2569,N_2093,N_2498);
or U2570 (N_2570,N_2486,N_2283);
nand U2571 (N_2571,N_2285,N_2242);
and U2572 (N_2572,N_2383,N_2013);
nor U2573 (N_2573,N_2032,N_2024);
and U2574 (N_2574,N_2118,N_2040);
nor U2575 (N_2575,N_2270,N_2100);
nor U2576 (N_2576,N_2198,N_2203);
and U2577 (N_2577,N_2150,N_2471);
and U2578 (N_2578,N_2154,N_2452);
nor U2579 (N_2579,N_2148,N_2419);
nor U2580 (N_2580,N_2494,N_2303);
and U2581 (N_2581,N_2252,N_2288);
nor U2582 (N_2582,N_2456,N_2431);
and U2583 (N_2583,N_2407,N_2477);
or U2584 (N_2584,N_2030,N_2006);
or U2585 (N_2585,N_2287,N_2379);
nor U2586 (N_2586,N_2404,N_2215);
nor U2587 (N_2587,N_2180,N_2192);
nand U2588 (N_2588,N_2469,N_2400);
or U2589 (N_2589,N_2239,N_2273);
nand U2590 (N_2590,N_2326,N_2152);
nand U2591 (N_2591,N_2476,N_2333);
and U2592 (N_2592,N_2279,N_2406);
or U2593 (N_2593,N_2359,N_2151);
and U2594 (N_2594,N_2245,N_2481);
and U2595 (N_2595,N_2134,N_2351);
or U2596 (N_2596,N_2393,N_2138);
or U2597 (N_2597,N_2384,N_2157);
and U2598 (N_2598,N_2212,N_2202);
nand U2599 (N_2599,N_2139,N_2329);
nand U2600 (N_2600,N_2193,N_2047);
or U2601 (N_2601,N_2137,N_2171);
nor U2602 (N_2602,N_2244,N_2336);
and U2603 (N_2603,N_2294,N_2307);
xor U2604 (N_2604,N_2022,N_2446);
nand U2605 (N_2605,N_2249,N_2440);
and U2606 (N_2606,N_2185,N_2349);
nor U2607 (N_2607,N_2416,N_2126);
and U2608 (N_2608,N_2339,N_2369);
and U2609 (N_2609,N_2052,N_2365);
and U2610 (N_2610,N_2291,N_2196);
and U2611 (N_2611,N_2344,N_2313);
nor U2612 (N_2612,N_2067,N_2489);
nand U2613 (N_2613,N_2050,N_2482);
and U2614 (N_2614,N_2485,N_2247);
or U2615 (N_2615,N_2464,N_2094);
or U2616 (N_2616,N_2465,N_2392);
or U2617 (N_2617,N_2061,N_2314);
nor U2618 (N_2618,N_2306,N_2257);
nor U2619 (N_2619,N_2309,N_2065);
nand U2620 (N_2620,N_2189,N_2223);
and U2621 (N_2621,N_2268,N_2132);
nor U2622 (N_2622,N_2271,N_2376);
or U2623 (N_2623,N_2216,N_2403);
or U2624 (N_2624,N_2290,N_2114);
nand U2625 (N_2625,N_2144,N_2281);
nor U2626 (N_2626,N_2099,N_2415);
nand U2627 (N_2627,N_2274,N_2101);
or U2628 (N_2628,N_2205,N_2248);
nand U2629 (N_2629,N_2163,N_2089);
or U2630 (N_2630,N_2278,N_2420);
nand U2631 (N_2631,N_2071,N_2097);
and U2632 (N_2632,N_2221,N_2327);
nand U2633 (N_2633,N_2428,N_2178);
xnor U2634 (N_2634,N_2229,N_2165);
or U2635 (N_2635,N_2430,N_2145);
nor U2636 (N_2636,N_2227,N_2226);
and U2637 (N_2637,N_2337,N_2475);
and U2638 (N_2638,N_2125,N_2079);
xor U2639 (N_2639,N_2317,N_2010);
nand U2640 (N_2640,N_2381,N_2352);
and U2641 (N_2641,N_2002,N_2348);
nand U2642 (N_2642,N_2077,N_2045);
nor U2643 (N_2643,N_2275,N_2391);
nor U2644 (N_2644,N_2373,N_2305);
nor U2645 (N_2645,N_2423,N_2461);
or U2646 (N_2646,N_2395,N_2058);
and U2647 (N_2647,N_2147,N_2241);
or U2648 (N_2648,N_2169,N_2473);
and U2649 (N_2649,N_2136,N_2479);
nor U2650 (N_2650,N_2260,N_2269);
nor U2651 (N_2651,N_2410,N_2412);
nand U2652 (N_2652,N_2368,N_2253);
or U2653 (N_2653,N_2394,N_2088);
nor U2654 (N_2654,N_2357,N_2117);
nor U2655 (N_2655,N_2445,N_2007);
nand U2656 (N_2656,N_2124,N_2116);
or U2657 (N_2657,N_2228,N_2049);
or U2658 (N_2658,N_2159,N_2302);
xor U2659 (N_2659,N_2462,N_2386);
nor U2660 (N_2660,N_2429,N_2033);
nand U2661 (N_2661,N_2312,N_2075);
nor U2662 (N_2662,N_2170,N_2167);
or U2663 (N_2663,N_2181,N_2451);
and U2664 (N_2664,N_2168,N_2340);
and U2665 (N_2665,N_2378,N_2289);
or U2666 (N_2666,N_2085,N_2054);
and U2667 (N_2667,N_2470,N_2350);
and U2668 (N_2668,N_2053,N_2036);
and U2669 (N_2669,N_2435,N_2266);
nor U2670 (N_2670,N_2078,N_2098);
nor U2671 (N_2671,N_2323,N_2254);
or U2672 (N_2672,N_2042,N_2095);
and U2673 (N_2673,N_2264,N_2194);
or U2674 (N_2674,N_2377,N_2204);
nand U2675 (N_2675,N_2310,N_2463);
or U2676 (N_2676,N_2236,N_2120);
nand U2677 (N_2677,N_2466,N_2405);
and U2678 (N_2678,N_2166,N_2316);
nor U2679 (N_2679,N_2214,N_2069);
or U2680 (N_2680,N_2018,N_2397);
nor U2681 (N_2681,N_2238,N_2041);
nand U2682 (N_2682,N_2343,N_2197);
and U2683 (N_2683,N_2090,N_2056);
nor U2684 (N_2684,N_2364,N_2454);
or U2685 (N_2685,N_2401,N_2360);
or U2686 (N_2686,N_2308,N_2103);
nor U2687 (N_2687,N_2459,N_2129);
and U2688 (N_2688,N_2358,N_2142);
xor U2689 (N_2689,N_2318,N_2076);
nor U2690 (N_2690,N_2443,N_2439);
and U2691 (N_2691,N_2390,N_2143);
nand U2692 (N_2692,N_2478,N_2107);
nor U2693 (N_2693,N_2276,N_2332);
nand U2694 (N_2694,N_2000,N_2367);
nor U2695 (N_2695,N_2155,N_2468);
and U2696 (N_2696,N_2038,N_2347);
nor U2697 (N_2697,N_2179,N_2282);
and U2698 (N_2698,N_2251,N_2421);
or U2699 (N_2699,N_2102,N_2237);
or U2700 (N_2700,N_2210,N_2297);
and U2701 (N_2701,N_2004,N_2491);
nand U2702 (N_2702,N_2073,N_2230);
nand U2703 (N_2703,N_2186,N_2200);
or U2704 (N_2704,N_2258,N_2450);
nand U2705 (N_2705,N_2434,N_2141);
or U2706 (N_2706,N_2025,N_2341);
and U2707 (N_2707,N_2493,N_2021);
nor U2708 (N_2708,N_2081,N_2201);
nand U2709 (N_2709,N_2418,N_2330);
and U2710 (N_2710,N_2361,N_2453);
nor U2711 (N_2711,N_2074,N_2195);
and U2712 (N_2712,N_2246,N_2023);
and U2713 (N_2713,N_2277,N_2322);
and U2714 (N_2714,N_2121,N_2255);
and U2715 (N_2715,N_2455,N_2424);
and U2716 (N_2716,N_2338,N_2020);
or U2717 (N_2717,N_2441,N_2388);
or U2718 (N_2718,N_2091,N_2436);
and U2719 (N_2719,N_2188,N_2387);
nand U2720 (N_2720,N_2012,N_2224);
or U2721 (N_2721,N_2109,N_2156);
nor U2722 (N_2722,N_2497,N_2262);
xor U2723 (N_2723,N_2447,N_2261);
nand U2724 (N_2724,N_2158,N_2222);
nor U2725 (N_2725,N_2072,N_2005);
or U2726 (N_2726,N_2346,N_2146);
or U2727 (N_2727,N_2174,N_2096);
or U2728 (N_2728,N_2084,N_2480);
nand U2729 (N_2729,N_2115,N_2111);
nor U2730 (N_2730,N_2133,N_2366);
nand U2731 (N_2731,N_2325,N_2286);
and U2732 (N_2732,N_2031,N_2304);
nand U2733 (N_2733,N_2335,N_2402);
or U2734 (N_2734,N_2355,N_2183);
or U2735 (N_2735,N_2014,N_2187);
or U2736 (N_2736,N_2009,N_2256);
nor U2737 (N_2737,N_2417,N_2034);
and U2738 (N_2738,N_2495,N_2345);
or U2739 (N_2739,N_2059,N_2008);
nor U2740 (N_2740,N_2301,N_2140);
nand U2741 (N_2741,N_2472,N_2128);
or U2742 (N_2742,N_2016,N_2371);
nor U2743 (N_2743,N_2295,N_2017);
nand U2744 (N_2744,N_2208,N_2026);
nand U2745 (N_2745,N_2105,N_2342);
nand U2746 (N_2746,N_2066,N_2191);
nand U2747 (N_2747,N_2382,N_2385);
nor U2748 (N_2748,N_2300,N_2176);
or U2749 (N_2749,N_2082,N_2160);
or U2750 (N_2750,N_2139,N_2220);
nand U2751 (N_2751,N_2004,N_2231);
and U2752 (N_2752,N_2212,N_2203);
nor U2753 (N_2753,N_2481,N_2212);
or U2754 (N_2754,N_2010,N_2100);
and U2755 (N_2755,N_2327,N_2453);
nand U2756 (N_2756,N_2363,N_2397);
or U2757 (N_2757,N_2205,N_2203);
nor U2758 (N_2758,N_2137,N_2453);
nor U2759 (N_2759,N_2261,N_2149);
and U2760 (N_2760,N_2484,N_2181);
or U2761 (N_2761,N_2410,N_2470);
and U2762 (N_2762,N_2417,N_2060);
and U2763 (N_2763,N_2330,N_2359);
nand U2764 (N_2764,N_2257,N_2240);
and U2765 (N_2765,N_2093,N_2029);
nor U2766 (N_2766,N_2380,N_2390);
nand U2767 (N_2767,N_2461,N_2169);
nand U2768 (N_2768,N_2083,N_2243);
or U2769 (N_2769,N_2269,N_2335);
nand U2770 (N_2770,N_2158,N_2172);
nor U2771 (N_2771,N_2032,N_2145);
nand U2772 (N_2772,N_2252,N_2172);
or U2773 (N_2773,N_2374,N_2224);
or U2774 (N_2774,N_2277,N_2330);
xnor U2775 (N_2775,N_2473,N_2266);
nor U2776 (N_2776,N_2306,N_2344);
nor U2777 (N_2777,N_2061,N_2374);
or U2778 (N_2778,N_2083,N_2161);
and U2779 (N_2779,N_2441,N_2369);
nor U2780 (N_2780,N_2255,N_2124);
and U2781 (N_2781,N_2273,N_2082);
and U2782 (N_2782,N_2209,N_2011);
nand U2783 (N_2783,N_2142,N_2053);
nor U2784 (N_2784,N_2443,N_2265);
and U2785 (N_2785,N_2140,N_2050);
nand U2786 (N_2786,N_2213,N_2367);
and U2787 (N_2787,N_2345,N_2419);
and U2788 (N_2788,N_2190,N_2301);
and U2789 (N_2789,N_2345,N_2016);
and U2790 (N_2790,N_2313,N_2037);
and U2791 (N_2791,N_2426,N_2321);
nand U2792 (N_2792,N_2118,N_2105);
and U2793 (N_2793,N_2354,N_2083);
nor U2794 (N_2794,N_2426,N_2342);
nand U2795 (N_2795,N_2397,N_2194);
nand U2796 (N_2796,N_2490,N_2275);
or U2797 (N_2797,N_2167,N_2081);
or U2798 (N_2798,N_2176,N_2327);
nand U2799 (N_2799,N_2355,N_2384);
and U2800 (N_2800,N_2442,N_2405);
or U2801 (N_2801,N_2097,N_2286);
or U2802 (N_2802,N_2490,N_2241);
nor U2803 (N_2803,N_2416,N_2303);
nor U2804 (N_2804,N_2247,N_2425);
nor U2805 (N_2805,N_2127,N_2107);
or U2806 (N_2806,N_2098,N_2461);
or U2807 (N_2807,N_2102,N_2135);
nand U2808 (N_2808,N_2000,N_2155);
nor U2809 (N_2809,N_2295,N_2413);
nor U2810 (N_2810,N_2115,N_2085);
nand U2811 (N_2811,N_2241,N_2025);
nor U2812 (N_2812,N_2124,N_2218);
or U2813 (N_2813,N_2343,N_2492);
xnor U2814 (N_2814,N_2178,N_2418);
or U2815 (N_2815,N_2385,N_2450);
or U2816 (N_2816,N_2483,N_2141);
nor U2817 (N_2817,N_2023,N_2019);
nand U2818 (N_2818,N_2025,N_2323);
nor U2819 (N_2819,N_2413,N_2448);
nand U2820 (N_2820,N_2299,N_2347);
and U2821 (N_2821,N_2406,N_2309);
and U2822 (N_2822,N_2473,N_2271);
or U2823 (N_2823,N_2372,N_2284);
and U2824 (N_2824,N_2166,N_2089);
nand U2825 (N_2825,N_2011,N_2136);
or U2826 (N_2826,N_2389,N_2068);
nand U2827 (N_2827,N_2087,N_2365);
nor U2828 (N_2828,N_2153,N_2429);
nor U2829 (N_2829,N_2384,N_2179);
nor U2830 (N_2830,N_2299,N_2113);
and U2831 (N_2831,N_2414,N_2092);
and U2832 (N_2832,N_2414,N_2310);
or U2833 (N_2833,N_2160,N_2005);
nand U2834 (N_2834,N_2367,N_2428);
and U2835 (N_2835,N_2335,N_2135);
or U2836 (N_2836,N_2074,N_2413);
nor U2837 (N_2837,N_2108,N_2399);
or U2838 (N_2838,N_2054,N_2091);
or U2839 (N_2839,N_2255,N_2380);
or U2840 (N_2840,N_2079,N_2268);
nor U2841 (N_2841,N_2392,N_2233);
nand U2842 (N_2842,N_2169,N_2464);
and U2843 (N_2843,N_2148,N_2128);
nand U2844 (N_2844,N_2232,N_2197);
or U2845 (N_2845,N_2176,N_2151);
nand U2846 (N_2846,N_2438,N_2162);
or U2847 (N_2847,N_2065,N_2381);
and U2848 (N_2848,N_2243,N_2392);
nand U2849 (N_2849,N_2407,N_2382);
or U2850 (N_2850,N_2090,N_2327);
nand U2851 (N_2851,N_2357,N_2092);
nor U2852 (N_2852,N_2353,N_2318);
and U2853 (N_2853,N_2305,N_2095);
nor U2854 (N_2854,N_2430,N_2283);
and U2855 (N_2855,N_2158,N_2033);
nand U2856 (N_2856,N_2087,N_2243);
and U2857 (N_2857,N_2079,N_2252);
nand U2858 (N_2858,N_2043,N_2107);
and U2859 (N_2859,N_2002,N_2092);
nand U2860 (N_2860,N_2433,N_2080);
and U2861 (N_2861,N_2405,N_2005);
or U2862 (N_2862,N_2101,N_2046);
nand U2863 (N_2863,N_2455,N_2466);
and U2864 (N_2864,N_2066,N_2186);
and U2865 (N_2865,N_2395,N_2319);
or U2866 (N_2866,N_2244,N_2464);
nand U2867 (N_2867,N_2011,N_2247);
or U2868 (N_2868,N_2090,N_2318);
nand U2869 (N_2869,N_2415,N_2427);
nor U2870 (N_2870,N_2270,N_2312);
and U2871 (N_2871,N_2353,N_2128);
nor U2872 (N_2872,N_2388,N_2107);
nor U2873 (N_2873,N_2247,N_2432);
nand U2874 (N_2874,N_2142,N_2071);
nor U2875 (N_2875,N_2183,N_2035);
and U2876 (N_2876,N_2324,N_2445);
nor U2877 (N_2877,N_2436,N_2189);
or U2878 (N_2878,N_2282,N_2204);
and U2879 (N_2879,N_2293,N_2419);
and U2880 (N_2880,N_2316,N_2081);
and U2881 (N_2881,N_2074,N_2217);
or U2882 (N_2882,N_2428,N_2097);
or U2883 (N_2883,N_2374,N_2383);
and U2884 (N_2884,N_2347,N_2067);
xnor U2885 (N_2885,N_2406,N_2187);
and U2886 (N_2886,N_2216,N_2251);
nand U2887 (N_2887,N_2233,N_2452);
or U2888 (N_2888,N_2120,N_2350);
nor U2889 (N_2889,N_2440,N_2285);
or U2890 (N_2890,N_2164,N_2186);
nor U2891 (N_2891,N_2364,N_2184);
nand U2892 (N_2892,N_2473,N_2494);
nand U2893 (N_2893,N_2091,N_2410);
or U2894 (N_2894,N_2012,N_2466);
and U2895 (N_2895,N_2021,N_2172);
and U2896 (N_2896,N_2382,N_2488);
or U2897 (N_2897,N_2150,N_2384);
nand U2898 (N_2898,N_2132,N_2139);
nand U2899 (N_2899,N_2120,N_2285);
or U2900 (N_2900,N_2425,N_2038);
nor U2901 (N_2901,N_2233,N_2220);
nor U2902 (N_2902,N_2072,N_2285);
and U2903 (N_2903,N_2178,N_2024);
or U2904 (N_2904,N_2333,N_2070);
xor U2905 (N_2905,N_2399,N_2122);
and U2906 (N_2906,N_2127,N_2376);
nand U2907 (N_2907,N_2394,N_2134);
or U2908 (N_2908,N_2040,N_2158);
nor U2909 (N_2909,N_2160,N_2104);
xnor U2910 (N_2910,N_2145,N_2341);
nor U2911 (N_2911,N_2320,N_2468);
nand U2912 (N_2912,N_2307,N_2441);
nor U2913 (N_2913,N_2171,N_2009);
nand U2914 (N_2914,N_2483,N_2495);
nand U2915 (N_2915,N_2274,N_2046);
nand U2916 (N_2916,N_2383,N_2071);
nand U2917 (N_2917,N_2043,N_2365);
and U2918 (N_2918,N_2317,N_2289);
nor U2919 (N_2919,N_2210,N_2119);
or U2920 (N_2920,N_2495,N_2312);
or U2921 (N_2921,N_2118,N_2113);
or U2922 (N_2922,N_2053,N_2191);
nor U2923 (N_2923,N_2052,N_2355);
nand U2924 (N_2924,N_2074,N_2172);
nand U2925 (N_2925,N_2327,N_2333);
and U2926 (N_2926,N_2252,N_2349);
or U2927 (N_2927,N_2111,N_2016);
nand U2928 (N_2928,N_2338,N_2279);
nand U2929 (N_2929,N_2301,N_2251);
nand U2930 (N_2930,N_2056,N_2148);
or U2931 (N_2931,N_2209,N_2082);
xnor U2932 (N_2932,N_2093,N_2021);
nand U2933 (N_2933,N_2273,N_2380);
and U2934 (N_2934,N_2207,N_2229);
nand U2935 (N_2935,N_2144,N_2184);
nor U2936 (N_2936,N_2308,N_2200);
nor U2937 (N_2937,N_2067,N_2311);
and U2938 (N_2938,N_2232,N_2270);
or U2939 (N_2939,N_2144,N_2031);
or U2940 (N_2940,N_2465,N_2365);
nor U2941 (N_2941,N_2231,N_2476);
or U2942 (N_2942,N_2011,N_2070);
nand U2943 (N_2943,N_2327,N_2321);
nor U2944 (N_2944,N_2475,N_2177);
or U2945 (N_2945,N_2284,N_2199);
or U2946 (N_2946,N_2498,N_2371);
nor U2947 (N_2947,N_2283,N_2285);
nor U2948 (N_2948,N_2344,N_2284);
and U2949 (N_2949,N_2011,N_2374);
xor U2950 (N_2950,N_2264,N_2277);
nor U2951 (N_2951,N_2423,N_2064);
and U2952 (N_2952,N_2250,N_2200);
nand U2953 (N_2953,N_2326,N_2437);
or U2954 (N_2954,N_2438,N_2222);
and U2955 (N_2955,N_2356,N_2445);
nor U2956 (N_2956,N_2467,N_2239);
nand U2957 (N_2957,N_2010,N_2399);
and U2958 (N_2958,N_2054,N_2088);
and U2959 (N_2959,N_2017,N_2164);
and U2960 (N_2960,N_2093,N_2409);
nor U2961 (N_2961,N_2144,N_2252);
and U2962 (N_2962,N_2172,N_2318);
or U2963 (N_2963,N_2370,N_2045);
nand U2964 (N_2964,N_2198,N_2072);
and U2965 (N_2965,N_2431,N_2336);
or U2966 (N_2966,N_2120,N_2219);
or U2967 (N_2967,N_2134,N_2036);
or U2968 (N_2968,N_2096,N_2100);
nand U2969 (N_2969,N_2168,N_2155);
or U2970 (N_2970,N_2339,N_2219);
nor U2971 (N_2971,N_2075,N_2287);
nand U2972 (N_2972,N_2451,N_2412);
or U2973 (N_2973,N_2098,N_2387);
nor U2974 (N_2974,N_2136,N_2161);
and U2975 (N_2975,N_2091,N_2215);
nand U2976 (N_2976,N_2409,N_2423);
nand U2977 (N_2977,N_2337,N_2352);
nor U2978 (N_2978,N_2375,N_2076);
nor U2979 (N_2979,N_2289,N_2285);
nand U2980 (N_2980,N_2434,N_2067);
and U2981 (N_2981,N_2322,N_2182);
nor U2982 (N_2982,N_2017,N_2340);
nor U2983 (N_2983,N_2020,N_2307);
nor U2984 (N_2984,N_2472,N_2151);
nor U2985 (N_2985,N_2304,N_2381);
nor U2986 (N_2986,N_2306,N_2266);
or U2987 (N_2987,N_2147,N_2329);
nand U2988 (N_2988,N_2475,N_2327);
nand U2989 (N_2989,N_2434,N_2317);
nor U2990 (N_2990,N_2304,N_2152);
nor U2991 (N_2991,N_2227,N_2459);
nor U2992 (N_2992,N_2102,N_2363);
nor U2993 (N_2993,N_2162,N_2261);
nor U2994 (N_2994,N_2118,N_2223);
or U2995 (N_2995,N_2262,N_2193);
and U2996 (N_2996,N_2313,N_2338);
and U2997 (N_2997,N_2111,N_2334);
or U2998 (N_2998,N_2221,N_2044);
or U2999 (N_2999,N_2318,N_2257);
and UO_0 (O_0,N_2522,N_2730);
or UO_1 (O_1,N_2885,N_2645);
nand UO_2 (O_2,N_2923,N_2672);
xor UO_3 (O_3,N_2664,N_2627);
nor UO_4 (O_4,N_2816,N_2783);
nor UO_5 (O_5,N_2750,N_2577);
nor UO_6 (O_6,N_2640,N_2813);
nand UO_7 (O_7,N_2858,N_2963);
nand UO_8 (O_8,N_2901,N_2796);
and UO_9 (O_9,N_2652,N_2504);
and UO_10 (O_10,N_2956,N_2597);
nand UO_11 (O_11,N_2596,N_2641);
nor UO_12 (O_12,N_2784,N_2543);
or UO_13 (O_13,N_2807,N_2836);
or UO_14 (O_14,N_2718,N_2926);
and UO_15 (O_15,N_2602,N_2630);
or UO_16 (O_16,N_2567,N_2920);
and UO_17 (O_17,N_2911,N_2969);
or UO_18 (O_18,N_2695,N_2592);
and UO_19 (O_19,N_2547,N_2966);
nand UO_20 (O_20,N_2982,N_2898);
nor UO_21 (O_21,N_2626,N_2835);
nor UO_22 (O_22,N_2929,N_2746);
nor UO_23 (O_23,N_2936,N_2518);
nand UO_24 (O_24,N_2669,N_2760);
nor UO_25 (O_25,N_2874,N_2600);
and UO_26 (O_26,N_2997,N_2955);
or UO_27 (O_27,N_2551,N_2872);
and UO_28 (O_28,N_2933,N_2741);
and UO_29 (O_29,N_2771,N_2698);
nand UO_30 (O_30,N_2992,N_2527);
and UO_31 (O_31,N_2801,N_2659);
or UO_32 (O_32,N_2788,N_2749);
or UO_33 (O_33,N_2615,N_2878);
and UO_34 (O_34,N_2799,N_2800);
nand UO_35 (O_35,N_2685,N_2945);
or UO_36 (O_36,N_2703,N_2941);
and UO_37 (O_37,N_2785,N_2675);
nor UO_38 (O_38,N_2908,N_2554);
and UO_39 (O_39,N_2891,N_2570);
and UO_40 (O_40,N_2976,N_2532);
nor UO_41 (O_41,N_2866,N_2793);
and UO_42 (O_42,N_2862,N_2819);
nor UO_43 (O_43,N_2530,N_2644);
xor UO_44 (O_44,N_2617,N_2721);
xor UO_45 (O_45,N_2795,N_2505);
and UO_46 (O_46,N_2715,N_2557);
or UO_47 (O_47,N_2893,N_2754);
or UO_48 (O_48,N_2841,N_2973);
and UO_49 (O_49,N_2538,N_2745);
and UO_50 (O_50,N_2553,N_2513);
or UO_51 (O_51,N_2914,N_2631);
or UO_52 (O_52,N_2759,N_2638);
and UO_53 (O_53,N_2734,N_2616);
or UO_54 (O_54,N_2556,N_2545);
nand UO_55 (O_55,N_2896,N_2516);
nor UO_56 (O_56,N_2736,N_2886);
or UO_57 (O_57,N_2740,N_2775);
and UO_58 (O_58,N_2993,N_2681);
nand UO_59 (O_59,N_2629,N_2578);
or UO_60 (O_60,N_2880,N_2820);
nand UO_61 (O_61,N_2687,N_2852);
and UO_62 (O_62,N_2620,N_2983);
and UO_63 (O_63,N_2931,N_2562);
nand UO_64 (O_64,N_2853,N_2821);
nor UO_65 (O_65,N_2743,N_2774);
or UO_66 (O_66,N_2894,N_2833);
or UO_67 (O_67,N_2937,N_2682);
nor UO_68 (O_68,N_2815,N_2934);
nand UO_69 (O_69,N_2628,N_2728);
nand UO_70 (O_70,N_2899,N_2716);
or UO_71 (O_71,N_2526,N_2710);
and UO_72 (O_72,N_2508,N_2671);
or UO_73 (O_73,N_2599,N_2890);
and UO_74 (O_74,N_2586,N_2634);
nor UO_75 (O_75,N_2909,N_2987);
and UO_76 (O_76,N_2732,N_2849);
and UO_77 (O_77,N_2704,N_2560);
nor UO_78 (O_78,N_2758,N_2674);
nand UO_79 (O_79,N_2613,N_2524);
or UO_80 (O_80,N_2737,N_2808);
nand UO_81 (O_81,N_2763,N_2738);
nand UO_82 (O_82,N_2739,N_2789);
nor UO_83 (O_83,N_2755,N_2731);
nor UO_84 (O_84,N_2762,N_2515);
or UO_85 (O_85,N_2947,N_2855);
or UO_86 (O_86,N_2511,N_2806);
nand UO_87 (O_87,N_2552,N_2848);
or UO_88 (O_88,N_2589,N_2921);
nor UO_89 (O_89,N_2531,N_2748);
nand UO_90 (O_90,N_2618,N_2946);
nor UO_91 (O_91,N_2861,N_2830);
nor UO_92 (O_92,N_2537,N_2870);
nand UO_93 (O_93,N_2561,N_2636);
nor UO_94 (O_94,N_2601,N_2940);
nand UO_95 (O_95,N_2677,N_2847);
or UO_96 (O_96,N_2814,N_2506);
and UO_97 (O_97,N_2679,N_2998);
nand UO_98 (O_98,N_2655,N_2590);
nor UO_99 (O_99,N_2905,N_2811);
nor UO_100 (O_100,N_2544,N_2883);
and UO_101 (O_101,N_2529,N_2954);
and UO_102 (O_102,N_2643,N_2585);
or UO_103 (O_103,N_2609,N_2573);
and UO_104 (O_104,N_2792,N_2591);
and UO_105 (O_105,N_2970,N_2794);
and UO_106 (O_106,N_2781,N_2717);
and UO_107 (O_107,N_2756,N_2888);
nor UO_108 (O_108,N_2536,N_2612);
nand UO_109 (O_109,N_2680,N_2844);
and UO_110 (O_110,N_2851,N_2935);
or UO_111 (O_111,N_2660,N_2533);
and UO_112 (O_112,N_2593,N_2803);
and UO_113 (O_113,N_2744,N_2810);
or UO_114 (O_114,N_2647,N_2753);
nor UO_115 (O_115,N_2882,N_2943);
nand UO_116 (O_116,N_2957,N_2779);
nor UO_117 (O_117,N_2777,N_2824);
or UO_118 (O_118,N_2942,N_2525);
nor UO_119 (O_119,N_2869,N_2509);
nand UO_120 (O_120,N_2773,N_2925);
nor UO_121 (O_121,N_2778,N_2694);
or UO_122 (O_122,N_2879,N_2850);
and UO_123 (O_123,N_2996,N_2632);
and UO_124 (O_124,N_2598,N_2767);
nor UO_125 (O_125,N_2772,N_2594);
nand UO_126 (O_126,N_2979,N_2770);
or UO_127 (O_127,N_2892,N_2708);
or UO_128 (O_128,N_2500,N_2507);
nor UO_129 (O_129,N_2757,N_2968);
nor UO_130 (O_130,N_2826,N_2633);
and UO_131 (O_131,N_2876,N_2521);
nand UO_132 (O_132,N_2904,N_2797);
nand UO_133 (O_133,N_2606,N_2678);
and UO_134 (O_134,N_2512,N_2765);
nand UO_135 (O_135,N_2692,N_2948);
and UO_136 (O_136,N_2610,N_2981);
and UO_137 (O_137,N_2877,N_2722);
nor UO_138 (O_138,N_2686,N_2607);
or UO_139 (O_139,N_2950,N_2747);
nand UO_140 (O_140,N_2802,N_2726);
nand UO_141 (O_141,N_2702,N_2584);
and UO_142 (O_142,N_2822,N_2729);
nand UO_143 (O_143,N_2699,N_2566);
and UO_144 (O_144,N_2667,N_2574);
nor UO_145 (O_145,N_2919,N_2614);
and UO_146 (O_146,N_2523,N_2579);
xor UO_147 (O_147,N_2534,N_2838);
or UO_148 (O_148,N_2501,N_2944);
nand UO_149 (O_149,N_2520,N_2907);
nand UO_150 (O_150,N_2915,N_2875);
or UO_151 (O_151,N_2622,N_2910);
and UO_152 (O_152,N_2846,N_2528);
nor UO_153 (O_153,N_2786,N_2798);
or UO_154 (O_154,N_2690,N_2913);
or UO_155 (O_155,N_2588,N_2952);
nand UO_156 (O_156,N_2502,N_2809);
xor UO_157 (O_157,N_2790,N_2724);
or UO_158 (O_158,N_2864,N_2546);
and UO_159 (O_159,N_2999,N_2571);
and UO_160 (O_160,N_2619,N_2707);
and UO_161 (O_161,N_2766,N_2549);
nor UO_162 (O_162,N_2658,N_2696);
and UO_163 (O_163,N_2563,N_2582);
nor UO_164 (O_164,N_2568,N_2697);
or UO_165 (O_165,N_2663,N_2666);
nor UO_166 (O_166,N_2889,N_2646);
and UO_167 (O_167,N_2719,N_2662);
nor UO_168 (O_168,N_2829,N_2902);
nor UO_169 (O_169,N_2927,N_2625);
nor UO_170 (O_170,N_2576,N_2980);
or UO_171 (O_171,N_2840,N_2949);
nor UO_172 (O_172,N_2959,N_2834);
nand UO_173 (O_173,N_2654,N_2791);
nand UO_174 (O_174,N_2906,N_2986);
or UO_175 (O_175,N_2825,N_2994);
nor UO_176 (O_176,N_2742,N_2651);
and UO_177 (O_177,N_2932,N_2510);
or UO_178 (O_178,N_2550,N_2503);
nand UO_179 (O_179,N_2871,N_2706);
nand UO_180 (O_180,N_2818,N_2608);
nor UO_181 (O_181,N_2924,N_2595);
nor UO_182 (O_182,N_2564,N_2649);
and UO_183 (O_183,N_2900,N_2860);
or UO_184 (O_184,N_2723,N_2583);
and UO_185 (O_185,N_2764,N_2832);
nand UO_186 (O_186,N_2656,N_2988);
nand UO_187 (O_187,N_2958,N_2916);
or UO_188 (O_188,N_2831,N_2960);
nand UO_189 (O_189,N_2548,N_2812);
and UO_190 (O_190,N_2845,N_2642);
or UO_191 (O_191,N_2751,N_2972);
nor UO_192 (O_192,N_2676,N_2558);
and UO_193 (O_193,N_2611,N_2857);
or UO_194 (O_194,N_2856,N_2542);
nand UO_195 (O_195,N_2565,N_2701);
xnor UO_196 (O_196,N_2922,N_2668);
or UO_197 (O_197,N_2637,N_2843);
and UO_198 (O_198,N_2985,N_2962);
nor UO_199 (O_199,N_2575,N_2863);
nor UO_200 (O_200,N_2868,N_2961);
and UO_201 (O_201,N_2733,N_2714);
nand UO_202 (O_202,N_2665,N_2572);
and UO_203 (O_203,N_2768,N_2938);
and UO_204 (O_204,N_2713,N_2657);
and UO_205 (O_205,N_2842,N_2727);
xor UO_206 (O_206,N_2918,N_2804);
nand UO_207 (O_207,N_2823,N_2965);
and UO_208 (O_208,N_2624,N_2683);
or UO_209 (O_209,N_2605,N_2917);
and UO_210 (O_210,N_2604,N_2873);
nand UO_211 (O_211,N_2653,N_2897);
nand UO_212 (O_212,N_2569,N_2684);
or UO_213 (O_213,N_2971,N_2635);
and UO_214 (O_214,N_2735,N_2650);
nand UO_215 (O_215,N_2700,N_2539);
nor UO_216 (O_216,N_2514,N_2555);
and UO_217 (O_217,N_2535,N_2978);
nor UO_218 (O_218,N_2991,N_2603);
and UO_219 (O_219,N_2540,N_2517);
nor UO_220 (O_220,N_2827,N_2623);
or UO_221 (O_221,N_2580,N_2688);
or UO_222 (O_222,N_2587,N_2903);
nor UO_223 (O_223,N_2776,N_2964);
nand UO_224 (O_224,N_2705,N_2661);
nand UO_225 (O_225,N_2951,N_2828);
nand UO_226 (O_226,N_2787,N_2648);
and UO_227 (O_227,N_2928,N_2673);
or UO_228 (O_228,N_2837,N_2712);
nand UO_229 (O_229,N_2621,N_2995);
nand UO_230 (O_230,N_2817,N_2805);
nor UO_231 (O_231,N_2693,N_2974);
and UO_232 (O_232,N_2782,N_2887);
nand UO_233 (O_233,N_2581,N_2725);
or UO_234 (O_234,N_2519,N_2884);
and UO_235 (O_235,N_2709,N_2881);
and UO_236 (O_236,N_2711,N_2761);
or UO_237 (O_237,N_2691,N_2967);
or UO_238 (O_238,N_2895,N_2930);
nand UO_239 (O_239,N_2977,N_2839);
nor UO_240 (O_240,N_2865,N_2854);
nor UO_241 (O_241,N_2670,N_2689);
nor UO_242 (O_242,N_2752,N_2541);
or UO_243 (O_243,N_2859,N_2720);
or UO_244 (O_244,N_2953,N_2867);
and UO_245 (O_245,N_2639,N_2939);
nor UO_246 (O_246,N_2990,N_2912);
or UO_247 (O_247,N_2769,N_2780);
nand UO_248 (O_248,N_2989,N_2559);
and UO_249 (O_249,N_2984,N_2975);
nand UO_250 (O_250,N_2563,N_2520);
and UO_251 (O_251,N_2683,N_2620);
and UO_252 (O_252,N_2917,N_2895);
or UO_253 (O_253,N_2605,N_2801);
nand UO_254 (O_254,N_2838,N_2503);
or UO_255 (O_255,N_2595,N_2518);
nand UO_256 (O_256,N_2862,N_2934);
or UO_257 (O_257,N_2940,N_2539);
nand UO_258 (O_258,N_2710,N_2661);
or UO_259 (O_259,N_2887,N_2777);
or UO_260 (O_260,N_2730,N_2773);
and UO_261 (O_261,N_2967,N_2687);
or UO_262 (O_262,N_2875,N_2520);
and UO_263 (O_263,N_2727,N_2591);
and UO_264 (O_264,N_2602,N_2694);
or UO_265 (O_265,N_2545,N_2611);
nor UO_266 (O_266,N_2828,N_2667);
nand UO_267 (O_267,N_2970,N_2869);
and UO_268 (O_268,N_2501,N_2518);
nor UO_269 (O_269,N_2763,N_2603);
and UO_270 (O_270,N_2796,N_2662);
nand UO_271 (O_271,N_2869,N_2600);
nand UO_272 (O_272,N_2955,N_2731);
nor UO_273 (O_273,N_2723,N_2685);
nor UO_274 (O_274,N_2735,N_2713);
or UO_275 (O_275,N_2873,N_2528);
or UO_276 (O_276,N_2944,N_2854);
nor UO_277 (O_277,N_2877,N_2761);
nand UO_278 (O_278,N_2686,N_2610);
nand UO_279 (O_279,N_2913,N_2604);
nand UO_280 (O_280,N_2578,N_2944);
nand UO_281 (O_281,N_2919,N_2564);
or UO_282 (O_282,N_2694,N_2800);
nand UO_283 (O_283,N_2951,N_2860);
and UO_284 (O_284,N_2607,N_2678);
and UO_285 (O_285,N_2602,N_2990);
nand UO_286 (O_286,N_2589,N_2622);
and UO_287 (O_287,N_2768,N_2926);
nor UO_288 (O_288,N_2761,N_2927);
nand UO_289 (O_289,N_2530,N_2505);
and UO_290 (O_290,N_2560,N_2568);
or UO_291 (O_291,N_2947,N_2876);
nor UO_292 (O_292,N_2928,N_2583);
nor UO_293 (O_293,N_2693,N_2678);
and UO_294 (O_294,N_2510,N_2854);
or UO_295 (O_295,N_2936,N_2956);
or UO_296 (O_296,N_2696,N_2924);
nor UO_297 (O_297,N_2540,N_2599);
and UO_298 (O_298,N_2939,N_2970);
and UO_299 (O_299,N_2742,N_2978);
nor UO_300 (O_300,N_2835,N_2896);
nor UO_301 (O_301,N_2717,N_2670);
nor UO_302 (O_302,N_2628,N_2906);
or UO_303 (O_303,N_2701,N_2815);
or UO_304 (O_304,N_2906,N_2595);
nand UO_305 (O_305,N_2515,N_2914);
nand UO_306 (O_306,N_2539,N_2706);
nand UO_307 (O_307,N_2659,N_2658);
and UO_308 (O_308,N_2594,N_2751);
and UO_309 (O_309,N_2672,N_2860);
and UO_310 (O_310,N_2772,N_2935);
nor UO_311 (O_311,N_2809,N_2831);
nor UO_312 (O_312,N_2953,N_2922);
and UO_313 (O_313,N_2811,N_2548);
or UO_314 (O_314,N_2918,N_2807);
nor UO_315 (O_315,N_2858,N_2559);
and UO_316 (O_316,N_2811,N_2832);
and UO_317 (O_317,N_2727,N_2610);
and UO_318 (O_318,N_2866,N_2620);
nor UO_319 (O_319,N_2857,N_2967);
or UO_320 (O_320,N_2526,N_2648);
nand UO_321 (O_321,N_2903,N_2752);
nor UO_322 (O_322,N_2821,N_2899);
or UO_323 (O_323,N_2544,N_2747);
or UO_324 (O_324,N_2624,N_2533);
nand UO_325 (O_325,N_2760,N_2618);
nand UO_326 (O_326,N_2709,N_2750);
nor UO_327 (O_327,N_2596,N_2586);
nand UO_328 (O_328,N_2560,N_2519);
and UO_329 (O_329,N_2925,N_2636);
nor UO_330 (O_330,N_2787,N_2774);
or UO_331 (O_331,N_2906,N_2575);
nor UO_332 (O_332,N_2510,N_2811);
and UO_333 (O_333,N_2709,N_2849);
nor UO_334 (O_334,N_2897,N_2650);
or UO_335 (O_335,N_2721,N_2694);
nor UO_336 (O_336,N_2618,N_2531);
nand UO_337 (O_337,N_2864,N_2537);
or UO_338 (O_338,N_2545,N_2940);
nand UO_339 (O_339,N_2968,N_2979);
nand UO_340 (O_340,N_2864,N_2821);
nor UO_341 (O_341,N_2735,N_2626);
and UO_342 (O_342,N_2633,N_2765);
nand UO_343 (O_343,N_2853,N_2574);
nand UO_344 (O_344,N_2513,N_2588);
and UO_345 (O_345,N_2791,N_2825);
and UO_346 (O_346,N_2995,N_2559);
or UO_347 (O_347,N_2861,N_2869);
and UO_348 (O_348,N_2632,N_2933);
xor UO_349 (O_349,N_2532,N_2533);
and UO_350 (O_350,N_2926,N_2852);
or UO_351 (O_351,N_2971,N_2531);
nor UO_352 (O_352,N_2751,N_2984);
or UO_353 (O_353,N_2897,N_2907);
or UO_354 (O_354,N_2945,N_2708);
nor UO_355 (O_355,N_2963,N_2726);
nand UO_356 (O_356,N_2821,N_2728);
nand UO_357 (O_357,N_2571,N_2785);
nor UO_358 (O_358,N_2813,N_2587);
nand UO_359 (O_359,N_2668,N_2909);
or UO_360 (O_360,N_2936,N_2874);
xor UO_361 (O_361,N_2640,N_2713);
or UO_362 (O_362,N_2890,N_2668);
nor UO_363 (O_363,N_2825,N_2726);
nor UO_364 (O_364,N_2631,N_2712);
nand UO_365 (O_365,N_2901,N_2536);
nand UO_366 (O_366,N_2955,N_2887);
nand UO_367 (O_367,N_2677,N_2531);
or UO_368 (O_368,N_2634,N_2621);
nand UO_369 (O_369,N_2578,N_2947);
nor UO_370 (O_370,N_2597,N_2767);
and UO_371 (O_371,N_2885,N_2586);
or UO_372 (O_372,N_2810,N_2858);
and UO_373 (O_373,N_2662,N_2813);
nor UO_374 (O_374,N_2752,N_2912);
and UO_375 (O_375,N_2894,N_2924);
nor UO_376 (O_376,N_2886,N_2937);
xor UO_377 (O_377,N_2538,N_2740);
and UO_378 (O_378,N_2974,N_2892);
and UO_379 (O_379,N_2997,N_2704);
nand UO_380 (O_380,N_2790,N_2585);
nor UO_381 (O_381,N_2919,N_2682);
nand UO_382 (O_382,N_2772,N_2644);
nor UO_383 (O_383,N_2844,N_2604);
or UO_384 (O_384,N_2942,N_2755);
and UO_385 (O_385,N_2874,N_2608);
and UO_386 (O_386,N_2748,N_2537);
xnor UO_387 (O_387,N_2948,N_2858);
or UO_388 (O_388,N_2610,N_2944);
or UO_389 (O_389,N_2650,N_2886);
or UO_390 (O_390,N_2707,N_2806);
nor UO_391 (O_391,N_2722,N_2580);
and UO_392 (O_392,N_2745,N_2929);
nor UO_393 (O_393,N_2797,N_2519);
nand UO_394 (O_394,N_2775,N_2530);
and UO_395 (O_395,N_2693,N_2524);
nand UO_396 (O_396,N_2938,N_2607);
nor UO_397 (O_397,N_2976,N_2723);
or UO_398 (O_398,N_2937,N_2510);
nor UO_399 (O_399,N_2809,N_2837);
and UO_400 (O_400,N_2638,N_2831);
or UO_401 (O_401,N_2833,N_2590);
xnor UO_402 (O_402,N_2866,N_2758);
nand UO_403 (O_403,N_2800,N_2512);
nor UO_404 (O_404,N_2696,N_2800);
nor UO_405 (O_405,N_2967,N_2982);
nor UO_406 (O_406,N_2677,N_2586);
and UO_407 (O_407,N_2858,N_2922);
or UO_408 (O_408,N_2792,N_2851);
nor UO_409 (O_409,N_2917,N_2724);
nand UO_410 (O_410,N_2977,N_2633);
and UO_411 (O_411,N_2521,N_2941);
and UO_412 (O_412,N_2782,N_2855);
and UO_413 (O_413,N_2615,N_2588);
nor UO_414 (O_414,N_2573,N_2833);
nand UO_415 (O_415,N_2767,N_2545);
nor UO_416 (O_416,N_2588,N_2733);
or UO_417 (O_417,N_2705,N_2552);
xnor UO_418 (O_418,N_2706,N_2613);
xor UO_419 (O_419,N_2594,N_2664);
and UO_420 (O_420,N_2547,N_2513);
and UO_421 (O_421,N_2861,N_2640);
or UO_422 (O_422,N_2602,N_2765);
nand UO_423 (O_423,N_2621,N_2618);
nor UO_424 (O_424,N_2984,N_2927);
nand UO_425 (O_425,N_2976,N_2635);
nand UO_426 (O_426,N_2935,N_2667);
or UO_427 (O_427,N_2576,N_2521);
nor UO_428 (O_428,N_2655,N_2927);
and UO_429 (O_429,N_2931,N_2875);
nand UO_430 (O_430,N_2538,N_2828);
and UO_431 (O_431,N_2796,N_2602);
nand UO_432 (O_432,N_2847,N_2954);
nand UO_433 (O_433,N_2959,N_2680);
or UO_434 (O_434,N_2600,N_2708);
nor UO_435 (O_435,N_2993,N_2728);
nor UO_436 (O_436,N_2867,N_2983);
nand UO_437 (O_437,N_2511,N_2861);
or UO_438 (O_438,N_2682,N_2540);
nor UO_439 (O_439,N_2890,N_2994);
xor UO_440 (O_440,N_2882,N_2784);
and UO_441 (O_441,N_2959,N_2850);
nor UO_442 (O_442,N_2585,N_2641);
and UO_443 (O_443,N_2636,N_2707);
nand UO_444 (O_444,N_2549,N_2655);
or UO_445 (O_445,N_2707,N_2755);
and UO_446 (O_446,N_2660,N_2600);
or UO_447 (O_447,N_2779,N_2572);
or UO_448 (O_448,N_2921,N_2976);
or UO_449 (O_449,N_2959,N_2516);
or UO_450 (O_450,N_2643,N_2839);
nor UO_451 (O_451,N_2800,N_2660);
nand UO_452 (O_452,N_2799,N_2544);
and UO_453 (O_453,N_2720,N_2740);
or UO_454 (O_454,N_2799,N_2744);
nor UO_455 (O_455,N_2729,N_2506);
nand UO_456 (O_456,N_2929,N_2891);
nor UO_457 (O_457,N_2683,N_2736);
xnor UO_458 (O_458,N_2710,N_2579);
or UO_459 (O_459,N_2635,N_2997);
nor UO_460 (O_460,N_2966,N_2935);
nor UO_461 (O_461,N_2811,N_2552);
or UO_462 (O_462,N_2942,N_2816);
or UO_463 (O_463,N_2564,N_2529);
nand UO_464 (O_464,N_2927,N_2544);
nand UO_465 (O_465,N_2950,N_2772);
nand UO_466 (O_466,N_2624,N_2646);
nor UO_467 (O_467,N_2558,N_2562);
nand UO_468 (O_468,N_2976,N_2770);
or UO_469 (O_469,N_2680,N_2822);
or UO_470 (O_470,N_2918,N_2695);
nand UO_471 (O_471,N_2886,N_2891);
or UO_472 (O_472,N_2777,N_2689);
or UO_473 (O_473,N_2521,N_2558);
nand UO_474 (O_474,N_2642,N_2662);
and UO_475 (O_475,N_2753,N_2663);
nor UO_476 (O_476,N_2999,N_2718);
or UO_477 (O_477,N_2769,N_2534);
or UO_478 (O_478,N_2765,N_2831);
nor UO_479 (O_479,N_2763,N_2911);
nand UO_480 (O_480,N_2761,N_2682);
or UO_481 (O_481,N_2532,N_2675);
nor UO_482 (O_482,N_2741,N_2579);
nor UO_483 (O_483,N_2986,N_2561);
and UO_484 (O_484,N_2565,N_2736);
and UO_485 (O_485,N_2746,N_2588);
or UO_486 (O_486,N_2934,N_2686);
or UO_487 (O_487,N_2896,N_2733);
nor UO_488 (O_488,N_2888,N_2567);
nor UO_489 (O_489,N_2607,N_2816);
and UO_490 (O_490,N_2788,N_2960);
or UO_491 (O_491,N_2563,N_2630);
xor UO_492 (O_492,N_2739,N_2787);
nand UO_493 (O_493,N_2571,N_2675);
and UO_494 (O_494,N_2658,N_2532);
or UO_495 (O_495,N_2553,N_2757);
or UO_496 (O_496,N_2732,N_2988);
and UO_497 (O_497,N_2879,N_2658);
and UO_498 (O_498,N_2898,N_2576);
or UO_499 (O_499,N_2894,N_2644);
endmodule