module basic_1000_10000_1500_100_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_741,In_324);
nor U1 (N_1,In_852,In_930);
nor U2 (N_2,In_829,In_855);
and U3 (N_3,In_670,In_86);
nand U4 (N_4,In_446,In_477);
nor U5 (N_5,In_864,In_76);
and U6 (N_6,In_912,In_158);
nor U7 (N_7,In_844,In_195);
or U8 (N_8,In_718,In_130);
or U9 (N_9,In_859,In_433);
nor U10 (N_10,In_419,In_574);
nor U11 (N_11,In_357,In_75);
xor U12 (N_12,In_915,In_811);
nand U13 (N_13,In_951,In_180);
xor U14 (N_14,In_84,In_385);
nor U15 (N_15,In_24,In_445);
nand U16 (N_16,In_560,In_918);
and U17 (N_17,In_427,In_914);
nor U18 (N_18,In_522,In_406);
nor U19 (N_19,In_408,In_422);
nand U20 (N_20,In_22,In_935);
nor U21 (N_21,In_671,In_801);
xor U22 (N_22,In_127,In_78);
and U23 (N_23,In_21,In_10);
or U24 (N_24,In_80,In_610);
or U25 (N_25,In_447,In_378);
xor U26 (N_26,In_582,In_182);
and U27 (N_27,In_628,In_299);
xor U28 (N_28,In_255,In_108);
nor U29 (N_29,In_339,In_579);
xor U30 (N_30,In_961,In_333);
nand U31 (N_31,In_536,In_424);
or U32 (N_32,In_364,In_744);
nand U33 (N_33,In_286,In_593);
and U34 (N_34,In_544,In_111);
nor U35 (N_35,In_767,In_420);
or U36 (N_36,In_97,In_649);
or U37 (N_37,In_463,In_92);
xor U38 (N_38,In_330,In_787);
xnor U39 (N_39,In_550,In_305);
and U40 (N_40,In_765,In_791);
xnor U41 (N_41,In_232,In_313);
and U42 (N_42,In_745,In_476);
nor U43 (N_43,In_7,In_224);
or U44 (N_44,In_486,In_191);
nand U45 (N_45,In_925,In_241);
and U46 (N_46,In_821,In_50);
and U47 (N_47,In_528,In_743);
xnor U48 (N_48,In_277,In_208);
nand U49 (N_49,In_329,In_250);
nor U50 (N_50,In_138,In_291);
or U51 (N_51,In_887,In_631);
or U52 (N_52,In_732,In_584);
nor U53 (N_53,In_203,In_387);
or U54 (N_54,In_350,In_518);
xor U55 (N_55,In_197,In_351);
and U56 (N_56,In_49,In_48);
and U57 (N_57,In_662,In_714);
or U58 (N_58,In_594,In_519);
nand U59 (N_59,In_828,In_673);
nand U60 (N_60,In_133,In_1);
nor U61 (N_61,In_166,In_966);
nand U62 (N_62,In_258,In_113);
and U63 (N_63,In_390,In_699);
or U64 (N_64,In_798,In_280);
xor U65 (N_65,In_805,In_386);
nor U66 (N_66,In_125,In_396);
and U67 (N_67,In_950,In_442);
or U68 (N_68,In_633,In_988);
and U69 (N_69,In_997,In_975);
xor U70 (N_70,In_894,In_356);
or U71 (N_71,In_660,In_465);
or U72 (N_72,In_939,In_140);
or U73 (N_73,In_168,In_938);
nor U74 (N_74,In_490,In_881);
nor U75 (N_75,In_395,In_459);
and U76 (N_76,In_60,In_481);
nor U77 (N_77,In_297,In_973);
nor U78 (N_78,In_306,In_622);
and U79 (N_79,In_268,In_581);
and U80 (N_80,In_399,In_440);
nand U81 (N_81,In_290,In_143);
xnor U82 (N_82,In_713,In_927);
and U83 (N_83,In_267,In_95);
and U84 (N_84,In_688,In_804);
nor U85 (N_85,In_728,In_615);
and U86 (N_86,In_30,In_300);
and U87 (N_87,In_61,In_82);
and U88 (N_88,In_690,In_81);
xor U89 (N_89,In_167,In_843);
nand U90 (N_90,In_318,In_704);
xnor U91 (N_91,In_851,In_776);
and U92 (N_92,In_205,In_611);
nand U93 (N_93,In_739,In_556);
xnor U94 (N_94,In_423,In_154);
nor U95 (N_95,In_149,In_293);
nand U96 (N_96,In_174,In_899);
nor U97 (N_97,In_984,In_421);
nor U98 (N_98,In_724,In_64);
and U99 (N_99,In_793,In_775);
xor U100 (N_100,In_188,In_994);
and U101 (N_101,In_900,In_58);
xnor U102 (N_102,N_18,In_948);
nor U103 (N_103,In_865,In_23);
and U104 (N_104,In_489,In_735);
nor U105 (N_105,In_555,In_678);
nor U106 (N_106,In_884,In_349);
xnor U107 (N_107,In_537,In_559);
or U108 (N_108,In_327,In_733);
or U109 (N_109,In_608,In_17);
and U110 (N_110,In_814,In_316);
or U111 (N_111,In_772,In_104);
nand U112 (N_112,In_756,In_837);
and U113 (N_113,In_659,In_897);
xnor U114 (N_114,N_88,In_261);
or U115 (N_115,In_100,In_681);
xor U116 (N_116,In_789,N_7);
or U117 (N_117,In_769,N_50);
or U118 (N_118,In_401,N_49);
and U119 (N_119,In_721,In_304);
nor U120 (N_120,In_353,N_69);
xor U121 (N_121,In_159,In_903);
nand U122 (N_122,N_29,In_53);
and U123 (N_123,In_856,In_507);
nand U124 (N_124,In_768,In_564);
or U125 (N_125,N_58,In_770);
and U126 (N_126,In_102,In_949);
nand U127 (N_127,In_359,In_664);
nand U128 (N_128,In_976,In_79);
xnor U129 (N_129,In_716,In_278);
or U130 (N_130,In_563,In_274);
or U131 (N_131,In_103,N_52);
or U132 (N_132,In_42,In_495);
xnor U133 (N_133,In_895,In_578);
nor U134 (N_134,In_230,In_591);
nor U135 (N_135,In_137,In_597);
xnor U136 (N_136,In_836,In_244);
and U137 (N_137,In_283,In_955);
nor U138 (N_138,In_114,In_840);
or U139 (N_139,In_693,In_527);
nand U140 (N_140,In_885,In_730);
and U141 (N_141,In_832,N_98);
nand U142 (N_142,In_242,In_566);
nor U143 (N_143,In_418,In_896);
and U144 (N_144,In_262,In_934);
nor U145 (N_145,In_219,In_691);
xor U146 (N_146,In_28,In_204);
nand U147 (N_147,In_347,In_485);
or U148 (N_148,In_956,In_431);
nand U149 (N_149,In_252,In_345);
and U150 (N_150,In_749,In_284);
or U151 (N_151,In_186,In_853);
xor U152 (N_152,In_971,In_797);
nand U153 (N_153,N_4,In_737);
nor U154 (N_154,In_783,In_193);
and U155 (N_155,In_14,In_876);
nor U156 (N_156,In_134,In_573);
or U157 (N_157,In_497,In_117);
xor U158 (N_158,In_157,In_947);
xnor U159 (N_159,In_107,In_389);
nor U160 (N_160,In_658,In_285);
nand U161 (N_161,In_746,In_227);
xnor U162 (N_162,In_405,In_668);
or U163 (N_163,In_263,In_554);
nor U164 (N_164,In_20,N_81);
xnor U165 (N_165,In_601,N_21);
xor U166 (N_166,In_57,In_128);
nor U167 (N_167,In_273,In_376);
or U168 (N_168,In_254,N_96);
or U169 (N_169,In_151,In_882);
and U170 (N_170,In_165,N_10);
or U171 (N_171,N_38,In_74);
nand U172 (N_172,In_707,In_806);
nand U173 (N_173,In_922,In_627);
or U174 (N_174,In_360,In_281);
or U175 (N_175,In_178,In_809);
xnor U176 (N_176,In_953,In_762);
nor U177 (N_177,In_786,In_407);
or U178 (N_178,N_55,In_785);
or U179 (N_179,In_220,In_669);
nand U180 (N_180,In_34,In_119);
xor U181 (N_181,In_334,In_484);
nand U182 (N_182,In_542,In_0);
nand U183 (N_183,In_478,In_501);
and U184 (N_184,N_0,In_583);
or U185 (N_185,In_637,In_500);
nor U186 (N_186,In_812,In_651);
or U187 (N_187,In_612,In_321);
xor U188 (N_188,In_910,In_298);
or U189 (N_189,In_229,In_27);
xor U190 (N_190,In_974,N_74);
nand U191 (N_191,In_392,In_474);
xnor U192 (N_192,In_531,In_319);
xnor U193 (N_193,In_546,In_525);
or U194 (N_194,In_513,In_512);
or U195 (N_195,In_99,In_845);
and U196 (N_196,In_600,In_818);
nor U197 (N_197,In_508,In_636);
and U198 (N_198,In_414,In_77);
and U199 (N_199,In_715,In_712);
xnor U200 (N_200,In_183,In_367);
and U201 (N_201,N_155,N_63);
nor U202 (N_202,In_368,In_585);
or U203 (N_203,In_838,In_701);
and U204 (N_204,In_901,In_993);
nor U205 (N_205,In_275,In_199);
nand U206 (N_206,N_31,In_264);
xor U207 (N_207,In_648,In_176);
nand U208 (N_208,N_171,In_210);
nand U209 (N_209,In_877,In_337);
or U210 (N_210,In_740,N_168);
nand U211 (N_211,In_842,In_247);
and U212 (N_212,In_39,In_609);
nor U213 (N_213,In_314,In_383);
xor U214 (N_214,In_943,In_626);
and U215 (N_215,N_78,In_443);
nand U216 (N_216,In_37,N_190);
xnor U217 (N_217,N_199,In_409);
and U218 (N_218,In_868,In_782);
and U219 (N_219,In_639,N_132);
or U220 (N_220,N_138,In_889);
and U221 (N_221,In_112,In_657);
or U222 (N_222,In_524,In_494);
nand U223 (N_223,In_549,In_67);
nor U224 (N_224,N_71,N_36);
nand U225 (N_225,In_482,In_857);
and U226 (N_226,In_553,In_514);
xor U227 (N_227,In_235,In_890);
nor U228 (N_228,In_36,In_216);
xnor U229 (N_229,In_985,In_799);
nand U230 (N_230,In_827,N_30);
nor U231 (N_231,In_187,In_25);
nor U232 (N_232,In_381,In_567);
and U233 (N_233,N_47,In_361);
and U234 (N_234,In_962,In_709);
nand U235 (N_235,In_439,In_945);
and U236 (N_236,N_19,In_120);
and U237 (N_237,In_995,In_121);
nand U238 (N_238,In_807,In_380);
xnor U239 (N_239,In_515,N_82);
nor U240 (N_240,In_924,In_764);
nor U241 (N_241,N_79,In_473);
nor U242 (N_242,In_342,In_365);
nand U243 (N_243,In_532,N_163);
nor U244 (N_244,In_619,In_603);
nand U245 (N_245,In_545,N_127);
xor U246 (N_246,In_652,In_9);
nand U247 (N_247,In_875,In_850);
or U248 (N_248,N_146,In_870);
nand U249 (N_249,N_147,In_605);
or U250 (N_250,In_136,In_116);
nand U251 (N_251,N_157,In_819);
nor U252 (N_252,N_193,In_906);
xnor U253 (N_253,In_63,In_592);
and U254 (N_254,In_867,N_135);
xor U255 (N_255,In_780,In_147);
nor U256 (N_256,In_238,In_12);
or U257 (N_257,In_251,In_35);
and U258 (N_258,In_687,In_589);
and U259 (N_259,In_717,In_279);
xnor U260 (N_260,In_31,In_982);
nand U261 (N_261,In_784,In_624);
nand U262 (N_262,In_547,In_509);
xnor U263 (N_263,In_282,In_675);
nor U264 (N_264,In_288,In_110);
xnor U265 (N_265,In_642,In_893);
nor U266 (N_266,N_152,In_908);
nand U267 (N_267,In_543,In_499);
xnor U268 (N_268,In_41,In_937);
and U269 (N_269,In_234,In_541);
nand U270 (N_270,In_808,In_779);
nand U271 (N_271,N_178,In_523);
nand U272 (N_272,In_335,In_833);
nor U273 (N_273,N_34,In_483);
or U274 (N_274,In_123,In_700);
or U275 (N_275,In_83,In_607);
and U276 (N_276,In_987,N_51);
nand U277 (N_277,In_503,N_112);
or U278 (N_278,In_276,In_469);
and U279 (N_279,In_343,In_667);
nor U280 (N_280,N_73,In_621);
nand U281 (N_281,In_511,In_972);
nor U282 (N_282,In_461,In_752);
xor U283 (N_283,In_978,In_587);
nand U284 (N_284,N_181,N_169);
xor U285 (N_285,In_352,In_144);
nand U286 (N_286,In_826,In_813);
or U287 (N_287,In_534,In_38);
and U288 (N_288,In_175,N_56);
and U289 (N_289,In_942,In_980);
and U290 (N_290,N_84,N_128);
xnor U291 (N_291,In_47,In_332);
or U292 (N_292,In_4,In_849);
nor U293 (N_293,In_70,In_944);
and U294 (N_294,In_986,N_14);
xor U295 (N_295,In_990,In_18);
nor U296 (N_296,N_93,In_222);
xnor U297 (N_297,In_417,In_43);
and U298 (N_298,In_795,In_634);
and U299 (N_299,In_432,In_246);
or U300 (N_300,In_548,In_835);
and U301 (N_301,In_348,N_172);
or U302 (N_302,N_247,N_218);
and U303 (N_303,In_3,In_727);
nor U304 (N_304,In_847,N_223);
or U305 (N_305,In_977,N_212);
or U306 (N_306,N_173,In_979);
xor U307 (N_307,In_320,In_493);
xnor U308 (N_308,N_153,In_822);
nand U309 (N_309,N_111,In_29);
xor U310 (N_310,In_931,In_854);
xor U311 (N_311,N_17,N_102);
xnor U312 (N_312,In_379,N_282);
xor U313 (N_313,N_6,N_123);
or U314 (N_314,In_653,In_954);
or U315 (N_315,In_757,N_228);
or U316 (N_316,In_689,In_710);
xnor U317 (N_317,In_702,N_13);
nand U318 (N_318,N_189,N_246);
or U319 (N_319,In_372,In_720);
nor U320 (N_320,N_184,N_270);
xnor U321 (N_321,In_317,N_225);
nand U322 (N_322,In_173,In_46);
nor U323 (N_323,In_362,In_923);
nand U324 (N_324,In_672,In_233);
and U325 (N_325,In_436,In_677);
or U326 (N_326,In_928,In_872);
nor U327 (N_327,In_16,N_261);
and U328 (N_328,N_149,N_120);
nand U329 (N_329,In_155,In_45);
or U330 (N_330,In_640,N_42);
nand U331 (N_331,In_748,N_264);
nand U332 (N_332,In_510,In_455);
xor U333 (N_333,In_646,N_260);
and U334 (N_334,In_598,N_241);
nand U335 (N_335,N_285,N_217);
nand U336 (N_336,In_212,N_105);
nand U337 (N_337,In_126,In_570);
or U338 (N_338,In_69,In_331);
or U339 (N_339,In_294,In_983);
or U340 (N_340,In_630,N_27);
nand U341 (N_341,In_338,N_242);
and U342 (N_342,In_635,N_195);
nor U343 (N_343,N_227,N_131);
or U344 (N_344,In_632,N_259);
and U345 (N_345,N_106,In_403);
nand U346 (N_346,In_620,N_253);
and U347 (N_347,In_94,In_572);
nand U348 (N_348,In_428,N_265);
nor U349 (N_349,N_254,In_302);
or U350 (N_350,N_295,In_415);
or U351 (N_351,In_802,In_839);
nor U352 (N_352,In_467,In_758);
xor U353 (N_353,N_215,N_283);
or U354 (N_354,N_272,N_243);
nor U355 (N_355,In_62,N_137);
nand U356 (N_356,In_11,In_878);
nor U357 (N_357,In_904,In_460);
xnor U358 (N_358,In_629,N_221);
and U359 (N_359,N_91,N_158);
and U360 (N_360,In_68,In_85);
or U361 (N_361,N_240,N_224);
or U362 (N_362,In_863,N_113);
or U363 (N_363,N_280,In_371);
nand U364 (N_364,In_109,N_211);
nand U365 (N_365,In_416,In_296);
and U366 (N_366,In_56,In_891);
nand U367 (N_367,N_142,In_400);
and U368 (N_368,In_480,In_655);
and U369 (N_369,In_450,In_861);
xnor U370 (N_370,N_257,In_231);
xnor U371 (N_371,In_142,In_596);
and U372 (N_372,In_604,In_645);
or U373 (N_373,In_911,N_216);
xnor U374 (N_374,N_290,In_115);
nor U375 (N_375,In_363,N_72);
nor U376 (N_376,In_370,In_736);
and U377 (N_377,In_245,In_464);
xor U378 (N_378,In_207,N_44);
and U379 (N_379,In_344,In_156);
nor U380 (N_380,N_35,N_286);
xor U381 (N_381,In_958,In_132);
or U382 (N_382,N_26,N_45);
xnor U383 (N_383,In_202,In_190);
nor U384 (N_384,In_516,In_265);
nand U385 (N_385,In_834,In_52);
and U386 (N_386,In_161,N_159);
or U387 (N_387,In_569,N_156);
and U388 (N_388,In_249,N_104);
xnor U389 (N_389,In_926,N_54);
and U390 (N_390,N_60,In_488);
nand U391 (N_391,N_239,In_462);
nor U392 (N_392,In_73,N_214);
and U393 (N_393,N_126,In_957);
and U394 (N_394,N_267,In_963);
nor U395 (N_395,In_124,In_434);
nand U396 (N_396,N_144,In_326);
xnor U397 (N_397,In_831,N_161);
xnor U398 (N_398,In_644,In_698);
and U399 (N_399,In_989,In_729);
nand U400 (N_400,N_385,N_380);
and U401 (N_401,In_919,N_145);
nor U402 (N_402,N_165,In_498);
and U403 (N_403,N_275,In_453);
nand U404 (N_404,In_153,In_451);
nand U405 (N_405,In_226,N_119);
or U406 (N_406,In_398,N_208);
nor U407 (N_407,In_101,N_20);
or U408 (N_408,N_32,N_396);
nor U409 (N_409,N_48,In_223);
and U410 (N_410,In_788,N_266);
nor U411 (N_411,In_917,In_858);
nand U412 (N_412,In_684,N_392);
nor U413 (N_413,In_412,N_330);
xor U414 (N_414,In_228,In_217);
nor U415 (N_415,N_278,In_369);
or U416 (N_416,In_456,In_883);
and U417 (N_417,N_174,In_169);
and U418 (N_418,N_256,In_529);
and U419 (N_419,In_613,In_269);
and U420 (N_420,In_270,N_133);
xor U421 (N_421,In_468,In_438);
xnor U422 (N_422,In_886,N_277);
xor U423 (N_423,In_391,N_373);
nand U424 (N_424,In_860,N_375);
nor U425 (N_425,In_921,N_298);
and U426 (N_426,N_357,In_694);
and U427 (N_427,In_181,In_152);
nor U428 (N_428,In_341,In_661);
and U429 (N_429,N_343,In_437);
and U430 (N_430,In_682,N_326);
and U431 (N_431,N_238,In_196);
nor U432 (N_432,N_309,In_773);
nand U433 (N_433,N_12,In_2);
nand U434 (N_434,N_170,In_763);
nor U435 (N_435,In_198,In_606);
or U436 (N_436,In_150,N_167);
or U437 (N_437,N_318,In_540);
nand U438 (N_438,N_176,In_201);
xnor U439 (N_439,In_747,N_316);
nand U440 (N_440,N_315,N_41);
nand U441 (N_441,In_708,In_663);
xnor U442 (N_442,N_2,In_71);
and U443 (N_443,In_685,In_384);
or U444 (N_444,N_255,In_706);
nor U445 (N_445,In_679,In_817);
xor U446 (N_446,In_616,In_410);
and U447 (N_447,N_95,In_96);
nor U448 (N_448,N_103,In_726);
nand U449 (N_449,N_268,In_236);
nor U450 (N_450,In_561,In_774);
nand U451 (N_451,N_139,In_665);
or U452 (N_452,N_334,N_3);
and U453 (N_453,N_207,In_841);
and U454 (N_454,In_239,In_129);
and U455 (N_455,In_830,In_404);
nand U456 (N_456,In_755,N_53);
nand U457 (N_457,N_9,N_370);
nand U458 (N_458,In_373,N_83);
or U459 (N_459,N_114,In_413);
xor U460 (N_460,In_580,In_457);
nand U461 (N_461,N_25,N_229);
and U462 (N_462,In_5,N_67);
and U463 (N_463,N_222,In_59);
nor U464 (N_464,N_303,N_397);
nor U465 (N_465,In_777,In_539);
xnor U466 (N_466,In_225,N_314);
xnor U467 (N_467,In_771,N_287);
nand U468 (N_468,N_379,In_625);
nand U469 (N_469,In_309,In_194);
xnor U470 (N_470,N_234,In_941);
and U471 (N_471,In_590,In_815);
xnor U472 (N_472,In_766,In_810);
xnor U473 (N_473,In_51,In_211);
and U474 (N_474,N_361,N_359);
nand U475 (N_475,N_335,In_444);
and U476 (N_476,N_205,In_595);
or U477 (N_477,N_230,In_394);
nand U478 (N_478,N_349,In_315);
and U479 (N_479,In_981,In_106);
nor U480 (N_480,In_308,In_271);
nor U481 (N_481,N_99,N_383);
and U482 (N_482,N_204,In_502);
nand U483 (N_483,N_46,In_54);
xor U484 (N_484,N_358,N_151);
or U485 (N_485,N_354,In_13);
nand U486 (N_486,N_324,In_575);
and U487 (N_487,In_599,In_172);
nand U488 (N_488,N_301,In_164);
or U489 (N_489,In_377,N_175);
or U490 (N_490,N_310,In_933);
xor U491 (N_491,In_90,N_179);
or U492 (N_492,In_683,N_24);
nor U493 (N_493,In_131,N_213);
or U494 (N_494,In_189,N_61);
and U495 (N_495,In_696,In_905);
and U496 (N_496,In_323,In_869);
nor U497 (N_497,N_92,In_435);
or U498 (N_498,N_399,In_577);
and U499 (N_499,N_107,N_244);
nor U500 (N_500,N_8,N_471);
xnor U501 (N_501,In_206,In_105);
nand U502 (N_502,N_446,In_761);
or U503 (N_503,N_450,In_122);
nor U504 (N_504,N_445,N_274);
nand U505 (N_505,N_395,N_140);
or U506 (N_506,N_121,In_55);
or U507 (N_507,N_485,In_656);
xor U508 (N_508,N_352,In_397);
nor U509 (N_509,N_365,In_824);
nor U510 (N_510,N_493,In_533);
xor U511 (N_511,In_848,In_192);
xnor U512 (N_512,In_719,N_39);
nor U513 (N_513,In_163,In_430);
and U514 (N_514,N_180,In_307);
nand U515 (N_515,N_443,N_143);
nor U516 (N_516,In_388,N_416);
nand U517 (N_517,N_23,N_339);
nand U518 (N_518,N_329,In_790);
and U519 (N_519,In_200,N_452);
nand U520 (N_520,N_430,N_220);
xor U521 (N_521,In_491,N_15);
xor U522 (N_522,N_360,N_109);
nand U523 (N_523,In_940,N_390);
and U524 (N_524,N_185,In_565);
nand U525 (N_525,In_209,N_474);
nor U526 (N_526,N_456,In_336);
nand U527 (N_527,In_162,In_898);
xor U528 (N_528,In_139,In_374);
and U529 (N_529,In_920,N_125);
or U530 (N_530,N_317,N_448);
or U531 (N_531,N_192,In_66);
nand U532 (N_532,N_164,In_325);
or U533 (N_533,N_321,In_676);
nor U534 (N_534,In_454,N_206);
nand U535 (N_535,N_368,N_403);
nand U536 (N_536,N_235,N_371);
and U537 (N_537,N_434,N_497);
nand U538 (N_538,In_778,N_65);
nand U539 (N_539,N_162,In_65);
and U540 (N_540,N_292,N_136);
nand U541 (N_541,In_521,N_304);
and U542 (N_542,N_245,In_145);
or U543 (N_543,N_182,N_362);
xor U544 (N_544,N_177,N_348);
nor U545 (N_545,N_372,In_98);
xor U546 (N_546,N_209,In_909);
and U547 (N_547,N_492,In_218);
nor U548 (N_548,N_391,N_364);
or U549 (N_549,N_141,N_384);
nand U550 (N_550,In_880,N_325);
xnor U551 (N_551,N_308,N_378);
nor U552 (N_552,N_263,N_101);
xor U553 (N_553,N_451,In_15);
and U554 (N_554,In_19,In_487);
xnor U555 (N_555,In_148,In_722);
xnor U556 (N_556,In_711,N_465);
nand U557 (N_557,N_76,In_32);
and U558 (N_558,In_289,In_479);
nand U559 (N_559,N_297,In_552);
xor U560 (N_560,In_253,N_464);
nor U561 (N_561,N_469,In_588);
or U562 (N_562,In_240,N_449);
or U563 (N_563,N_294,N_442);
or U564 (N_564,In_340,In_393);
xnor U565 (N_565,N_322,N_386);
xor U566 (N_566,In_301,N_89);
nand U567 (N_567,N_342,In_970);
and U568 (N_568,N_289,In_40);
and U569 (N_569,In_402,In_742);
and U570 (N_570,In_322,In_471);
xor U571 (N_571,In_866,N_475);
xnor U572 (N_572,N_484,N_332);
xor U573 (N_573,In_557,N_337);
nand U574 (N_574,N_377,N_404);
nand U575 (N_575,N_134,N_414);
xnor U576 (N_576,In_411,N_408);
or U577 (N_577,N_226,In_551);
nand U578 (N_578,N_75,N_85);
nand U579 (N_579,N_350,N_202);
and U580 (N_580,N_70,In_358);
nor U581 (N_581,In_697,N_398);
xnor U582 (N_582,N_305,In_759);
xnor U583 (N_583,N_115,N_409);
and U584 (N_584,In_731,N_210);
xor U585 (N_585,In_879,In_602);
nor U586 (N_586,In_179,In_520);
or U587 (N_587,In_825,N_300);
nand U588 (N_588,N_498,N_415);
nand U589 (N_589,In_91,In_259);
or U590 (N_590,N_249,N_478);
nand U591 (N_591,N_288,N_400);
or U592 (N_592,In_674,In_506);
nand U593 (N_593,In_530,In_87);
or U594 (N_594,In_171,N_435);
or U595 (N_595,In_862,In_647);
nand U596 (N_596,N_296,N_495);
and U597 (N_597,N_381,N_401);
nor U598 (N_598,N_87,N_436);
nand U599 (N_599,N_453,N_299);
xor U600 (N_600,In_734,In_562);
nor U601 (N_601,N_33,N_307);
nor U602 (N_602,In_256,N_470);
nor U603 (N_603,In_871,N_312);
and U604 (N_604,In_213,N_406);
or U605 (N_605,In_458,N_355);
or U606 (N_606,N_477,N_501);
nor U607 (N_607,N_271,N_571);
nand U608 (N_608,N_586,N_411);
nor U609 (N_609,In_586,In_969);
nor U610 (N_610,In_623,In_846);
and U611 (N_611,N_319,In_781);
nand U612 (N_612,N_486,N_594);
and U613 (N_613,In_816,N_596);
nand U614 (N_614,N_80,N_203);
or U615 (N_615,In_526,In_754);
or U616 (N_616,N_467,N_510);
nand U617 (N_617,N_338,N_540);
or U618 (N_618,In_243,N_328);
xnor U619 (N_619,In_72,N_539);
nor U620 (N_620,N_468,N_437);
and U621 (N_621,In_643,N_573);
or U622 (N_622,N_547,In_170);
nand U623 (N_623,In_185,N_565);
xor U624 (N_624,N_555,In_141);
nor U625 (N_625,N_592,N_550);
xnor U626 (N_626,N_518,N_320);
or U627 (N_627,N_412,In_425);
and U628 (N_628,N_545,N_524);
nor U629 (N_629,N_503,N_447);
nand U630 (N_630,In_492,N_461);
or U631 (N_631,In_214,N_422);
and U632 (N_632,N_351,In_820);
nand U633 (N_633,In_650,N_347);
and U634 (N_634,N_237,N_194);
nor U635 (N_635,N_363,In_504);
xnor U636 (N_636,N_463,N_410);
or U637 (N_637,In_558,N_419);
nor U638 (N_638,N_129,N_595);
nor U639 (N_639,N_440,N_302);
and U640 (N_640,In_967,N_198);
nand U641 (N_641,N_580,In_452);
and U642 (N_642,N_311,In_965);
nor U643 (N_643,N_559,N_97);
or U644 (N_644,N_489,N_252);
xnor U645 (N_645,In_221,N_534);
and U646 (N_646,N_116,In_705);
xor U647 (N_647,N_582,N_425);
xnor U648 (N_648,N_191,N_344);
and U649 (N_649,In_666,N_94);
nor U650 (N_650,N_513,N_533);
xnor U651 (N_651,N_483,N_327);
or U652 (N_652,In_6,N_346);
and U653 (N_653,N_64,N_490);
or U654 (N_654,N_313,N_472);
and U655 (N_655,N_507,N_90);
nand U656 (N_656,In_873,N_557);
xnor U657 (N_657,In_466,N_460);
and U658 (N_658,N_454,In_686);
nand U659 (N_659,N_585,In_792);
xor U660 (N_660,N_231,N_269);
nand U661 (N_661,In_538,In_366);
nor U662 (N_662,N_481,N_487);
nand U663 (N_663,N_438,N_196);
or U664 (N_664,N_567,N_522);
xnor U665 (N_665,N_405,N_457);
or U666 (N_666,In_725,In_160);
nand U667 (N_667,In_751,In_936);
nor U668 (N_668,N_100,In_311);
nand U669 (N_669,N_186,In_800);
or U670 (N_670,N_232,In_874);
nor U671 (N_671,N_553,N_528);
and U672 (N_672,N_200,In_248);
xnor U673 (N_673,N_572,N_323);
xor U674 (N_674,N_291,N_462);
and U675 (N_675,N_394,N_166);
or U676 (N_676,N_541,N_554);
xnor U677 (N_677,N_546,N_331);
and U678 (N_678,N_480,N_563);
nand U679 (N_679,N_581,N_366);
and U680 (N_680,N_598,N_542);
nor U681 (N_681,N_262,In_88);
nand U682 (N_682,N_16,N_521);
nor U683 (N_683,N_588,N_482);
nand U684 (N_684,N_421,In_641);
nor U685 (N_685,N_599,N_426);
nand U686 (N_686,In_888,In_272);
and U687 (N_687,N_505,N_62);
nor U688 (N_688,In_260,N_543);
nor U689 (N_689,In_932,In_568);
and U690 (N_690,In_292,N_532);
nor U691 (N_691,N_511,N_479);
xnor U692 (N_692,N_509,N_560);
xor U693 (N_693,In_441,N_576);
nor U694 (N_694,N_504,N_529);
nor U695 (N_695,In_952,N_433);
xnor U696 (N_696,In_916,N_154);
and U697 (N_697,N_236,N_110);
or U698 (N_698,N_11,In_803);
nor U699 (N_699,N_1,In_496);
nor U700 (N_700,N_219,N_642);
nor U701 (N_701,N_691,In_449);
xnor U702 (N_702,N_494,N_387);
nand U703 (N_703,N_686,N_611);
nand U704 (N_704,In_738,N_197);
xnor U705 (N_705,N_431,N_650);
xnor U706 (N_706,N_306,In_237);
nand U707 (N_707,N_148,In_26);
nand U708 (N_708,N_459,In_354);
and U709 (N_709,N_466,N_376);
xor U710 (N_710,N_613,N_680);
nor U711 (N_711,N_685,N_516);
nand U712 (N_712,N_679,N_428);
or U713 (N_713,N_637,In_753);
xor U714 (N_714,N_458,N_625);
nand U715 (N_715,N_556,N_694);
and U716 (N_716,N_699,N_696);
and U717 (N_717,N_160,N_659);
or U718 (N_718,N_616,N_671);
and U719 (N_719,N_692,N_626);
xnor U720 (N_720,N_336,N_284);
xor U721 (N_721,N_669,N_183);
or U722 (N_722,N_427,N_622);
nand U723 (N_723,N_356,N_640);
nor U724 (N_724,N_549,N_604);
nand U725 (N_725,N_612,N_551);
nand U726 (N_726,In_576,In_571);
xnor U727 (N_727,In_426,N_657);
xnor U728 (N_728,N_620,N_629);
nand U729 (N_729,In_638,In_429);
nand U730 (N_730,In_328,N_636);
or U731 (N_731,N_618,N_500);
nand U732 (N_732,In_295,In_760);
nand U733 (N_733,N_608,N_248);
and U734 (N_734,In_902,N_628);
or U735 (N_735,In_794,N_634);
nand U736 (N_736,N_677,N_77);
nand U737 (N_737,N_584,N_353);
or U738 (N_738,In_470,N_644);
nor U739 (N_739,N_108,N_597);
nand U740 (N_740,N_662,N_601);
xor U741 (N_741,N_647,N_369);
xnor U742 (N_742,N_402,N_279);
or U743 (N_743,N_651,N_670);
nand U744 (N_744,N_418,N_258);
and U745 (N_745,N_488,N_698);
nand U746 (N_746,N_491,N_499);
and U747 (N_747,In_382,N_544);
or U748 (N_748,N_345,N_523);
nand U749 (N_749,N_630,N_668);
or U750 (N_750,N_5,N_579);
xor U751 (N_751,In_184,In_448);
or U752 (N_752,N_37,N_664);
nor U753 (N_753,N_639,N_658);
nand U754 (N_754,In_991,N_537);
nand U755 (N_755,N_382,N_473);
xnor U756 (N_756,N_496,N_610);
or U757 (N_757,N_250,N_517);
nand U758 (N_758,N_59,N_43);
nand U759 (N_759,N_538,N_506);
nand U760 (N_760,N_393,N_432);
or U761 (N_761,N_624,N_623);
and U762 (N_762,In_355,N_643);
nor U763 (N_763,In_146,N_631);
xor U764 (N_764,In_892,In_215);
nor U765 (N_765,N_661,N_407);
or U766 (N_766,N_439,In_472);
xor U767 (N_767,N_519,In_618);
xor U768 (N_768,N_388,N_530);
nand U769 (N_769,N_649,N_281);
and U770 (N_770,In_654,In_907);
nand U771 (N_771,In_93,N_593);
and U772 (N_772,N_693,In_964);
nor U773 (N_773,In_257,N_86);
xor U774 (N_774,N_676,N_591);
nand U775 (N_775,In_999,N_600);
or U776 (N_776,N_455,N_577);
nand U777 (N_777,N_690,N_645);
or U778 (N_778,In_266,N_251);
nand U779 (N_779,N_333,N_564);
nand U780 (N_780,N_28,N_632);
or U781 (N_781,N_590,In_505);
xnor U782 (N_782,N_589,N_655);
nand U783 (N_783,N_688,N_68);
nand U784 (N_784,N_635,N_660);
xor U785 (N_785,N_117,N_389);
and U786 (N_786,N_201,N_374);
or U787 (N_787,N_672,N_535);
nand U788 (N_788,N_627,N_602);
nor U789 (N_789,N_675,In_929);
xnor U790 (N_790,N_525,N_609);
and U791 (N_791,N_646,N_276);
nand U792 (N_792,In_177,In_992);
and U793 (N_793,In_692,N_531);
xor U794 (N_794,N_341,N_648);
xnor U795 (N_795,N_621,N_566);
nor U796 (N_796,In_703,N_633);
nand U797 (N_797,N_673,In_8);
or U798 (N_798,N_683,In_996);
nand U799 (N_799,N_429,In_968);
nand U800 (N_800,In_695,In_33);
nand U801 (N_801,N_667,N_652);
and U802 (N_802,N_687,N_561);
nor U803 (N_803,In_998,N_420);
nand U804 (N_804,N_705,N_124);
nor U805 (N_805,N_757,N_697);
and U806 (N_806,N_707,N_723);
nor U807 (N_807,N_663,N_770);
nand U808 (N_808,N_558,N_799);
or U809 (N_809,N_767,In_135);
and U810 (N_810,N_714,N_780);
and U811 (N_811,In_823,N_721);
nand U812 (N_812,N_66,N_764);
nor U813 (N_813,In_375,N_740);
nand U814 (N_814,N_656,N_340);
xor U815 (N_815,N_605,N_796);
xor U816 (N_816,In_614,In_303);
nand U817 (N_817,N_562,N_750);
xnor U818 (N_818,N_737,N_653);
and U819 (N_819,N_57,N_797);
nand U820 (N_820,N_717,N_674);
nand U821 (N_821,N_575,N_666);
and U822 (N_822,N_733,N_731);
nand U823 (N_823,In_959,N_614);
xor U824 (N_824,N_735,N_752);
nand U825 (N_825,N_761,N_570);
or U826 (N_826,N_700,N_689);
nand U827 (N_827,N_715,N_794);
or U828 (N_828,N_730,N_710);
xor U829 (N_829,N_606,N_552);
nor U830 (N_830,N_413,N_768);
nor U831 (N_831,N_441,N_712);
nor U832 (N_832,N_782,N_744);
nand U833 (N_833,In_312,In_346);
or U834 (N_834,In_475,In_617);
and U835 (N_835,N_743,N_568);
nor U836 (N_836,N_751,N_756);
or U837 (N_837,N_512,N_367);
and U838 (N_838,N_615,N_40);
nand U839 (N_839,N_781,N_759);
nor U840 (N_840,In_287,N_607);
xnor U841 (N_841,N_417,N_130);
and U842 (N_842,N_118,N_654);
and U843 (N_843,N_709,N_726);
nor U844 (N_844,N_695,N_776);
or U845 (N_845,N_758,N_703);
and U846 (N_846,N_748,N_792);
nor U847 (N_847,N_773,N_520);
and U848 (N_848,In_89,N_187);
and U849 (N_849,N_587,N_548);
nand U850 (N_850,N_514,N_787);
nor U851 (N_851,N_641,N_619);
xnor U852 (N_852,N_746,In_960);
nor U853 (N_853,N_738,N_719);
xnor U854 (N_854,N_728,N_766);
nand U855 (N_855,N_777,N_769);
xnor U856 (N_856,In_750,N_795);
and U857 (N_857,N_760,N_502);
nor U858 (N_858,N_745,N_617);
or U859 (N_859,N_578,N_739);
or U860 (N_860,N_763,N_783);
and U861 (N_861,In_796,N_775);
nand U862 (N_862,N_716,N_708);
or U863 (N_863,N_790,N_702);
xor U864 (N_864,In_680,N_749);
xor U865 (N_865,In_913,N_765);
nor U866 (N_866,N_526,N_720);
nor U867 (N_867,N_536,N_678);
and U868 (N_868,N_772,N_755);
nand U869 (N_869,N_574,N_150);
and U870 (N_870,N_681,N_747);
and U871 (N_871,N_774,N_583);
and U872 (N_872,N_122,N_718);
and U873 (N_873,N_785,N_684);
xor U874 (N_874,N_444,N_423);
xnor U875 (N_875,N_569,N_704);
nor U876 (N_876,N_508,N_273);
nand U877 (N_877,N_638,N_725);
nand U878 (N_878,N_791,N_476);
nor U879 (N_879,N_424,N_701);
and U880 (N_880,N_682,In_517);
or U881 (N_881,In_723,In_118);
nand U882 (N_882,N_729,In_946);
or U883 (N_883,N_188,N_293);
and U884 (N_884,N_665,N_786);
and U885 (N_885,N_753,N_741);
and U886 (N_886,N_734,N_762);
xnor U887 (N_887,N_706,N_724);
and U888 (N_888,N_713,In_310);
nor U889 (N_889,N_771,N_788);
xnor U890 (N_890,N_732,N_727);
and U891 (N_891,N_742,N_798);
xnor U892 (N_892,N_711,N_233);
or U893 (N_893,N_778,N_736);
and U894 (N_894,In_535,N_22);
and U895 (N_895,In_44,N_779);
nor U896 (N_896,N_527,N_789);
and U897 (N_897,N_603,N_784);
and U898 (N_898,N_722,N_793);
xor U899 (N_899,N_754,N_515);
nor U900 (N_900,N_839,N_814);
nor U901 (N_901,N_858,N_837);
or U902 (N_902,N_800,N_877);
nand U903 (N_903,N_809,N_822);
or U904 (N_904,N_844,N_891);
nand U905 (N_905,N_855,N_817);
and U906 (N_906,N_813,N_876);
nand U907 (N_907,N_888,N_848);
nor U908 (N_908,N_856,N_854);
xor U909 (N_909,N_845,N_886);
xnor U910 (N_910,N_818,N_860);
and U911 (N_911,N_820,N_898);
and U912 (N_912,N_881,N_849);
nor U913 (N_913,N_892,N_893);
or U914 (N_914,N_806,N_808);
or U915 (N_915,N_834,N_897);
nand U916 (N_916,N_842,N_804);
and U917 (N_917,N_843,N_824);
xnor U918 (N_918,N_887,N_801);
nor U919 (N_919,N_884,N_852);
xor U920 (N_920,N_851,N_835);
or U921 (N_921,N_811,N_873);
or U922 (N_922,N_825,N_863);
or U923 (N_923,N_870,N_869);
xnor U924 (N_924,N_831,N_826);
nand U925 (N_925,N_857,N_819);
or U926 (N_926,N_815,N_846);
or U927 (N_927,N_866,N_803);
nor U928 (N_928,N_828,N_807);
nand U929 (N_929,N_840,N_868);
and U930 (N_930,N_875,N_841);
nand U931 (N_931,N_890,N_878);
nor U932 (N_932,N_805,N_867);
and U933 (N_933,N_823,N_895);
nor U934 (N_934,N_872,N_874);
nand U935 (N_935,N_885,N_821);
or U936 (N_936,N_864,N_832);
xnor U937 (N_937,N_889,N_879);
and U938 (N_938,N_896,N_833);
nand U939 (N_939,N_836,N_882);
nor U940 (N_940,N_861,N_865);
nand U941 (N_941,N_894,N_802);
nand U942 (N_942,N_827,N_830);
xnor U943 (N_943,N_850,N_883);
and U944 (N_944,N_859,N_862);
nor U945 (N_945,N_829,N_810);
nand U946 (N_946,N_812,N_899);
nand U947 (N_947,N_838,N_816);
xnor U948 (N_948,N_847,N_853);
nor U949 (N_949,N_880,N_871);
and U950 (N_950,N_842,N_852);
nor U951 (N_951,N_849,N_877);
and U952 (N_952,N_819,N_814);
or U953 (N_953,N_830,N_864);
and U954 (N_954,N_802,N_855);
nor U955 (N_955,N_870,N_897);
nor U956 (N_956,N_890,N_807);
xor U957 (N_957,N_821,N_870);
nor U958 (N_958,N_865,N_856);
xor U959 (N_959,N_830,N_884);
nor U960 (N_960,N_813,N_814);
or U961 (N_961,N_811,N_870);
xnor U962 (N_962,N_868,N_883);
nor U963 (N_963,N_866,N_818);
nor U964 (N_964,N_896,N_805);
nor U965 (N_965,N_847,N_881);
xor U966 (N_966,N_881,N_870);
nor U967 (N_967,N_884,N_819);
nand U968 (N_968,N_892,N_813);
nand U969 (N_969,N_833,N_878);
and U970 (N_970,N_809,N_828);
or U971 (N_971,N_891,N_863);
and U972 (N_972,N_804,N_810);
nand U973 (N_973,N_882,N_871);
or U974 (N_974,N_850,N_806);
nand U975 (N_975,N_881,N_878);
or U976 (N_976,N_898,N_866);
and U977 (N_977,N_885,N_850);
and U978 (N_978,N_894,N_883);
and U979 (N_979,N_846,N_814);
or U980 (N_980,N_869,N_823);
and U981 (N_981,N_873,N_806);
nor U982 (N_982,N_847,N_891);
or U983 (N_983,N_866,N_884);
and U984 (N_984,N_856,N_858);
nor U985 (N_985,N_863,N_816);
or U986 (N_986,N_860,N_811);
or U987 (N_987,N_885,N_855);
xor U988 (N_988,N_878,N_837);
xor U989 (N_989,N_801,N_884);
nor U990 (N_990,N_844,N_882);
nor U991 (N_991,N_817,N_868);
xnor U992 (N_992,N_874,N_870);
nor U993 (N_993,N_855,N_878);
nand U994 (N_994,N_876,N_837);
nand U995 (N_995,N_852,N_882);
or U996 (N_996,N_815,N_887);
nor U997 (N_997,N_897,N_859);
xor U998 (N_998,N_865,N_854);
and U999 (N_999,N_849,N_815);
nand U1000 (N_1000,N_922,N_962);
nand U1001 (N_1001,N_917,N_992);
nor U1002 (N_1002,N_932,N_925);
nor U1003 (N_1003,N_915,N_985);
xor U1004 (N_1004,N_901,N_995);
and U1005 (N_1005,N_928,N_984);
and U1006 (N_1006,N_940,N_904);
or U1007 (N_1007,N_946,N_909);
nor U1008 (N_1008,N_971,N_938);
or U1009 (N_1009,N_957,N_907);
nor U1010 (N_1010,N_951,N_961);
nand U1011 (N_1011,N_979,N_916);
xor U1012 (N_1012,N_934,N_980);
nand U1013 (N_1013,N_903,N_983);
and U1014 (N_1014,N_949,N_989);
or U1015 (N_1015,N_996,N_997);
and U1016 (N_1016,N_906,N_923);
xnor U1017 (N_1017,N_935,N_943);
and U1018 (N_1018,N_994,N_913);
xor U1019 (N_1019,N_924,N_937);
and U1020 (N_1020,N_999,N_921);
xor U1021 (N_1021,N_988,N_965);
nand U1022 (N_1022,N_941,N_958);
nor U1023 (N_1023,N_975,N_919);
xor U1024 (N_1024,N_977,N_974);
and U1025 (N_1025,N_948,N_926);
and U1026 (N_1026,N_929,N_954);
and U1027 (N_1027,N_952,N_933);
or U1028 (N_1028,N_978,N_936);
or U1029 (N_1029,N_912,N_945);
xor U1030 (N_1030,N_993,N_953);
and U1031 (N_1031,N_960,N_987);
nand U1032 (N_1032,N_973,N_950);
nand U1033 (N_1033,N_931,N_900);
and U1034 (N_1034,N_905,N_902);
nand U1035 (N_1035,N_908,N_967);
xnor U1036 (N_1036,N_944,N_963);
nor U1037 (N_1037,N_914,N_959);
or U1038 (N_1038,N_976,N_972);
nor U1039 (N_1039,N_955,N_930);
xnor U1040 (N_1040,N_966,N_911);
and U1041 (N_1041,N_927,N_964);
nand U1042 (N_1042,N_920,N_939);
nor U1043 (N_1043,N_942,N_981);
nand U1044 (N_1044,N_910,N_990);
nor U1045 (N_1045,N_986,N_969);
xor U1046 (N_1046,N_991,N_918);
and U1047 (N_1047,N_956,N_998);
and U1048 (N_1048,N_968,N_947);
or U1049 (N_1049,N_982,N_970);
nand U1050 (N_1050,N_959,N_905);
or U1051 (N_1051,N_908,N_907);
or U1052 (N_1052,N_965,N_953);
nand U1053 (N_1053,N_930,N_941);
and U1054 (N_1054,N_944,N_955);
or U1055 (N_1055,N_991,N_982);
nand U1056 (N_1056,N_979,N_955);
nand U1057 (N_1057,N_959,N_906);
and U1058 (N_1058,N_922,N_940);
and U1059 (N_1059,N_901,N_952);
xnor U1060 (N_1060,N_905,N_991);
nand U1061 (N_1061,N_978,N_964);
nand U1062 (N_1062,N_919,N_970);
xor U1063 (N_1063,N_980,N_981);
and U1064 (N_1064,N_941,N_909);
nor U1065 (N_1065,N_956,N_942);
and U1066 (N_1066,N_922,N_969);
and U1067 (N_1067,N_933,N_901);
and U1068 (N_1068,N_997,N_934);
or U1069 (N_1069,N_978,N_920);
nand U1070 (N_1070,N_940,N_943);
and U1071 (N_1071,N_947,N_985);
nor U1072 (N_1072,N_975,N_973);
nand U1073 (N_1073,N_966,N_958);
or U1074 (N_1074,N_989,N_929);
and U1075 (N_1075,N_974,N_901);
nand U1076 (N_1076,N_904,N_981);
nand U1077 (N_1077,N_978,N_981);
or U1078 (N_1078,N_926,N_958);
and U1079 (N_1079,N_902,N_924);
nor U1080 (N_1080,N_966,N_946);
xor U1081 (N_1081,N_901,N_900);
nand U1082 (N_1082,N_936,N_944);
and U1083 (N_1083,N_943,N_988);
nand U1084 (N_1084,N_913,N_931);
nor U1085 (N_1085,N_983,N_912);
and U1086 (N_1086,N_991,N_976);
xnor U1087 (N_1087,N_921,N_994);
nor U1088 (N_1088,N_957,N_956);
and U1089 (N_1089,N_903,N_975);
nor U1090 (N_1090,N_987,N_945);
nand U1091 (N_1091,N_966,N_986);
or U1092 (N_1092,N_902,N_989);
or U1093 (N_1093,N_931,N_970);
or U1094 (N_1094,N_910,N_923);
and U1095 (N_1095,N_973,N_913);
nand U1096 (N_1096,N_964,N_934);
xnor U1097 (N_1097,N_970,N_983);
or U1098 (N_1098,N_995,N_907);
nand U1099 (N_1099,N_945,N_931);
xor U1100 (N_1100,N_1028,N_1062);
nand U1101 (N_1101,N_1079,N_1021);
or U1102 (N_1102,N_1092,N_1074);
xnor U1103 (N_1103,N_1097,N_1076);
xnor U1104 (N_1104,N_1098,N_1068);
or U1105 (N_1105,N_1063,N_1096);
and U1106 (N_1106,N_1038,N_1009);
nand U1107 (N_1107,N_1016,N_1040);
xor U1108 (N_1108,N_1069,N_1057);
nand U1109 (N_1109,N_1019,N_1078);
or U1110 (N_1110,N_1060,N_1032);
or U1111 (N_1111,N_1071,N_1056);
nor U1112 (N_1112,N_1031,N_1067);
nor U1113 (N_1113,N_1089,N_1084);
nand U1114 (N_1114,N_1030,N_1025);
and U1115 (N_1115,N_1011,N_1029);
nor U1116 (N_1116,N_1070,N_1020);
nand U1117 (N_1117,N_1035,N_1000);
nor U1118 (N_1118,N_1023,N_1039);
xnor U1119 (N_1119,N_1099,N_1042);
nor U1120 (N_1120,N_1027,N_1059);
or U1121 (N_1121,N_1066,N_1018);
or U1122 (N_1122,N_1075,N_1045);
and U1123 (N_1123,N_1087,N_1061);
nand U1124 (N_1124,N_1002,N_1065);
or U1125 (N_1125,N_1041,N_1017);
and U1126 (N_1126,N_1014,N_1033);
nand U1127 (N_1127,N_1094,N_1093);
xnor U1128 (N_1128,N_1095,N_1004);
and U1129 (N_1129,N_1001,N_1055);
nand U1130 (N_1130,N_1044,N_1026);
and U1131 (N_1131,N_1037,N_1048);
xor U1132 (N_1132,N_1007,N_1072);
nor U1133 (N_1133,N_1081,N_1013);
nor U1134 (N_1134,N_1080,N_1008);
nand U1135 (N_1135,N_1010,N_1064);
or U1136 (N_1136,N_1049,N_1088);
nor U1137 (N_1137,N_1046,N_1091);
and U1138 (N_1138,N_1024,N_1083);
nand U1139 (N_1139,N_1012,N_1015);
xnor U1140 (N_1140,N_1051,N_1054);
nor U1141 (N_1141,N_1003,N_1006);
or U1142 (N_1142,N_1034,N_1090);
nor U1143 (N_1143,N_1053,N_1043);
nor U1144 (N_1144,N_1086,N_1085);
or U1145 (N_1145,N_1073,N_1052);
nor U1146 (N_1146,N_1036,N_1005);
and U1147 (N_1147,N_1047,N_1077);
nand U1148 (N_1148,N_1058,N_1082);
and U1149 (N_1149,N_1050,N_1022);
and U1150 (N_1150,N_1049,N_1091);
and U1151 (N_1151,N_1071,N_1083);
nand U1152 (N_1152,N_1054,N_1096);
nand U1153 (N_1153,N_1062,N_1027);
nor U1154 (N_1154,N_1054,N_1020);
nand U1155 (N_1155,N_1082,N_1085);
or U1156 (N_1156,N_1033,N_1001);
xor U1157 (N_1157,N_1080,N_1052);
nor U1158 (N_1158,N_1031,N_1082);
nor U1159 (N_1159,N_1016,N_1037);
nor U1160 (N_1160,N_1099,N_1000);
or U1161 (N_1161,N_1024,N_1000);
nand U1162 (N_1162,N_1002,N_1095);
nor U1163 (N_1163,N_1089,N_1025);
nor U1164 (N_1164,N_1004,N_1033);
xnor U1165 (N_1165,N_1050,N_1042);
xnor U1166 (N_1166,N_1082,N_1067);
xnor U1167 (N_1167,N_1010,N_1069);
nor U1168 (N_1168,N_1088,N_1032);
xnor U1169 (N_1169,N_1095,N_1001);
nand U1170 (N_1170,N_1056,N_1000);
or U1171 (N_1171,N_1037,N_1059);
nor U1172 (N_1172,N_1005,N_1050);
and U1173 (N_1173,N_1037,N_1011);
and U1174 (N_1174,N_1053,N_1050);
or U1175 (N_1175,N_1045,N_1093);
xor U1176 (N_1176,N_1016,N_1043);
nor U1177 (N_1177,N_1053,N_1065);
or U1178 (N_1178,N_1028,N_1013);
xor U1179 (N_1179,N_1069,N_1068);
nand U1180 (N_1180,N_1099,N_1064);
nor U1181 (N_1181,N_1084,N_1012);
and U1182 (N_1182,N_1022,N_1000);
or U1183 (N_1183,N_1012,N_1020);
and U1184 (N_1184,N_1044,N_1027);
or U1185 (N_1185,N_1063,N_1036);
and U1186 (N_1186,N_1075,N_1014);
nor U1187 (N_1187,N_1066,N_1028);
and U1188 (N_1188,N_1055,N_1084);
xor U1189 (N_1189,N_1083,N_1054);
nand U1190 (N_1190,N_1033,N_1053);
xor U1191 (N_1191,N_1064,N_1094);
or U1192 (N_1192,N_1072,N_1040);
xnor U1193 (N_1193,N_1022,N_1059);
xor U1194 (N_1194,N_1061,N_1038);
nor U1195 (N_1195,N_1092,N_1023);
and U1196 (N_1196,N_1064,N_1051);
and U1197 (N_1197,N_1055,N_1088);
xnor U1198 (N_1198,N_1075,N_1089);
or U1199 (N_1199,N_1072,N_1003);
nor U1200 (N_1200,N_1108,N_1155);
xor U1201 (N_1201,N_1197,N_1148);
and U1202 (N_1202,N_1123,N_1178);
or U1203 (N_1203,N_1102,N_1149);
nand U1204 (N_1204,N_1147,N_1100);
xnor U1205 (N_1205,N_1135,N_1183);
or U1206 (N_1206,N_1112,N_1189);
and U1207 (N_1207,N_1177,N_1156);
xor U1208 (N_1208,N_1185,N_1113);
nor U1209 (N_1209,N_1193,N_1157);
or U1210 (N_1210,N_1184,N_1158);
nor U1211 (N_1211,N_1124,N_1103);
or U1212 (N_1212,N_1139,N_1136);
or U1213 (N_1213,N_1145,N_1152);
nand U1214 (N_1214,N_1180,N_1137);
nand U1215 (N_1215,N_1132,N_1118);
xor U1216 (N_1216,N_1162,N_1150);
nand U1217 (N_1217,N_1170,N_1126);
xnor U1218 (N_1218,N_1138,N_1153);
xor U1219 (N_1219,N_1168,N_1161);
nor U1220 (N_1220,N_1171,N_1111);
nand U1221 (N_1221,N_1172,N_1194);
nor U1222 (N_1222,N_1131,N_1169);
nand U1223 (N_1223,N_1179,N_1173);
nand U1224 (N_1224,N_1167,N_1106);
nor U1225 (N_1225,N_1129,N_1159);
nand U1226 (N_1226,N_1186,N_1176);
and U1227 (N_1227,N_1195,N_1174);
or U1228 (N_1228,N_1120,N_1119);
nor U1229 (N_1229,N_1154,N_1181);
nor U1230 (N_1230,N_1122,N_1107);
nand U1231 (N_1231,N_1140,N_1166);
and U1232 (N_1232,N_1192,N_1105);
xor U1233 (N_1233,N_1175,N_1104);
and U1234 (N_1234,N_1109,N_1190);
nor U1235 (N_1235,N_1198,N_1187);
xor U1236 (N_1236,N_1163,N_1117);
or U1237 (N_1237,N_1165,N_1144);
and U1238 (N_1238,N_1133,N_1146);
nor U1239 (N_1239,N_1196,N_1160);
and U1240 (N_1240,N_1114,N_1101);
and U1241 (N_1241,N_1164,N_1191);
nor U1242 (N_1242,N_1151,N_1115);
nor U1243 (N_1243,N_1110,N_1116);
nand U1244 (N_1244,N_1141,N_1134);
nor U1245 (N_1245,N_1199,N_1142);
or U1246 (N_1246,N_1127,N_1182);
nor U1247 (N_1247,N_1143,N_1128);
or U1248 (N_1248,N_1130,N_1125);
or U1249 (N_1249,N_1188,N_1121);
xor U1250 (N_1250,N_1175,N_1134);
or U1251 (N_1251,N_1104,N_1134);
and U1252 (N_1252,N_1197,N_1167);
xor U1253 (N_1253,N_1144,N_1113);
xnor U1254 (N_1254,N_1189,N_1129);
or U1255 (N_1255,N_1119,N_1180);
xnor U1256 (N_1256,N_1114,N_1109);
and U1257 (N_1257,N_1115,N_1177);
nand U1258 (N_1258,N_1146,N_1155);
or U1259 (N_1259,N_1173,N_1107);
or U1260 (N_1260,N_1185,N_1198);
nor U1261 (N_1261,N_1149,N_1178);
nor U1262 (N_1262,N_1179,N_1176);
nand U1263 (N_1263,N_1118,N_1174);
nand U1264 (N_1264,N_1196,N_1178);
or U1265 (N_1265,N_1106,N_1130);
xor U1266 (N_1266,N_1194,N_1153);
or U1267 (N_1267,N_1189,N_1185);
nor U1268 (N_1268,N_1175,N_1192);
xor U1269 (N_1269,N_1112,N_1124);
nand U1270 (N_1270,N_1169,N_1182);
nor U1271 (N_1271,N_1152,N_1185);
and U1272 (N_1272,N_1161,N_1175);
xnor U1273 (N_1273,N_1112,N_1173);
nand U1274 (N_1274,N_1135,N_1111);
nand U1275 (N_1275,N_1139,N_1123);
and U1276 (N_1276,N_1185,N_1165);
nand U1277 (N_1277,N_1141,N_1184);
nor U1278 (N_1278,N_1187,N_1111);
nand U1279 (N_1279,N_1175,N_1108);
xnor U1280 (N_1280,N_1130,N_1167);
nor U1281 (N_1281,N_1152,N_1122);
and U1282 (N_1282,N_1197,N_1119);
nor U1283 (N_1283,N_1110,N_1141);
or U1284 (N_1284,N_1150,N_1167);
or U1285 (N_1285,N_1127,N_1192);
nor U1286 (N_1286,N_1154,N_1149);
and U1287 (N_1287,N_1148,N_1145);
xnor U1288 (N_1288,N_1102,N_1106);
xnor U1289 (N_1289,N_1103,N_1131);
xnor U1290 (N_1290,N_1140,N_1159);
and U1291 (N_1291,N_1164,N_1162);
xnor U1292 (N_1292,N_1186,N_1164);
nor U1293 (N_1293,N_1190,N_1142);
or U1294 (N_1294,N_1108,N_1183);
or U1295 (N_1295,N_1189,N_1175);
nand U1296 (N_1296,N_1155,N_1157);
nand U1297 (N_1297,N_1147,N_1123);
nand U1298 (N_1298,N_1156,N_1129);
and U1299 (N_1299,N_1181,N_1174);
nand U1300 (N_1300,N_1260,N_1293);
nand U1301 (N_1301,N_1259,N_1243);
and U1302 (N_1302,N_1237,N_1251);
nor U1303 (N_1303,N_1223,N_1235);
xnor U1304 (N_1304,N_1275,N_1230);
nor U1305 (N_1305,N_1288,N_1278);
and U1306 (N_1306,N_1201,N_1234);
or U1307 (N_1307,N_1200,N_1219);
and U1308 (N_1308,N_1244,N_1282);
nand U1309 (N_1309,N_1232,N_1286);
nor U1310 (N_1310,N_1202,N_1218);
nor U1311 (N_1311,N_1250,N_1265);
nand U1312 (N_1312,N_1285,N_1297);
nor U1313 (N_1313,N_1258,N_1209);
nor U1314 (N_1314,N_1225,N_1240);
nand U1315 (N_1315,N_1221,N_1248);
and U1316 (N_1316,N_1203,N_1277);
and U1317 (N_1317,N_1222,N_1247);
nor U1318 (N_1318,N_1255,N_1211);
and U1319 (N_1319,N_1231,N_1249);
xnor U1320 (N_1320,N_1287,N_1252);
nor U1321 (N_1321,N_1273,N_1204);
or U1322 (N_1322,N_1279,N_1229);
nand U1323 (N_1323,N_1276,N_1292);
or U1324 (N_1324,N_1207,N_1215);
nor U1325 (N_1325,N_1274,N_1228);
xnor U1326 (N_1326,N_1269,N_1220);
nor U1327 (N_1327,N_1257,N_1296);
and U1328 (N_1328,N_1216,N_1246);
xnor U1329 (N_1329,N_1270,N_1266);
xnor U1330 (N_1330,N_1289,N_1281);
xor U1331 (N_1331,N_1208,N_1290);
xor U1332 (N_1332,N_1262,N_1242);
xor U1333 (N_1333,N_1238,N_1236);
and U1334 (N_1334,N_1214,N_1227);
and U1335 (N_1335,N_1245,N_1261);
and U1336 (N_1336,N_1268,N_1212);
xnor U1337 (N_1337,N_1291,N_1256);
nand U1338 (N_1338,N_1298,N_1226);
and U1339 (N_1339,N_1271,N_1224);
and U1340 (N_1340,N_1241,N_1299);
nand U1341 (N_1341,N_1283,N_1213);
or U1342 (N_1342,N_1294,N_1267);
xnor U1343 (N_1343,N_1210,N_1206);
nand U1344 (N_1344,N_1264,N_1295);
nor U1345 (N_1345,N_1217,N_1280);
xnor U1346 (N_1346,N_1205,N_1263);
and U1347 (N_1347,N_1272,N_1284);
or U1348 (N_1348,N_1253,N_1233);
and U1349 (N_1349,N_1254,N_1239);
nand U1350 (N_1350,N_1286,N_1265);
xor U1351 (N_1351,N_1284,N_1214);
and U1352 (N_1352,N_1202,N_1214);
or U1353 (N_1353,N_1252,N_1296);
nand U1354 (N_1354,N_1239,N_1275);
nand U1355 (N_1355,N_1201,N_1206);
or U1356 (N_1356,N_1277,N_1200);
nand U1357 (N_1357,N_1283,N_1230);
xnor U1358 (N_1358,N_1226,N_1217);
or U1359 (N_1359,N_1297,N_1223);
and U1360 (N_1360,N_1245,N_1217);
nor U1361 (N_1361,N_1206,N_1231);
nor U1362 (N_1362,N_1201,N_1277);
nor U1363 (N_1363,N_1225,N_1263);
nand U1364 (N_1364,N_1203,N_1211);
and U1365 (N_1365,N_1299,N_1282);
or U1366 (N_1366,N_1206,N_1237);
nor U1367 (N_1367,N_1254,N_1236);
or U1368 (N_1368,N_1259,N_1264);
xor U1369 (N_1369,N_1224,N_1254);
and U1370 (N_1370,N_1274,N_1270);
or U1371 (N_1371,N_1281,N_1269);
nand U1372 (N_1372,N_1278,N_1295);
xnor U1373 (N_1373,N_1204,N_1240);
nand U1374 (N_1374,N_1291,N_1222);
and U1375 (N_1375,N_1273,N_1229);
or U1376 (N_1376,N_1232,N_1201);
or U1377 (N_1377,N_1246,N_1207);
xor U1378 (N_1378,N_1286,N_1235);
or U1379 (N_1379,N_1225,N_1258);
nand U1380 (N_1380,N_1212,N_1232);
nor U1381 (N_1381,N_1254,N_1268);
and U1382 (N_1382,N_1290,N_1209);
and U1383 (N_1383,N_1270,N_1275);
nor U1384 (N_1384,N_1293,N_1233);
or U1385 (N_1385,N_1209,N_1210);
nor U1386 (N_1386,N_1295,N_1267);
xnor U1387 (N_1387,N_1210,N_1256);
xnor U1388 (N_1388,N_1292,N_1249);
or U1389 (N_1389,N_1212,N_1279);
nand U1390 (N_1390,N_1241,N_1209);
nor U1391 (N_1391,N_1233,N_1201);
xor U1392 (N_1392,N_1294,N_1231);
nand U1393 (N_1393,N_1251,N_1243);
nand U1394 (N_1394,N_1210,N_1233);
nor U1395 (N_1395,N_1264,N_1225);
nor U1396 (N_1396,N_1234,N_1219);
xor U1397 (N_1397,N_1238,N_1248);
xnor U1398 (N_1398,N_1269,N_1205);
nor U1399 (N_1399,N_1241,N_1293);
or U1400 (N_1400,N_1346,N_1325);
nor U1401 (N_1401,N_1360,N_1351);
nor U1402 (N_1402,N_1344,N_1320);
nor U1403 (N_1403,N_1334,N_1340);
nor U1404 (N_1404,N_1338,N_1318);
or U1405 (N_1405,N_1376,N_1308);
xnor U1406 (N_1406,N_1337,N_1397);
nand U1407 (N_1407,N_1326,N_1390);
nor U1408 (N_1408,N_1301,N_1389);
xor U1409 (N_1409,N_1356,N_1367);
nand U1410 (N_1410,N_1342,N_1336);
nand U1411 (N_1411,N_1317,N_1328);
nor U1412 (N_1412,N_1302,N_1324);
or U1413 (N_1413,N_1387,N_1385);
and U1414 (N_1414,N_1363,N_1357);
or U1415 (N_1415,N_1312,N_1330);
nand U1416 (N_1416,N_1372,N_1394);
nand U1417 (N_1417,N_1381,N_1322);
nand U1418 (N_1418,N_1348,N_1379);
and U1419 (N_1419,N_1349,N_1306);
xor U1420 (N_1420,N_1332,N_1369);
nand U1421 (N_1421,N_1362,N_1316);
and U1422 (N_1422,N_1392,N_1321);
and U1423 (N_1423,N_1359,N_1345);
nor U1424 (N_1424,N_1366,N_1364);
or U1425 (N_1425,N_1377,N_1352);
nor U1426 (N_1426,N_1395,N_1341);
or U1427 (N_1427,N_1365,N_1309);
nand U1428 (N_1428,N_1339,N_1391);
or U1429 (N_1429,N_1361,N_1343);
or U1430 (N_1430,N_1313,N_1375);
nand U1431 (N_1431,N_1384,N_1393);
and U1432 (N_1432,N_1380,N_1374);
xnor U1433 (N_1433,N_1327,N_1319);
or U1434 (N_1434,N_1399,N_1303);
or U1435 (N_1435,N_1311,N_1307);
or U1436 (N_1436,N_1314,N_1333);
and U1437 (N_1437,N_1350,N_1398);
nand U1438 (N_1438,N_1323,N_1347);
and U1439 (N_1439,N_1370,N_1335);
xnor U1440 (N_1440,N_1368,N_1378);
xor U1441 (N_1441,N_1386,N_1382);
nor U1442 (N_1442,N_1300,N_1383);
nor U1443 (N_1443,N_1331,N_1371);
nand U1444 (N_1444,N_1396,N_1329);
xnor U1445 (N_1445,N_1315,N_1310);
xnor U1446 (N_1446,N_1388,N_1305);
and U1447 (N_1447,N_1355,N_1353);
or U1448 (N_1448,N_1373,N_1358);
nor U1449 (N_1449,N_1354,N_1304);
nor U1450 (N_1450,N_1374,N_1328);
and U1451 (N_1451,N_1359,N_1392);
nor U1452 (N_1452,N_1338,N_1352);
xnor U1453 (N_1453,N_1329,N_1365);
nor U1454 (N_1454,N_1383,N_1354);
xnor U1455 (N_1455,N_1394,N_1349);
or U1456 (N_1456,N_1371,N_1383);
xnor U1457 (N_1457,N_1331,N_1385);
and U1458 (N_1458,N_1370,N_1351);
xnor U1459 (N_1459,N_1368,N_1395);
and U1460 (N_1460,N_1309,N_1368);
nor U1461 (N_1461,N_1347,N_1360);
and U1462 (N_1462,N_1354,N_1322);
nor U1463 (N_1463,N_1337,N_1368);
nor U1464 (N_1464,N_1391,N_1326);
xor U1465 (N_1465,N_1355,N_1388);
or U1466 (N_1466,N_1337,N_1328);
xor U1467 (N_1467,N_1317,N_1366);
nand U1468 (N_1468,N_1323,N_1338);
xor U1469 (N_1469,N_1335,N_1353);
xor U1470 (N_1470,N_1370,N_1303);
nor U1471 (N_1471,N_1359,N_1328);
and U1472 (N_1472,N_1374,N_1398);
xnor U1473 (N_1473,N_1309,N_1302);
and U1474 (N_1474,N_1334,N_1304);
xnor U1475 (N_1475,N_1377,N_1303);
nor U1476 (N_1476,N_1350,N_1332);
xnor U1477 (N_1477,N_1380,N_1339);
and U1478 (N_1478,N_1380,N_1355);
nand U1479 (N_1479,N_1332,N_1306);
or U1480 (N_1480,N_1361,N_1337);
nand U1481 (N_1481,N_1380,N_1384);
nand U1482 (N_1482,N_1345,N_1364);
and U1483 (N_1483,N_1358,N_1312);
or U1484 (N_1484,N_1323,N_1356);
or U1485 (N_1485,N_1376,N_1383);
nor U1486 (N_1486,N_1371,N_1339);
nand U1487 (N_1487,N_1314,N_1373);
nand U1488 (N_1488,N_1366,N_1333);
nand U1489 (N_1489,N_1306,N_1309);
xnor U1490 (N_1490,N_1309,N_1391);
nand U1491 (N_1491,N_1319,N_1341);
xnor U1492 (N_1492,N_1319,N_1381);
or U1493 (N_1493,N_1367,N_1338);
xor U1494 (N_1494,N_1343,N_1342);
or U1495 (N_1495,N_1354,N_1371);
or U1496 (N_1496,N_1310,N_1321);
and U1497 (N_1497,N_1354,N_1316);
xor U1498 (N_1498,N_1336,N_1330);
or U1499 (N_1499,N_1384,N_1335);
and U1500 (N_1500,N_1494,N_1462);
xnor U1501 (N_1501,N_1402,N_1434);
or U1502 (N_1502,N_1468,N_1475);
nand U1503 (N_1503,N_1430,N_1441);
and U1504 (N_1504,N_1435,N_1471);
and U1505 (N_1505,N_1440,N_1493);
and U1506 (N_1506,N_1458,N_1443);
xor U1507 (N_1507,N_1477,N_1470);
and U1508 (N_1508,N_1433,N_1428);
nand U1509 (N_1509,N_1474,N_1465);
and U1510 (N_1510,N_1446,N_1424);
xor U1511 (N_1511,N_1452,N_1469);
and U1512 (N_1512,N_1429,N_1419);
and U1513 (N_1513,N_1448,N_1490);
or U1514 (N_1514,N_1454,N_1412);
nand U1515 (N_1515,N_1410,N_1400);
nor U1516 (N_1516,N_1455,N_1489);
nor U1517 (N_1517,N_1464,N_1449);
xnor U1518 (N_1518,N_1413,N_1467);
nor U1519 (N_1519,N_1406,N_1431);
nor U1520 (N_1520,N_1492,N_1438);
xor U1521 (N_1521,N_1444,N_1451);
nor U1522 (N_1522,N_1417,N_1463);
or U1523 (N_1523,N_1450,N_1495);
xor U1524 (N_1524,N_1445,N_1457);
or U1525 (N_1525,N_1447,N_1423);
or U1526 (N_1526,N_1486,N_1411);
and U1527 (N_1527,N_1487,N_1432);
nand U1528 (N_1528,N_1460,N_1491);
xor U1529 (N_1529,N_1425,N_1426);
nor U1530 (N_1530,N_1427,N_1415);
and U1531 (N_1531,N_1403,N_1421);
nand U1532 (N_1532,N_1422,N_1401);
nor U1533 (N_1533,N_1482,N_1456);
or U1534 (N_1534,N_1418,N_1436);
nor U1535 (N_1535,N_1442,N_1488);
and U1536 (N_1536,N_1416,N_1437);
nor U1537 (N_1537,N_1461,N_1466);
nand U1538 (N_1538,N_1481,N_1414);
or U1539 (N_1539,N_1484,N_1405);
xor U1540 (N_1540,N_1498,N_1499);
nor U1541 (N_1541,N_1478,N_1407);
xor U1542 (N_1542,N_1496,N_1453);
nor U1543 (N_1543,N_1404,N_1497);
xnor U1544 (N_1544,N_1480,N_1409);
nor U1545 (N_1545,N_1439,N_1476);
xor U1546 (N_1546,N_1420,N_1472);
nand U1547 (N_1547,N_1459,N_1408);
and U1548 (N_1548,N_1485,N_1483);
nor U1549 (N_1549,N_1473,N_1479);
xnor U1550 (N_1550,N_1433,N_1474);
nor U1551 (N_1551,N_1466,N_1419);
and U1552 (N_1552,N_1438,N_1498);
nor U1553 (N_1553,N_1472,N_1413);
nor U1554 (N_1554,N_1492,N_1465);
nand U1555 (N_1555,N_1498,N_1476);
nor U1556 (N_1556,N_1463,N_1434);
nand U1557 (N_1557,N_1419,N_1483);
xnor U1558 (N_1558,N_1431,N_1498);
and U1559 (N_1559,N_1404,N_1418);
and U1560 (N_1560,N_1428,N_1437);
xnor U1561 (N_1561,N_1456,N_1493);
or U1562 (N_1562,N_1459,N_1484);
nor U1563 (N_1563,N_1450,N_1421);
xnor U1564 (N_1564,N_1475,N_1451);
and U1565 (N_1565,N_1448,N_1474);
nor U1566 (N_1566,N_1413,N_1409);
xor U1567 (N_1567,N_1421,N_1491);
nand U1568 (N_1568,N_1454,N_1430);
or U1569 (N_1569,N_1485,N_1436);
nor U1570 (N_1570,N_1440,N_1485);
and U1571 (N_1571,N_1438,N_1400);
or U1572 (N_1572,N_1438,N_1455);
nor U1573 (N_1573,N_1480,N_1493);
and U1574 (N_1574,N_1460,N_1408);
nor U1575 (N_1575,N_1442,N_1496);
nand U1576 (N_1576,N_1455,N_1495);
and U1577 (N_1577,N_1445,N_1425);
or U1578 (N_1578,N_1435,N_1446);
nand U1579 (N_1579,N_1488,N_1496);
or U1580 (N_1580,N_1465,N_1461);
and U1581 (N_1581,N_1461,N_1431);
or U1582 (N_1582,N_1444,N_1454);
nor U1583 (N_1583,N_1487,N_1433);
nor U1584 (N_1584,N_1401,N_1400);
nor U1585 (N_1585,N_1448,N_1492);
nor U1586 (N_1586,N_1413,N_1451);
and U1587 (N_1587,N_1427,N_1474);
and U1588 (N_1588,N_1459,N_1458);
xor U1589 (N_1589,N_1496,N_1443);
nand U1590 (N_1590,N_1444,N_1402);
nor U1591 (N_1591,N_1478,N_1438);
or U1592 (N_1592,N_1450,N_1420);
or U1593 (N_1593,N_1430,N_1491);
nor U1594 (N_1594,N_1488,N_1478);
nor U1595 (N_1595,N_1427,N_1448);
nor U1596 (N_1596,N_1487,N_1454);
or U1597 (N_1597,N_1435,N_1444);
and U1598 (N_1598,N_1411,N_1419);
and U1599 (N_1599,N_1445,N_1458);
xnor U1600 (N_1600,N_1543,N_1528);
nand U1601 (N_1601,N_1595,N_1504);
nand U1602 (N_1602,N_1514,N_1570);
or U1603 (N_1603,N_1574,N_1555);
nand U1604 (N_1604,N_1524,N_1538);
xor U1605 (N_1605,N_1580,N_1591);
nand U1606 (N_1606,N_1507,N_1596);
nor U1607 (N_1607,N_1590,N_1508);
or U1608 (N_1608,N_1513,N_1581);
or U1609 (N_1609,N_1573,N_1522);
xnor U1610 (N_1610,N_1536,N_1537);
nor U1611 (N_1611,N_1586,N_1558);
nand U1612 (N_1612,N_1523,N_1568);
nand U1613 (N_1613,N_1593,N_1525);
xnor U1614 (N_1614,N_1566,N_1561);
or U1615 (N_1615,N_1547,N_1521);
or U1616 (N_1616,N_1571,N_1501);
and U1617 (N_1617,N_1535,N_1518);
and U1618 (N_1618,N_1510,N_1577);
and U1619 (N_1619,N_1526,N_1585);
xnor U1620 (N_1620,N_1506,N_1515);
and U1621 (N_1621,N_1592,N_1562);
and U1622 (N_1622,N_1587,N_1544);
nand U1623 (N_1623,N_1563,N_1503);
nand U1624 (N_1624,N_1519,N_1589);
nor U1625 (N_1625,N_1541,N_1545);
xnor U1626 (N_1626,N_1575,N_1505);
xnor U1627 (N_1627,N_1540,N_1549);
and U1628 (N_1628,N_1552,N_1530);
xor U1629 (N_1629,N_1527,N_1582);
xor U1630 (N_1630,N_1557,N_1516);
nor U1631 (N_1631,N_1567,N_1583);
or U1632 (N_1632,N_1532,N_1546);
and U1633 (N_1633,N_1529,N_1500);
nor U1634 (N_1634,N_1539,N_1578);
nand U1635 (N_1635,N_1559,N_1550);
xnor U1636 (N_1636,N_1548,N_1564);
and U1637 (N_1637,N_1531,N_1576);
or U1638 (N_1638,N_1511,N_1569);
or U1639 (N_1639,N_1597,N_1560);
and U1640 (N_1640,N_1553,N_1551);
nor U1641 (N_1641,N_1509,N_1598);
nor U1642 (N_1642,N_1579,N_1554);
xnor U1643 (N_1643,N_1542,N_1517);
nor U1644 (N_1644,N_1520,N_1572);
nor U1645 (N_1645,N_1565,N_1594);
xnor U1646 (N_1646,N_1534,N_1599);
and U1647 (N_1647,N_1512,N_1556);
or U1648 (N_1648,N_1533,N_1502);
nor U1649 (N_1649,N_1584,N_1588);
xor U1650 (N_1650,N_1523,N_1552);
nand U1651 (N_1651,N_1519,N_1555);
nor U1652 (N_1652,N_1548,N_1560);
or U1653 (N_1653,N_1518,N_1573);
or U1654 (N_1654,N_1511,N_1531);
xor U1655 (N_1655,N_1506,N_1580);
or U1656 (N_1656,N_1574,N_1590);
and U1657 (N_1657,N_1545,N_1578);
xnor U1658 (N_1658,N_1561,N_1505);
and U1659 (N_1659,N_1511,N_1550);
nor U1660 (N_1660,N_1527,N_1517);
or U1661 (N_1661,N_1544,N_1534);
and U1662 (N_1662,N_1553,N_1597);
nand U1663 (N_1663,N_1545,N_1546);
nand U1664 (N_1664,N_1570,N_1582);
and U1665 (N_1665,N_1545,N_1534);
nand U1666 (N_1666,N_1506,N_1586);
and U1667 (N_1667,N_1564,N_1540);
or U1668 (N_1668,N_1570,N_1501);
xnor U1669 (N_1669,N_1563,N_1584);
or U1670 (N_1670,N_1524,N_1585);
and U1671 (N_1671,N_1553,N_1546);
or U1672 (N_1672,N_1538,N_1597);
nor U1673 (N_1673,N_1552,N_1541);
nand U1674 (N_1674,N_1594,N_1532);
and U1675 (N_1675,N_1528,N_1555);
and U1676 (N_1676,N_1598,N_1520);
and U1677 (N_1677,N_1599,N_1585);
and U1678 (N_1678,N_1579,N_1544);
xnor U1679 (N_1679,N_1585,N_1562);
and U1680 (N_1680,N_1560,N_1526);
xnor U1681 (N_1681,N_1573,N_1509);
nand U1682 (N_1682,N_1518,N_1586);
nor U1683 (N_1683,N_1548,N_1580);
xor U1684 (N_1684,N_1590,N_1592);
xor U1685 (N_1685,N_1549,N_1527);
xnor U1686 (N_1686,N_1580,N_1577);
or U1687 (N_1687,N_1578,N_1533);
or U1688 (N_1688,N_1523,N_1555);
and U1689 (N_1689,N_1575,N_1522);
xor U1690 (N_1690,N_1591,N_1597);
and U1691 (N_1691,N_1519,N_1561);
nand U1692 (N_1692,N_1589,N_1576);
nor U1693 (N_1693,N_1506,N_1579);
xnor U1694 (N_1694,N_1518,N_1502);
or U1695 (N_1695,N_1572,N_1592);
or U1696 (N_1696,N_1591,N_1535);
and U1697 (N_1697,N_1554,N_1552);
xnor U1698 (N_1698,N_1507,N_1566);
xnor U1699 (N_1699,N_1532,N_1595);
nand U1700 (N_1700,N_1670,N_1696);
xor U1701 (N_1701,N_1629,N_1638);
xnor U1702 (N_1702,N_1664,N_1648);
nand U1703 (N_1703,N_1627,N_1693);
xor U1704 (N_1704,N_1600,N_1640);
or U1705 (N_1705,N_1657,N_1605);
and U1706 (N_1706,N_1612,N_1667);
and U1707 (N_1707,N_1609,N_1675);
nand U1708 (N_1708,N_1635,N_1634);
and U1709 (N_1709,N_1613,N_1681);
nor U1710 (N_1710,N_1644,N_1677);
nand U1711 (N_1711,N_1689,N_1669);
and U1712 (N_1712,N_1645,N_1652);
xor U1713 (N_1713,N_1687,N_1625);
nand U1714 (N_1714,N_1630,N_1617);
nand U1715 (N_1715,N_1653,N_1606);
and U1716 (N_1716,N_1695,N_1643);
nand U1717 (N_1717,N_1619,N_1622);
or U1718 (N_1718,N_1694,N_1685);
nand U1719 (N_1719,N_1679,N_1607);
or U1720 (N_1720,N_1697,N_1632);
and U1721 (N_1721,N_1647,N_1671);
or U1722 (N_1722,N_1601,N_1688);
nor U1723 (N_1723,N_1610,N_1608);
and U1724 (N_1724,N_1639,N_1641);
nor U1725 (N_1725,N_1626,N_1650);
nor U1726 (N_1726,N_1649,N_1642);
xor U1727 (N_1727,N_1680,N_1656);
nand U1728 (N_1728,N_1623,N_1690);
nor U1729 (N_1729,N_1651,N_1691);
or U1730 (N_1730,N_1633,N_1646);
nor U1731 (N_1731,N_1662,N_1660);
nand U1732 (N_1732,N_1673,N_1628);
nor U1733 (N_1733,N_1676,N_1668);
xnor U1734 (N_1734,N_1636,N_1659);
and U1735 (N_1735,N_1616,N_1637);
or U1736 (N_1736,N_1611,N_1604);
or U1737 (N_1737,N_1603,N_1682);
and U1738 (N_1738,N_1699,N_1684);
nand U1739 (N_1739,N_1683,N_1624);
nand U1740 (N_1740,N_1621,N_1672);
and U1741 (N_1741,N_1666,N_1655);
or U1742 (N_1742,N_1674,N_1620);
xnor U1743 (N_1743,N_1678,N_1654);
xor U1744 (N_1744,N_1631,N_1686);
nand U1745 (N_1745,N_1615,N_1665);
nand U1746 (N_1746,N_1692,N_1661);
nand U1747 (N_1747,N_1663,N_1698);
or U1748 (N_1748,N_1614,N_1618);
nor U1749 (N_1749,N_1602,N_1658);
nand U1750 (N_1750,N_1638,N_1687);
xor U1751 (N_1751,N_1619,N_1621);
nand U1752 (N_1752,N_1674,N_1688);
and U1753 (N_1753,N_1690,N_1603);
or U1754 (N_1754,N_1655,N_1605);
or U1755 (N_1755,N_1668,N_1614);
and U1756 (N_1756,N_1601,N_1637);
xor U1757 (N_1757,N_1659,N_1656);
xor U1758 (N_1758,N_1644,N_1652);
nor U1759 (N_1759,N_1680,N_1686);
and U1760 (N_1760,N_1638,N_1686);
xor U1761 (N_1761,N_1696,N_1665);
xor U1762 (N_1762,N_1650,N_1645);
or U1763 (N_1763,N_1644,N_1689);
nand U1764 (N_1764,N_1634,N_1698);
or U1765 (N_1765,N_1655,N_1626);
xnor U1766 (N_1766,N_1624,N_1623);
nand U1767 (N_1767,N_1661,N_1681);
or U1768 (N_1768,N_1649,N_1677);
nand U1769 (N_1769,N_1644,N_1653);
or U1770 (N_1770,N_1650,N_1641);
nor U1771 (N_1771,N_1656,N_1679);
xor U1772 (N_1772,N_1621,N_1648);
and U1773 (N_1773,N_1626,N_1654);
and U1774 (N_1774,N_1621,N_1631);
and U1775 (N_1775,N_1659,N_1613);
nand U1776 (N_1776,N_1612,N_1681);
and U1777 (N_1777,N_1605,N_1614);
xor U1778 (N_1778,N_1672,N_1605);
and U1779 (N_1779,N_1686,N_1634);
or U1780 (N_1780,N_1692,N_1694);
xor U1781 (N_1781,N_1634,N_1626);
and U1782 (N_1782,N_1681,N_1699);
nand U1783 (N_1783,N_1691,N_1601);
nor U1784 (N_1784,N_1699,N_1604);
nor U1785 (N_1785,N_1627,N_1694);
and U1786 (N_1786,N_1614,N_1675);
nor U1787 (N_1787,N_1611,N_1659);
or U1788 (N_1788,N_1681,N_1651);
nand U1789 (N_1789,N_1686,N_1690);
and U1790 (N_1790,N_1668,N_1691);
nand U1791 (N_1791,N_1668,N_1661);
nor U1792 (N_1792,N_1625,N_1654);
xnor U1793 (N_1793,N_1646,N_1665);
xnor U1794 (N_1794,N_1640,N_1660);
or U1795 (N_1795,N_1639,N_1687);
nor U1796 (N_1796,N_1607,N_1604);
nor U1797 (N_1797,N_1690,N_1667);
nor U1798 (N_1798,N_1624,N_1640);
or U1799 (N_1799,N_1640,N_1634);
and U1800 (N_1800,N_1729,N_1739);
xnor U1801 (N_1801,N_1709,N_1789);
xnor U1802 (N_1802,N_1771,N_1732);
nor U1803 (N_1803,N_1795,N_1715);
xor U1804 (N_1804,N_1767,N_1720);
nor U1805 (N_1805,N_1755,N_1722);
or U1806 (N_1806,N_1791,N_1716);
and U1807 (N_1807,N_1714,N_1758);
or U1808 (N_1808,N_1798,N_1718);
nor U1809 (N_1809,N_1770,N_1799);
and U1810 (N_1810,N_1701,N_1785);
or U1811 (N_1811,N_1766,N_1719);
xor U1812 (N_1812,N_1700,N_1752);
nand U1813 (N_1813,N_1743,N_1703);
nor U1814 (N_1814,N_1759,N_1733);
nand U1815 (N_1815,N_1749,N_1708);
nor U1816 (N_1816,N_1778,N_1757);
nand U1817 (N_1817,N_1737,N_1765);
or U1818 (N_1818,N_1727,N_1774);
xor U1819 (N_1819,N_1702,N_1721);
xor U1820 (N_1820,N_1777,N_1797);
nand U1821 (N_1821,N_1787,N_1736);
and U1822 (N_1822,N_1753,N_1741);
xor U1823 (N_1823,N_1760,N_1745);
nor U1824 (N_1824,N_1713,N_1779);
and U1825 (N_1825,N_1790,N_1761);
and U1826 (N_1826,N_1772,N_1705);
or U1827 (N_1827,N_1738,N_1768);
or U1828 (N_1828,N_1746,N_1762);
or U1829 (N_1829,N_1792,N_1784);
nand U1830 (N_1830,N_1794,N_1751);
or U1831 (N_1831,N_1782,N_1756);
or U1832 (N_1832,N_1740,N_1724);
xnor U1833 (N_1833,N_1728,N_1735);
xnor U1834 (N_1834,N_1734,N_1747);
nor U1835 (N_1835,N_1780,N_1744);
xnor U1836 (N_1836,N_1754,N_1730);
and U1837 (N_1837,N_1786,N_1764);
or U1838 (N_1838,N_1748,N_1726);
or U1839 (N_1839,N_1710,N_1711);
and U1840 (N_1840,N_1796,N_1717);
nand U1841 (N_1841,N_1723,N_1707);
or U1842 (N_1842,N_1775,N_1750);
xor U1843 (N_1843,N_1773,N_1781);
or U1844 (N_1844,N_1704,N_1725);
xnor U1845 (N_1845,N_1776,N_1793);
nand U1846 (N_1846,N_1783,N_1706);
xnor U1847 (N_1847,N_1788,N_1769);
or U1848 (N_1848,N_1742,N_1712);
xnor U1849 (N_1849,N_1763,N_1731);
and U1850 (N_1850,N_1768,N_1764);
xor U1851 (N_1851,N_1777,N_1781);
nand U1852 (N_1852,N_1704,N_1753);
and U1853 (N_1853,N_1788,N_1727);
or U1854 (N_1854,N_1702,N_1775);
nor U1855 (N_1855,N_1772,N_1717);
nor U1856 (N_1856,N_1793,N_1732);
xnor U1857 (N_1857,N_1721,N_1778);
and U1858 (N_1858,N_1734,N_1766);
or U1859 (N_1859,N_1780,N_1705);
nand U1860 (N_1860,N_1784,N_1706);
xor U1861 (N_1861,N_1760,N_1722);
or U1862 (N_1862,N_1752,N_1769);
or U1863 (N_1863,N_1788,N_1749);
or U1864 (N_1864,N_1787,N_1784);
and U1865 (N_1865,N_1790,N_1749);
nor U1866 (N_1866,N_1714,N_1708);
nor U1867 (N_1867,N_1791,N_1759);
nand U1868 (N_1868,N_1791,N_1740);
or U1869 (N_1869,N_1797,N_1776);
nand U1870 (N_1870,N_1790,N_1799);
or U1871 (N_1871,N_1798,N_1745);
nor U1872 (N_1872,N_1763,N_1771);
or U1873 (N_1873,N_1726,N_1783);
or U1874 (N_1874,N_1784,N_1704);
or U1875 (N_1875,N_1764,N_1780);
or U1876 (N_1876,N_1789,N_1705);
and U1877 (N_1877,N_1786,N_1758);
nor U1878 (N_1878,N_1788,N_1723);
nor U1879 (N_1879,N_1768,N_1749);
nand U1880 (N_1880,N_1743,N_1715);
nor U1881 (N_1881,N_1738,N_1796);
and U1882 (N_1882,N_1718,N_1776);
nand U1883 (N_1883,N_1774,N_1741);
xor U1884 (N_1884,N_1713,N_1702);
nor U1885 (N_1885,N_1772,N_1724);
xnor U1886 (N_1886,N_1756,N_1751);
nand U1887 (N_1887,N_1709,N_1707);
xor U1888 (N_1888,N_1763,N_1786);
nand U1889 (N_1889,N_1758,N_1797);
nand U1890 (N_1890,N_1762,N_1711);
nand U1891 (N_1891,N_1737,N_1775);
nor U1892 (N_1892,N_1709,N_1726);
nand U1893 (N_1893,N_1703,N_1772);
or U1894 (N_1894,N_1707,N_1733);
xnor U1895 (N_1895,N_1799,N_1760);
xor U1896 (N_1896,N_1767,N_1719);
nand U1897 (N_1897,N_1780,N_1799);
and U1898 (N_1898,N_1772,N_1745);
xor U1899 (N_1899,N_1793,N_1756);
and U1900 (N_1900,N_1840,N_1874);
nor U1901 (N_1901,N_1882,N_1841);
and U1902 (N_1902,N_1839,N_1848);
nor U1903 (N_1903,N_1867,N_1887);
xor U1904 (N_1904,N_1827,N_1842);
nand U1905 (N_1905,N_1833,N_1844);
or U1906 (N_1906,N_1801,N_1828);
xnor U1907 (N_1907,N_1823,N_1829);
and U1908 (N_1908,N_1845,N_1805);
or U1909 (N_1909,N_1885,N_1895);
or U1910 (N_1910,N_1836,N_1821);
or U1911 (N_1911,N_1822,N_1806);
or U1912 (N_1912,N_1859,N_1809);
xor U1913 (N_1913,N_1877,N_1897);
or U1914 (N_1914,N_1866,N_1824);
and U1915 (N_1915,N_1883,N_1888);
nor U1916 (N_1916,N_1818,N_1856);
nand U1917 (N_1917,N_1868,N_1802);
or U1918 (N_1918,N_1872,N_1855);
nand U1919 (N_1919,N_1870,N_1843);
xor U1920 (N_1920,N_1826,N_1837);
xor U1921 (N_1921,N_1832,N_1814);
or U1922 (N_1922,N_1862,N_1871);
nor U1923 (N_1923,N_1854,N_1876);
xnor U1924 (N_1924,N_1899,N_1830);
nand U1925 (N_1925,N_1834,N_1811);
or U1926 (N_1926,N_1820,N_1890);
xor U1927 (N_1927,N_1891,N_1861);
or U1928 (N_1928,N_1803,N_1851);
and U1929 (N_1929,N_1879,N_1847);
or U1930 (N_1930,N_1860,N_1800);
xnor U1931 (N_1931,N_1863,N_1894);
nor U1932 (N_1932,N_1857,N_1804);
nand U1933 (N_1933,N_1869,N_1853);
and U1934 (N_1934,N_1846,N_1884);
and U1935 (N_1935,N_1849,N_1808);
or U1936 (N_1936,N_1807,N_1865);
and U1937 (N_1937,N_1813,N_1893);
and U1938 (N_1938,N_1875,N_1815);
nand U1939 (N_1939,N_1810,N_1873);
nor U1940 (N_1940,N_1898,N_1819);
or U1941 (N_1941,N_1881,N_1817);
nand U1942 (N_1942,N_1880,N_1878);
xnor U1943 (N_1943,N_1850,N_1838);
or U1944 (N_1944,N_1892,N_1858);
and U1945 (N_1945,N_1852,N_1812);
and U1946 (N_1946,N_1896,N_1889);
xnor U1947 (N_1947,N_1886,N_1825);
nor U1948 (N_1948,N_1831,N_1864);
nand U1949 (N_1949,N_1835,N_1816);
nor U1950 (N_1950,N_1824,N_1811);
or U1951 (N_1951,N_1854,N_1857);
and U1952 (N_1952,N_1890,N_1896);
nand U1953 (N_1953,N_1875,N_1840);
nand U1954 (N_1954,N_1890,N_1883);
xnor U1955 (N_1955,N_1827,N_1808);
and U1956 (N_1956,N_1856,N_1860);
and U1957 (N_1957,N_1878,N_1871);
or U1958 (N_1958,N_1800,N_1806);
xnor U1959 (N_1959,N_1892,N_1831);
or U1960 (N_1960,N_1880,N_1821);
and U1961 (N_1961,N_1884,N_1819);
nor U1962 (N_1962,N_1843,N_1858);
nor U1963 (N_1963,N_1807,N_1826);
or U1964 (N_1964,N_1873,N_1842);
or U1965 (N_1965,N_1854,N_1858);
nand U1966 (N_1966,N_1862,N_1882);
and U1967 (N_1967,N_1844,N_1875);
xnor U1968 (N_1968,N_1844,N_1807);
nand U1969 (N_1969,N_1823,N_1899);
nor U1970 (N_1970,N_1879,N_1807);
xor U1971 (N_1971,N_1857,N_1894);
nand U1972 (N_1972,N_1804,N_1824);
nand U1973 (N_1973,N_1811,N_1879);
nand U1974 (N_1974,N_1831,N_1865);
nand U1975 (N_1975,N_1849,N_1840);
and U1976 (N_1976,N_1824,N_1801);
nor U1977 (N_1977,N_1836,N_1876);
or U1978 (N_1978,N_1862,N_1816);
nand U1979 (N_1979,N_1863,N_1812);
nand U1980 (N_1980,N_1811,N_1817);
xnor U1981 (N_1981,N_1818,N_1870);
or U1982 (N_1982,N_1839,N_1860);
nand U1983 (N_1983,N_1878,N_1888);
or U1984 (N_1984,N_1884,N_1806);
or U1985 (N_1985,N_1837,N_1813);
or U1986 (N_1986,N_1858,N_1830);
nand U1987 (N_1987,N_1829,N_1815);
nor U1988 (N_1988,N_1898,N_1833);
and U1989 (N_1989,N_1853,N_1873);
and U1990 (N_1990,N_1896,N_1837);
nand U1991 (N_1991,N_1871,N_1803);
and U1992 (N_1992,N_1881,N_1847);
nor U1993 (N_1993,N_1830,N_1804);
nand U1994 (N_1994,N_1871,N_1844);
or U1995 (N_1995,N_1869,N_1804);
nor U1996 (N_1996,N_1867,N_1818);
nand U1997 (N_1997,N_1850,N_1842);
nor U1998 (N_1998,N_1847,N_1831);
nand U1999 (N_1999,N_1816,N_1883);
xnor U2000 (N_2000,N_1947,N_1905);
and U2001 (N_2001,N_1954,N_1964);
xor U2002 (N_2002,N_1911,N_1993);
nor U2003 (N_2003,N_1961,N_1910);
xnor U2004 (N_2004,N_1935,N_1968);
and U2005 (N_2005,N_1907,N_1986);
xor U2006 (N_2006,N_1999,N_1976);
nor U2007 (N_2007,N_1920,N_1943);
nand U2008 (N_2008,N_1962,N_1927);
nor U2009 (N_2009,N_1966,N_1909);
nand U2010 (N_2010,N_1984,N_1938);
or U2011 (N_2011,N_1967,N_1924);
and U2012 (N_2012,N_1987,N_1979);
or U2013 (N_2013,N_1992,N_1958);
xor U2014 (N_2014,N_1914,N_1973);
and U2015 (N_2015,N_1931,N_1998);
xor U2016 (N_2016,N_1952,N_1974);
and U2017 (N_2017,N_1906,N_1980);
nor U2018 (N_2018,N_1903,N_1960);
or U2019 (N_2019,N_1955,N_1915);
xnor U2020 (N_2020,N_1957,N_1971);
nand U2021 (N_2021,N_1946,N_1941);
nand U2022 (N_2022,N_1983,N_1939);
nand U2023 (N_2023,N_1995,N_1975);
nor U2024 (N_2024,N_1990,N_1908);
nor U2025 (N_2025,N_1940,N_1919);
nor U2026 (N_2026,N_1949,N_1944);
xnor U2027 (N_2027,N_1922,N_1997);
nor U2028 (N_2028,N_1965,N_1948);
or U2029 (N_2029,N_1972,N_1932);
nand U2030 (N_2030,N_1937,N_1981);
nand U2031 (N_2031,N_1928,N_1977);
nand U2032 (N_2032,N_1913,N_1978);
and U2033 (N_2033,N_1916,N_1982);
xor U2034 (N_2034,N_1951,N_1989);
xnor U2035 (N_2035,N_1963,N_1900);
or U2036 (N_2036,N_1917,N_1959);
and U2037 (N_2037,N_1969,N_1912);
nand U2038 (N_2038,N_1936,N_1934);
xnor U2039 (N_2039,N_1923,N_1901);
nand U2040 (N_2040,N_1902,N_1970);
nand U2041 (N_2041,N_1996,N_1933);
or U2042 (N_2042,N_1953,N_1988);
nor U2043 (N_2043,N_1929,N_1925);
xor U2044 (N_2044,N_1985,N_1926);
or U2045 (N_2045,N_1994,N_1950);
and U2046 (N_2046,N_1918,N_1942);
and U2047 (N_2047,N_1945,N_1930);
nand U2048 (N_2048,N_1921,N_1956);
nand U2049 (N_2049,N_1991,N_1904);
and U2050 (N_2050,N_1989,N_1941);
or U2051 (N_2051,N_1912,N_1993);
or U2052 (N_2052,N_1900,N_1924);
xor U2053 (N_2053,N_1963,N_1913);
nor U2054 (N_2054,N_1951,N_1995);
nor U2055 (N_2055,N_1996,N_1925);
xor U2056 (N_2056,N_1969,N_1988);
nand U2057 (N_2057,N_1937,N_1948);
nor U2058 (N_2058,N_1964,N_1942);
xor U2059 (N_2059,N_1943,N_1953);
nand U2060 (N_2060,N_1981,N_1985);
nor U2061 (N_2061,N_1982,N_1984);
or U2062 (N_2062,N_1961,N_1990);
or U2063 (N_2063,N_1968,N_1947);
nand U2064 (N_2064,N_1968,N_1921);
or U2065 (N_2065,N_1989,N_1920);
nor U2066 (N_2066,N_1918,N_1995);
xnor U2067 (N_2067,N_1907,N_1904);
nand U2068 (N_2068,N_1999,N_1923);
or U2069 (N_2069,N_1997,N_1968);
and U2070 (N_2070,N_1959,N_1924);
and U2071 (N_2071,N_1936,N_1961);
nand U2072 (N_2072,N_1993,N_1927);
nand U2073 (N_2073,N_1950,N_1908);
nand U2074 (N_2074,N_1900,N_1983);
or U2075 (N_2075,N_1905,N_1931);
xnor U2076 (N_2076,N_1977,N_1999);
nor U2077 (N_2077,N_1968,N_1928);
or U2078 (N_2078,N_1918,N_1917);
or U2079 (N_2079,N_1956,N_1971);
or U2080 (N_2080,N_1943,N_1967);
nor U2081 (N_2081,N_1985,N_1921);
nor U2082 (N_2082,N_1904,N_1914);
and U2083 (N_2083,N_1978,N_1995);
or U2084 (N_2084,N_1970,N_1999);
or U2085 (N_2085,N_1956,N_1979);
or U2086 (N_2086,N_1906,N_1996);
nor U2087 (N_2087,N_1933,N_1952);
nand U2088 (N_2088,N_1965,N_1931);
nand U2089 (N_2089,N_1930,N_1942);
nand U2090 (N_2090,N_1944,N_1998);
nor U2091 (N_2091,N_1960,N_1995);
or U2092 (N_2092,N_1972,N_1915);
nand U2093 (N_2093,N_1913,N_1911);
and U2094 (N_2094,N_1907,N_1970);
xor U2095 (N_2095,N_1926,N_1986);
and U2096 (N_2096,N_1960,N_1984);
nor U2097 (N_2097,N_1940,N_1964);
nand U2098 (N_2098,N_1976,N_1956);
nor U2099 (N_2099,N_1903,N_1936);
or U2100 (N_2100,N_2052,N_2051);
and U2101 (N_2101,N_2065,N_2079);
and U2102 (N_2102,N_2000,N_2070);
and U2103 (N_2103,N_2064,N_2087);
or U2104 (N_2104,N_2057,N_2032);
nor U2105 (N_2105,N_2068,N_2080);
or U2106 (N_2106,N_2004,N_2010);
and U2107 (N_2107,N_2003,N_2069);
or U2108 (N_2108,N_2088,N_2085);
nor U2109 (N_2109,N_2055,N_2029);
or U2110 (N_2110,N_2031,N_2047);
and U2111 (N_2111,N_2006,N_2098);
and U2112 (N_2112,N_2063,N_2053);
nor U2113 (N_2113,N_2081,N_2027);
nand U2114 (N_2114,N_2019,N_2048);
nor U2115 (N_2115,N_2056,N_2038);
nor U2116 (N_2116,N_2015,N_2062);
nor U2117 (N_2117,N_2086,N_2084);
or U2118 (N_2118,N_2016,N_2049);
nand U2119 (N_2119,N_2024,N_2090);
xnor U2120 (N_2120,N_2075,N_2060);
nand U2121 (N_2121,N_2037,N_2005);
nand U2122 (N_2122,N_2040,N_2092);
nor U2123 (N_2123,N_2041,N_2091);
nor U2124 (N_2124,N_2007,N_2046);
or U2125 (N_2125,N_2061,N_2073);
nand U2126 (N_2126,N_2059,N_2009);
or U2127 (N_2127,N_2012,N_2039);
nand U2128 (N_2128,N_2023,N_2001);
nand U2129 (N_2129,N_2026,N_2066);
and U2130 (N_2130,N_2067,N_2028);
nand U2131 (N_2131,N_2021,N_2089);
and U2132 (N_2132,N_2017,N_2044);
nor U2133 (N_2133,N_2008,N_2022);
nor U2134 (N_2134,N_2045,N_2025);
or U2135 (N_2135,N_2095,N_2076);
nand U2136 (N_2136,N_2034,N_2050);
nand U2137 (N_2137,N_2042,N_2018);
and U2138 (N_2138,N_2097,N_2096);
or U2139 (N_2139,N_2035,N_2077);
nor U2140 (N_2140,N_2071,N_2013);
and U2141 (N_2141,N_2074,N_2082);
or U2142 (N_2142,N_2014,N_2020);
or U2143 (N_2143,N_2043,N_2058);
and U2144 (N_2144,N_2054,N_2036);
nor U2145 (N_2145,N_2078,N_2002);
xor U2146 (N_2146,N_2083,N_2099);
and U2147 (N_2147,N_2094,N_2030);
or U2148 (N_2148,N_2072,N_2093);
nor U2149 (N_2149,N_2033,N_2011);
nand U2150 (N_2150,N_2034,N_2059);
nand U2151 (N_2151,N_2022,N_2046);
xor U2152 (N_2152,N_2097,N_2066);
nand U2153 (N_2153,N_2079,N_2017);
and U2154 (N_2154,N_2020,N_2096);
xnor U2155 (N_2155,N_2031,N_2008);
and U2156 (N_2156,N_2031,N_2053);
and U2157 (N_2157,N_2052,N_2033);
and U2158 (N_2158,N_2065,N_2039);
and U2159 (N_2159,N_2048,N_2035);
nand U2160 (N_2160,N_2053,N_2012);
nor U2161 (N_2161,N_2083,N_2021);
xor U2162 (N_2162,N_2010,N_2085);
nor U2163 (N_2163,N_2010,N_2092);
or U2164 (N_2164,N_2029,N_2046);
xor U2165 (N_2165,N_2011,N_2044);
xor U2166 (N_2166,N_2060,N_2051);
xnor U2167 (N_2167,N_2054,N_2053);
nand U2168 (N_2168,N_2027,N_2057);
and U2169 (N_2169,N_2091,N_2037);
nand U2170 (N_2170,N_2059,N_2017);
nor U2171 (N_2171,N_2079,N_2037);
nor U2172 (N_2172,N_2053,N_2011);
nor U2173 (N_2173,N_2060,N_2037);
or U2174 (N_2174,N_2021,N_2024);
xor U2175 (N_2175,N_2050,N_2031);
and U2176 (N_2176,N_2017,N_2040);
nor U2177 (N_2177,N_2088,N_2084);
nor U2178 (N_2178,N_2077,N_2002);
or U2179 (N_2179,N_2093,N_2017);
nand U2180 (N_2180,N_2028,N_2015);
and U2181 (N_2181,N_2003,N_2013);
or U2182 (N_2182,N_2030,N_2056);
xor U2183 (N_2183,N_2014,N_2092);
xnor U2184 (N_2184,N_2037,N_2047);
or U2185 (N_2185,N_2007,N_2087);
nand U2186 (N_2186,N_2081,N_2021);
and U2187 (N_2187,N_2044,N_2081);
nor U2188 (N_2188,N_2046,N_2064);
or U2189 (N_2189,N_2089,N_2030);
and U2190 (N_2190,N_2044,N_2028);
nand U2191 (N_2191,N_2031,N_2017);
xnor U2192 (N_2192,N_2036,N_2057);
nor U2193 (N_2193,N_2040,N_2002);
xnor U2194 (N_2194,N_2045,N_2091);
xor U2195 (N_2195,N_2022,N_2010);
nand U2196 (N_2196,N_2078,N_2036);
nand U2197 (N_2197,N_2039,N_2031);
xor U2198 (N_2198,N_2019,N_2057);
nor U2199 (N_2199,N_2050,N_2074);
nand U2200 (N_2200,N_2139,N_2127);
and U2201 (N_2201,N_2136,N_2133);
xnor U2202 (N_2202,N_2166,N_2143);
nor U2203 (N_2203,N_2104,N_2162);
xor U2204 (N_2204,N_2171,N_2101);
nand U2205 (N_2205,N_2117,N_2113);
xnor U2206 (N_2206,N_2181,N_2187);
or U2207 (N_2207,N_2114,N_2158);
xnor U2208 (N_2208,N_2174,N_2107);
or U2209 (N_2209,N_2157,N_2147);
nand U2210 (N_2210,N_2149,N_2120);
or U2211 (N_2211,N_2184,N_2154);
or U2212 (N_2212,N_2160,N_2126);
and U2213 (N_2213,N_2148,N_2137);
nor U2214 (N_2214,N_2173,N_2138);
nor U2215 (N_2215,N_2130,N_2168);
xnor U2216 (N_2216,N_2188,N_2196);
nand U2217 (N_2217,N_2183,N_2194);
nand U2218 (N_2218,N_2146,N_2161);
nand U2219 (N_2219,N_2105,N_2185);
and U2220 (N_2220,N_2134,N_2145);
and U2221 (N_2221,N_2108,N_2155);
xor U2222 (N_2222,N_2132,N_2182);
nor U2223 (N_2223,N_2150,N_2110);
xor U2224 (N_2224,N_2189,N_2169);
nand U2225 (N_2225,N_2170,N_2152);
or U2226 (N_2226,N_2167,N_2192);
nor U2227 (N_2227,N_2163,N_2135);
xor U2228 (N_2228,N_2124,N_2122);
nand U2229 (N_2229,N_2179,N_2131);
nand U2230 (N_2230,N_2156,N_2193);
nand U2231 (N_2231,N_2109,N_2165);
xnor U2232 (N_2232,N_2125,N_2178);
nand U2233 (N_2233,N_2112,N_2128);
or U2234 (N_2234,N_2197,N_2159);
or U2235 (N_2235,N_2119,N_2115);
nand U2236 (N_2236,N_2176,N_2144);
and U2237 (N_2237,N_2199,N_2175);
xnor U2238 (N_2238,N_2142,N_2172);
nor U2239 (N_2239,N_2153,N_2116);
nor U2240 (N_2240,N_2140,N_2102);
xnor U2241 (N_2241,N_2106,N_2190);
xor U2242 (N_2242,N_2103,N_2198);
and U2243 (N_2243,N_2123,N_2141);
or U2244 (N_2244,N_2118,N_2121);
xor U2245 (N_2245,N_2100,N_2129);
xnor U2246 (N_2246,N_2186,N_2180);
or U2247 (N_2247,N_2195,N_2177);
or U2248 (N_2248,N_2191,N_2164);
nand U2249 (N_2249,N_2151,N_2111);
nor U2250 (N_2250,N_2112,N_2143);
nand U2251 (N_2251,N_2101,N_2106);
xnor U2252 (N_2252,N_2150,N_2128);
nand U2253 (N_2253,N_2100,N_2124);
nand U2254 (N_2254,N_2106,N_2126);
nor U2255 (N_2255,N_2107,N_2115);
nand U2256 (N_2256,N_2151,N_2184);
nor U2257 (N_2257,N_2121,N_2147);
xnor U2258 (N_2258,N_2100,N_2160);
nand U2259 (N_2259,N_2112,N_2168);
or U2260 (N_2260,N_2141,N_2176);
xor U2261 (N_2261,N_2149,N_2126);
nand U2262 (N_2262,N_2193,N_2135);
nand U2263 (N_2263,N_2104,N_2122);
or U2264 (N_2264,N_2131,N_2150);
nor U2265 (N_2265,N_2174,N_2152);
or U2266 (N_2266,N_2101,N_2174);
and U2267 (N_2267,N_2166,N_2145);
nor U2268 (N_2268,N_2119,N_2176);
nor U2269 (N_2269,N_2103,N_2110);
xnor U2270 (N_2270,N_2178,N_2193);
xnor U2271 (N_2271,N_2125,N_2128);
and U2272 (N_2272,N_2108,N_2137);
xor U2273 (N_2273,N_2108,N_2193);
nand U2274 (N_2274,N_2156,N_2122);
nand U2275 (N_2275,N_2130,N_2185);
nor U2276 (N_2276,N_2165,N_2121);
nand U2277 (N_2277,N_2109,N_2162);
nor U2278 (N_2278,N_2193,N_2192);
or U2279 (N_2279,N_2115,N_2164);
and U2280 (N_2280,N_2191,N_2182);
xnor U2281 (N_2281,N_2128,N_2191);
or U2282 (N_2282,N_2153,N_2169);
xnor U2283 (N_2283,N_2115,N_2158);
nand U2284 (N_2284,N_2142,N_2162);
and U2285 (N_2285,N_2108,N_2132);
or U2286 (N_2286,N_2145,N_2173);
nand U2287 (N_2287,N_2131,N_2108);
and U2288 (N_2288,N_2106,N_2139);
xor U2289 (N_2289,N_2118,N_2102);
xnor U2290 (N_2290,N_2152,N_2113);
nor U2291 (N_2291,N_2195,N_2105);
nor U2292 (N_2292,N_2199,N_2146);
and U2293 (N_2293,N_2188,N_2184);
nor U2294 (N_2294,N_2192,N_2101);
nor U2295 (N_2295,N_2177,N_2126);
xnor U2296 (N_2296,N_2181,N_2110);
and U2297 (N_2297,N_2130,N_2188);
xor U2298 (N_2298,N_2142,N_2156);
nand U2299 (N_2299,N_2174,N_2100);
nand U2300 (N_2300,N_2215,N_2246);
and U2301 (N_2301,N_2249,N_2245);
xnor U2302 (N_2302,N_2232,N_2243);
nand U2303 (N_2303,N_2258,N_2201);
nor U2304 (N_2304,N_2286,N_2298);
xnor U2305 (N_2305,N_2223,N_2204);
and U2306 (N_2306,N_2296,N_2269);
xnor U2307 (N_2307,N_2202,N_2214);
and U2308 (N_2308,N_2282,N_2250);
or U2309 (N_2309,N_2244,N_2285);
nand U2310 (N_2310,N_2239,N_2275);
or U2311 (N_2311,N_2255,N_2231);
xnor U2312 (N_2312,N_2272,N_2236);
or U2313 (N_2313,N_2252,N_2206);
or U2314 (N_2314,N_2284,N_2222);
or U2315 (N_2315,N_2292,N_2248);
or U2316 (N_2316,N_2253,N_2268);
or U2317 (N_2317,N_2256,N_2230);
xnor U2318 (N_2318,N_2221,N_2277);
nand U2319 (N_2319,N_2290,N_2208);
xnor U2320 (N_2320,N_2287,N_2234);
and U2321 (N_2321,N_2218,N_2210);
or U2322 (N_2322,N_2288,N_2281);
and U2323 (N_2323,N_2293,N_2226);
xor U2324 (N_2324,N_2254,N_2264);
nor U2325 (N_2325,N_2247,N_2278);
or U2326 (N_2326,N_2203,N_2240);
nor U2327 (N_2327,N_2237,N_2228);
nand U2328 (N_2328,N_2213,N_2270);
or U2329 (N_2329,N_2283,N_2219);
xor U2330 (N_2330,N_2205,N_2242);
xor U2331 (N_2331,N_2251,N_2224);
xnor U2332 (N_2332,N_2276,N_2297);
and U2333 (N_2333,N_2279,N_2257);
or U2334 (N_2334,N_2265,N_2217);
nor U2335 (N_2335,N_2261,N_2262);
nor U2336 (N_2336,N_2207,N_2216);
xnor U2337 (N_2337,N_2294,N_2200);
xor U2338 (N_2338,N_2263,N_2211);
and U2339 (N_2339,N_2241,N_2273);
nand U2340 (N_2340,N_2274,N_2229);
xnor U2341 (N_2341,N_2227,N_2233);
nand U2342 (N_2342,N_2259,N_2267);
and U2343 (N_2343,N_2220,N_2225);
or U2344 (N_2344,N_2209,N_2260);
and U2345 (N_2345,N_2212,N_2271);
xnor U2346 (N_2346,N_2289,N_2280);
nand U2347 (N_2347,N_2235,N_2299);
xor U2348 (N_2348,N_2238,N_2295);
and U2349 (N_2349,N_2291,N_2266);
xor U2350 (N_2350,N_2283,N_2234);
or U2351 (N_2351,N_2295,N_2232);
and U2352 (N_2352,N_2210,N_2235);
and U2353 (N_2353,N_2238,N_2294);
nand U2354 (N_2354,N_2267,N_2228);
xor U2355 (N_2355,N_2251,N_2226);
and U2356 (N_2356,N_2267,N_2272);
and U2357 (N_2357,N_2275,N_2237);
and U2358 (N_2358,N_2290,N_2288);
and U2359 (N_2359,N_2249,N_2251);
and U2360 (N_2360,N_2243,N_2268);
xnor U2361 (N_2361,N_2265,N_2210);
or U2362 (N_2362,N_2299,N_2249);
or U2363 (N_2363,N_2266,N_2240);
nand U2364 (N_2364,N_2265,N_2276);
and U2365 (N_2365,N_2225,N_2294);
xor U2366 (N_2366,N_2248,N_2274);
nand U2367 (N_2367,N_2229,N_2221);
and U2368 (N_2368,N_2297,N_2284);
nor U2369 (N_2369,N_2296,N_2271);
and U2370 (N_2370,N_2260,N_2211);
nand U2371 (N_2371,N_2243,N_2204);
xnor U2372 (N_2372,N_2260,N_2274);
nand U2373 (N_2373,N_2234,N_2294);
xnor U2374 (N_2374,N_2206,N_2233);
nand U2375 (N_2375,N_2299,N_2263);
xor U2376 (N_2376,N_2202,N_2230);
xor U2377 (N_2377,N_2268,N_2212);
and U2378 (N_2378,N_2284,N_2263);
or U2379 (N_2379,N_2275,N_2214);
nor U2380 (N_2380,N_2252,N_2235);
xnor U2381 (N_2381,N_2202,N_2298);
xor U2382 (N_2382,N_2282,N_2271);
or U2383 (N_2383,N_2280,N_2291);
nor U2384 (N_2384,N_2294,N_2227);
xnor U2385 (N_2385,N_2285,N_2241);
and U2386 (N_2386,N_2244,N_2233);
nand U2387 (N_2387,N_2208,N_2297);
or U2388 (N_2388,N_2286,N_2201);
nand U2389 (N_2389,N_2246,N_2264);
nor U2390 (N_2390,N_2260,N_2235);
nor U2391 (N_2391,N_2216,N_2252);
nor U2392 (N_2392,N_2284,N_2287);
xnor U2393 (N_2393,N_2252,N_2203);
or U2394 (N_2394,N_2284,N_2295);
or U2395 (N_2395,N_2285,N_2288);
nand U2396 (N_2396,N_2205,N_2275);
nand U2397 (N_2397,N_2253,N_2266);
or U2398 (N_2398,N_2238,N_2227);
nor U2399 (N_2399,N_2215,N_2276);
or U2400 (N_2400,N_2303,N_2316);
nor U2401 (N_2401,N_2317,N_2311);
and U2402 (N_2402,N_2399,N_2359);
nand U2403 (N_2403,N_2319,N_2326);
nand U2404 (N_2404,N_2304,N_2349);
nor U2405 (N_2405,N_2324,N_2356);
nor U2406 (N_2406,N_2395,N_2367);
nand U2407 (N_2407,N_2363,N_2364);
and U2408 (N_2408,N_2348,N_2385);
and U2409 (N_2409,N_2362,N_2315);
or U2410 (N_2410,N_2333,N_2375);
nand U2411 (N_2411,N_2308,N_2355);
nor U2412 (N_2412,N_2378,N_2314);
nand U2413 (N_2413,N_2320,N_2387);
xor U2414 (N_2414,N_2340,N_2394);
or U2415 (N_2415,N_2325,N_2382);
nand U2416 (N_2416,N_2306,N_2390);
and U2417 (N_2417,N_2309,N_2376);
or U2418 (N_2418,N_2383,N_2336);
xor U2419 (N_2419,N_2300,N_2370);
xor U2420 (N_2420,N_2369,N_2353);
or U2421 (N_2421,N_2358,N_2374);
xnor U2422 (N_2422,N_2380,N_2313);
nor U2423 (N_2423,N_2328,N_2384);
or U2424 (N_2424,N_2346,N_2305);
xnor U2425 (N_2425,N_2379,N_2366);
and U2426 (N_2426,N_2357,N_2377);
nor U2427 (N_2427,N_2334,N_2307);
xor U2428 (N_2428,N_2396,N_2329);
nand U2429 (N_2429,N_2360,N_2388);
and U2430 (N_2430,N_2397,N_2332);
nand U2431 (N_2431,N_2302,N_2312);
and U2432 (N_2432,N_2343,N_2354);
xor U2433 (N_2433,N_2391,N_2361);
xor U2434 (N_2434,N_2368,N_2350);
and U2435 (N_2435,N_2338,N_2322);
and U2436 (N_2436,N_2301,N_2372);
xor U2437 (N_2437,N_2389,N_2347);
nand U2438 (N_2438,N_2310,N_2323);
nor U2439 (N_2439,N_2335,N_2365);
nand U2440 (N_2440,N_2321,N_2331);
nand U2441 (N_2441,N_2327,N_2393);
xor U2442 (N_2442,N_2381,N_2339);
and U2443 (N_2443,N_2386,N_2344);
and U2444 (N_2444,N_2351,N_2318);
nand U2445 (N_2445,N_2341,N_2330);
nand U2446 (N_2446,N_2373,N_2392);
xor U2447 (N_2447,N_2371,N_2342);
nor U2448 (N_2448,N_2352,N_2337);
nor U2449 (N_2449,N_2398,N_2345);
xor U2450 (N_2450,N_2340,N_2347);
and U2451 (N_2451,N_2384,N_2361);
nor U2452 (N_2452,N_2363,N_2339);
or U2453 (N_2453,N_2361,N_2377);
nor U2454 (N_2454,N_2375,N_2304);
nor U2455 (N_2455,N_2355,N_2318);
nor U2456 (N_2456,N_2341,N_2389);
nor U2457 (N_2457,N_2330,N_2316);
nand U2458 (N_2458,N_2325,N_2399);
and U2459 (N_2459,N_2387,N_2317);
xor U2460 (N_2460,N_2392,N_2344);
or U2461 (N_2461,N_2347,N_2305);
or U2462 (N_2462,N_2313,N_2364);
and U2463 (N_2463,N_2306,N_2332);
nor U2464 (N_2464,N_2330,N_2351);
and U2465 (N_2465,N_2336,N_2379);
nor U2466 (N_2466,N_2303,N_2341);
or U2467 (N_2467,N_2353,N_2343);
nor U2468 (N_2468,N_2314,N_2355);
xor U2469 (N_2469,N_2323,N_2338);
and U2470 (N_2470,N_2312,N_2316);
or U2471 (N_2471,N_2358,N_2327);
xor U2472 (N_2472,N_2385,N_2395);
nand U2473 (N_2473,N_2365,N_2340);
nand U2474 (N_2474,N_2381,N_2377);
nand U2475 (N_2475,N_2385,N_2397);
xnor U2476 (N_2476,N_2336,N_2376);
and U2477 (N_2477,N_2389,N_2301);
nand U2478 (N_2478,N_2398,N_2316);
and U2479 (N_2479,N_2310,N_2311);
and U2480 (N_2480,N_2323,N_2318);
or U2481 (N_2481,N_2394,N_2335);
nor U2482 (N_2482,N_2339,N_2326);
xnor U2483 (N_2483,N_2394,N_2306);
xnor U2484 (N_2484,N_2363,N_2377);
nand U2485 (N_2485,N_2335,N_2348);
or U2486 (N_2486,N_2320,N_2391);
or U2487 (N_2487,N_2394,N_2327);
or U2488 (N_2488,N_2367,N_2382);
xor U2489 (N_2489,N_2349,N_2335);
nor U2490 (N_2490,N_2336,N_2388);
nor U2491 (N_2491,N_2358,N_2369);
or U2492 (N_2492,N_2330,N_2361);
xor U2493 (N_2493,N_2393,N_2335);
xnor U2494 (N_2494,N_2354,N_2347);
and U2495 (N_2495,N_2300,N_2359);
and U2496 (N_2496,N_2393,N_2350);
and U2497 (N_2497,N_2356,N_2351);
or U2498 (N_2498,N_2309,N_2331);
and U2499 (N_2499,N_2386,N_2329);
nor U2500 (N_2500,N_2497,N_2476);
nor U2501 (N_2501,N_2436,N_2428);
nor U2502 (N_2502,N_2448,N_2408);
or U2503 (N_2503,N_2480,N_2432);
nand U2504 (N_2504,N_2493,N_2469);
xor U2505 (N_2505,N_2456,N_2470);
nand U2506 (N_2506,N_2417,N_2430);
or U2507 (N_2507,N_2423,N_2479);
nand U2508 (N_2508,N_2486,N_2429);
nor U2509 (N_2509,N_2473,N_2405);
nand U2510 (N_2510,N_2441,N_2488);
or U2511 (N_2511,N_2450,N_2466);
or U2512 (N_2512,N_2403,N_2478);
nand U2513 (N_2513,N_2459,N_2481);
nand U2514 (N_2514,N_2485,N_2421);
or U2515 (N_2515,N_2484,N_2435);
xor U2516 (N_2516,N_2451,N_2444);
xor U2517 (N_2517,N_2402,N_2406);
and U2518 (N_2518,N_2462,N_2461);
or U2519 (N_2519,N_2427,N_2491);
and U2520 (N_2520,N_2460,N_2415);
xnor U2521 (N_2521,N_2410,N_2433);
xor U2522 (N_2522,N_2453,N_2487);
or U2523 (N_2523,N_2496,N_2422);
nand U2524 (N_2524,N_2437,N_2426);
xor U2525 (N_2525,N_2463,N_2438);
and U2526 (N_2526,N_2455,N_2424);
xnor U2527 (N_2527,N_2449,N_2425);
and U2528 (N_2528,N_2477,N_2464);
and U2529 (N_2529,N_2401,N_2442);
nor U2530 (N_2530,N_2409,N_2471);
nor U2531 (N_2531,N_2467,N_2414);
nor U2532 (N_2532,N_2468,N_2418);
xor U2533 (N_2533,N_2407,N_2431);
nor U2534 (N_2534,N_2475,N_2452);
nand U2535 (N_2535,N_2416,N_2434);
or U2536 (N_2536,N_2400,N_2412);
nor U2537 (N_2537,N_2419,N_2465);
and U2538 (N_2538,N_2420,N_2482);
nand U2539 (N_2539,N_2495,N_2413);
or U2540 (N_2540,N_2490,N_2454);
or U2541 (N_2541,N_2439,N_2447);
xnor U2542 (N_2542,N_2494,N_2472);
and U2543 (N_2543,N_2440,N_2411);
nor U2544 (N_2544,N_2457,N_2498);
and U2545 (N_2545,N_2443,N_2499);
nor U2546 (N_2546,N_2445,N_2446);
xnor U2547 (N_2547,N_2489,N_2474);
or U2548 (N_2548,N_2483,N_2492);
nand U2549 (N_2549,N_2404,N_2458);
nand U2550 (N_2550,N_2415,N_2463);
nand U2551 (N_2551,N_2473,N_2486);
nor U2552 (N_2552,N_2467,N_2422);
xor U2553 (N_2553,N_2488,N_2470);
nand U2554 (N_2554,N_2469,N_2448);
xor U2555 (N_2555,N_2466,N_2417);
and U2556 (N_2556,N_2460,N_2414);
nand U2557 (N_2557,N_2449,N_2409);
and U2558 (N_2558,N_2476,N_2491);
nand U2559 (N_2559,N_2487,N_2431);
xor U2560 (N_2560,N_2483,N_2414);
or U2561 (N_2561,N_2452,N_2457);
nand U2562 (N_2562,N_2408,N_2471);
nor U2563 (N_2563,N_2454,N_2496);
nand U2564 (N_2564,N_2474,N_2420);
and U2565 (N_2565,N_2449,N_2461);
xnor U2566 (N_2566,N_2425,N_2415);
or U2567 (N_2567,N_2482,N_2433);
nand U2568 (N_2568,N_2498,N_2424);
xor U2569 (N_2569,N_2423,N_2425);
and U2570 (N_2570,N_2438,N_2443);
and U2571 (N_2571,N_2415,N_2420);
or U2572 (N_2572,N_2483,N_2437);
nor U2573 (N_2573,N_2440,N_2417);
or U2574 (N_2574,N_2487,N_2457);
nand U2575 (N_2575,N_2402,N_2412);
and U2576 (N_2576,N_2424,N_2431);
nor U2577 (N_2577,N_2473,N_2409);
nor U2578 (N_2578,N_2431,N_2446);
or U2579 (N_2579,N_2488,N_2497);
nand U2580 (N_2580,N_2471,N_2460);
xnor U2581 (N_2581,N_2479,N_2436);
and U2582 (N_2582,N_2447,N_2493);
or U2583 (N_2583,N_2490,N_2402);
nor U2584 (N_2584,N_2487,N_2436);
nor U2585 (N_2585,N_2488,N_2468);
nor U2586 (N_2586,N_2492,N_2432);
and U2587 (N_2587,N_2466,N_2491);
nor U2588 (N_2588,N_2462,N_2466);
nand U2589 (N_2589,N_2444,N_2477);
and U2590 (N_2590,N_2401,N_2494);
and U2591 (N_2591,N_2456,N_2497);
or U2592 (N_2592,N_2487,N_2401);
and U2593 (N_2593,N_2417,N_2426);
and U2594 (N_2594,N_2418,N_2451);
nand U2595 (N_2595,N_2434,N_2473);
nor U2596 (N_2596,N_2431,N_2436);
nand U2597 (N_2597,N_2420,N_2410);
xnor U2598 (N_2598,N_2404,N_2452);
xnor U2599 (N_2599,N_2460,N_2450);
xnor U2600 (N_2600,N_2592,N_2524);
nand U2601 (N_2601,N_2593,N_2576);
or U2602 (N_2602,N_2581,N_2507);
nand U2603 (N_2603,N_2565,N_2521);
nand U2604 (N_2604,N_2505,N_2549);
nor U2605 (N_2605,N_2587,N_2558);
nor U2606 (N_2606,N_2582,N_2503);
nor U2607 (N_2607,N_2546,N_2577);
and U2608 (N_2608,N_2514,N_2595);
or U2609 (N_2609,N_2541,N_2537);
nand U2610 (N_2610,N_2562,N_2566);
xor U2611 (N_2611,N_2536,N_2580);
nor U2612 (N_2612,N_2552,N_2515);
and U2613 (N_2613,N_2548,N_2538);
or U2614 (N_2614,N_2500,N_2554);
or U2615 (N_2615,N_2573,N_2520);
nand U2616 (N_2616,N_2534,N_2584);
or U2617 (N_2617,N_2528,N_2532);
nand U2618 (N_2618,N_2510,N_2544);
and U2619 (N_2619,N_2530,N_2559);
nor U2620 (N_2620,N_2570,N_2572);
nor U2621 (N_2621,N_2523,N_2535);
or U2622 (N_2622,N_2589,N_2588);
nor U2623 (N_2623,N_2560,N_2512);
or U2624 (N_2624,N_2501,N_2556);
xnor U2625 (N_2625,N_2553,N_2519);
nand U2626 (N_2626,N_2502,N_2578);
and U2627 (N_2627,N_2563,N_2511);
xor U2628 (N_2628,N_2555,N_2575);
or U2629 (N_2629,N_2547,N_2586);
or U2630 (N_2630,N_2567,N_2590);
nor U2631 (N_2631,N_2508,N_2518);
xnor U2632 (N_2632,N_2591,N_2571);
nand U2633 (N_2633,N_2533,N_2545);
xnor U2634 (N_2634,N_2540,N_2583);
xor U2635 (N_2635,N_2513,N_2594);
nor U2636 (N_2636,N_2531,N_2585);
nor U2637 (N_2637,N_2568,N_2557);
and U2638 (N_2638,N_2551,N_2509);
nor U2639 (N_2639,N_2569,N_2516);
xnor U2640 (N_2640,N_2529,N_2539);
and U2641 (N_2641,N_2527,N_2522);
and U2642 (N_2642,N_2564,N_2599);
or U2643 (N_2643,N_2525,N_2579);
nor U2644 (N_2644,N_2596,N_2574);
and U2645 (N_2645,N_2542,N_2504);
or U2646 (N_2646,N_2543,N_2526);
and U2647 (N_2647,N_2561,N_2597);
or U2648 (N_2648,N_2506,N_2598);
and U2649 (N_2649,N_2517,N_2550);
nand U2650 (N_2650,N_2531,N_2574);
nand U2651 (N_2651,N_2535,N_2532);
xnor U2652 (N_2652,N_2590,N_2578);
and U2653 (N_2653,N_2591,N_2512);
nor U2654 (N_2654,N_2540,N_2596);
or U2655 (N_2655,N_2526,N_2589);
xnor U2656 (N_2656,N_2578,N_2540);
nor U2657 (N_2657,N_2543,N_2594);
xor U2658 (N_2658,N_2518,N_2572);
xnor U2659 (N_2659,N_2596,N_2519);
nand U2660 (N_2660,N_2512,N_2550);
nand U2661 (N_2661,N_2555,N_2573);
nor U2662 (N_2662,N_2521,N_2503);
nor U2663 (N_2663,N_2582,N_2595);
or U2664 (N_2664,N_2541,N_2584);
nand U2665 (N_2665,N_2558,N_2532);
nor U2666 (N_2666,N_2563,N_2576);
nand U2667 (N_2667,N_2583,N_2516);
xor U2668 (N_2668,N_2585,N_2569);
and U2669 (N_2669,N_2507,N_2516);
or U2670 (N_2670,N_2509,N_2521);
nor U2671 (N_2671,N_2514,N_2520);
and U2672 (N_2672,N_2595,N_2568);
nor U2673 (N_2673,N_2580,N_2543);
xnor U2674 (N_2674,N_2575,N_2556);
and U2675 (N_2675,N_2507,N_2575);
nor U2676 (N_2676,N_2575,N_2598);
nand U2677 (N_2677,N_2591,N_2502);
nand U2678 (N_2678,N_2540,N_2556);
or U2679 (N_2679,N_2565,N_2577);
nor U2680 (N_2680,N_2570,N_2500);
or U2681 (N_2681,N_2511,N_2539);
or U2682 (N_2682,N_2544,N_2526);
xor U2683 (N_2683,N_2570,N_2516);
nand U2684 (N_2684,N_2514,N_2534);
xor U2685 (N_2685,N_2579,N_2589);
and U2686 (N_2686,N_2524,N_2534);
and U2687 (N_2687,N_2573,N_2540);
nand U2688 (N_2688,N_2550,N_2547);
and U2689 (N_2689,N_2503,N_2504);
or U2690 (N_2690,N_2561,N_2578);
nand U2691 (N_2691,N_2508,N_2580);
nor U2692 (N_2692,N_2593,N_2517);
or U2693 (N_2693,N_2554,N_2510);
xnor U2694 (N_2694,N_2571,N_2537);
nand U2695 (N_2695,N_2513,N_2567);
xnor U2696 (N_2696,N_2597,N_2558);
xor U2697 (N_2697,N_2579,N_2576);
nor U2698 (N_2698,N_2598,N_2511);
nor U2699 (N_2699,N_2571,N_2584);
nor U2700 (N_2700,N_2696,N_2620);
nor U2701 (N_2701,N_2687,N_2630);
nor U2702 (N_2702,N_2665,N_2609);
nor U2703 (N_2703,N_2675,N_2610);
or U2704 (N_2704,N_2672,N_2690);
nor U2705 (N_2705,N_2680,N_2639);
or U2706 (N_2706,N_2691,N_2684);
nor U2707 (N_2707,N_2683,N_2602);
nand U2708 (N_2708,N_2657,N_2625);
and U2709 (N_2709,N_2640,N_2699);
xnor U2710 (N_2710,N_2634,N_2613);
xor U2711 (N_2711,N_2662,N_2621);
or U2712 (N_2712,N_2693,N_2611);
or U2713 (N_2713,N_2681,N_2661);
or U2714 (N_2714,N_2612,N_2695);
or U2715 (N_2715,N_2679,N_2607);
xnor U2716 (N_2716,N_2604,N_2647);
or U2717 (N_2717,N_2646,N_2605);
nand U2718 (N_2718,N_2641,N_2631);
nand U2719 (N_2719,N_2678,N_2669);
xor U2720 (N_2720,N_2660,N_2624);
and U2721 (N_2721,N_2663,N_2682);
or U2722 (N_2722,N_2653,N_2619);
and U2723 (N_2723,N_2673,N_2664);
and U2724 (N_2724,N_2688,N_2622);
nand U2725 (N_2725,N_2697,N_2668);
xor U2726 (N_2726,N_2685,N_2676);
nand U2727 (N_2727,N_2626,N_2648);
or U2728 (N_2728,N_2603,N_2628);
and U2729 (N_2729,N_2632,N_2698);
nand U2730 (N_2730,N_2650,N_2615);
xor U2731 (N_2731,N_2627,N_2674);
and U2732 (N_2732,N_2671,N_2633);
or U2733 (N_2733,N_2642,N_2677);
or U2734 (N_2734,N_2670,N_2643);
nand U2735 (N_2735,N_2654,N_2659);
xor U2736 (N_2736,N_2608,N_2645);
nor U2737 (N_2737,N_2689,N_2651);
nand U2738 (N_2738,N_2617,N_2649);
and U2739 (N_2739,N_2616,N_2666);
and U2740 (N_2740,N_2629,N_2655);
xnor U2741 (N_2741,N_2637,N_2652);
nor U2742 (N_2742,N_2623,N_2638);
and U2743 (N_2743,N_2694,N_2635);
and U2744 (N_2744,N_2658,N_2636);
or U2745 (N_2745,N_2667,N_2614);
nand U2746 (N_2746,N_2692,N_2686);
or U2747 (N_2747,N_2618,N_2600);
xor U2748 (N_2748,N_2656,N_2644);
and U2749 (N_2749,N_2601,N_2606);
nor U2750 (N_2750,N_2661,N_2692);
nand U2751 (N_2751,N_2695,N_2601);
nor U2752 (N_2752,N_2669,N_2654);
xor U2753 (N_2753,N_2663,N_2609);
or U2754 (N_2754,N_2667,N_2686);
or U2755 (N_2755,N_2624,N_2697);
and U2756 (N_2756,N_2698,N_2679);
and U2757 (N_2757,N_2622,N_2653);
and U2758 (N_2758,N_2631,N_2608);
nand U2759 (N_2759,N_2657,N_2674);
or U2760 (N_2760,N_2655,N_2650);
nor U2761 (N_2761,N_2642,N_2644);
nand U2762 (N_2762,N_2662,N_2698);
nor U2763 (N_2763,N_2630,N_2648);
and U2764 (N_2764,N_2628,N_2694);
nand U2765 (N_2765,N_2660,N_2646);
nand U2766 (N_2766,N_2616,N_2675);
nand U2767 (N_2767,N_2671,N_2658);
nand U2768 (N_2768,N_2682,N_2649);
and U2769 (N_2769,N_2668,N_2629);
xor U2770 (N_2770,N_2667,N_2629);
nand U2771 (N_2771,N_2636,N_2650);
xnor U2772 (N_2772,N_2606,N_2662);
nand U2773 (N_2773,N_2637,N_2612);
and U2774 (N_2774,N_2619,N_2611);
nor U2775 (N_2775,N_2677,N_2641);
nor U2776 (N_2776,N_2632,N_2670);
nand U2777 (N_2777,N_2667,N_2605);
xnor U2778 (N_2778,N_2616,N_2645);
xor U2779 (N_2779,N_2642,N_2626);
or U2780 (N_2780,N_2678,N_2646);
nand U2781 (N_2781,N_2600,N_2647);
and U2782 (N_2782,N_2643,N_2623);
xnor U2783 (N_2783,N_2616,N_2613);
nand U2784 (N_2784,N_2648,N_2652);
nand U2785 (N_2785,N_2621,N_2687);
nor U2786 (N_2786,N_2660,N_2652);
nor U2787 (N_2787,N_2624,N_2673);
nor U2788 (N_2788,N_2690,N_2669);
and U2789 (N_2789,N_2645,N_2614);
and U2790 (N_2790,N_2658,N_2675);
nand U2791 (N_2791,N_2694,N_2632);
xor U2792 (N_2792,N_2622,N_2659);
or U2793 (N_2793,N_2650,N_2691);
nand U2794 (N_2794,N_2617,N_2686);
nor U2795 (N_2795,N_2682,N_2684);
nand U2796 (N_2796,N_2681,N_2696);
xor U2797 (N_2797,N_2619,N_2648);
and U2798 (N_2798,N_2636,N_2620);
nor U2799 (N_2799,N_2668,N_2605);
xnor U2800 (N_2800,N_2787,N_2711);
xnor U2801 (N_2801,N_2783,N_2747);
and U2802 (N_2802,N_2788,N_2793);
xnor U2803 (N_2803,N_2738,N_2704);
nand U2804 (N_2804,N_2717,N_2708);
nand U2805 (N_2805,N_2745,N_2731);
or U2806 (N_2806,N_2718,N_2706);
xor U2807 (N_2807,N_2746,N_2784);
nor U2808 (N_2808,N_2781,N_2749);
nor U2809 (N_2809,N_2796,N_2712);
xor U2810 (N_2810,N_2730,N_2715);
nand U2811 (N_2811,N_2792,N_2786);
nor U2812 (N_2812,N_2765,N_2739);
nand U2813 (N_2813,N_2703,N_2709);
nor U2814 (N_2814,N_2754,N_2727);
nor U2815 (N_2815,N_2737,N_2756);
nand U2816 (N_2816,N_2764,N_2753);
nand U2817 (N_2817,N_2759,N_2728);
and U2818 (N_2818,N_2725,N_2757);
nand U2819 (N_2819,N_2760,N_2732);
nor U2820 (N_2820,N_2751,N_2799);
and U2821 (N_2821,N_2752,N_2729);
nor U2822 (N_2822,N_2733,N_2726);
nand U2823 (N_2823,N_2789,N_2798);
xor U2824 (N_2824,N_2742,N_2797);
xor U2825 (N_2825,N_2776,N_2775);
nor U2826 (N_2826,N_2770,N_2741);
or U2827 (N_2827,N_2701,N_2707);
or U2828 (N_2828,N_2769,N_2710);
nand U2829 (N_2829,N_2755,N_2705);
or U2830 (N_2830,N_2763,N_2748);
xor U2831 (N_2831,N_2734,N_2721);
nand U2832 (N_2832,N_2702,N_2744);
nor U2833 (N_2833,N_2719,N_2716);
xnor U2834 (N_2834,N_2723,N_2791);
nand U2835 (N_2835,N_2785,N_2735);
xor U2836 (N_2836,N_2743,N_2782);
xnor U2837 (N_2837,N_2774,N_2761);
and U2838 (N_2838,N_2700,N_2795);
nor U2839 (N_2839,N_2766,N_2780);
xor U2840 (N_2840,N_2779,N_2714);
and U2841 (N_2841,N_2713,N_2772);
xor U2842 (N_2842,N_2750,N_2778);
nand U2843 (N_2843,N_2740,N_2758);
or U2844 (N_2844,N_2722,N_2768);
nor U2845 (N_2845,N_2794,N_2790);
nand U2846 (N_2846,N_2767,N_2720);
nor U2847 (N_2847,N_2777,N_2771);
and U2848 (N_2848,N_2724,N_2762);
or U2849 (N_2849,N_2773,N_2736);
nor U2850 (N_2850,N_2714,N_2738);
and U2851 (N_2851,N_2765,N_2763);
and U2852 (N_2852,N_2754,N_2794);
nand U2853 (N_2853,N_2731,N_2720);
and U2854 (N_2854,N_2774,N_2775);
nor U2855 (N_2855,N_2709,N_2726);
xor U2856 (N_2856,N_2715,N_2794);
nor U2857 (N_2857,N_2714,N_2763);
nand U2858 (N_2858,N_2772,N_2715);
nand U2859 (N_2859,N_2701,N_2740);
or U2860 (N_2860,N_2709,N_2797);
and U2861 (N_2861,N_2772,N_2766);
or U2862 (N_2862,N_2752,N_2713);
and U2863 (N_2863,N_2755,N_2710);
and U2864 (N_2864,N_2701,N_2749);
or U2865 (N_2865,N_2700,N_2703);
nand U2866 (N_2866,N_2726,N_2738);
nor U2867 (N_2867,N_2772,N_2711);
nor U2868 (N_2868,N_2769,N_2717);
nor U2869 (N_2869,N_2733,N_2727);
and U2870 (N_2870,N_2719,N_2751);
or U2871 (N_2871,N_2726,N_2740);
or U2872 (N_2872,N_2742,N_2769);
nand U2873 (N_2873,N_2777,N_2752);
or U2874 (N_2874,N_2753,N_2745);
nand U2875 (N_2875,N_2777,N_2784);
nand U2876 (N_2876,N_2704,N_2726);
xnor U2877 (N_2877,N_2796,N_2771);
nand U2878 (N_2878,N_2746,N_2783);
nor U2879 (N_2879,N_2757,N_2748);
nor U2880 (N_2880,N_2727,N_2710);
nand U2881 (N_2881,N_2715,N_2763);
and U2882 (N_2882,N_2787,N_2768);
nor U2883 (N_2883,N_2756,N_2761);
nand U2884 (N_2884,N_2795,N_2775);
or U2885 (N_2885,N_2761,N_2702);
nor U2886 (N_2886,N_2793,N_2717);
and U2887 (N_2887,N_2783,N_2708);
or U2888 (N_2888,N_2740,N_2735);
nor U2889 (N_2889,N_2758,N_2784);
xnor U2890 (N_2890,N_2774,N_2781);
and U2891 (N_2891,N_2785,N_2752);
xnor U2892 (N_2892,N_2766,N_2769);
or U2893 (N_2893,N_2771,N_2762);
nor U2894 (N_2894,N_2729,N_2750);
nand U2895 (N_2895,N_2778,N_2722);
xor U2896 (N_2896,N_2735,N_2750);
xnor U2897 (N_2897,N_2731,N_2789);
xor U2898 (N_2898,N_2797,N_2773);
xnor U2899 (N_2899,N_2737,N_2708);
nor U2900 (N_2900,N_2803,N_2889);
and U2901 (N_2901,N_2860,N_2899);
or U2902 (N_2902,N_2830,N_2804);
xnor U2903 (N_2903,N_2845,N_2813);
or U2904 (N_2904,N_2868,N_2844);
nor U2905 (N_2905,N_2896,N_2802);
nor U2906 (N_2906,N_2823,N_2861);
and U2907 (N_2907,N_2837,N_2892);
or U2908 (N_2908,N_2834,N_2819);
nor U2909 (N_2909,N_2820,N_2859);
nand U2910 (N_2910,N_2851,N_2824);
xor U2911 (N_2911,N_2875,N_2843);
and U2912 (N_2912,N_2831,N_2895);
nand U2913 (N_2913,N_2815,N_2878);
nand U2914 (N_2914,N_2810,N_2857);
or U2915 (N_2915,N_2849,N_2808);
nand U2916 (N_2916,N_2876,N_2882);
xor U2917 (N_2917,N_2829,N_2847);
or U2918 (N_2918,N_2855,N_2806);
or U2919 (N_2919,N_2872,N_2801);
nor U2920 (N_2920,N_2826,N_2856);
or U2921 (N_2921,N_2852,N_2864);
or U2922 (N_2922,N_2898,N_2807);
or U2923 (N_2923,N_2805,N_2866);
and U2924 (N_2924,N_2888,N_2893);
nand U2925 (N_2925,N_2825,N_2867);
xor U2926 (N_2926,N_2809,N_2842);
or U2927 (N_2927,N_2880,N_2816);
nand U2928 (N_2928,N_2877,N_2817);
nand U2929 (N_2929,N_2848,N_2894);
or U2930 (N_2930,N_2832,N_2836);
and U2931 (N_2931,N_2897,N_2858);
or U2932 (N_2932,N_2874,N_2891);
and U2933 (N_2933,N_2873,N_2800);
or U2934 (N_2934,N_2863,N_2818);
or U2935 (N_2935,N_2883,N_2884);
nor U2936 (N_2936,N_2835,N_2812);
and U2937 (N_2937,N_2887,N_2881);
and U2938 (N_2938,N_2885,N_2886);
or U2939 (N_2939,N_2854,N_2828);
nor U2940 (N_2940,N_2865,N_2870);
nor U2941 (N_2941,N_2833,N_2871);
and U2942 (N_2942,N_2821,N_2838);
nor U2943 (N_2943,N_2850,N_2890);
nor U2944 (N_2944,N_2822,N_2853);
or U2945 (N_2945,N_2814,N_2811);
xor U2946 (N_2946,N_2879,N_2846);
and U2947 (N_2947,N_2827,N_2862);
or U2948 (N_2948,N_2841,N_2869);
nor U2949 (N_2949,N_2840,N_2839);
and U2950 (N_2950,N_2818,N_2837);
and U2951 (N_2951,N_2858,N_2862);
xnor U2952 (N_2952,N_2871,N_2837);
xnor U2953 (N_2953,N_2862,N_2841);
or U2954 (N_2954,N_2812,N_2822);
xnor U2955 (N_2955,N_2856,N_2802);
and U2956 (N_2956,N_2816,N_2877);
and U2957 (N_2957,N_2809,N_2879);
xnor U2958 (N_2958,N_2842,N_2851);
nor U2959 (N_2959,N_2835,N_2876);
and U2960 (N_2960,N_2828,N_2873);
and U2961 (N_2961,N_2814,N_2883);
nand U2962 (N_2962,N_2839,N_2844);
xor U2963 (N_2963,N_2815,N_2859);
and U2964 (N_2964,N_2806,N_2824);
nand U2965 (N_2965,N_2806,N_2841);
xnor U2966 (N_2966,N_2852,N_2875);
xnor U2967 (N_2967,N_2821,N_2886);
and U2968 (N_2968,N_2811,N_2815);
xnor U2969 (N_2969,N_2804,N_2832);
and U2970 (N_2970,N_2831,N_2878);
xnor U2971 (N_2971,N_2850,N_2894);
nand U2972 (N_2972,N_2841,N_2890);
or U2973 (N_2973,N_2861,N_2867);
nand U2974 (N_2974,N_2812,N_2825);
nand U2975 (N_2975,N_2864,N_2821);
or U2976 (N_2976,N_2833,N_2838);
nand U2977 (N_2977,N_2839,N_2858);
and U2978 (N_2978,N_2882,N_2855);
nor U2979 (N_2979,N_2820,N_2846);
xor U2980 (N_2980,N_2832,N_2801);
nand U2981 (N_2981,N_2856,N_2888);
nand U2982 (N_2982,N_2854,N_2891);
xnor U2983 (N_2983,N_2825,N_2882);
nand U2984 (N_2984,N_2800,N_2874);
xor U2985 (N_2985,N_2880,N_2821);
and U2986 (N_2986,N_2823,N_2894);
nor U2987 (N_2987,N_2847,N_2851);
xnor U2988 (N_2988,N_2800,N_2876);
nor U2989 (N_2989,N_2898,N_2851);
or U2990 (N_2990,N_2878,N_2863);
nand U2991 (N_2991,N_2807,N_2810);
nand U2992 (N_2992,N_2883,N_2813);
xnor U2993 (N_2993,N_2887,N_2825);
nor U2994 (N_2994,N_2867,N_2801);
xor U2995 (N_2995,N_2858,N_2826);
xor U2996 (N_2996,N_2846,N_2832);
nor U2997 (N_2997,N_2873,N_2822);
and U2998 (N_2998,N_2895,N_2845);
or U2999 (N_2999,N_2828,N_2821);
xor U3000 (N_3000,N_2988,N_2934);
and U3001 (N_3001,N_2936,N_2907);
xnor U3002 (N_3002,N_2954,N_2921);
and U3003 (N_3003,N_2906,N_2933);
xnor U3004 (N_3004,N_2904,N_2952);
xor U3005 (N_3005,N_2966,N_2944);
xnor U3006 (N_3006,N_2985,N_2983);
or U3007 (N_3007,N_2975,N_2957);
or U3008 (N_3008,N_2901,N_2996);
or U3009 (N_3009,N_2964,N_2908);
nand U3010 (N_3010,N_2949,N_2915);
nand U3011 (N_3011,N_2972,N_2984);
xnor U3012 (N_3012,N_2974,N_2951);
nand U3013 (N_3013,N_2962,N_2958);
nor U3014 (N_3014,N_2919,N_2910);
nor U3015 (N_3015,N_2947,N_2955);
xor U3016 (N_3016,N_2913,N_2994);
nand U3017 (N_3017,N_2997,N_2969);
and U3018 (N_3018,N_2909,N_2940);
xor U3019 (N_3019,N_2967,N_2905);
xor U3020 (N_3020,N_2953,N_2978);
nor U3021 (N_3021,N_2939,N_2937);
nor U3022 (N_3022,N_2981,N_2923);
or U3023 (N_3023,N_2943,N_2941);
xor U3024 (N_3024,N_2920,N_2938);
and U3025 (N_3025,N_2965,N_2989);
xor U3026 (N_3026,N_2970,N_2995);
and U3027 (N_3027,N_2950,N_2917);
xnor U3028 (N_3028,N_2986,N_2956);
or U3029 (N_3029,N_2977,N_2992);
nand U3030 (N_3030,N_2900,N_2929);
or U3031 (N_3031,N_2980,N_2948);
nor U3032 (N_3032,N_2946,N_2926);
nor U3033 (N_3033,N_2932,N_2911);
xor U3034 (N_3034,N_2902,N_2903);
xor U3035 (N_3035,N_2918,N_2942);
xnor U3036 (N_3036,N_2961,N_2930);
or U3037 (N_3037,N_2914,N_2924);
or U3038 (N_3038,N_2999,N_2931);
and U3039 (N_3039,N_2976,N_2945);
nand U3040 (N_3040,N_2987,N_2963);
nand U3041 (N_3041,N_2927,N_2928);
or U3042 (N_3042,N_2991,N_2968);
and U3043 (N_3043,N_2990,N_2973);
nor U3044 (N_3044,N_2935,N_2922);
or U3045 (N_3045,N_2959,N_2993);
xnor U3046 (N_3046,N_2971,N_2916);
and U3047 (N_3047,N_2979,N_2912);
or U3048 (N_3048,N_2960,N_2982);
xnor U3049 (N_3049,N_2998,N_2925);
or U3050 (N_3050,N_2968,N_2969);
or U3051 (N_3051,N_2950,N_2990);
nor U3052 (N_3052,N_2927,N_2994);
xnor U3053 (N_3053,N_2927,N_2924);
and U3054 (N_3054,N_2985,N_2911);
xor U3055 (N_3055,N_2988,N_2938);
nor U3056 (N_3056,N_2900,N_2969);
nand U3057 (N_3057,N_2998,N_2920);
xnor U3058 (N_3058,N_2917,N_2911);
or U3059 (N_3059,N_2942,N_2957);
and U3060 (N_3060,N_2923,N_2958);
or U3061 (N_3061,N_2951,N_2964);
xor U3062 (N_3062,N_2964,N_2984);
nand U3063 (N_3063,N_2972,N_2937);
or U3064 (N_3064,N_2936,N_2925);
or U3065 (N_3065,N_2956,N_2921);
nor U3066 (N_3066,N_2962,N_2941);
and U3067 (N_3067,N_2910,N_2927);
nand U3068 (N_3068,N_2936,N_2973);
nand U3069 (N_3069,N_2961,N_2931);
nor U3070 (N_3070,N_2993,N_2943);
or U3071 (N_3071,N_2989,N_2947);
and U3072 (N_3072,N_2915,N_2918);
nand U3073 (N_3073,N_2948,N_2983);
and U3074 (N_3074,N_2956,N_2954);
xor U3075 (N_3075,N_2931,N_2980);
and U3076 (N_3076,N_2943,N_2972);
nand U3077 (N_3077,N_2918,N_2986);
xor U3078 (N_3078,N_2951,N_2907);
nand U3079 (N_3079,N_2922,N_2901);
and U3080 (N_3080,N_2944,N_2976);
nor U3081 (N_3081,N_2948,N_2929);
nor U3082 (N_3082,N_2983,N_2902);
nand U3083 (N_3083,N_2956,N_2969);
nand U3084 (N_3084,N_2908,N_2939);
xnor U3085 (N_3085,N_2949,N_2966);
nor U3086 (N_3086,N_2928,N_2963);
nor U3087 (N_3087,N_2930,N_2916);
xor U3088 (N_3088,N_2998,N_2911);
and U3089 (N_3089,N_2931,N_2969);
xnor U3090 (N_3090,N_2908,N_2998);
or U3091 (N_3091,N_2952,N_2995);
and U3092 (N_3092,N_2938,N_2916);
or U3093 (N_3093,N_2989,N_2986);
or U3094 (N_3094,N_2939,N_2999);
xor U3095 (N_3095,N_2937,N_2960);
or U3096 (N_3096,N_2935,N_2909);
and U3097 (N_3097,N_2923,N_2985);
xnor U3098 (N_3098,N_2941,N_2985);
nor U3099 (N_3099,N_2920,N_2949);
and U3100 (N_3100,N_3090,N_3019);
nor U3101 (N_3101,N_3055,N_3096);
and U3102 (N_3102,N_3094,N_3056);
and U3103 (N_3103,N_3065,N_3004);
and U3104 (N_3104,N_3032,N_3041);
nand U3105 (N_3105,N_3040,N_3000);
or U3106 (N_3106,N_3050,N_3011);
and U3107 (N_3107,N_3010,N_3084);
or U3108 (N_3108,N_3060,N_3097);
nor U3109 (N_3109,N_3043,N_3051);
xnor U3110 (N_3110,N_3037,N_3088);
and U3111 (N_3111,N_3068,N_3008);
and U3112 (N_3112,N_3069,N_3009);
xnor U3113 (N_3113,N_3017,N_3045);
or U3114 (N_3114,N_3007,N_3074);
and U3115 (N_3115,N_3039,N_3076);
xor U3116 (N_3116,N_3033,N_3062);
or U3117 (N_3117,N_3072,N_3075);
xnor U3118 (N_3118,N_3083,N_3058);
and U3119 (N_3119,N_3052,N_3093);
or U3120 (N_3120,N_3024,N_3036);
xor U3121 (N_3121,N_3070,N_3034);
xor U3122 (N_3122,N_3042,N_3013);
nor U3123 (N_3123,N_3029,N_3054);
nor U3124 (N_3124,N_3005,N_3073);
nor U3125 (N_3125,N_3016,N_3026);
nor U3126 (N_3126,N_3092,N_3089);
xor U3127 (N_3127,N_3081,N_3085);
nor U3128 (N_3128,N_3001,N_3048);
xnor U3129 (N_3129,N_3099,N_3079);
and U3130 (N_3130,N_3022,N_3014);
and U3131 (N_3131,N_3057,N_3095);
nand U3132 (N_3132,N_3071,N_3086);
and U3133 (N_3133,N_3063,N_3020);
nand U3134 (N_3134,N_3047,N_3059);
or U3135 (N_3135,N_3023,N_3035);
nand U3136 (N_3136,N_3098,N_3067);
nand U3137 (N_3137,N_3002,N_3038);
xor U3138 (N_3138,N_3087,N_3049);
or U3139 (N_3139,N_3015,N_3012);
and U3140 (N_3140,N_3077,N_3025);
nor U3141 (N_3141,N_3053,N_3061);
or U3142 (N_3142,N_3018,N_3066);
or U3143 (N_3143,N_3030,N_3082);
nor U3144 (N_3144,N_3028,N_3064);
and U3145 (N_3145,N_3006,N_3078);
xnor U3146 (N_3146,N_3044,N_3046);
nor U3147 (N_3147,N_3091,N_3080);
and U3148 (N_3148,N_3021,N_3003);
nor U3149 (N_3149,N_3027,N_3031);
nor U3150 (N_3150,N_3027,N_3003);
nor U3151 (N_3151,N_3070,N_3030);
and U3152 (N_3152,N_3060,N_3073);
or U3153 (N_3153,N_3005,N_3081);
and U3154 (N_3154,N_3003,N_3009);
or U3155 (N_3155,N_3069,N_3016);
nor U3156 (N_3156,N_3059,N_3030);
and U3157 (N_3157,N_3016,N_3063);
or U3158 (N_3158,N_3024,N_3099);
xor U3159 (N_3159,N_3023,N_3053);
or U3160 (N_3160,N_3093,N_3022);
and U3161 (N_3161,N_3084,N_3012);
nor U3162 (N_3162,N_3038,N_3013);
nand U3163 (N_3163,N_3067,N_3043);
or U3164 (N_3164,N_3046,N_3099);
and U3165 (N_3165,N_3030,N_3084);
and U3166 (N_3166,N_3056,N_3012);
and U3167 (N_3167,N_3085,N_3089);
and U3168 (N_3168,N_3087,N_3051);
xnor U3169 (N_3169,N_3056,N_3039);
and U3170 (N_3170,N_3040,N_3080);
nor U3171 (N_3171,N_3064,N_3075);
nor U3172 (N_3172,N_3048,N_3034);
nor U3173 (N_3173,N_3071,N_3036);
xor U3174 (N_3174,N_3053,N_3088);
xor U3175 (N_3175,N_3063,N_3055);
or U3176 (N_3176,N_3002,N_3089);
and U3177 (N_3177,N_3059,N_3055);
nand U3178 (N_3178,N_3071,N_3025);
or U3179 (N_3179,N_3020,N_3027);
and U3180 (N_3180,N_3059,N_3021);
xor U3181 (N_3181,N_3062,N_3037);
nor U3182 (N_3182,N_3028,N_3072);
nor U3183 (N_3183,N_3085,N_3046);
nor U3184 (N_3184,N_3055,N_3086);
and U3185 (N_3185,N_3030,N_3093);
or U3186 (N_3186,N_3078,N_3087);
nand U3187 (N_3187,N_3020,N_3058);
nand U3188 (N_3188,N_3028,N_3029);
or U3189 (N_3189,N_3045,N_3088);
xor U3190 (N_3190,N_3073,N_3047);
xnor U3191 (N_3191,N_3074,N_3059);
xnor U3192 (N_3192,N_3022,N_3054);
or U3193 (N_3193,N_3061,N_3076);
and U3194 (N_3194,N_3090,N_3078);
nand U3195 (N_3195,N_3034,N_3038);
or U3196 (N_3196,N_3054,N_3096);
or U3197 (N_3197,N_3004,N_3074);
or U3198 (N_3198,N_3012,N_3076);
or U3199 (N_3199,N_3001,N_3068);
nor U3200 (N_3200,N_3106,N_3167);
nand U3201 (N_3201,N_3145,N_3159);
xor U3202 (N_3202,N_3165,N_3119);
and U3203 (N_3203,N_3132,N_3120);
and U3204 (N_3204,N_3155,N_3125);
nor U3205 (N_3205,N_3104,N_3148);
xnor U3206 (N_3206,N_3156,N_3107);
and U3207 (N_3207,N_3142,N_3112);
nand U3208 (N_3208,N_3193,N_3110);
nor U3209 (N_3209,N_3188,N_3138);
or U3210 (N_3210,N_3134,N_3151);
and U3211 (N_3211,N_3121,N_3131);
xor U3212 (N_3212,N_3164,N_3111);
xnor U3213 (N_3213,N_3105,N_3103);
or U3214 (N_3214,N_3170,N_3190);
and U3215 (N_3215,N_3181,N_3189);
or U3216 (N_3216,N_3137,N_3197);
xor U3217 (N_3217,N_3128,N_3113);
nand U3218 (N_3218,N_3146,N_3123);
or U3219 (N_3219,N_3143,N_3160);
nor U3220 (N_3220,N_3173,N_3109);
or U3221 (N_3221,N_3144,N_3169);
nor U3222 (N_3222,N_3147,N_3135);
xnor U3223 (N_3223,N_3184,N_3194);
xor U3224 (N_3224,N_3154,N_3136);
nand U3225 (N_3225,N_3122,N_3161);
and U3226 (N_3226,N_3126,N_3130);
or U3227 (N_3227,N_3162,N_3185);
or U3228 (N_3228,N_3139,N_3166);
or U3229 (N_3229,N_3192,N_3195);
nand U3230 (N_3230,N_3191,N_3101);
nand U3231 (N_3231,N_3118,N_3149);
nor U3232 (N_3232,N_3176,N_3171);
xnor U3233 (N_3233,N_3177,N_3127);
xor U3234 (N_3234,N_3153,N_3152);
nor U3235 (N_3235,N_3157,N_3168);
and U3236 (N_3236,N_3133,N_3129);
nand U3237 (N_3237,N_3141,N_3150);
xnor U3238 (N_3238,N_3100,N_3108);
and U3239 (N_3239,N_3199,N_3182);
or U3240 (N_3240,N_3198,N_3172);
or U3241 (N_3241,N_3179,N_3178);
nand U3242 (N_3242,N_3187,N_3102);
nor U3243 (N_3243,N_3140,N_3117);
xor U3244 (N_3244,N_3163,N_3183);
xnor U3245 (N_3245,N_3114,N_3186);
nor U3246 (N_3246,N_3158,N_3180);
and U3247 (N_3247,N_3196,N_3175);
xnor U3248 (N_3248,N_3115,N_3174);
xor U3249 (N_3249,N_3116,N_3124);
nor U3250 (N_3250,N_3174,N_3141);
nand U3251 (N_3251,N_3174,N_3195);
and U3252 (N_3252,N_3134,N_3114);
nor U3253 (N_3253,N_3157,N_3154);
or U3254 (N_3254,N_3149,N_3107);
nand U3255 (N_3255,N_3193,N_3169);
xnor U3256 (N_3256,N_3177,N_3111);
or U3257 (N_3257,N_3137,N_3152);
nand U3258 (N_3258,N_3147,N_3106);
xnor U3259 (N_3259,N_3170,N_3122);
and U3260 (N_3260,N_3172,N_3161);
or U3261 (N_3261,N_3152,N_3142);
xnor U3262 (N_3262,N_3196,N_3101);
xnor U3263 (N_3263,N_3192,N_3117);
and U3264 (N_3264,N_3138,N_3104);
and U3265 (N_3265,N_3152,N_3155);
nand U3266 (N_3266,N_3140,N_3195);
and U3267 (N_3267,N_3157,N_3145);
and U3268 (N_3268,N_3134,N_3187);
xnor U3269 (N_3269,N_3152,N_3182);
xnor U3270 (N_3270,N_3108,N_3199);
and U3271 (N_3271,N_3183,N_3138);
and U3272 (N_3272,N_3161,N_3164);
or U3273 (N_3273,N_3116,N_3176);
xnor U3274 (N_3274,N_3160,N_3149);
xor U3275 (N_3275,N_3160,N_3123);
or U3276 (N_3276,N_3177,N_3114);
xor U3277 (N_3277,N_3133,N_3120);
xor U3278 (N_3278,N_3119,N_3160);
or U3279 (N_3279,N_3199,N_3174);
or U3280 (N_3280,N_3163,N_3123);
nand U3281 (N_3281,N_3167,N_3183);
nor U3282 (N_3282,N_3126,N_3176);
or U3283 (N_3283,N_3120,N_3138);
nor U3284 (N_3284,N_3175,N_3131);
and U3285 (N_3285,N_3105,N_3172);
nand U3286 (N_3286,N_3178,N_3160);
xor U3287 (N_3287,N_3102,N_3105);
and U3288 (N_3288,N_3147,N_3179);
or U3289 (N_3289,N_3186,N_3140);
and U3290 (N_3290,N_3120,N_3198);
nor U3291 (N_3291,N_3159,N_3121);
nand U3292 (N_3292,N_3181,N_3113);
and U3293 (N_3293,N_3145,N_3103);
and U3294 (N_3294,N_3157,N_3199);
and U3295 (N_3295,N_3110,N_3114);
xor U3296 (N_3296,N_3185,N_3184);
and U3297 (N_3297,N_3151,N_3142);
nand U3298 (N_3298,N_3113,N_3138);
nor U3299 (N_3299,N_3190,N_3186);
and U3300 (N_3300,N_3242,N_3250);
xnor U3301 (N_3301,N_3263,N_3280);
and U3302 (N_3302,N_3287,N_3217);
nand U3303 (N_3303,N_3256,N_3241);
nor U3304 (N_3304,N_3254,N_3282);
nand U3305 (N_3305,N_3227,N_3215);
nand U3306 (N_3306,N_3258,N_3286);
or U3307 (N_3307,N_3204,N_3234);
xor U3308 (N_3308,N_3294,N_3213);
nor U3309 (N_3309,N_3216,N_3210);
nor U3310 (N_3310,N_3226,N_3253);
nand U3311 (N_3311,N_3221,N_3291);
nand U3312 (N_3312,N_3247,N_3285);
and U3313 (N_3313,N_3235,N_3249);
or U3314 (N_3314,N_3293,N_3262);
or U3315 (N_3315,N_3274,N_3224);
and U3316 (N_3316,N_3231,N_3205);
nor U3317 (N_3317,N_3246,N_3207);
nand U3318 (N_3318,N_3223,N_3270);
and U3319 (N_3319,N_3232,N_3260);
nor U3320 (N_3320,N_3261,N_3279);
xnor U3321 (N_3321,N_3230,N_3218);
and U3322 (N_3322,N_3219,N_3267);
nand U3323 (N_3323,N_3292,N_3278);
nor U3324 (N_3324,N_3203,N_3212);
xnor U3325 (N_3325,N_3271,N_3211);
xor U3326 (N_3326,N_3259,N_3295);
nor U3327 (N_3327,N_3265,N_3272);
or U3328 (N_3328,N_3200,N_3284);
and U3329 (N_3329,N_3251,N_3229);
nand U3330 (N_3330,N_3289,N_3233);
or U3331 (N_3331,N_3206,N_3209);
nand U3332 (N_3332,N_3288,N_3236);
or U3333 (N_3333,N_3248,N_3208);
xor U3334 (N_3334,N_3225,N_3275);
xor U3335 (N_3335,N_3255,N_3283);
nand U3336 (N_3336,N_3268,N_3220);
and U3337 (N_3337,N_3202,N_3297);
nor U3338 (N_3338,N_3298,N_3201);
nor U3339 (N_3339,N_3269,N_3238);
xnor U3340 (N_3340,N_3237,N_3281);
nor U3341 (N_3341,N_3257,N_3276);
xor U3342 (N_3342,N_3266,N_3239);
xnor U3343 (N_3343,N_3244,N_3214);
and U3344 (N_3344,N_3252,N_3245);
nand U3345 (N_3345,N_3290,N_3296);
and U3346 (N_3346,N_3240,N_3277);
xor U3347 (N_3347,N_3299,N_3273);
nand U3348 (N_3348,N_3264,N_3228);
and U3349 (N_3349,N_3243,N_3222);
or U3350 (N_3350,N_3238,N_3226);
or U3351 (N_3351,N_3295,N_3287);
and U3352 (N_3352,N_3200,N_3218);
and U3353 (N_3353,N_3229,N_3222);
or U3354 (N_3354,N_3267,N_3221);
or U3355 (N_3355,N_3297,N_3281);
or U3356 (N_3356,N_3295,N_3208);
or U3357 (N_3357,N_3224,N_3226);
nor U3358 (N_3358,N_3232,N_3219);
nand U3359 (N_3359,N_3221,N_3255);
xor U3360 (N_3360,N_3296,N_3263);
and U3361 (N_3361,N_3235,N_3230);
nor U3362 (N_3362,N_3234,N_3224);
xor U3363 (N_3363,N_3254,N_3202);
or U3364 (N_3364,N_3205,N_3245);
or U3365 (N_3365,N_3285,N_3204);
and U3366 (N_3366,N_3291,N_3278);
xnor U3367 (N_3367,N_3235,N_3242);
or U3368 (N_3368,N_3225,N_3228);
nand U3369 (N_3369,N_3258,N_3270);
nand U3370 (N_3370,N_3285,N_3289);
nor U3371 (N_3371,N_3269,N_3207);
or U3372 (N_3372,N_3255,N_3256);
nor U3373 (N_3373,N_3296,N_3271);
or U3374 (N_3374,N_3207,N_3239);
xnor U3375 (N_3375,N_3257,N_3254);
nand U3376 (N_3376,N_3248,N_3223);
and U3377 (N_3377,N_3204,N_3291);
nand U3378 (N_3378,N_3262,N_3235);
or U3379 (N_3379,N_3229,N_3234);
nand U3380 (N_3380,N_3205,N_3274);
nand U3381 (N_3381,N_3255,N_3224);
or U3382 (N_3382,N_3219,N_3286);
or U3383 (N_3383,N_3287,N_3265);
or U3384 (N_3384,N_3292,N_3256);
nor U3385 (N_3385,N_3213,N_3271);
and U3386 (N_3386,N_3266,N_3229);
and U3387 (N_3387,N_3257,N_3256);
nor U3388 (N_3388,N_3293,N_3265);
nand U3389 (N_3389,N_3285,N_3267);
or U3390 (N_3390,N_3209,N_3267);
nand U3391 (N_3391,N_3210,N_3238);
xnor U3392 (N_3392,N_3269,N_3227);
nor U3393 (N_3393,N_3274,N_3276);
or U3394 (N_3394,N_3289,N_3263);
nor U3395 (N_3395,N_3223,N_3285);
xor U3396 (N_3396,N_3220,N_3221);
or U3397 (N_3397,N_3211,N_3287);
and U3398 (N_3398,N_3240,N_3257);
and U3399 (N_3399,N_3205,N_3259);
and U3400 (N_3400,N_3347,N_3330);
xnor U3401 (N_3401,N_3323,N_3340);
xor U3402 (N_3402,N_3392,N_3328);
nand U3403 (N_3403,N_3332,N_3377);
and U3404 (N_3404,N_3367,N_3353);
nor U3405 (N_3405,N_3354,N_3379);
or U3406 (N_3406,N_3318,N_3351);
xnor U3407 (N_3407,N_3344,N_3343);
and U3408 (N_3408,N_3324,N_3338);
or U3409 (N_3409,N_3365,N_3325);
or U3410 (N_3410,N_3384,N_3305);
or U3411 (N_3411,N_3382,N_3319);
nor U3412 (N_3412,N_3301,N_3300);
nor U3413 (N_3413,N_3322,N_3363);
and U3414 (N_3414,N_3375,N_3333);
or U3415 (N_3415,N_3394,N_3398);
nand U3416 (N_3416,N_3397,N_3372);
or U3417 (N_3417,N_3371,N_3321);
or U3418 (N_3418,N_3378,N_3381);
nand U3419 (N_3419,N_3306,N_3356);
and U3420 (N_3420,N_3390,N_3337);
nand U3421 (N_3421,N_3316,N_3352);
xnor U3422 (N_3422,N_3303,N_3311);
nor U3423 (N_3423,N_3385,N_3395);
xor U3424 (N_3424,N_3369,N_3327);
or U3425 (N_3425,N_3334,N_3345);
or U3426 (N_3426,N_3335,N_3309);
nor U3427 (N_3427,N_3387,N_3331);
nor U3428 (N_3428,N_3368,N_3302);
nand U3429 (N_3429,N_3304,N_3399);
or U3430 (N_3430,N_3341,N_3396);
or U3431 (N_3431,N_3310,N_3383);
nand U3432 (N_3432,N_3359,N_3366);
and U3433 (N_3433,N_3370,N_3308);
and U3434 (N_3434,N_3391,N_3307);
xnor U3435 (N_3435,N_3373,N_3362);
and U3436 (N_3436,N_3393,N_3358);
xor U3437 (N_3437,N_3374,N_3361);
nor U3438 (N_3438,N_3346,N_3355);
and U3439 (N_3439,N_3329,N_3339);
nand U3440 (N_3440,N_3313,N_3360);
xor U3441 (N_3441,N_3388,N_3342);
nor U3442 (N_3442,N_3314,N_3312);
xor U3443 (N_3443,N_3350,N_3317);
xnor U3444 (N_3444,N_3386,N_3364);
xnor U3445 (N_3445,N_3326,N_3349);
xnor U3446 (N_3446,N_3357,N_3389);
nand U3447 (N_3447,N_3380,N_3320);
xor U3448 (N_3448,N_3336,N_3376);
and U3449 (N_3449,N_3315,N_3348);
and U3450 (N_3450,N_3363,N_3344);
xnor U3451 (N_3451,N_3314,N_3363);
nor U3452 (N_3452,N_3349,N_3383);
and U3453 (N_3453,N_3361,N_3399);
or U3454 (N_3454,N_3308,N_3361);
nand U3455 (N_3455,N_3323,N_3398);
and U3456 (N_3456,N_3320,N_3369);
nand U3457 (N_3457,N_3305,N_3368);
nor U3458 (N_3458,N_3353,N_3314);
and U3459 (N_3459,N_3355,N_3329);
or U3460 (N_3460,N_3318,N_3386);
and U3461 (N_3461,N_3318,N_3322);
nand U3462 (N_3462,N_3343,N_3353);
and U3463 (N_3463,N_3386,N_3394);
and U3464 (N_3464,N_3337,N_3322);
and U3465 (N_3465,N_3306,N_3341);
xnor U3466 (N_3466,N_3337,N_3328);
and U3467 (N_3467,N_3374,N_3395);
nand U3468 (N_3468,N_3300,N_3353);
nor U3469 (N_3469,N_3367,N_3362);
xor U3470 (N_3470,N_3352,N_3303);
nand U3471 (N_3471,N_3352,N_3326);
nor U3472 (N_3472,N_3368,N_3380);
nand U3473 (N_3473,N_3347,N_3380);
nor U3474 (N_3474,N_3378,N_3365);
xnor U3475 (N_3475,N_3382,N_3312);
or U3476 (N_3476,N_3370,N_3337);
nor U3477 (N_3477,N_3336,N_3342);
nand U3478 (N_3478,N_3325,N_3314);
or U3479 (N_3479,N_3384,N_3391);
xor U3480 (N_3480,N_3318,N_3359);
or U3481 (N_3481,N_3371,N_3332);
nor U3482 (N_3482,N_3359,N_3330);
and U3483 (N_3483,N_3338,N_3323);
and U3484 (N_3484,N_3316,N_3353);
nand U3485 (N_3485,N_3351,N_3331);
and U3486 (N_3486,N_3359,N_3354);
and U3487 (N_3487,N_3383,N_3338);
nor U3488 (N_3488,N_3315,N_3339);
and U3489 (N_3489,N_3374,N_3306);
or U3490 (N_3490,N_3354,N_3357);
xor U3491 (N_3491,N_3302,N_3374);
or U3492 (N_3492,N_3377,N_3371);
nor U3493 (N_3493,N_3395,N_3347);
xor U3494 (N_3494,N_3358,N_3354);
or U3495 (N_3495,N_3352,N_3370);
nand U3496 (N_3496,N_3333,N_3332);
or U3497 (N_3497,N_3345,N_3352);
or U3498 (N_3498,N_3389,N_3380);
nand U3499 (N_3499,N_3357,N_3328);
and U3500 (N_3500,N_3430,N_3413);
nor U3501 (N_3501,N_3487,N_3494);
nand U3502 (N_3502,N_3421,N_3450);
xor U3503 (N_3503,N_3414,N_3474);
xnor U3504 (N_3504,N_3493,N_3417);
nor U3505 (N_3505,N_3495,N_3400);
nand U3506 (N_3506,N_3441,N_3463);
and U3507 (N_3507,N_3490,N_3419);
xor U3508 (N_3508,N_3468,N_3447);
or U3509 (N_3509,N_3428,N_3458);
nand U3510 (N_3510,N_3451,N_3457);
or U3511 (N_3511,N_3401,N_3435);
xor U3512 (N_3512,N_3431,N_3489);
or U3513 (N_3513,N_3406,N_3498);
and U3514 (N_3514,N_3433,N_3470);
nor U3515 (N_3515,N_3403,N_3461);
or U3516 (N_3516,N_3473,N_3437);
or U3517 (N_3517,N_3454,N_3476);
and U3518 (N_3518,N_3464,N_3411);
nand U3519 (N_3519,N_3492,N_3480);
nor U3520 (N_3520,N_3424,N_3496);
or U3521 (N_3521,N_3405,N_3442);
xnor U3522 (N_3522,N_3416,N_3481);
xor U3523 (N_3523,N_3491,N_3499);
xnor U3524 (N_3524,N_3408,N_3434);
xor U3525 (N_3525,N_3484,N_3409);
xor U3526 (N_3526,N_3427,N_3436);
nand U3527 (N_3527,N_3475,N_3443);
and U3528 (N_3528,N_3467,N_3456);
nand U3529 (N_3529,N_3483,N_3477);
nor U3530 (N_3530,N_3438,N_3478);
nand U3531 (N_3531,N_3459,N_3440);
nor U3532 (N_3532,N_3448,N_3425);
nand U3533 (N_3533,N_3423,N_3472);
nor U3534 (N_3534,N_3404,N_3453);
and U3535 (N_3535,N_3486,N_3452);
nor U3536 (N_3536,N_3446,N_3469);
or U3537 (N_3537,N_3418,N_3445);
xnor U3538 (N_3538,N_3465,N_3462);
xor U3539 (N_3539,N_3426,N_3482);
or U3540 (N_3540,N_3402,N_3485);
nor U3541 (N_3541,N_3449,N_3412);
or U3542 (N_3542,N_3407,N_3432);
or U3543 (N_3543,N_3420,N_3497);
or U3544 (N_3544,N_3422,N_3466);
xnor U3545 (N_3545,N_3455,N_3444);
or U3546 (N_3546,N_3410,N_3488);
and U3547 (N_3547,N_3429,N_3479);
xnor U3548 (N_3548,N_3415,N_3460);
nor U3549 (N_3549,N_3471,N_3439);
or U3550 (N_3550,N_3412,N_3486);
and U3551 (N_3551,N_3482,N_3437);
nor U3552 (N_3552,N_3440,N_3428);
nand U3553 (N_3553,N_3454,N_3464);
nand U3554 (N_3554,N_3486,N_3477);
xor U3555 (N_3555,N_3485,N_3401);
and U3556 (N_3556,N_3401,N_3429);
xnor U3557 (N_3557,N_3460,N_3499);
xnor U3558 (N_3558,N_3497,N_3400);
or U3559 (N_3559,N_3403,N_3441);
xnor U3560 (N_3560,N_3455,N_3415);
and U3561 (N_3561,N_3403,N_3467);
nand U3562 (N_3562,N_3472,N_3467);
nor U3563 (N_3563,N_3465,N_3444);
or U3564 (N_3564,N_3461,N_3490);
or U3565 (N_3565,N_3459,N_3453);
xnor U3566 (N_3566,N_3494,N_3483);
xnor U3567 (N_3567,N_3405,N_3478);
xor U3568 (N_3568,N_3478,N_3481);
nand U3569 (N_3569,N_3461,N_3426);
nor U3570 (N_3570,N_3442,N_3483);
nand U3571 (N_3571,N_3467,N_3402);
nand U3572 (N_3572,N_3460,N_3401);
xnor U3573 (N_3573,N_3421,N_3448);
xnor U3574 (N_3574,N_3480,N_3440);
nand U3575 (N_3575,N_3493,N_3463);
nor U3576 (N_3576,N_3456,N_3400);
xnor U3577 (N_3577,N_3468,N_3403);
nor U3578 (N_3578,N_3457,N_3476);
and U3579 (N_3579,N_3408,N_3407);
nand U3580 (N_3580,N_3495,N_3408);
and U3581 (N_3581,N_3434,N_3444);
or U3582 (N_3582,N_3415,N_3494);
or U3583 (N_3583,N_3454,N_3489);
xnor U3584 (N_3584,N_3433,N_3447);
or U3585 (N_3585,N_3499,N_3459);
xor U3586 (N_3586,N_3409,N_3434);
nor U3587 (N_3587,N_3414,N_3489);
nand U3588 (N_3588,N_3474,N_3433);
nand U3589 (N_3589,N_3486,N_3444);
nand U3590 (N_3590,N_3419,N_3473);
nand U3591 (N_3591,N_3480,N_3423);
and U3592 (N_3592,N_3439,N_3433);
and U3593 (N_3593,N_3412,N_3497);
or U3594 (N_3594,N_3427,N_3400);
xnor U3595 (N_3595,N_3486,N_3450);
nand U3596 (N_3596,N_3443,N_3427);
or U3597 (N_3597,N_3464,N_3410);
or U3598 (N_3598,N_3404,N_3444);
or U3599 (N_3599,N_3473,N_3458);
or U3600 (N_3600,N_3559,N_3574);
xor U3601 (N_3601,N_3579,N_3589);
nand U3602 (N_3602,N_3503,N_3592);
and U3603 (N_3603,N_3542,N_3583);
nor U3604 (N_3604,N_3537,N_3523);
nor U3605 (N_3605,N_3599,N_3518);
nor U3606 (N_3606,N_3560,N_3540);
and U3607 (N_3607,N_3564,N_3538);
nor U3608 (N_3608,N_3590,N_3507);
or U3609 (N_3609,N_3511,N_3500);
nor U3610 (N_3610,N_3570,N_3598);
xnor U3611 (N_3611,N_3515,N_3575);
or U3612 (N_3612,N_3534,N_3584);
nand U3613 (N_3613,N_3525,N_3571);
nor U3614 (N_3614,N_3551,N_3562);
xnor U3615 (N_3615,N_3550,N_3508);
xnor U3616 (N_3616,N_3544,N_3580);
or U3617 (N_3617,N_3545,N_3530);
or U3618 (N_3618,N_3506,N_3597);
nand U3619 (N_3619,N_3568,N_3594);
nor U3620 (N_3620,N_3533,N_3581);
nand U3621 (N_3621,N_3576,N_3573);
or U3622 (N_3622,N_3595,N_3536);
xnor U3623 (N_3623,N_3539,N_3578);
and U3624 (N_3624,N_3529,N_3566);
nand U3625 (N_3625,N_3524,N_3557);
and U3626 (N_3626,N_3563,N_3510);
and U3627 (N_3627,N_3521,N_3519);
and U3628 (N_3628,N_3505,N_3561);
and U3629 (N_3629,N_3554,N_3543);
or U3630 (N_3630,N_3531,N_3582);
or U3631 (N_3631,N_3586,N_3547);
nor U3632 (N_3632,N_3516,N_3577);
and U3633 (N_3633,N_3549,N_3527);
xor U3634 (N_3634,N_3555,N_3517);
nor U3635 (N_3635,N_3567,N_3588);
nand U3636 (N_3636,N_3526,N_3553);
nand U3637 (N_3637,N_3528,N_3514);
xnor U3638 (N_3638,N_3569,N_3596);
or U3639 (N_3639,N_3520,N_3532);
xnor U3640 (N_3640,N_3558,N_3585);
or U3641 (N_3641,N_3504,N_3502);
nand U3642 (N_3642,N_3556,N_3565);
nand U3643 (N_3643,N_3541,N_3513);
and U3644 (N_3644,N_3522,N_3591);
nor U3645 (N_3645,N_3501,N_3572);
nand U3646 (N_3646,N_3535,N_3552);
xor U3647 (N_3647,N_3509,N_3512);
nand U3648 (N_3648,N_3548,N_3587);
or U3649 (N_3649,N_3546,N_3593);
xnor U3650 (N_3650,N_3526,N_3521);
xor U3651 (N_3651,N_3586,N_3599);
nand U3652 (N_3652,N_3544,N_3542);
xor U3653 (N_3653,N_3576,N_3543);
nor U3654 (N_3654,N_3581,N_3555);
and U3655 (N_3655,N_3503,N_3506);
and U3656 (N_3656,N_3595,N_3569);
xor U3657 (N_3657,N_3578,N_3571);
nor U3658 (N_3658,N_3512,N_3572);
nand U3659 (N_3659,N_3569,N_3538);
or U3660 (N_3660,N_3576,N_3541);
nor U3661 (N_3661,N_3517,N_3590);
xnor U3662 (N_3662,N_3549,N_3568);
nor U3663 (N_3663,N_3547,N_3575);
xor U3664 (N_3664,N_3504,N_3539);
xnor U3665 (N_3665,N_3524,N_3533);
nand U3666 (N_3666,N_3511,N_3582);
nor U3667 (N_3667,N_3545,N_3514);
xnor U3668 (N_3668,N_3573,N_3588);
xor U3669 (N_3669,N_3555,N_3599);
xnor U3670 (N_3670,N_3549,N_3516);
or U3671 (N_3671,N_3596,N_3513);
nor U3672 (N_3672,N_3590,N_3536);
nor U3673 (N_3673,N_3557,N_3504);
nor U3674 (N_3674,N_3513,N_3572);
nor U3675 (N_3675,N_3556,N_3574);
nor U3676 (N_3676,N_3545,N_3560);
and U3677 (N_3677,N_3565,N_3524);
nand U3678 (N_3678,N_3560,N_3589);
xnor U3679 (N_3679,N_3557,N_3560);
or U3680 (N_3680,N_3507,N_3593);
nand U3681 (N_3681,N_3545,N_3572);
and U3682 (N_3682,N_3556,N_3505);
nor U3683 (N_3683,N_3558,N_3536);
nor U3684 (N_3684,N_3541,N_3506);
and U3685 (N_3685,N_3517,N_3508);
or U3686 (N_3686,N_3592,N_3583);
xnor U3687 (N_3687,N_3557,N_3558);
nor U3688 (N_3688,N_3510,N_3524);
nor U3689 (N_3689,N_3591,N_3509);
and U3690 (N_3690,N_3514,N_3552);
and U3691 (N_3691,N_3544,N_3591);
or U3692 (N_3692,N_3557,N_3501);
nor U3693 (N_3693,N_3528,N_3523);
or U3694 (N_3694,N_3551,N_3541);
nand U3695 (N_3695,N_3500,N_3595);
nor U3696 (N_3696,N_3598,N_3592);
nand U3697 (N_3697,N_3534,N_3559);
nand U3698 (N_3698,N_3534,N_3514);
nor U3699 (N_3699,N_3561,N_3597);
nand U3700 (N_3700,N_3691,N_3616);
or U3701 (N_3701,N_3615,N_3694);
nand U3702 (N_3702,N_3630,N_3699);
or U3703 (N_3703,N_3660,N_3614);
xor U3704 (N_3704,N_3679,N_3650);
nand U3705 (N_3705,N_3675,N_3669);
xnor U3706 (N_3706,N_3662,N_3611);
nand U3707 (N_3707,N_3684,N_3620);
and U3708 (N_3708,N_3693,N_3631);
and U3709 (N_3709,N_3641,N_3653);
xnor U3710 (N_3710,N_3692,N_3685);
and U3711 (N_3711,N_3647,N_3666);
nand U3712 (N_3712,N_3689,N_3678);
nand U3713 (N_3713,N_3636,N_3651);
nand U3714 (N_3714,N_3655,N_3658);
nor U3715 (N_3715,N_3610,N_3613);
nand U3716 (N_3716,N_3686,N_3668);
or U3717 (N_3717,N_3628,N_3639);
and U3718 (N_3718,N_3607,N_3665);
or U3719 (N_3719,N_3626,N_3652);
nand U3720 (N_3720,N_3635,N_3663);
nand U3721 (N_3721,N_3671,N_3648);
and U3722 (N_3722,N_3698,N_3600);
xor U3723 (N_3723,N_3608,N_3623);
nor U3724 (N_3724,N_3622,N_3609);
and U3725 (N_3725,N_3672,N_3612);
nand U3726 (N_3726,N_3659,N_3643);
xor U3727 (N_3727,N_3645,N_3633);
nand U3728 (N_3728,N_3618,N_3627);
and U3729 (N_3729,N_3603,N_3619);
nand U3730 (N_3730,N_3602,N_3632);
nor U3731 (N_3731,N_3601,N_3682);
or U3732 (N_3732,N_3690,N_3661);
xnor U3733 (N_3733,N_3625,N_3629);
and U3734 (N_3734,N_3674,N_3617);
xor U3735 (N_3735,N_3683,N_3657);
nor U3736 (N_3736,N_3604,N_3681);
nand U3737 (N_3737,N_3637,N_3644);
nor U3738 (N_3738,N_3688,N_3670);
or U3739 (N_3739,N_3677,N_3664);
xnor U3740 (N_3740,N_3654,N_3640);
xor U3741 (N_3741,N_3667,N_3642);
and U3742 (N_3742,N_3696,N_3673);
or U3743 (N_3743,N_3606,N_3649);
nand U3744 (N_3744,N_3634,N_3695);
xor U3745 (N_3745,N_3680,N_3605);
nor U3746 (N_3746,N_3646,N_3676);
nand U3747 (N_3747,N_3621,N_3638);
xor U3748 (N_3748,N_3624,N_3656);
nand U3749 (N_3749,N_3687,N_3697);
nor U3750 (N_3750,N_3604,N_3623);
nand U3751 (N_3751,N_3610,N_3664);
nand U3752 (N_3752,N_3683,N_3617);
nand U3753 (N_3753,N_3696,N_3620);
or U3754 (N_3754,N_3695,N_3606);
nand U3755 (N_3755,N_3608,N_3621);
nand U3756 (N_3756,N_3656,N_3674);
xnor U3757 (N_3757,N_3608,N_3640);
and U3758 (N_3758,N_3635,N_3632);
nand U3759 (N_3759,N_3682,N_3695);
or U3760 (N_3760,N_3697,N_3606);
nor U3761 (N_3761,N_3612,N_3658);
xnor U3762 (N_3762,N_3642,N_3621);
or U3763 (N_3763,N_3660,N_3696);
and U3764 (N_3764,N_3608,N_3675);
nand U3765 (N_3765,N_3699,N_3621);
and U3766 (N_3766,N_3671,N_3634);
nand U3767 (N_3767,N_3639,N_3611);
xor U3768 (N_3768,N_3611,N_3638);
nand U3769 (N_3769,N_3608,N_3665);
nand U3770 (N_3770,N_3622,N_3652);
nand U3771 (N_3771,N_3647,N_3672);
nor U3772 (N_3772,N_3644,N_3685);
xor U3773 (N_3773,N_3605,N_3622);
nand U3774 (N_3774,N_3620,N_3679);
or U3775 (N_3775,N_3664,N_3695);
or U3776 (N_3776,N_3626,N_3633);
or U3777 (N_3777,N_3658,N_3683);
nand U3778 (N_3778,N_3604,N_3638);
and U3779 (N_3779,N_3645,N_3627);
or U3780 (N_3780,N_3607,N_3611);
nand U3781 (N_3781,N_3624,N_3642);
nand U3782 (N_3782,N_3642,N_3650);
or U3783 (N_3783,N_3630,N_3633);
xor U3784 (N_3784,N_3698,N_3613);
nor U3785 (N_3785,N_3697,N_3681);
or U3786 (N_3786,N_3638,N_3679);
nor U3787 (N_3787,N_3676,N_3623);
and U3788 (N_3788,N_3623,N_3673);
and U3789 (N_3789,N_3603,N_3695);
nand U3790 (N_3790,N_3635,N_3687);
and U3791 (N_3791,N_3694,N_3649);
and U3792 (N_3792,N_3668,N_3698);
and U3793 (N_3793,N_3663,N_3667);
nor U3794 (N_3794,N_3698,N_3637);
and U3795 (N_3795,N_3649,N_3608);
nor U3796 (N_3796,N_3644,N_3666);
or U3797 (N_3797,N_3642,N_3669);
nand U3798 (N_3798,N_3687,N_3612);
nand U3799 (N_3799,N_3619,N_3611);
or U3800 (N_3800,N_3776,N_3705);
nand U3801 (N_3801,N_3789,N_3796);
or U3802 (N_3802,N_3773,N_3713);
or U3803 (N_3803,N_3766,N_3791);
nand U3804 (N_3804,N_3786,N_3711);
or U3805 (N_3805,N_3715,N_3721);
xnor U3806 (N_3806,N_3746,N_3726);
nor U3807 (N_3807,N_3701,N_3748);
and U3808 (N_3808,N_3774,N_3775);
and U3809 (N_3809,N_3798,N_3722);
nand U3810 (N_3810,N_3708,N_3743);
xor U3811 (N_3811,N_3744,N_3717);
nand U3812 (N_3812,N_3757,N_3700);
xnor U3813 (N_3813,N_3771,N_3797);
xor U3814 (N_3814,N_3799,N_3707);
nand U3815 (N_3815,N_3735,N_3730);
or U3816 (N_3816,N_3706,N_3778);
nand U3817 (N_3817,N_3709,N_3759);
xnor U3818 (N_3818,N_3731,N_3741);
nand U3819 (N_3819,N_3781,N_3742);
nor U3820 (N_3820,N_3779,N_3763);
nand U3821 (N_3821,N_3732,N_3783);
or U3822 (N_3822,N_3758,N_3734);
or U3823 (N_3823,N_3790,N_3740);
nor U3824 (N_3824,N_3792,N_3787);
nor U3825 (N_3825,N_3764,N_3780);
or U3826 (N_3826,N_3794,N_3749);
and U3827 (N_3827,N_3719,N_3752);
nor U3828 (N_3828,N_3736,N_3712);
nor U3829 (N_3829,N_3751,N_3777);
xor U3830 (N_3830,N_3702,N_3765);
and U3831 (N_3831,N_3785,N_3737);
and U3832 (N_3832,N_3703,N_3788);
nand U3833 (N_3833,N_3782,N_3770);
nor U3834 (N_3834,N_3724,N_3733);
xor U3835 (N_3835,N_3755,N_3784);
and U3836 (N_3836,N_3772,N_3714);
nor U3837 (N_3837,N_3750,N_3745);
nor U3838 (N_3838,N_3718,N_3725);
nor U3839 (N_3839,N_3728,N_3768);
xnor U3840 (N_3840,N_3729,N_3767);
nand U3841 (N_3841,N_3756,N_3738);
nand U3842 (N_3842,N_3747,N_3739);
and U3843 (N_3843,N_3710,N_3769);
nand U3844 (N_3844,N_3760,N_3761);
nand U3845 (N_3845,N_3704,N_3727);
xor U3846 (N_3846,N_3762,N_3754);
xor U3847 (N_3847,N_3795,N_3723);
and U3848 (N_3848,N_3753,N_3793);
xnor U3849 (N_3849,N_3720,N_3716);
or U3850 (N_3850,N_3765,N_3720);
nand U3851 (N_3851,N_3790,N_3747);
and U3852 (N_3852,N_3770,N_3779);
or U3853 (N_3853,N_3785,N_3739);
nor U3854 (N_3854,N_3730,N_3765);
nand U3855 (N_3855,N_3734,N_3738);
nand U3856 (N_3856,N_3738,N_3754);
nand U3857 (N_3857,N_3791,N_3723);
and U3858 (N_3858,N_3786,N_3712);
nor U3859 (N_3859,N_3783,N_3799);
and U3860 (N_3860,N_3757,N_3723);
nand U3861 (N_3861,N_3726,N_3708);
xor U3862 (N_3862,N_3797,N_3786);
nor U3863 (N_3863,N_3718,N_3733);
or U3864 (N_3864,N_3716,N_3728);
nor U3865 (N_3865,N_3738,N_3726);
or U3866 (N_3866,N_3779,N_3785);
xor U3867 (N_3867,N_3706,N_3747);
nor U3868 (N_3868,N_3762,N_3718);
xnor U3869 (N_3869,N_3774,N_3794);
xor U3870 (N_3870,N_3781,N_3764);
nor U3871 (N_3871,N_3778,N_3742);
nor U3872 (N_3872,N_3714,N_3777);
or U3873 (N_3873,N_3738,N_3777);
or U3874 (N_3874,N_3792,N_3715);
nand U3875 (N_3875,N_3784,N_3785);
or U3876 (N_3876,N_3739,N_3796);
nor U3877 (N_3877,N_3708,N_3751);
xnor U3878 (N_3878,N_3775,N_3786);
and U3879 (N_3879,N_3745,N_3739);
nor U3880 (N_3880,N_3771,N_3769);
and U3881 (N_3881,N_3703,N_3770);
nor U3882 (N_3882,N_3751,N_3786);
or U3883 (N_3883,N_3774,N_3751);
nor U3884 (N_3884,N_3733,N_3782);
and U3885 (N_3885,N_3771,N_3700);
nand U3886 (N_3886,N_3718,N_3784);
xnor U3887 (N_3887,N_3782,N_3747);
xor U3888 (N_3888,N_3764,N_3775);
and U3889 (N_3889,N_3700,N_3772);
xnor U3890 (N_3890,N_3780,N_3756);
xnor U3891 (N_3891,N_3726,N_3751);
or U3892 (N_3892,N_3769,N_3755);
or U3893 (N_3893,N_3704,N_3737);
nand U3894 (N_3894,N_3792,N_3754);
xnor U3895 (N_3895,N_3738,N_3769);
nor U3896 (N_3896,N_3739,N_3753);
and U3897 (N_3897,N_3773,N_3708);
nor U3898 (N_3898,N_3719,N_3768);
and U3899 (N_3899,N_3712,N_3758);
xor U3900 (N_3900,N_3804,N_3889);
and U3901 (N_3901,N_3841,N_3885);
xor U3902 (N_3902,N_3878,N_3849);
nor U3903 (N_3903,N_3896,N_3869);
nor U3904 (N_3904,N_3887,N_3846);
xor U3905 (N_3905,N_3882,N_3897);
xnor U3906 (N_3906,N_3823,N_3864);
nand U3907 (N_3907,N_3845,N_3873);
xnor U3908 (N_3908,N_3862,N_3812);
nand U3909 (N_3909,N_3847,N_3839);
xor U3910 (N_3910,N_3874,N_3868);
nand U3911 (N_3911,N_3805,N_3827);
xnor U3912 (N_3912,N_3892,N_3884);
xnor U3913 (N_3913,N_3809,N_3848);
and U3914 (N_3914,N_3871,N_3818);
or U3915 (N_3915,N_3894,N_3837);
or U3916 (N_3916,N_3854,N_3899);
and U3917 (N_3917,N_3824,N_3880);
xnor U3918 (N_3918,N_3816,N_3815);
nand U3919 (N_3919,N_3829,N_3886);
nand U3920 (N_3920,N_3875,N_3851);
nand U3921 (N_3921,N_3852,N_3821);
xnor U3922 (N_3922,N_3822,N_3858);
or U3923 (N_3923,N_3881,N_3866);
nor U3924 (N_3924,N_3870,N_3876);
nor U3925 (N_3925,N_3800,N_3861);
or U3926 (N_3926,N_3883,N_3835);
nor U3927 (N_3927,N_3853,N_3828);
xor U3928 (N_3928,N_3893,N_3820);
and U3929 (N_3929,N_3898,N_3850);
nand U3930 (N_3930,N_3831,N_3819);
nand U3931 (N_3931,N_3860,N_3840);
xnor U3932 (N_3932,N_3836,N_3801);
and U3933 (N_3933,N_3863,N_3888);
xnor U3934 (N_3934,N_3855,N_3867);
and U3935 (N_3935,N_3879,N_3877);
nand U3936 (N_3936,N_3808,N_3802);
and U3937 (N_3937,N_3842,N_3806);
xnor U3938 (N_3938,N_3810,N_3859);
xnor U3939 (N_3939,N_3844,N_3814);
and U3940 (N_3940,N_3857,N_3895);
nor U3941 (N_3941,N_3834,N_3807);
or U3942 (N_3942,N_3813,N_3803);
xnor U3943 (N_3943,N_3832,N_3825);
xnor U3944 (N_3944,N_3830,N_3838);
nor U3945 (N_3945,N_3826,N_3890);
nor U3946 (N_3946,N_3856,N_3833);
nor U3947 (N_3947,N_3843,N_3891);
nand U3948 (N_3948,N_3811,N_3872);
nand U3949 (N_3949,N_3865,N_3817);
or U3950 (N_3950,N_3810,N_3868);
nand U3951 (N_3951,N_3832,N_3807);
xor U3952 (N_3952,N_3838,N_3852);
xnor U3953 (N_3953,N_3862,N_3868);
xor U3954 (N_3954,N_3886,N_3807);
nand U3955 (N_3955,N_3887,N_3879);
nor U3956 (N_3956,N_3893,N_3852);
or U3957 (N_3957,N_3801,N_3898);
nor U3958 (N_3958,N_3872,N_3803);
nor U3959 (N_3959,N_3888,N_3839);
xnor U3960 (N_3960,N_3866,N_3864);
or U3961 (N_3961,N_3801,N_3868);
xnor U3962 (N_3962,N_3896,N_3892);
nor U3963 (N_3963,N_3827,N_3872);
nand U3964 (N_3964,N_3820,N_3815);
nand U3965 (N_3965,N_3811,N_3864);
nand U3966 (N_3966,N_3884,N_3896);
nor U3967 (N_3967,N_3898,N_3872);
nor U3968 (N_3968,N_3872,N_3820);
nand U3969 (N_3969,N_3851,N_3870);
xnor U3970 (N_3970,N_3806,N_3824);
nor U3971 (N_3971,N_3864,N_3892);
and U3972 (N_3972,N_3833,N_3842);
and U3973 (N_3973,N_3823,N_3879);
and U3974 (N_3974,N_3879,N_3868);
nor U3975 (N_3975,N_3827,N_3885);
or U3976 (N_3976,N_3880,N_3875);
and U3977 (N_3977,N_3840,N_3802);
and U3978 (N_3978,N_3868,N_3870);
xnor U3979 (N_3979,N_3855,N_3857);
xor U3980 (N_3980,N_3802,N_3863);
nand U3981 (N_3981,N_3815,N_3854);
xnor U3982 (N_3982,N_3889,N_3873);
or U3983 (N_3983,N_3849,N_3819);
or U3984 (N_3984,N_3835,N_3893);
nor U3985 (N_3985,N_3805,N_3828);
nor U3986 (N_3986,N_3869,N_3868);
xnor U3987 (N_3987,N_3822,N_3861);
and U3988 (N_3988,N_3807,N_3862);
nor U3989 (N_3989,N_3852,N_3860);
or U3990 (N_3990,N_3818,N_3823);
xnor U3991 (N_3991,N_3840,N_3893);
or U3992 (N_3992,N_3880,N_3866);
nand U3993 (N_3993,N_3809,N_3820);
xnor U3994 (N_3994,N_3828,N_3877);
nor U3995 (N_3995,N_3817,N_3841);
nand U3996 (N_3996,N_3805,N_3898);
or U3997 (N_3997,N_3860,N_3833);
nand U3998 (N_3998,N_3877,N_3855);
and U3999 (N_3999,N_3809,N_3824);
and U4000 (N_4000,N_3901,N_3993);
or U4001 (N_4001,N_3900,N_3947);
and U4002 (N_4002,N_3974,N_3957);
nor U4003 (N_4003,N_3976,N_3991);
or U4004 (N_4004,N_3915,N_3917);
nand U4005 (N_4005,N_3966,N_3926);
nor U4006 (N_4006,N_3943,N_3909);
nand U4007 (N_4007,N_3902,N_3972);
nand U4008 (N_4008,N_3911,N_3994);
xnor U4009 (N_4009,N_3980,N_3914);
and U4010 (N_4010,N_3983,N_3903);
and U4011 (N_4011,N_3951,N_3969);
or U4012 (N_4012,N_3973,N_3977);
xor U4013 (N_4013,N_3989,N_3986);
nor U4014 (N_4014,N_3998,N_3941);
nand U4015 (N_4015,N_3921,N_3931);
xnor U4016 (N_4016,N_3950,N_3952);
nor U4017 (N_4017,N_3913,N_3912);
xnor U4018 (N_4018,N_3963,N_3970);
nor U4019 (N_4019,N_3999,N_3982);
and U4020 (N_4020,N_3928,N_3933);
xor U4021 (N_4021,N_3916,N_3955);
nor U4022 (N_4022,N_3927,N_3924);
nor U4023 (N_4023,N_3946,N_3925);
and U4024 (N_4024,N_3995,N_3988);
xor U4025 (N_4025,N_3904,N_3979);
xor U4026 (N_4026,N_3919,N_3932);
nor U4027 (N_4027,N_3985,N_3945);
nor U4028 (N_4028,N_3960,N_3949);
xnor U4029 (N_4029,N_3975,N_3910);
nand U4030 (N_4030,N_3918,N_3923);
nor U4031 (N_4031,N_3997,N_3987);
and U4032 (N_4032,N_3939,N_3940);
nor U4033 (N_4033,N_3906,N_3938);
nand U4034 (N_4034,N_3962,N_3992);
and U4035 (N_4035,N_3936,N_3942);
and U4036 (N_4036,N_3956,N_3920);
and U4037 (N_4037,N_3953,N_3930);
and U4038 (N_4038,N_3961,N_3967);
or U4039 (N_4039,N_3981,N_3959);
nand U4040 (N_4040,N_3905,N_3984);
xnor U4041 (N_4041,N_3935,N_3958);
nor U4042 (N_4042,N_3937,N_3978);
xnor U4043 (N_4043,N_3907,N_3990);
xor U4044 (N_4044,N_3954,N_3968);
or U4045 (N_4045,N_3971,N_3934);
and U4046 (N_4046,N_3922,N_3948);
nor U4047 (N_4047,N_3996,N_3964);
nand U4048 (N_4048,N_3944,N_3965);
xor U4049 (N_4049,N_3908,N_3929);
nor U4050 (N_4050,N_3992,N_3934);
nor U4051 (N_4051,N_3952,N_3921);
nand U4052 (N_4052,N_3940,N_3997);
xor U4053 (N_4053,N_3954,N_3962);
and U4054 (N_4054,N_3980,N_3948);
or U4055 (N_4055,N_3947,N_3951);
xnor U4056 (N_4056,N_3974,N_3915);
or U4057 (N_4057,N_3937,N_3985);
or U4058 (N_4058,N_3945,N_3942);
xnor U4059 (N_4059,N_3986,N_3945);
nand U4060 (N_4060,N_3953,N_3968);
xor U4061 (N_4061,N_3913,N_3953);
nand U4062 (N_4062,N_3900,N_3925);
or U4063 (N_4063,N_3961,N_3902);
or U4064 (N_4064,N_3975,N_3920);
nor U4065 (N_4065,N_3909,N_3937);
nor U4066 (N_4066,N_3914,N_3964);
xor U4067 (N_4067,N_3971,N_3933);
nand U4068 (N_4068,N_3910,N_3974);
and U4069 (N_4069,N_3985,N_3977);
nand U4070 (N_4070,N_3903,N_3933);
xor U4071 (N_4071,N_3940,N_3933);
nand U4072 (N_4072,N_3955,N_3992);
nand U4073 (N_4073,N_3999,N_3969);
and U4074 (N_4074,N_3950,N_3906);
xor U4075 (N_4075,N_3926,N_3987);
and U4076 (N_4076,N_3984,N_3972);
xnor U4077 (N_4077,N_3925,N_3987);
nand U4078 (N_4078,N_3924,N_3975);
or U4079 (N_4079,N_3910,N_3983);
xnor U4080 (N_4080,N_3956,N_3983);
nand U4081 (N_4081,N_3928,N_3940);
or U4082 (N_4082,N_3999,N_3905);
xnor U4083 (N_4083,N_3928,N_3975);
and U4084 (N_4084,N_3902,N_3920);
nor U4085 (N_4085,N_3942,N_3941);
or U4086 (N_4086,N_3951,N_3975);
nand U4087 (N_4087,N_3911,N_3903);
and U4088 (N_4088,N_3976,N_3973);
xnor U4089 (N_4089,N_3928,N_3963);
nand U4090 (N_4090,N_3966,N_3967);
nor U4091 (N_4091,N_3935,N_3981);
nor U4092 (N_4092,N_3947,N_3942);
xnor U4093 (N_4093,N_3922,N_3960);
or U4094 (N_4094,N_3997,N_3945);
and U4095 (N_4095,N_3983,N_3984);
and U4096 (N_4096,N_3987,N_3958);
and U4097 (N_4097,N_3929,N_3981);
nor U4098 (N_4098,N_3958,N_3994);
xor U4099 (N_4099,N_3902,N_3921);
nor U4100 (N_4100,N_4086,N_4066);
or U4101 (N_4101,N_4059,N_4037);
nand U4102 (N_4102,N_4014,N_4009);
xnor U4103 (N_4103,N_4032,N_4052);
and U4104 (N_4104,N_4060,N_4062);
xor U4105 (N_4105,N_4007,N_4018);
nor U4106 (N_4106,N_4077,N_4004);
nor U4107 (N_4107,N_4024,N_4000);
xor U4108 (N_4108,N_4053,N_4061);
xor U4109 (N_4109,N_4039,N_4033);
or U4110 (N_4110,N_4003,N_4098);
nand U4111 (N_4111,N_4076,N_4038);
nor U4112 (N_4112,N_4011,N_4022);
or U4113 (N_4113,N_4088,N_4015);
nand U4114 (N_4114,N_4051,N_4075);
and U4115 (N_4115,N_4064,N_4031);
and U4116 (N_4116,N_4092,N_4005);
nor U4117 (N_4117,N_4002,N_4069);
or U4118 (N_4118,N_4068,N_4072);
and U4119 (N_4119,N_4023,N_4028);
nand U4120 (N_4120,N_4044,N_4041);
or U4121 (N_4121,N_4089,N_4049);
xnor U4122 (N_4122,N_4035,N_4047);
or U4123 (N_4123,N_4067,N_4006);
xor U4124 (N_4124,N_4095,N_4016);
and U4125 (N_4125,N_4082,N_4073);
and U4126 (N_4126,N_4099,N_4097);
nor U4127 (N_4127,N_4034,N_4074);
xnor U4128 (N_4128,N_4094,N_4096);
nor U4129 (N_4129,N_4029,N_4090);
nor U4130 (N_4130,N_4054,N_4057);
xor U4131 (N_4131,N_4036,N_4025);
nor U4132 (N_4132,N_4085,N_4084);
nor U4133 (N_4133,N_4027,N_4081);
nand U4134 (N_4134,N_4021,N_4078);
or U4135 (N_4135,N_4055,N_4026);
and U4136 (N_4136,N_4050,N_4042);
nor U4137 (N_4137,N_4020,N_4079);
or U4138 (N_4138,N_4048,N_4019);
nand U4139 (N_4139,N_4043,N_4017);
xor U4140 (N_4140,N_4013,N_4001);
xor U4141 (N_4141,N_4071,N_4070);
and U4142 (N_4142,N_4093,N_4056);
or U4143 (N_4143,N_4065,N_4030);
or U4144 (N_4144,N_4040,N_4091);
xor U4145 (N_4145,N_4012,N_4010);
nand U4146 (N_4146,N_4045,N_4087);
nand U4147 (N_4147,N_4008,N_4046);
nor U4148 (N_4148,N_4063,N_4083);
and U4149 (N_4149,N_4058,N_4080);
and U4150 (N_4150,N_4039,N_4064);
xnor U4151 (N_4151,N_4063,N_4088);
xnor U4152 (N_4152,N_4029,N_4000);
nor U4153 (N_4153,N_4082,N_4052);
xnor U4154 (N_4154,N_4087,N_4010);
and U4155 (N_4155,N_4008,N_4003);
or U4156 (N_4156,N_4078,N_4050);
or U4157 (N_4157,N_4074,N_4000);
and U4158 (N_4158,N_4062,N_4025);
nand U4159 (N_4159,N_4056,N_4079);
or U4160 (N_4160,N_4028,N_4079);
nand U4161 (N_4161,N_4034,N_4017);
or U4162 (N_4162,N_4054,N_4076);
xor U4163 (N_4163,N_4062,N_4068);
nor U4164 (N_4164,N_4087,N_4026);
nor U4165 (N_4165,N_4099,N_4083);
nand U4166 (N_4166,N_4029,N_4011);
or U4167 (N_4167,N_4040,N_4047);
xor U4168 (N_4168,N_4082,N_4015);
and U4169 (N_4169,N_4055,N_4040);
and U4170 (N_4170,N_4067,N_4004);
nand U4171 (N_4171,N_4051,N_4061);
nor U4172 (N_4172,N_4009,N_4036);
nand U4173 (N_4173,N_4097,N_4033);
xor U4174 (N_4174,N_4043,N_4044);
and U4175 (N_4175,N_4021,N_4056);
nor U4176 (N_4176,N_4080,N_4091);
nor U4177 (N_4177,N_4027,N_4019);
xnor U4178 (N_4178,N_4002,N_4057);
and U4179 (N_4179,N_4048,N_4008);
nor U4180 (N_4180,N_4081,N_4091);
nor U4181 (N_4181,N_4048,N_4080);
nand U4182 (N_4182,N_4043,N_4094);
or U4183 (N_4183,N_4006,N_4088);
and U4184 (N_4184,N_4009,N_4019);
nand U4185 (N_4185,N_4086,N_4019);
nor U4186 (N_4186,N_4038,N_4072);
or U4187 (N_4187,N_4074,N_4047);
nand U4188 (N_4188,N_4097,N_4028);
and U4189 (N_4189,N_4001,N_4073);
or U4190 (N_4190,N_4018,N_4098);
and U4191 (N_4191,N_4062,N_4043);
or U4192 (N_4192,N_4062,N_4019);
or U4193 (N_4193,N_4021,N_4070);
and U4194 (N_4194,N_4027,N_4005);
xnor U4195 (N_4195,N_4053,N_4016);
xor U4196 (N_4196,N_4031,N_4018);
xor U4197 (N_4197,N_4085,N_4019);
nor U4198 (N_4198,N_4088,N_4062);
nand U4199 (N_4199,N_4038,N_4050);
nor U4200 (N_4200,N_4139,N_4107);
xnor U4201 (N_4201,N_4137,N_4145);
or U4202 (N_4202,N_4163,N_4160);
xor U4203 (N_4203,N_4136,N_4186);
nor U4204 (N_4204,N_4164,N_4184);
and U4205 (N_4205,N_4121,N_4115);
or U4206 (N_4206,N_4191,N_4178);
nand U4207 (N_4207,N_4124,N_4170);
nor U4208 (N_4208,N_4157,N_4106);
nand U4209 (N_4209,N_4150,N_4132);
and U4210 (N_4210,N_4140,N_4158);
nor U4211 (N_4211,N_4138,N_4126);
nor U4212 (N_4212,N_4189,N_4143);
nor U4213 (N_4213,N_4188,N_4176);
nand U4214 (N_4214,N_4125,N_4195);
nor U4215 (N_4215,N_4120,N_4154);
nand U4216 (N_4216,N_4182,N_4117);
and U4217 (N_4217,N_4172,N_4197);
xor U4218 (N_4218,N_4173,N_4190);
and U4219 (N_4219,N_4179,N_4165);
or U4220 (N_4220,N_4109,N_4131);
nand U4221 (N_4221,N_4100,N_4108);
nor U4222 (N_4222,N_4198,N_4133);
or U4223 (N_4223,N_4104,N_4159);
nand U4224 (N_4224,N_4185,N_4180);
xor U4225 (N_4225,N_4166,N_4141);
nor U4226 (N_4226,N_4114,N_4144);
and U4227 (N_4227,N_4128,N_4153);
and U4228 (N_4228,N_4127,N_4123);
and U4229 (N_4229,N_4101,N_4129);
nand U4230 (N_4230,N_4199,N_4167);
and U4231 (N_4231,N_4111,N_4102);
or U4232 (N_4232,N_4193,N_4156);
and U4233 (N_4233,N_4152,N_4113);
nand U4234 (N_4234,N_4119,N_4134);
nor U4235 (N_4235,N_4149,N_4171);
nor U4236 (N_4236,N_4155,N_4105);
or U4237 (N_4237,N_4196,N_4142);
nand U4238 (N_4238,N_4151,N_4116);
or U4239 (N_4239,N_4103,N_4181);
nand U4240 (N_4240,N_4130,N_4162);
nor U4241 (N_4241,N_4122,N_4147);
xor U4242 (N_4242,N_4175,N_4135);
and U4243 (N_4243,N_4148,N_4168);
and U4244 (N_4244,N_4177,N_4169);
and U4245 (N_4245,N_4183,N_4174);
xnor U4246 (N_4246,N_4192,N_4146);
nand U4247 (N_4247,N_4118,N_4112);
nand U4248 (N_4248,N_4187,N_4110);
nand U4249 (N_4249,N_4194,N_4161);
xnor U4250 (N_4250,N_4177,N_4168);
and U4251 (N_4251,N_4143,N_4159);
xnor U4252 (N_4252,N_4171,N_4173);
or U4253 (N_4253,N_4158,N_4193);
xnor U4254 (N_4254,N_4122,N_4153);
or U4255 (N_4255,N_4183,N_4166);
and U4256 (N_4256,N_4149,N_4196);
and U4257 (N_4257,N_4193,N_4163);
or U4258 (N_4258,N_4179,N_4180);
nand U4259 (N_4259,N_4199,N_4193);
nand U4260 (N_4260,N_4148,N_4175);
nor U4261 (N_4261,N_4164,N_4179);
nor U4262 (N_4262,N_4143,N_4114);
or U4263 (N_4263,N_4174,N_4147);
nor U4264 (N_4264,N_4122,N_4198);
nor U4265 (N_4265,N_4180,N_4188);
nor U4266 (N_4266,N_4175,N_4193);
xor U4267 (N_4267,N_4122,N_4170);
and U4268 (N_4268,N_4142,N_4101);
and U4269 (N_4269,N_4115,N_4186);
nand U4270 (N_4270,N_4183,N_4139);
nor U4271 (N_4271,N_4135,N_4150);
or U4272 (N_4272,N_4199,N_4140);
or U4273 (N_4273,N_4181,N_4171);
and U4274 (N_4274,N_4118,N_4185);
xnor U4275 (N_4275,N_4195,N_4114);
or U4276 (N_4276,N_4147,N_4157);
nor U4277 (N_4277,N_4189,N_4167);
xnor U4278 (N_4278,N_4175,N_4124);
and U4279 (N_4279,N_4166,N_4152);
nor U4280 (N_4280,N_4155,N_4191);
nor U4281 (N_4281,N_4162,N_4167);
or U4282 (N_4282,N_4197,N_4114);
nor U4283 (N_4283,N_4126,N_4193);
nand U4284 (N_4284,N_4157,N_4137);
or U4285 (N_4285,N_4129,N_4109);
and U4286 (N_4286,N_4181,N_4175);
and U4287 (N_4287,N_4108,N_4178);
nor U4288 (N_4288,N_4160,N_4113);
or U4289 (N_4289,N_4135,N_4120);
or U4290 (N_4290,N_4157,N_4154);
or U4291 (N_4291,N_4111,N_4176);
or U4292 (N_4292,N_4186,N_4108);
nand U4293 (N_4293,N_4159,N_4174);
and U4294 (N_4294,N_4106,N_4156);
nor U4295 (N_4295,N_4143,N_4146);
xor U4296 (N_4296,N_4132,N_4169);
and U4297 (N_4297,N_4160,N_4102);
or U4298 (N_4298,N_4183,N_4165);
nor U4299 (N_4299,N_4144,N_4124);
and U4300 (N_4300,N_4289,N_4284);
and U4301 (N_4301,N_4209,N_4249);
nand U4302 (N_4302,N_4272,N_4220);
nand U4303 (N_4303,N_4237,N_4288);
and U4304 (N_4304,N_4299,N_4269);
nand U4305 (N_4305,N_4265,N_4231);
xor U4306 (N_4306,N_4287,N_4222);
nor U4307 (N_4307,N_4219,N_4238);
nand U4308 (N_4308,N_4282,N_4201);
xnor U4309 (N_4309,N_4273,N_4202);
or U4310 (N_4310,N_4240,N_4295);
nand U4311 (N_4311,N_4258,N_4217);
and U4312 (N_4312,N_4277,N_4234);
nand U4313 (N_4313,N_4216,N_4276);
or U4314 (N_4314,N_4256,N_4211);
nor U4315 (N_4315,N_4253,N_4227);
nand U4316 (N_4316,N_4260,N_4248);
nor U4317 (N_4317,N_4278,N_4213);
nand U4318 (N_4318,N_4228,N_4212);
xnor U4319 (N_4319,N_4236,N_4210);
xor U4320 (N_4320,N_4298,N_4233);
nand U4321 (N_4321,N_4266,N_4244);
nor U4322 (N_4322,N_4224,N_4291);
or U4323 (N_4323,N_4251,N_4286);
nand U4324 (N_4324,N_4207,N_4208);
nand U4325 (N_4325,N_4221,N_4200);
nor U4326 (N_4326,N_4206,N_4270);
nor U4327 (N_4327,N_4232,N_4205);
nor U4328 (N_4328,N_4297,N_4274);
or U4329 (N_4329,N_4241,N_4242);
nor U4330 (N_4330,N_4243,N_4215);
xor U4331 (N_4331,N_4226,N_4280);
and U4332 (N_4332,N_4271,N_4261);
and U4333 (N_4333,N_4294,N_4262);
nor U4334 (N_4334,N_4225,N_4263);
nand U4335 (N_4335,N_4259,N_4204);
xnor U4336 (N_4336,N_4252,N_4292);
or U4337 (N_4337,N_4246,N_4293);
xnor U4338 (N_4338,N_4285,N_4296);
or U4339 (N_4339,N_4267,N_4275);
nor U4340 (N_4340,N_4247,N_4214);
nand U4341 (N_4341,N_4250,N_4268);
and U4342 (N_4342,N_4230,N_4254);
and U4343 (N_4343,N_4290,N_4235);
or U4344 (N_4344,N_4281,N_4255);
xnor U4345 (N_4345,N_4218,N_4203);
nor U4346 (N_4346,N_4239,N_4283);
and U4347 (N_4347,N_4229,N_4264);
nor U4348 (N_4348,N_4257,N_4223);
or U4349 (N_4349,N_4245,N_4279);
xor U4350 (N_4350,N_4242,N_4274);
or U4351 (N_4351,N_4277,N_4226);
nand U4352 (N_4352,N_4278,N_4206);
nand U4353 (N_4353,N_4260,N_4289);
and U4354 (N_4354,N_4260,N_4296);
or U4355 (N_4355,N_4275,N_4282);
xnor U4356 (N_4356,N_4241,N_4270);
nand U4357 (N_4357,N_4237,N_4245);
nand U4358 (N_4358,N_4217,N_4210);
or U4359 (N_4359,N_4217,N_4276);
nand U4360 (N_4360,N_4205,N_4231);
or U4361 (N_4361,N_4294,N_4200);
and U4362 (N_4362,N_4258,N_4235);
nor U4363 (N_4363,N_4298,N_4277);
nand U4364 (N_4364,N_4273,N_4245);
nor U4365 (N_4365,N_4241,N_4244);
nand U4366 (N_4366,N_4205,N_4212);
or U4367 (N_4367,N_4262,N_4236);
nor U4368 (N_4368,N_4213,N_4281);
nor U4369 (N_4369,N_4246,N_4271);
xor U4370 (N_4370,N_4211,N_4204);
or U4371 (N_4371,N_4280,N_4242);
nor U4372 (N_4372,N_4227,N_4225);
nor U4373 (N_4373,N_4239,N_4284);
and U4374 (N_4374,N_4292,N_4248);
nor U4375 (N_4375,N_4274,N_4265);
nor U4376 (N_4376,N_4272,N_4226);
or U4377 (N_4377,N_4221,N_4261);
xor U4378 (N_4378,N_4276,N_4270);
nor U4379 (N_4379,N_4287,N_4200);
xor U4380 (N_4380,N_4228,N_4257);
nand U4381 (N_4381,N_4219,N_4239);
and U4382 (N_4382,N_4289,N_4228);
xor U4383 (N_4383,N_4294,N_4257);
nor U4384 (N_4384,N_4240,N_4237);
nor U4385 (N_4385,N_4231,N_4290);
xnor U4386 (N_4386,N_4251,N_4262);
xnor U4387 (N_4387,N_4257,N_4244);
or U4388 (N_4388,N_4215,N_4229);
and U4389 (N_4389,N_4298,N_4240);
nand U4390 (N_4390,N_4294,N_4243);
and U4391 (N_4391,N_4289,N_4285);
or U4392 (N_4392,N_4296,N_4268);
xor U4393 (N_4393,N_4291,N_4221);
nor U4394 (N_4394,N_4251,N_4276);
nor U4395 (N_4395,N_4244,N_4233);
nand U4396 (N_4396,N_4242,N_4227);
nand U4397 (N_4397,N_4274,N_4211);
and U4398 (N_4398,N_4293,N_4206);
nand U4399 (N_4399,N_4266,N_4285);
and U4400 (N_4400,N_4302,N_4324);
nand U4401 (N_4401,N_4303,N_4333);
nand U4402 (N_4402,N_4336,N_4364);
nand U4403 (N_4403,N_4323,N_4371);
and U4404 (N_4404,N_4389,N_4308);
nor U4405 (N_4405,N_4376,N_4366);
and U4406 (N_4406,N_4352,N_4317);
xnor U4407 (N_4407,N_4332,N_4343);
nor U4408 (N_4408,N_4397,N_4355);
or U4409 (N_4409,N_4348,N_4320);
nor U4410 (N_4410,N_4318,N_4354);
or U4411 (N_4411,N_4313,N_4375);
nand U4412 (N_4412,N_4382,N_4329);
xor U4413 (N_4413,N_4306,N_4351);
and U4414 (N_4414,N_4307,N_4331);
or U4415 (N_4415,N_4368,N_4315);
nand U4416 (N_4416,N_4321,N_4350);
nor U4417 (N_4417,N_4305,N_4345);
and U4418 (N_4418,N_4378,N_4353);
and U4419 (N_4419,N_4398,N_4341);
nor U4420 (N_4420,N_4328,N_4349);
nand U4421 (N_4421,N_4370,N_4386);
or U4422 (N_4422,N_4337,N_4340);
xor U4423 (N_4423,N_4361,N_4309);
and U4424 (N_4424,N_4338,N_4393);
nor U4425 (N_4425,N_4322,N_4396);
nand U4426 (N_4426,N_4316,N_4356);
or U4427 (N_4427,N_4374,N_4377);
xor U4428 (N_4428,N_4373,N_4325);
and U4429 (N_4429,N_4384,N_4330);
or U4430 (N_4430,N_4358,N_4387);
or U4431 (N_4431,N_4326,N_4342);
nor U4432 (N_4432,N_4380,N_4312);
and U4433 (N_4433,N_4304,N_4347);
and U4434 (N_4434,N_4327,N_4311);
or U4435 (N_4435,N_4319,N_4394);
xnor U4436 (N_4436,N_4392,N_4391);
nor U4437 (N_4437,N_4362,N_4372);
or U4438 (N_4438,N_4367,N_4381);
and U4439 (N_4439,N_4388,N_4385);
and U4440 (N_4440,N_4360,N_4357);
or U4441 (N_4441,N_4346,N_4310);
or U4442 (N_4442,N_4369,N_4359);
nor U4443 (N_4443,N_4300,N_4363);
nor U4444 (N_4444,N_4335,N_4379);
nand U4445 (N_4445,N_4334,N_4390);
and U4446 (N_4446,N_4301,N_4344);
nand U4447 (N_4447,N_4383,N_4365);
or U4448 (N_4448,N_4339,N_4399);
and U4449 (N_4449,N_4314,N_4395);
nor U4450 (N_4450,N_4335,N_4343);
nand U4451 (N_4451,N_4361,N_4383);
xor U4452 (N_4452,N_4381,N_4314);
xnor U4453 (N_4453,N_4335,N_4324);
and U4454 (N_4454,N_4339,N_4353);
and U4455 (N_4455,N_4336,N_4391);
xnor U4456 (N_4456,N_4328,N_4319);
xnor U4457 (N_4457,N_4324,N_4323);
or U4458 (N_4458,N_4311,N_4315);
xor U4459 (N_4459,N_4378,N_4315);
or U4460 (N_4460,N_4300,N_4313);
or U4461 (N_4461,N_4344,N_4345);
xor U4462 (N_4462,N_4372,N_4369);
xor U4463 (N_4463,N_4396,N_4369);
or U4464 (N_4464,N_4390,N_4346);
or U4465 (N_4465,N_4375,N_4344);
nor U4466 (N_4466,N_4322,N_4312);
or U4467 (N_4467,N_4342,N_4316);
nor U4468 (N_4468,N_4392,N_4306);
xor U4469 (N_4469,N_4305,N_4350);
xor U4470 (N_4470,N_4347,N_4398);
and U4471 (N_4471,N_4301,N_4388);
and U4472 (N_4472,N_4362,N_4300);
and U4473 (N_4473,N_4389,N_4303);
xor U4474 (N_4474,N_4308,N_4338);
nor U4475 (N_4475,N_4320,N_4363);
and U4476 (N_4476,N_4326,N_4339);
xor U4477 (N_4477,N_4333,N_4321);
nand U4478 (N_4478,N_4332,N_4315);
nand U4479 (N_4479,N_4354,N_4324);
or U4480 (N_4480,N_4327,N_4324);
or U4481 (N_4481,N_4389,N_4383);
nand U4482 (N_4482,N_4395,N_4363);
and U4483 (N_4483,N_4377,N_4380);
and U4484 (N_4484,N_4342,N_4387);
nor U4485 (N_4485,N_4366,N_4337);
nand U4486 (N_4486,N_4371,N_4361);
nand U4487 (N_4487,N_4391,N_4360);
or U4488 (N_4488,N_4337,N_4345);
nor U4489 (N_4489,N_4344,N_4335);
or U4490 (N_4490,N_4316,N_4300);
nor U4491 (N_4491,N_4391,N_4335);
nor U4492 (N_4492,N_4327,N_4332);
and U4493 (N_4493,N_4340,N_4341);
or U4494 (N_4494,N_4332,N_4394);
nand U4495 (N_4495,N_4332,N_4388);
or U4496 (N_4496,N_4397,N_4313);
nand U4497 (N_4497,N_4387,N_4317);
nand U4498 (N_4498,N_4364,N_4398);
xnor U4499 (N_4499,N_4376,N_4352);
or U4500 (N_4500,N_4480,N_4428);
nor U4501 (N_4501,N_4445,N_4446);
xor U4502 (N_4502,N_4458,N_4450);
or U4503 (N_4503,N_4481,N_4433);
nand U4504 (N_4504,N_4464,N_4484);
and U4505 (N_4505,N_4494,N_4475);
nor U4506 (N_4506,N_4460,N_4442);
or U4507 (N_4507,N_4470,N_4430);
and U4508 (N_4508,N_4491,N_4496);
and U4509 (N_4509,N_4474,N_4472);
xor U4510 (N_4510,N_4449,N_4465);
or U4511 (N_4511,N_4463,N_4486);
nand U4512 (N_4512,N_4416,N_4462);
nor U4513 (N_4513,N_4448,N_4498);
and U4514 (N_4514,N_4432,N_4437);
xor U4515 (N_4515,N_4495,N_4400);
or U4516 (N_4516,N_4492,N_4473);
xnor U4517 (N_4517,N_4412,N_4439);
xor U4518 (N_4518,N_4434,N_4483);
nand U4519 (N_4519,N_4461,N_4485);
nor U4520 (N_4520,N_4443,N_4440);
and U4521 (N_4521,N_4468,N_4489);
nand U4522 (N_4522,N_4420,N_4493);
or U4523 (N_4523,N_4452,N_4431);
or U4524 (N_4524,N_4487,N_4424);
and U4525 (N_4525,N_4459,N_4438);
or U4526 (N_4526,N_4418,N_4411);
xnor U4527 (N_4527,N_4456,N_4415);
or U4528 (N_4528,N_4447,N_4401);
or U4529 (N_4529,N_4478,N_4423);
or U4530 (N_4530,N_4441,N_4409);
xor U4531 (N_4531,N_4451,N_4407);
xor U4532 (N_4532,N_4469,N_4467);
or U4533 (N_4533,N_4427,N_4414);
xor U4534 (N_4534,N_4406,N_4413);
nor U4535 (N_4535,N_4455,N_4405);
or U4536 (N_4536,N_4477,N_4476);
nor U4537 (N_4537,N_4403,N_4402);
and U4538 (N_4538,N_4466,N_4425);
or U4539 (N_4539,N_4421,N_4408);
xor U4540 (N_4540,N_4436,N_4419);
nand U4541 (N_4541,N_4429,N_4404);
or U4542 (N_4542,N_4457,N_4454);
nand U4543 (N_4543,N_4426,N_4497);
nor U4544 (N_4544,N_4488,N_4444);
or U4545 (N_4545,N_4422,N_4471);
nor U4546 (N_4546,N_4417,N_4453);
nor U4547 (N_4547,N_4479,N_4410);
xor U4548 (N_4548,N_4499,N_4435);
nand U4549 (N_4549,N_4490,N_4482);
and U4550 (N_4550,N_4415,N_4463);
or U4551 (N_4551,N_4421,N_4422);
xnor U4552 (N_4552,N_4480,N_4441);
and U4553 (N_4553,N_4408,N_4486);
nor U4554 (N_4554,N_4472,N_4441);
and U4555 (N_4555,N_4467,N_4416);
nor U4556 (N_4556,N_4451,N_4409);
nand U4557 (N_4557,N_4409,N_4499);
nor U4558 (N_4558,N_4481,N_4466);
xor U4559 (N_4559,N_4460,N_4477);
or U4560 (N_4560,N_4482,N_4408);
or U4561 (N_4561,N_4412,N_4478);
nor U4562 (N_4562,N_4422,N_4473);
and U4563 (N_4563,N_4443,N_4417);
nor U4564 (N_4564,N_4462,N_4489);
xor U4565 (N_4565,N_4454,N_4488);
nand U4566 (N_4566,N_4485,N_4426);
nor U4567 (N_4567,N_4486,N_4475);
xnor U4568 (N_4568,N_4492,N_4478);
and U4569 (N_4569,N_4482,N_4493);
nand U4570 (N_4570,N_4474,N_4434);
and U4571 (N_4571,N_4424,N_4483);
xnor U4572 (N_4572,N_4488,N_4401);
nor U4573 (N_4573,N_4426,N_4444);
or U4574 (N_4574,N_4423,N_4481);
or U4575 (N_4575,N_4434,N_4445);
and U4576 (N_4576,N_4485,N_4443);
xnor U4577 (N_4577,N_4498,N_4447);
or U4578 (N_4578,N_4429,N_4434);
and U4579 (N_4579,N_4470,N_4434);
nand U4580 (N_4580,N_4491,N_4402);
nor U4581 (N_4581,N_4465,N_4436);
and U4582 (N_4582,N_4453,N_4495);
nor U4583 (N_4583,N_4427,N_4493);
nor U4584 (N_4584,N_4433,N_4442);
or U4585 (N_4585,N_4433,N_4465);
xnor U4586 (N_4586,N_4468,N_4476);
nand U4587 (N_4587,N_4486,N_4433);
nor U4588 (N_4588,N_4407,N_4403);
and U4589 (N_4589,N_4488,N_4407);
or U4590 (N_4590,N_4428,N_4430);
and U4591 (N_4591,N_4437,N_4457);
xor U4592 (N_4592,N_4451,N_4491);
xor U4593 (N_4593,N_4421,N_4461);
nand U4594 (N_4594,N_4443,N_4469);
xor U4595 (N_4595,N_4442,N_4467);
nand U4596 (N_4596,N_4462,N_4402);
xnor U4597 (N_4597,N_4429,N_4492);
or U4598 (N_4598,N_4431,N_4477);
nor U4599 (N_4599,N_4431,N_4475);
nor U4600 (N_4600,N_4525,N_4515);
xor U4601 (N_4601,N_4594,N_4532);
or U4602 (N_4602,N_4531,N_4550);
xnor U4603 (N_4603,N_4506,N_4510);
or U4604 (N_4604,N_4545,N_4568);
nand U4605 (N_4605,N_4500,N_4556);
nor U4606 (N_4606,N_4570,N_4501);
xnor U4607 (N_4607,N_4599,N_4582);
or U4608 (N_4608,N_4520,N_4580);
nor U4609 (N_4609,N_4585,N_4551);
or U4610 (N_4610,N_4565,N_4535);
nand U4611 (N_4611,N_4575,N_4591);
xor U4612 (N_4612,N_4566,N_4597);
or U4613 (N_4613,N_4567,N_4559);
nand U4614 (N_4614,N_4543,N_4589);
nand U4615 (N_4615,N_4598,N_4564);
xor U4616 (N_4616,N_4562,N_4584);
and U4617 (N_4617,N_4523,N_4563);
xnor U4618 (N_4618,N_4513,N_4554);
or U4619 (N_4619,N_4504,N_4519);
and U4620 (N_4620,N_4524,N_4511);
or U4621 (N_4621,N_4507,N_4553);
or U4622 (N_4622,N_4546,N_4536);
nand U4623 (N_4623,N_4583,N_4505);
xor U4624 (N_4624,N_4561,N_4569);
nor U4625 (N_4625,N_4539,N_4541);
xnor U4626 (N_4626,N_4529,N_4538);
nand U4627 (N_4627,N_4558,N_4560);
nor U4628 (N_4628,N_4548,N_4527);
or U4629 (N_4629,N_4521,N_4512);
xor U4630 (N_4630,N_4576,N_4574);
nor U4631 (N_4631,N_4542,N_4537);
nand U4632 (N_4632,N_4593,N_4516);
xor U4633 (N_4633,N_4588,N_4572);
nor U4634 (N_4634,N_4573,N_4540);
or U4635 (N_4635,N_4552,N_4586);
nor U4636 (N_4636,N_4579,N_4581);
xnor U4637 (N_4637,N_4544,N_4555);
or U4638 (N_4638,N_4530,N_4508);
xor U4639 (N_4639,N_4514,N_4578);
nor U4640 (N_4640,N_4509,N_4557);
or U4641 (N_4641,N_4534,N_4528);
xor U4642 (N_4642,N_4502,N_4587);
nand U4643 (N_4643,N_4592,N_4518);
or U4644 (N_4644,N_4577,N_4517);
and U4645 (N_4645,N_4522,N_4503);
xnor U4646 (N_4646,N_4595,N_4549);
xor U4647 (N_4647,N_4590,N_4571);
xor U4648 (N_4648,N_4596,N_4526);
or U4649 (N_4649,N_4533,N_4547);
nor U4650 (N_4650,N_4533,N_4561);
xor U4651 (N_4651,N_4537,N_4501);
and U4652 (N_4652,N_4585,N_4508);
nor U4653 (N_4653,N_4567,N_4550);
xor U4654 (N_4654,N_4529,N_4586);
xnor U4655 (N_4655,N_4537,N_4583);
nand U4656 (N_4656,N_4508,N_4535);
nor U4657 (N_4657,N_4528,N_4571);
nor U4658 (N_4658,N_4586,N_4520);
nor U4659 (N_4659,N_4505,N_4556);
nor U4660 (N_4660,N_4559,N_4571);
xnor U4661 (N_4661,N_4594,N_4599);
and U4662 (N_4662,N_4504,N_4546);
and U4663 (N_4663,N_4587,N_4517);
xor U4664 (N_4664,N_4525,N_4537);
nor U4665 (N_4665,N_4506,N_4590);
nand U4666 (N_4666,N_4538,N_4599);
nor U4667 (N_4667,N_4554,N_4519);
and U4668 (N_4668,N_4542,N_4532);
or U4669 (N_4669,N_4548,N_4521);
or U4670 (N_4670,N_4551,N_4579);
nor U4671 (N_4671,N_4502,N_4549);
or U4672 (N_4672,N_4533,N_4538);
or U4673 (N_4673,N_4537,N_4503);
or U4674 (N_4674,N_4554,N_4551);
xnor U4675 (N_4675,N_4517,N_4596);
xor U4676 (N_4676,N_4520,N_4518);
and U4677 (N_4677,N_4500,N_4559);
and U4678 (N_4678,N_4566,N_4560);
xor U4679 (N_4679,N_4519,N_4563);
or U4680 (N_4680,N_4557,N_4550);
and U4681 (N_4681,N_4586,N_4580);
nand U4682 (N_4682,N_4557,N_4523);
or U4683 (N_4683,N_4517,N_4533);
xnor U4684 (N_4684,N_4523,N_4502);
nand U4685 (N_4685,N_4508,N_4586);
nand U4686 (N_4686,N_4571,N_4525);
nand U4687 (N_4687,N_4515,N_4599);
xnor U4688 (N_4688,N_4519,N_4580);
xnor U4689 (N_4689,N_4539,N_4519);
and U4690 (N_4690,N_4575,N_4577);
nor U4691 (N_4691,N_4539,N_4544);
nor U4692 (N_4692,N_4500,N_4591);
and U4693 (N_4693,N_4556,N_4589);
or U4694 (N_4694,N_4574,N_4571);
nand U4695 (N_4695,N_4503,N_4526);
xnor U4696 (N_4696,N_4589,N_4505);
or U4697 (N_4697,N_4557,N_4581);
or U4698 (N_4698,N_4558,N_4579);
nand U4699 (N_4699,N_4557,N_4522);
nor U4700 (N_4700,N_4651,N_4653);
nor U4701 (N_4701,N_4673,N_4655);
and U4702 (N_4702,N_4641,N_4686);
and U4703 (N_4703,N_4642,N_4603);
nand U4704 (N_4704,N_4637,N_4645);
and U4705 (N_4705,N_4665,N_4654);
or U4706 (N_4706,N_4685,N_4663);
or U4707 (N_4707,N_4695,N_4696);
or U4708 (N_4708,N_4676,N_4616);
nor U4709 (N_4709,N_4648,N_4638);
xnor U4710 (N_4710,N_4602,N_4659);
xor U4711 (N_4711,N_4631,N_4680);
xnor U4712 (N_4712,N_4687,N_4683);
and U4713 (N_4713,N_4636,N_4626);
nor U4714 (N_4714,N_4620,N_4605);
and U4715 (N_4715,N_4691,N_4618);
nand U4716 (N_4716,N_4647,N_4632);
nor U4717 (N_4717,N_4617,N_4610);
or U4718 (N_4718,N_4657,N_4698);
nand U4719 (N_4719,N_4664,N_4639);
xor U4720 (N_4720,N_4604,N_4677);
nand U4721 (N_4721,N_4660,N_4678);
or U4722 (N_4722,N_4633,N_4615);
xnor U4723 (N_4723,N_4611,N_4608);
xnor U4724 (N_4724,N_4670,N_4630);
nand U4725 (N_4725,N_4697,N_4601);
and U4726 (N_4726,N_4606,N_4684);
nand U4727 (N_4727,N_4643,N_4609);
nand U4728 (N_4728,N_4693,N_4646);
nor U4729 (N_4729,N_4694,N_4672);
xnor U4730 (N_4730,N_4689,N_4649);
or U4731 (N_4731,N_4668,N_4635);
and U4732 (N_4732,N_4644,N_4640);
xor U4733 (N_4733,N_4671,N_4625);
xor U4734 (N_4734,N_4692,N_4669);
and U4735 (N_4735,N_4622,N_4662);
xnor U4736 (N_4736,N_4607,N_4675);
xor U4737 (N_4737,N_4628,N_4679);
or U4738 (N_4738,N_4612,N_4699);
or U4739 (N_4739,N_4627,N_4656);
or U4740 (N_4740,N_4674,N_4621);
or U4741 (N_4741,N_4614,N_4600);
nand U4742 (N_4742,N_4661,N_4623);
nor U4743 (N_4743,N_4619,N_4688);
and U4744 (N_4744,N_4629,N_4650);
nand U4745 (N_4745,N_4613,N_4624);
or U4746 (N_4746,N_4652,N_4667);
and U4747 (N_4747,N_4634,N_4690);
and U4748 (N_4748,N_4681,N_4658);
xnor U4749 (N_4749,N_4666,N_4682);
nor U4750 (N_4750,N_4627,N_4603);
xor U4751 (N_4751,N_4600,N_4658);
xnor U4752 (N_4752,N_4657,N_4623);
nand U4753 (N_4753,N_4606,N_4628);
nand U4754 (N_4754,N_4670,N_4616);
nand U4755 (N_4755,N_4686,N_4629);
nand U4756 (N_4756,N_4608,N_4635);
xor U4757 (N_4757,N_4656,N_4688);
xnor U4758 (N_4758,N_4685,N_4647);
xnor U4759 (N_4759,N_4657,N_4667);
nand U4760 (N_4760,N_4623,N_4659);
xnor U4761 (N_4761,N_4651,N_4696);
nor U4762 (N_4762,N_4635,N_4679);
or U4763 (N_4763,N_4642,N_4672);
nor U4764 (N_4764,N_4688,N_4666);
nor U4765 (N_4765,N_4660,N_4689);
nand U4766 (N_4766,N_4674,N_4629);
xor U4767 (N_4767,N_4646,N_4670);
xor U4768 (N_4768,N_4654,N_4634);
nor U4769 (N_4769,N_4667,N_4622);
or U4770 (N_4770,N_4614,N_4663);
and U4771 (N_4771,N_4656,N_4648);
nor U4772 (N_4772,N_4616,N_4673);
nand U4773 (N_4773,N_4653,N_4656);
nand U4774 (N_4774,N_4614,N_4628);
nor U4775 (N_4775,N_4694,N_4607);
or U4776 (N_4776,N_4668,N_4682);
nor U4777 (N_4777,N_4604,N_4607);
nor U4778 (N_4778,N_4636,N_4630);
and U4779 (N_4779,N_4647,N_4680);
nor U4780 (N_4780,N_4612,N_4608);
nand U4781 (N_4781,N_4685,N_4677);
or U4782 (N_4782,N_4644,N_4641);
xnor U4783 (N_4783,N_4636,N_4648);
nand U4784 (N_4784,N_4635,N_4666);
and U4785 (N_4785,N_4640,N_4611);
nor U4786 (N_4786,N_4615,N_4647);
nor U4787 (N_4787,N_4601,N_4600);
nor U4788 (N_4788,N_4617,N_4687);
nor U4789 (N_4789,N_4656,N_4678);
xor U4790 (N_4790,N_4685,N_4600);
xor U4791 (N_4791,N_4653,N_4633);
xor U4792 (N_4792,N_4628,N_4681);
nand U4793 (N_4793,N_4651,N_4602);
nand U4794 (N_4794,N_4687,N_4659);
or U4795 (N_4795,N_4637,N_4622);
xor U4796 (N_4796,N_4606,N_4685);
xnor U4797 (N_4797,N_4653,N_4607);
nor U4798 (N_4798,N_4664,N_4698);
xor U4799 (N_4799,N_4667,N_4691);
nand U4800 (N_4800,N_4724,N_4737);
nor U4801 (N_4801,N_4735,N_4779);
and U4802 (N_4802,N_4716,N_4715);
and U4803 (N_4803,N_4750,N_4767);
nor U4804 (N_4804,N_4706,N_4705);
and U4805 (N_4805,N_4728,N_4784);
or U4806 (N_4806,N_4701,N_4703);
nor U4807 (N_4807,N_4773,N_4792);
or U4808 (N_4808,N_4789,N_4770);
and U4809 (N_4809,N_4730,N_4748);
nand U4810 (N_4810,N_4726,N_4761);
or U4811 (N_4811,N_4788,N_4714);
and U4812 (N_4812,N_4700,N_4744);
xor U4813 (N_4813,N_4711,N_4790);
nand U4814 (N_4814,N_4783,N_4739);
or U4815 (N_4815,N_4754,N_4766);
and U4816 (N_4816,N_4787,N_4719);
nand U4817 (N_4817,N_4718,N_4702);
and U4818 (N_4818,N_4776,N_4762);
and U4819 (N_4819,N_4771,N_4743);
and U4820 (N_4820,N_4785,N_4778);
and U4821 (N_4821,N_4791,N_4768);
and U4822 (N_4822,N_4759,N_4774);
nand U4823 (N_4823,N_4721,N_4745);
or U4824 (N_4824,N_4738,N_4749);
xor U4825 (N_4825,N_4707,N_4758);
xor U4826 (N_4826,N_4764,N_4712);
nand U4827 (N_4827,N_4799,N_4713);
nor U4828 (N_4828,N_4732,N_4710);
or U4829 (N_4829,N_4765,N_4751);
nor U4830 (N_4830,N_4777,N_4775);
nor U4831 (N_4831,N_4746,N_4722);
nand U4832 (N_4832,N_4793,N_4752);
or U4833 (N_4833,N_4796,N_4723);
nor U4834 (N_4834,N_4772,N_4786);
nand U4835 (N_4835,N_4740,N_4720);
and U4836 (N_4836,N_4780,N_4727);
nor U4837 (N_4837,N_4797,N_4755);
nand U4838 (N_4838,N_4763,N_4734);
xnor U4839 (N_4839,N_4742,N_4725);
and U4840 (N_4840,N_4753,N_4708);
and U4841 (N_4841,N_4731,N_4704);
or U4842 (N_4842,N_4747,N_4717);
xnor U4843 (N_4843,N_4782,N_4795);
and U4844 (N_4844,N_4741,N_4769);
xnor U4845 (N_4845,N_4756,N_4733);
or U4846 (N_4846,N_4798,N_4729);
and U4847 (N_4847,N_4736,N_4757);
and U4848 (N_4848,N_4709,N_4781);
xor U4849 (N_4849,N_4760,N_4794);
nor U4850 (N_4850,N_4791,N_4798);
nor U4851 (N_4851,N_4712,N_4773);
nor U4852 (N_4852,N_4708,N_4796);
xnor U4853 (N_4853,N_4700,N_4751);
nor U4854 (N_4854,N_4775,N_4729);
and U4855 (N_4855,N_4761,N_4728);
and U4856 (N_4856,N_4776,N_4724);
or U4857 (N_4857,N_4715,N_4750);
xnor U4858 (N_4858,N_4744,N_4756);
nor U4859 (N_4859,N_4728,N_4786);
xnor U4860 (N_4860,N_4790,N_4754);
nor U4861 (N_4861,N_4784,N_4745);
and U4862 (N_4862,N_4744,N_4790);
or U4863 (N_4863,N_4763,N_4747);
xor U4864 (N_4864,N_4749,N_4793);
or U4865 (N_4865,N_4755,N_4747);
or U4866 (N_4866,N_4728,N_4705);
and U4867 (N_4867,N_4759,N_4744);
nor U4868 (N_4868,N_4720,N_4748);
nand U4869 (N_4869,N_4721,N_4706);
or U4870 (N_4870,N_4757,N_4763);
nor U4871 (N_4871,N_4746,N_4721);
xor U4872 (N_4872,N_4724,N_4741);
nor U4873 (N_4873,N_4709,N_4744);
or U4874 (N_4874,N_4747,N_4725);
xor U4875 (N_4875,N_4789,N_4787);
or U4876 (N_4876,N_4714,N_4777);
xor U4877 (N_4877,N_4727,N_4713);
nand U4878 (N_4878,N_4761,N_4720);
and U4879 (N_4879,N_4755,N_4792);
or U4880 (N_4880,N_4783,N_4735);
nand U4881 (N_4881,N_4703,N_4700);
xnor U4882 (N_4882,N_4769,N_4756);
or U4883 (N_4883,N_4794,N_4739);
or U4884 (N_4884,N_4745,N_4737);
or U4885 (N_4885,N_4794,N_4780);
nand U4886 (N_4886,N_4725,N_4775);
or U4887 (N_4887,N_4702,N_4777);
nor U4888 (N_4888,N_4752,N_4740);
nor U4889 (N_4889,N_4769,N_4726);
or U4890 (N_4890,N_4754,N_4707);
or U4891 (N_4891,N_4714,N_4740);
and U4892 (N_4892,N_4717,N_4712);
nor U4893 (N_4893,N_4746,N_4799);
xor U4894 (N_4894,N_4727,N_4733);
and U4895 (N_4895,N_4716,N_4769);
nand U4896 (N_4896,N_4747,N_4744);
xor U4897 (N_4897,N_4794,N_4776);
xor U4898 (N_4898,N_4725,N_4735);
nor U4899 (N_4899,N_4737,N_4719);
or U4900 (N_4900,N_4843,N_4800);
nand U4901 (N_4901,N_4879,N_4822);
nand U4902 (N_4902,N_4827,N_4808);
xnor U4903 (N_4903,N_4845,N_4841);
and U4904 (N_4904,N_4807,N_4844);
or U4905 (N_4905,N_4878,N_4893);
xnor U4906 (N_4906,N_4890,N_4829);
nand U4907 (N_4907,N_4860,N_4864);
xor U4908 (N_4908,N_4828,N_4872);
nor U4909 (N_4909,N_4820,N_4876);
nor U4910 (N_4910,N_4850,N_4838);
nor U4911 (N_4911,N_4881,N_4870);
or U4912 (N_4912,N_4839,N_4812);
and U4913 (N_4913,N_4896,N_4892);
or U4914 (N_4914,N_4867,N_4847);
nand U4915 (N_4915,N_4809,N_4819);
xor U4916 (N_4916,N_4857,N_4817);
nand U4917 (N_4917,N_4855,N_4802);
xor U4918 (N_4918,N_4814,N_4891);
xnor U4919 (N_4919,N_4883,N_4889);
xnor U4920 (N_4920,N_4853,N_4863);
and U4921 (N_4921,N_4842,N_4804);
nor U4922 (N_4922,N_4859,N_4833);
or U4923 (N_4923,N_4869,N_4813);
xnor U4924 (N_4924,N_4811,N_4810);
xor U4925 (N_4925,N_4803,N_4873);
and U4926 (N_4926,N_4825,N_4880);
or U4927 (N_4927,N_4801,N_4806);
and U4928 (N_4928,N_4815,N_4836);
xnor U4929 (N_4929,N_4885,N_4898);
nor U4930 (N_4930,N_4824,N_4852);
xor U4931 (N_4931,N_4899,N_4866);
and U4932 (N_4932,N_4816,N_4862);
xor U4933 (N_4933,N_4830,N_4871);
nand U4934 (N_4934,N_4888,N_4851);
or U4935 (N_4935,N_4877,N_4856);
nand U4936 (N_4936,N_4831,N_4832);
xor U4937 (N_4937,N_4874,N_4840);
nor U4938 (N_4938,N_4868,N_4887);
or U4939 (N_4939,N_4886,N_4826);
and U4940 (N_4940,N_4835,N_4834);
nor U4941 (N_4941,N_4894,N_4882);
xnor U4942 (N_4942,N_4849,N_4823);
xor U4943 (N_4943,N_4805,N_4865);
nor U4944 (N_4944,N_4875,N_4821);
xnor U4945 (N_4945,N_4858,N_4895);
or U4946 (N_4946,N_4854,N_4846);
nand U4947 (N_4947,N_4848,N_4897);
xnor U4948 (N_4948,N_4818,N_4837);
or U4949 (N_4949,N_4861,N_4884);
and U4950 (N_4950,N_4801,N_4850);
nor U4951 (N_4951,N_4827,N_4825);
and U4952 (N_4952,N_4803,N_4888);
nor U4953 (N_4953,N_4847,N_4862);
nand U4954 (N_4954,N_4808,N_4847);
nand U4955 (N_4955,N_4865,N_4880);
nand U4956 (N_4956,N_4821,N_4884);
or U4957 (N_4957,N_4892,N_4870);
nand U4958 (N_4958,N_4823,N_4876);
nor U4959 (N_4959,N_4812,N_4885);
and U4960 (N_4960,N_4861,N_4854);
xnor U4961 (N_4961,N_4873,N_4817);
xnor U4962 (N_4962,N_4818,N_4865);
nor U4963 (N_4963,N_4880,N_4889);
or U4964 (N_4964,N_4844,N_4873);
xnor U4965 (N_4965,N_4866,N_4820);
nor U4966 (N_4966,N_4898,N_4894);
or U4967 (N_4967,N_4896,N_4875);
nor U4968 (N_4968,N_4809,N_4829);
nand U4969 (N_4969,N_4863,N_4832);
and U4970 (N_4970,N_4846,N_4894);
or U4971 (N_4971,N_4852,N_4830);
nor U4972 (N_4972,N_4864,N_4816);
xnor U4973 (N_4973,N_4818,N_4853);
and U4974 (N_4974,N_4846,N_4825);
nand U4975 (N_4975,N_4823,N_4847);
and U4976 (N_4976,N_4813,N_4810);
nor U4977 (N_4977,N_4889,N_4810);
or U4978 (N_4978,N_4811,N_4884);
and U4979 (N_4979,N_4810,N_4877);
and U4980 (N_4980,N_4829,N_4875);
and U4981 (N_4981,N_4849,N_4807);
or U4982 (N_4982,N_4832,N_4817);
or U4983 (N_4983,N_4847,N_4869);
xor U4984 (N_4984,N_4841,N_4811);
nand U4985 (N_4985,N_4854,N_4879);
nand U4986 (N_4986,N_4807,N_4821);
and U4987 (N_4987,N_4858,N_4818);
or U4988 (N_4988,N_4856,N_4814);
or U4989 (N_4989,N_4807,N_4805);
xnor U4990 (N_4990,N_4845,N_4843);
and U4991 (N_4991,N_4814,N_4828);
nor U4992 (N_4992,N_4827,N_4838);
or U4993 (N_4993,N_4861,N_4853);
nor U4994 (N_4994,N_4817,N_4833);
and U4995 (N_4995,N_4862,N_4878);
xnor U4996 (N_4996,N_4831,N_4836);
nand U4997 (N_4997,N_4826,N_4853);
or U4998 (N_4998,N_4864,N_4834);
nor U4999 (N_4999,N_4815,N_4866);
and U5000 (N_5000,N_4994,N_4944);
xnor U5001 (N_5001,N_4979,N_4951);
or U5002 (N_5002,N_4912,N_4959);
nor U5003 (N_5003,N_4972,N_4992);
and U5004 (N_5004,N_4999,N_4901);
or U5005 (N_5005,N_4995,N_4993);
or U5006 (N_5006,N_4996,N_4903);
nand U5007 (N_5007,N_4920,N_4905);
or U5008 (N_5008,N_4960,N_4990);
nor U5009 (N_5009,N_4982,N_4984);
nand U5010 (N_5010,N_4991,N_4954);
or U5011 (N_5011,N_4987,N_4929);
nand U5012 (N_5012,N_4986,N_4919);
or U5013 (N_5013,N_4936,N_4989);
or U5014 (N_5014,N_4997,N_4956);
xnor U5015 (N_5015,N_4930,N_4917);
and U5016 (N_5016,N_4964,N_4914);
nor U5017 (N_5017,N_4934,N_4910);
nor U5018 (N_5018,N_4950,N_4907);
nor U5019 (N_5019,N_4943,N_4967);
nor U5020 (N_5020,N_4941,N_4922);
nor U5021 (N_5021,N_4970,N_4916);
or U5022 (N_5022,N_4980,N_4949);
and U5023 (N_5023,N_4939,N_4966);
nor U5024 (N_5024,N_4942,N_4975);
or U5025 (N_5025,N_4958,N_4974);
or U5026 (N_5026,N_4981,N_4918);
nor U5027 (N_5027,N_4969,N_4926);
nand U5028 (N_5028,N_4945,N_4953);
nand U5029 (N_5029,N_4940,N_4955);
or U5030 (N_5030,N_4937,N_4957);
and U5031 (N_5031,N_4947,N_4978);
nand U5032 (N_5032,N_4988,N_4977);
nor U5033 (N_5033,N_4925,N_4931);
xnor U5034 (N_5034,N_4928,N_4924);
nor U5035 (N_5035,N_4973,N_4985);
and U5036 (N_5036,N_4952,N_4915);
or U5037 (N_5037,N_4961,N_4921);
xnor U5038 (N_5038,N_4983,N_4998);
nor U5039 (N_5039,N_4913,N_4976);
and U5040 (N_5040,N_4935,N_4904);
and U5041 (N_5041,N_4948,N_4909);
xnor U5042 (N_5042,N_4968,N_4946);
xor U5043 (N_5043,N_4900,N_4932);
nand U5044 (N_5044,N_4971,N_4965);
nor U5045 (N_5045,N_4906,N_4927);
xnor U5046 (N_5046,N_4963,N_4933);
xnor U5047 (N_5047,N_4902,N_4938);
xnor U5048 (N_5048,N_4923,N_4908);
nand U5049 (N_5049,N_4962,N_4911);
nor U5050 (N_5050,N_4950,N_4972);
or U5051 (N_5051,N_4963,N_4971);
nand U5052 (N_5052,N_4901,N_4915);
xor U5053 (N_5053,N_4960,N_4982);
and U5054 (N_5054,N_4974,N_4948);
xor U5055 (N_5055,N_4979,N_4956);
nor U5056 (N_5056,N_4924,N_4949);
nand U5057 (N_5057,N_4996,N_4933);
nand U5058 (N_5058,N_4983,N_4985);
nor U5059 (N_5059,N_4932,N_4929);
and U5060 (N_5060,N_4969,N_4983);
nor U5061 (N_5061,N_4961,N_4963);
and U5062 (N_5062,N_4966,N_4957);
nor U5063 (N_5063,N_4959,N_4913);
nor U5064 (N_5064,N_4981,N_4973);
or U5065 (N_5065,N_4967,N_4927);
nand U5066 (N_5066,N_4952,N_4973);
or U5067 (N_5067,N_4989,N_4990);
or U5068 (N_5068,N_4922,N_4968);
or U5069 (N_5069,N_4959,N_4991);
nand U5070 (N_5070,N_4968,N_4989);
nor U5071 (N_5071,N_4910,N_4904);
and U5072 (N_5072,N_4988,N_4929);
or U5073 (N_5073,N_4939,N_4931);
and U5074 (N_5074,N_4964,N_4975);
xnor U5075 (N_5075,N_4927,N_4988);
nand U5076 (N_5076,N_4991,N_4946);
and U5077 (N_5077,N_4968,N_4945);
and U5078 (N_5078,N_4904,N_4924);
nor U5079 (N_5079,N_4917,N_4964);
nand U5080 (N_5080,N_4915,N_4958);
or U5081 (N_5081,N_4968,N_4908);
or U5082 (N_5082,N_4974,N_4936);
or U5083 (N_5083,N_4927,N_4937);
xor U5084 (N_5084,N_4990,N_4930);
and U5085 (N_5085,N_4925,N_4952);
and U5086 (N_5086,N_4906,N_4930);
or U5087 (N_5087,N_4939,N_4949);
xnor U5088 (N_5088,N_4977,N_4904);
nand U5089 (N_5089,N_4999,N_4916);
or U5090 (N_5090,N_4947,N_4929);
nor U5091 (N_5091,N_4965,N_4913);
nand U5092 (N_5092,N_4972,N_4981);
xnor U5093 (N_5093,N_4960,N_4971);
nor U5094 (N_5094,N_4981,N_4909);
xor U5095 (N_5095,N_4952,N_4956);
nand U5096 (N_5096,N_4950,N_4974);
xor U5097 (N_5097,N_4901,N_4929);
nor U5098 (N_5098,N_4994,N_4942);
nor U5099 (N_5099,N_4925,N_4902);
or U5100 (N_5100,N_5007,N_5081);
nor U5101 (N_5101,N_5098,N_5008);
nor U5102 (N_5102,N_5078,N_5084);
xor U5103 (N_5103,N_5097,N_5045);
or U5104 (N_5104,N_5095,N_5009);
and U5105 (N_5105,N_5018,N_5069);
or U5106 (N_5106,N_5052,N_5051);
nand U5107 (N_5107,N_5023,N_5074);
nand U5108 (N_5108,N_5082,N_5031);
xnor U5109 (N_5109,N_5041,N_5089);
and U5110 (N_5110,N_5040,N_5032);
nand U5111 (N_5111,N_5072,N_5096);
nor U5112 (N_5112,N_5014,N_5060);
and U5113 (N_5113,N_5063,N_5071);
and U5114 (N_5114,N_5010,N_5001);
and U5115 (N_5115,N_5017,N_5046);
nand U5116 (N_5116,N_5061,N_5004);
nor U5117 (N_5117,N_5044,N_5058);
and U5118 (N_5118,N_5073,N_5062);
xnor U5119 (N_5119,N_5085,N_5019);
nand U5120 (N_5120,N_5083,N_5021);
nor U5121 (N_5121,N_5038,N_5012);
nor U5122 (N_5122,N_5070,N_5090);
and U5123 (N_5123,N_5077,N_5016);
nand U5124 (N_5124,N_5066,N_5056);
and U5125 (N_5125,N_5067,N_5025);
xor U5126 (N_5126,N_5011,N_5053);
and U5127 (N_5127,N_5030,N_5035);
or U5128 (N_5128,N_5022,N_5036);
or U5129 (N_5129,N_5065,N_5005);
and U5130 (N_5130,N_5003,N_5000);
xor U5131 (N_5131,N_5050,N_5002);
nor U5132 (N_5132,N_5047,N_5076);
xor U5133 (N_5133,N_5028,N_5093);
xnor U5134 (N_5134,N_5059,N_5034);
nand U5135 (N_5135,N_5006,N_5094);
nand U5136 (N_5136,N_5057,N_5087);
or U5137 (N_5137,N_5099,N_5049);
nand U5138 (N_5138,N_5043,N_5029);
xnor U5139 (N_5139,N_5092,N_5054);
nor U5140 (N_5140,N_5048,N_5068);
nand U5141 (N_5141,N_5079,N_5020);
nor U5142 (N_5142,N_5026,N_5075);
nand U5143 (N_5143,N_5091,N_5086);
nor U5144 (N_5144,N_5013,N_5088);
or U5145 (N_5145,N_5042,N_5080);
xnor U5146 (N_5146,N_5064,N_5024);
xor U5147 (N_5147,N_5055,N_5027);
nor U5148 (N_5148,N_5033,N_5039);
nor U5149 (N_5149,N_5037,N_5015);
nand U5150 (N_5150,N_5080,N_5027);
nor U5151 (N_5151,N_5060,N_5049);
nor U5152 (N_5152,N_5054,N_5093);
or U5153 (N_5153,N_5067,N_5001);
nor U5154 (N_5154,N_5008,N_5022);
xnor U5155 (N_5155,N_5091,N_5018);
nor U5156 (N_5156,N_5035,N_5072);
nand U5157 (N_5157,N_5070,N_5075);
or U5158 (N_5158,N_5093,N_5042);
nor U5159 (N_5159,N_5092,N_5013);
nand U5160 (N_5160,N_5062,N_5014);
nand U5161 (N_5161,N_5028,N_5011);
or U5162 (N_5162,N_5037,N_5063);
nand U5163 (N_5163,N_5014,N_5083);
or U5164 (N_5164,N_5089,N_5016);
and U5165 (N_5165,N_5052,N_5065);
or U5166 (N_5166,N_5023,N_5038);
nand U5167 (N_5167,N_5098,N_5032);
xnor U5168 (N_5168,N_5011,N_5022);
or U5169 (N_5169,N_5004,N_5010);
or U5170 (N_5170,N_5034,N_5050);
xor U5171 (N_5171,N_5079,N_5095);
nand U5172 (N_5172,N_5001,N_5045);
nand U5173 (N_5173,N_5002,N_5035);
nand U5174 (N_5174,N_5023,N_5013);
xnor U5175 (N_5175,N_5048,N_5011);
and U5176 (N_5176,N_5070,N_5085);
or U5177 (N_5177,N_5009,N_5072);
or U5178 (N_5178,N_5079,N_5069);
nand U5179 (N_5179,N_5094,N_5032);
or U5180 (N_5180,N_5033,N_5029);
nor U5181 (N_5181,N_5040,N_5072);
and U5182 (N_5182,N_5048,N_5035);
nor U5183 (N_5183,N_5068,N_5000);
and U5184 (N_5184,N_5061,N_5092);
and U5185 (N_5185,N_5077,N_5021);
nor U5186 (N_5186,N_5046,N_5024);
xor U5187 (N_5187,N_5050,N_5071);
xor U5188 (N_5188,N_5017,N_5058);
nor U5189 (N_5189,N_5041,N_5000);
and U5190 (N_5190,N_5011,N_5065);
nor U5191 (N_5191,N_5059,N_5001);
xor U5192 (N_5192,N_5021,N_5059);
nor U5193 (N_5193,N_5084,N_5033);
xor U5194 (N_5194,N_5063,N_5013);
and U5195 (N_5195,N_5077,N_5088);
or U5196 (N_5196,N_5024,N_5061);
nand U5197 (N_5197,N_5088,N_5031);
xnor U5198 (N_5198,N_5032,N_5050);
xor U5199 (N_5199,N_5079,N_5077);
xnor U5200 (N_5200,N_5103,N_5128);
or U5201 (N_5201,N_5135,N_5175);
and U5202 (N_5202,N_5102,N_5113);
or U5203 (N_5203,N_5196,N_5198);
and U5204 (N_5204,N_5114,N_5144);
or U5205 (N_5205,N_5122,N_5165);
xor U5206 (N_5206,N_5140,N_5130);
nand U5207 (N_5207,N_5171,N_5146);
nor U5208 (N_5208,N_5189,N_5156);
xnor U5209 (N_5209,N_5187,N_5125);
xor U5210 (N_5210,N_5121,N_5134);
or U5211 (N_5211,N_5149,N_5127);
xor U5212 (N_5212,N_5104,N_5172);
or U5213 (N_5213,N_5184,N_5166);
nor U5214 (N_5214,N_5126,N_5139);
and U5215 (N_5215,N_5162,N_5163);
nor U5216 (N_5216,N_5193,N_5117);
or U5217 (N_5217,N_5164,N_5194);
nor U5218 (N_5218,N_5143,N_5112);
or U5219 (N_5219,N_5111,N_5105);
nor U5220 (N_5220,N_5138,N_5168);
nor U5221 (N_5221,N_5199,N_5160);
and U5222 (N_5222,N_5137,N_5176);
nor U5223 (N_5223,N_5174,N_5150);
or U5224 (N_5224,N_5129,N_5157);
and U5225 (N_5225,N_5183,N_5115);
xor U5226 (N_5226,N_5186,N_5148);
xor U5227 (N_5227,N_5120,N_5188);
and U5228 (N_5228,N_5132,N_5100);
nand U5229 (N_5229,N_5158,N_5116);
and U5230 (N_5230,N_5154,N_5142);
nand U5231 (N_5231,N_5169,N_5182);
or U5232 (N_5232,N_5133,N_5153);
nand U5233 (N_5233,N_5177,N_5141);
nor U5234 (N_5234,N_5192,N_5123);
and U5235 (N_5235,N_5109,N_5124);
nor U5236 (N_5236,N_5190,N_5191);
nor U5237 (N_5237,N_5195,N_5181);
xnor U5238 (N_5238,N_5108,N_5159);
or U5239 (N_5239,N_5155,N_5136);
nor U5240 (N_5240,N_5145,N_5178);
nor U5241 (N_5241,N_5118,N_5170);
or U5242 (N_5242,N_5185,N_5173);
or U5243 (N_5243,N_5167,N_5197);
nor U5244 (N_5244,N_5106,N_5131);
and U5245 (N_5245,N_5147,N_5110);
and U5246 (N_5246,N_5119,N_5152);
nand U5247 (N_5247,N_5180,N_5151);
nor U5248 (N_5248,N_5107,N_5161);
xnor U5249 (N_5249,N_5101,N_5179);
and U5250 (N_5250,N_5196,N_5195);
nor U5251 (N_5251,N_5188,N_5113);
xnor U5252 (N_5252,N_5111,N_5133);
nand U5253 (N_5253,N_5134,N_5160);
nand U5254 (N_5254,N_5152,N_5155);
nand U5255 (N_5255,N_5108,N_5118);
or U5256 (N_5256,N_5181,N_5141);
nor U5257 (N_5257,N_5128,N_5188);
nor U5258 (N_5258,N_5137,N_5164);
xor U5259 (N_5259,N_5108,N_5101);
or U5260 (N_5260,N_5145,N_5158);
or U5261 (N_5261,N_5100,N_5147);
or U5262 (N_5262,N_5145,N_5128);
xnor U5263 (N_5263,N_5174,N_5179);
nor U5264 (N_5264,N_5127,N_5109);
nand U5265 (N_5265,N_5152,N_5172);
nand U5266 (N_5266,N_5109,N_5154);
nand U5267 (N_5267,N_5135,N_5160);
or U5268 (N_5268,N_5107,N_5176);
nor U5269 (N_5269,N_5174,N_5103);
nand U5270 (N_5270,N_5115,N_5195);
xnor U5271 (N_5271,N_5104,N_5122);
and U5272 (N_5272,N_5115,N_5174);
or U5273 (N_5273,N_5180,N_5126);
nand U5274 (N_5274,N_5191,N_5195);
nand U5275 (N_5275,N_5123,N_5151);
and U5276 (N_5276,N_5169,N_5164);
and U5277 (N_5277,N_5131,N_5111);
nand U5278 (N_5278,N_5127,N_5123);
or U5279 (N_5279,N_5167,N_5142);
nand U5280 (N_5280,N_5142,N_5199);
nor U5281 (N_5281,N_5193,N_5168);
nor U5282 (N_5282,N_5162,N_5127);
and U5283 (N_5283,N_5140,N_5132);
and U5284 (N_5284,N_5100,N_5126);
and U5285 (N_5285,N_5194,N_5147);
and U5286 (N_5286,N_5115,N_5163);
nor U5287 (N_5287,N_5138,N_5137);
and U5288 (N_5288,N_5186,N_5118);
nand U5289 (N_5289,N_5124,N_5155);
xnor U5290 (N_5290,N_5177,N_5104);
and U5291 (N_5291,N_5173,N_5109);
and U5292 (N_5292,N_5150,N_5159);
xor U5293 (N_5293,N_5140,N_5103);
nand U5294 (N_5294,N_5161,N_5101);
xor U5295 (N_5295,N_5108,N_5148);
nor U5296 (N_5296,N_5154,N_5121);
and U5297 (N_5297,N_5142,N_5146);
or U5298 (N_5298,N_5112,N_5154);
nand U5299 (N_5299,N_5156,N_5168);
or U5300 (N_5300,N_5205,N_5216);
nor U5301 (N_5301,N_5221,N_5249);
xnor U5302 (N_5302,N_5264,N_5233);
xnor U5303 (N_5303,N_5258,N_5232);
nor U5304 (N_5304,N_5272,N_5291);
or U5305 (N_5305,N_5247,N_5227);
nand U5306 (N_5306,N_5244,N_5203);
or U5307 (N_5307,N_5288,N_5235);
nor U5308 (N_5308,N_5220,N_5222);
and U5309 (N_5309,N_5229,N_5200);
xnor U5310 (N_5310,N_5231,N_5211);
or U5311 (N_5311,N_5289,N_5283);
nand U5312 (N_5312,N_5275,N_5278);
nor U5313 (N_5313,N_5255,N_5267);
or U5314 (N_5314,N_5210,N_5202);
nand U5315 (N_5315,N_5271,N_5274);
nand U5316 (N_5316,N_5269,N_5242);
and U5317 (N_5317,N_5273,N_5295);
nor U5318 (N_5318,N_5270,N_5223);
nand U5319 (N_5319,N_5296,N_5230);
and U5320 (N_5320,N_5241,N_5245);
or U5321 (N_5321,N_5236,N_5265);
xnor U5322 (N_5322,N_5292,N_5293);
or U5323 (N_5323,N_5282,N_5243);
nand U5324 (N_5324,N_5204,N_5259);
nand U5325 (N_5325,N_5239,N_5248);
or U5326 (N_5326,N_5212,N_5226);
or U5327 (N_5327,N_5240,N_5234);
or U5328 (N_5328,N_5208,N_5268);
xnor U5329 (N_5329,N_5266,N_5252);
and U5330 (N_5330,N_5218,N_5281);
nand U5331 (N_5331,N_5286,N_5253);
nor U5332 (N_5332,N_5224,N_5280);
xor U5333 (N_5333,N_5257,N_5251);
or U5334 (N_5334,N_5215,N_5284);
xnor U5335 (N_5335,N_5213,N_5209);
or U5336 (N_5336,N_5254,N_5201);
and U5337 (N_5337,N_5228,N_5206);
nand U5338 (N_5338,N_5285,N_5207);
nor U5339 (N_5339,N_5250,N_5238);
and U5340 (N_5340,N_5214,N_5298);
or U5341 (N_5341,N_5261,N_5276);
xnor U5342 (N_5342,N_5263,N_5217);
and U5343 (N_5343,N_5262,N_5219);
or U5344 (N_5344,N_5260,N_5225);
xnor U5345 (N_5345,N_5237,N_5297);
nor U5346 (N_5346,N_5279,N_5256);
nor U5347 (N_5347,N_5277,N_5294);
nand U5348 (N_5348,N_5246,N_5299);
and U5349 (N_5349,N_5290,N_5287);
nand U5350 (N_5350,N_5204,N_5215);
xor U5351 (N_5351,N_5264,N_5261);
nor U5352 (N_5352,N_5250,N_5270);
or U5353 (N_5353,N_5214,N_5282);
nand U5354 (N_5354,N_5236,N_5217);
nor U5355 (N_5355,N_5286,N_5205);
or U5356 (N_5356,N_5293,N_5297);
nand U5357 (N_5357,N_5284,N_5212);
and U5358 (N_5358,N_5244,N_5260);
nor U5359 (N_5359,N_5201,N_5240);
or U5360 (N_5360,N_5273,N_5209);
nor U5361 (N_5361,N_5253,N_5257);
nor U5362 (N_5362,N_5239,N_5204);
and U5363 (N_5363,N_5239,N_5253);
nand U5364 (N_5364,N_5287,N_5292);
nand U5365 (N_5365,N_5221,N_5229);
or U5366 (N_5366,N_5272,N_5256);
nor U5367 (N_5367,N_5278,N_5213);
and U5368 (N_5368,N_5294,N_5276);
and U5369 (N_5369,N_5250,N_5251);
nor U5370 (N_5370,N_5231,N_5286);
or U5371 (N_5371,N_5287,N_5214);
or U5372 (N_5372,N_5246,N_5200);
or U5373 (N_5373,N_5280,N_5279);
and U5374 (N_5374,N_5259,N_5262);
xnor U5375 (N_5375,N_5292,N_5212);
nand U5376 (N_5376,N_5274,N_5237);
and U5377 (N_5377,N_5262,N_5288);
nor U5378 (N_5378,N_5228,N_5214);
and U5379 (N_5379,N_5228,N_5229);
or U5380 (N_5380,N_5247,N_5241);
nor U5381 (N_5381,N_5214,N_5211);
nand U5382 (N_5382,N_5202,N_5216);
or U5383 (N_5383,N_5215,N_5219);
and U5384 (N_5384,N_5222,N_5234);
nand U5385 (N_5385,N_5277,N_5223);
xnor U5386 (N_5386,N_5204,N_5233);
xnor U5387 (N_5387,N_5264,N_5207);
or U5388 (N_5388,N_5287,N_5260);
nand U5389 (N_5389,N_5233,N_5286);
nor U5390 (N_5390,N_5237,N_5239);
nand U5391 (N_5391,N_5292,N_5296);
and U5392 (N_5392,N_5276,N_5239);
nor U5393 (N_5393,N_5204,N_5269);
or U5394 (N_5394,N_5225,N_5211);
and U5395 (N_5395,N_5268,N_5231);
or U5396 (N_5396,N_5234,N_5285);
or U5397 (N_5397,N_5291,N_5202);
nor U5398 (N_5398,N_5271,N_5299);
or U5399 (N_5399,N_5293,N_5245);
nand U5400 (N_5400,N_5350,N_5372);
or U5401 (N_5401,N_5344,N_5316);
or U5402 (N_5402,N_5390,N_5332);
or U5403 (N_5403,N_5318,N_5374);
nand U5404 (N_5404,N_5309,N_5365);
or U5405 (N_5405,N_5343,N_5361);
nand U5406 (N_5406,N_5333,N_5364);
xnor U5407 (N_5407,N_5337,N_5305);
or U5408 (N_5408,N_5381,N_5347);
and U5409 (N_5409,N_5330,N_5363);
and U5410 (N_5410,N_5304,N_5395);
nand U5411 (N_5411,N_5398,N_5338);
xor U5412 (N_5412,N_5306,N_5302);
or U5413 (N_5413,N_5368,N_5303);
nand U5414 (N_5414,N_5353,N_5360);
and U5415 (N_5415,N_5382,N_5311);
and U5416 (N_5416,N_5342,N_5308);
nor U5417 (N_5417,N_5329,N_5315);
or U5418 (N_5418,N_5339,N_5393);
and U5419 (N_5419,N_5352,N_5307);
or U5420 (N_5420,N_5387,N_5325);
and U5421 (N_5421,N_5392,N_5322);
xor U5422 (N_5422,N_5383,N_5379);
nand U5423 (N_5423,N_5335,N_5351);
xnor U5424 (N_5424,N_5328,N_5336);
nand U5425 (N_5425,N_5385,N_5327);
nand U5426 (N_5426,N_5378,N_5384);
and U5427 (N_5427,N_5386,N_5321);
nand U5428 (N_5428,N_5312,N_5313);
and U5429 (N_5429,N_5346,N_5341);
nor U5430 (N_5430,N_5399,N_5396);
or U5431 (N_5431,N_5391,N_5356);
xor U5432 (N_5432,N_5357,N_5388);
or U5433 (N_5433,N_5320,N_5310);
and U5434 (N_5434,N_5371,N_5359);
or U5435 (N_5435,N_5345,N_5375);
xnor U5436 (N_5436,N_5362,N_5366);
nor U5437 (N_5437,N_5348,N_5394);
xor U5438 (N_5438,N_5377,N_5370);
nor U5439 (N_5439,N_5324,N_5334);
nor U5440 (N_5440,N_5380,N_5354);
nor U5441 (N_5441,N_5355,N_5331);
or U5442 (N_5442,N_5319,N_5314);
nand U5443 (N_5443,N_5317,N_5367);
xor U5444 (N_5444,N_5301,N_5358);
or U5445 (N_5445,N_5376,N_5397);
and U5446 (N_5446,N_5323,N_5326);
nor U5447 (N_5447,N_5389,N_5369);
or U5448 (N_5448,N_5300,N_5349);
xor U5449 (N_5449,N_5340,N_5373);
xor U5450 (N_5450,N_5301,N_5322);
or U5451 (N_5451,N_5392,N_5389);
nand U5452 (N_5452,N_5315,N_5352);
nand U5453 (N_5453,N_5363,N_5332);
nor U5454 (N_5454,N_5387,N_5354);
nor U5455 (N_5455,N_5388,N_5364);
xor U5456 (N_5456,N_5332,N_5322);
nand U5457 (N_5457,N_5305,N_5399);
nand U5458 (N_5458,N_5325,N_5336);
or U5459 (N_5459,N_5317,N_5356);
xor U5460 (N_5460,N_5310,N_5367);
or U5461 (N_5461,N_5361,N_5362);
nand U5462 (N_5462,N_5307,N_5331);
and U5463 (N_5463,N_5371,N_5310);
and U5464 (N_5464,N_5387,N_5362);
nor U5465 (N_5465,N_5362,N_5392);
or U5466 (N_5466,N_5321,N_5342);
xnor U5467 (N_5467,N_5356,N_5376);
xor U5468 (N_5468,N_5319,N_5369);
or U5469 (N_5469,N_5392,N_5357);
nand U5470 (N_5470,N_5364,N_5348);
nand U5471 (N_5471,N_5303,N_5346);
and U5472 (N_5472,N_5313,N_5322);
or U5473 (N_5473,N_5333,N_5309);
or U5474 (N_5474,N_5323,N_5333);
nand U5475 (N_5475,N_5362,N_5379);
nand U5476 (N_5476,N_5333,N_5310);
nor U5477 (N_5477,N_5351,N_5389);
and U5478 (N_5478,N_5350,N_5336);
nand U5479 (N_5479,N_5355,N_5332);
xnor U5480 (N_5480,N_5358,N_5374);
and U5481 (N_5481,N_5313,N_5369);
nand U5482 (N_5482,N_5384,N_5389);
or U5483 (N_5483,N_5396,N_5380);
nand U5484 (N_5484,N_5309,N_5303);
or U5485 (N_5485,N_5370,N_5301);
or U5486 (N_5486,N_5302,N_5386);
or U5487 (N_5487,N_5347,N_5326);
xnor U5488 (N_5488,N_5327,N_5304);
xnor U5489 (N_5489,N_5308,N_5334);
nand U5490 (N_5490,N_5390,N_5323);
nand U5491 (N_5491,N_5383,N_5303);
nor U5492 (N_5492,N_5394,N_5384);
nor U5493 (N_5493,N_5385,N_5338);
or U5494 (N_5494,N_5394,N_5397);
xnor U5495 (N_5495,N_5346,N_5371);
nand U5496 (N_5496,N_5332,N_5364);
and U5497 (N_5497,N_5349,N_5325);
and U5498 (N_5498,N_5351,N_5352);
or U5499 (N_5499,N_5386,N_5319);
and U5500 (N_5500,N_5407,N_5454);
nand U5501 (N_5501,N_5475,N_5440);
xnor U5502 (N_5502,N_5473,N_5447);
and U5503 (N_5503,N_5481,N_5487);
and U5504 (N_5504,N_5439,N_5404);
xnor U5505 (N_5505,N_5409,N_5457);
nor U5506 (N_5506,N_5460,N_5412);
nor U5507 (N_5507,N_5490,N_5437);
xor U5508 (N_5508,N_5483,N_5482);
nand U5509 (N_5509,N_5418,N_5430);
xor U5510 (N_5510,N_5452,N_5456);
and U5511 (N_5511,N_5428,N_5444);
xor U5512 (N_5512,N_5484,N_5497);
nor U5513 (N_5513,N_5403,N_5486);
or U5514 (N_5514,N_5491,N_5435);
xor U5515 (N_5515,N_5474,N_5410);
and U5516 (N_5516,N_5498,N_5489);
xor U5517 (N_5517,N_5461,N_5419);
and U5518 (N_5518,N_5431,N_5406);
nand U5519 (N_5519,N_5496,N_5413);
nor U5520 (N_5520,N_5408,N_5425);
nor U5521 (N_5521,N_5469,N_5459);
or U5522 (N_5522,N_5417,N_5400);
and U5523 (N_5523,N_5468,N_5401);
nor U5524 (N_5524,N_5485,N_5415);
xor U5525 (N_5525,N_5488,N_5480);
nand U5526 (N_5526,N_5464,N_5436);
nor U5527 (N_5527,N_5438,N_5402);
nor U5528 (N_5528,N_5443,N_5449);
nand U5529 (N_5529,N_5479,N_5495);
xor U5530 (N_5530,N_5427,N_5445);
nand U5531 (N_5531,N_5432,N_5458);
and U5532 (N_5532,N_5446,N_5453);
or U5533 (N_5533,N_5421,N_5462);
or U5534 (N_5534,N_5470,N_5472);
nor U5535 (N_5535,N_5494,N_5499);
nor U5536 (N_5536,N_5467,N_5448);
xnor U5537 (N_5537,N_5416,N_5476);
nor U5538 (N_5538,N_5405,N_5463);
xor U5539 (N_5539,N_5434,N_5426);
and U5540 (N_5540,N_5422,N_5471);
or U5541 (N_5541,N_5429,N_5450);
or U5542 (N_5542,N_5442,N_5465);
and U5543 (N_5543,N_5477,N_5411);
and U5544 (N_5544,N_5466,N_5420);
or U5545 (N_5545,N_5451,N_5433);
nor U5546 (N_5546,N_5414,N_5441);
and U5547 (N_5547,N_5424,N_5455);
and U5548 (N_5548,N_5423,N_5478);
and U5549 (N_5549,N_5493,N_5492);
or U5550 (N_5550,N_5464,N_5408);
or U5551 (N_5551,N_5427,N_5474);
and U5552 (N_5552,N_5438,N_5434);
nand U5553 (N_5553,N_5435,N_5450);
and U5554 (N_5554,N_5426,N_5465);
or U5555 (N_5555,N_5404,N_5440);
nand U5556 (N_5556,N_5425,N_5426);
and U5557 (N_5557,N_5472,N_5499);
xor U5558 (N_5558,N_5409,N_5433);
nand U5559 (N_5559,N_5400,N_5469);
xnor U5560 (N_5560,N_5429,N_5483);
or U5561 (N_5561,N_5402,N_5465);
or U5562 (N_5562,N_5469,N_5436);
nand U5563 (N_5563,N_5438,N_5483);
or U5564 (N_5564,N_5476,N_5466);
nor U5565 (N_5565,N_5487,N_5409);
and U5566 (N_5566,N_5407,N_5492);
xor U5567 (N_5567,N_5436,N_5405);
xnor U5568 (N_5568,N_5436,N_5471);
or U5569 (N_5569,N_5438,N_5471);
nor U5570 (N_5570,N_5416,N_5424);
or U5571 (N_5571,N_5458,N_5465);
xnor U5572 (N_5572,N_5496,N_5420);
or U5573 (N_5573,N_5418,N_5410);
nand U5574 (N_5574,N_5442,N_5493);
xor U5575 (N_5575,N_5417,N_5449);
nor U5576 (N_5576,N_5486,N_5423);
or U5577 (N_5577,N_5415,N_5418);
nor U5578 (N_5578,N_5418,N_5432);
nand U5579 (N_5579,N_5499,N_5414);
and U5580 (N_5580,N_5418,N_5491);
or U5581 (N_5581,N_5430,N_5428);
or U5582 (N_5582,N_5490,N_5406);
xor U5583 (N_5583,N_5406,N_5443);
xnor U5584 (N_5584,N_5442,N_5434);
nand U5585 (N_5585,N_5480,N_5430);
nor U5586 (N_5586,N_5410,N_5409);
nor U5587 (N_5587,N_5409,N_5463);
or U5588 (N_5588,N_5449,N_5405);
nand U5589 (N_5589,N_5450,N_5480);
nor U5590 (N_5590,N_5463,N_5499);
nand U5591 (N_5591,N_5448,N_5494);
nor U5592 (N_5592,N_5423,N_5487);
or U5593 (N_5593,N_5405,N_5429);
nand U5594 (N_5594,N_5401,N_5451);
or U5595 (N_5595,N_5401,N_5495);
nand U5596 (N_5596,N_5441,N_5435);
nand U5597 (N_5597,N_5491,N_5472);
xnor U5598 (N_5598,N_5405,N_5431);
nand U5599 (N_5599,N_5468,N_5461);
nand U5600 (N_5600,N_5570,N_5522);
xnor U5601 (N_5601,N_5576,N_5533);
nand U5602 (N_5602,N_5578,N_5527);
nor U5603 (N_5603,N_5586,N_5568);
nand U5604 (N_5604,N_5560,N_5591);
xor U5605 (N_5605,N_5577,N_5582);
and U5606 (N_5606,N_5548,N_5553);
nor U5607 (N_5607,N_5564,N_5510);
and U5608 (N_5608,N_5585,N_5538);
xnor U5609 (N_5609,N_5539,N_5589);
or U5610 (N_5610,N_5542,N_5580);
nand U5611 (N_5611,N_5562,N_5505);
nor U5612 (N_5612,N_5536,N_5583);
or U5613 (N_5613,N_5509,N_5599);
and U5614 (N_5614,N_5501,N_5588);
and U5615 (N_5615,N_5540,N_5561);
nand U5616 (N_5616,N_5550,N_5547);
and U5617 (N_5617,N_5514,N_5584);
or U5618 (N_5618,N_5513,N_5594);
xor U5619 (N_5619,N_5504,N_5529);
xnor U5620 (N_5620,N_5579,N_5556);
xnor U5621 (N_5621,N_5537,N_5511);
or U5622 (N_5622,N_5515,N_5587);
or U5623 (N_5623,N_5544,N_5546);
nand U5624 (N_5624,N_5518,N_5549);
nand U5625 (N_5625,N_5598,N_5558);
xor U5626 (N_5626,N_5552,N_5535);
nor U5627 (N_5627,N_5503,N_5559);
xnor U5628 (N_5628,N_5526,N_5574);
and U5629 (N_5629,N_5521,N_5508);
or U5630 (N_5630,N_5534,N_5519);
nor U5631 (N_5631,N_5525,N_5545);
xnor U5632 (N_5632,N_5563,N_5500);
nand U5633 (N_5633,N_5596,N_5507);
xor U5634 (N_5634,N_5520,N_5592);
or U5635 (N_5635,N_5569,N_5530);
xor U5636 (N_5636,N_5543,N_5502);
and U5637 (N_5637,N_5554,N_5595);
and U5638 (N_5638,N_5512,N_5532);
and U5639 (N_5639,N_5565,N_5557);
nand U5640 (N_5640,N_5506,N_5593);
and U5641 (N_5641,N_5528,N_5581);
xor U5642 (N_5642,N_5573,N_5572);
nor U5643 (N_5643,N_5516,N_5567);
and U5644 (N_5644,N_5597,N_5541);
or U5645 (N_5645,N_5531,N_5555);
or U5646 (N_5646,N_5551,N_5566);
nor U5647 (N_5647,N_5517,N_5524);
nand U5648 (N_5648,N_5590,N_5571);
nand U5649 (N_5649,N_5575,N_5523);
nand U5650 (N_5650,N_5507,N_5550);
xor U5651 (N_5651,N_5593,N_5539);
and U5652 (N_5652,N_5541,N_5531);
xor U5653 (N_5653,N_5534,N_5568);
or U5654 (N_5654,N_5506,N_5553);
and U5655 (N_5655,N_5583,N_5596);
nor U5656 (N_5656,N_5557,N_5528);
nand U5657 (N_5657,N_5596,N_5539);
nor U5658 (N_5658,N_5505,N_5530);
xnor U5659 (N_5659,N_5581,N_5505);
or U5660 (N_5660,N_5532,N_5531);
xnor U5661 (N_5661,N_5574,N_5529);
and U5662 (N_5662,N_5528,N_5538);
and U5663 (N_5663,N_5596,N_5565);
or U5664 (N_5664,N_5532,N_5539);
and U5665 (N_5665,N_5525,N_5536);
nor U5666 (N_5666,N_5506,N_5530);
or U5667 (N_5667,N_5525,N_5553);
and U5668 (N_5668,N_5584,N_5507);
xnor U5669 (N_5669,N_5508,N_5524);
nor U5670 (N_5670,N_5538,N_5583);
nand U5671 (N_5671,N_5597,N_5584);
nor U5672 (N_5672,N_5536,N_5581);
or U5673 (N_5673,N_5556,N_5520);
nor U5674 (N_5674,N_5565,N_5522);
nand U5675 (N_5675,N_5537,N_5571);
nand U5676 (N_5676,N_5520,N_5583);
xor U5677 (N_5677,N_5590,N_5510);
xnor U5678 (N_5678,N_5568,N_5510);
and U5679 (N_5679,N_5598,N_5521);
nor U5680 (N_5680,N_5584,N_5508);
nor U5681 (N_5681,N_5578,N_5502);
nor U5682 (N_5682,N_5541,N_5573);
or U5683 (N_5683,N_5511,N_5546);
nand U5684 (N_5684,N_5598,N_5506);
and U5685 (N_5685,N_5540,N_5539);
or U5686 (N_5686,N_5545,N_5591);
nor U5687 (N_5687,N_5544,N_5591);
xor U5688 (N_5688,N_5501,N_5515);
and U5689 (N_5689,N_5510,N_5596);
or U5690 (N_5690,N_5564,N_5583);
and U5691 (N_5691,N_5577,N_5501);
nand U5692 (N_5692,N_5545,N_5520);
or U5693 (N_5693,N_5526,N_5564);
nand U5694 (N_5694,N_5598,N_5504);
and U5695 (N_5695,N_5599,N_5587);
or U5696 (N_5696,N_5562,N_5500);
xor U5697 (N_5697,N_5538,N_5562);
nor U5698 (N_5698,N_5533,N_5545);
nor U5699 (N_5699,N_5595,N_5519);
and U5700 (N_5700,N_5625,N_5677);
and U5701 (N_5701,N_5652,N_5671);
or U5702 (N_5702,N_5660,N_5675);
xor U5703 (N_5703,N_5664,N_5608);
and U5704 (N_5704,N_5692,N_5680);
or U5705 (N_5705,N_5629,N_5684);
nand U5706 (N_5706,N_5602,N_5670);
and U5707 (N_5707,N_5637,N_5687);
and U5708 (N_5708,N_5678,N_5667);
nor U5709 (N_5709,N_5647,N_5605);
xor U5710 (N_5710,N_5632,N_5663);
xnor U5711 (N_5711,N_5679,N_5607);
xor U5712 (N_5712,N_5657,N_5611);
nor U5713 (N_5713,N_5666,N_5658);
nand U5714 (N_5714,N_5691,N_5600);
xor U5715 (N_5715,N_5699,N_5601);
nor U5716 (N_5716,N_5610,N_5643);
nor U5717 (N_5717,N_5686,N_5688);
nor U5718 (N_5718,N_5615,N_5682);
nor U5719 (N_5719,N_5673,N_5634);
or U5720 (N_5720,N_5639,N_5676);
and U5721 (N_5721,N_5622,N_5623);
and U5722 (N_5722,N_5683,N_5656);
or U5723 (N_5723,N_5613,N_5644);
nand U5724 (N_5724,N_5640,N_5638);
nor U5725 (N_5725,N_5650,N_5662);
and U5726 (N_5726,N_5626,N_5618);
nor U5727 (N_5727,N_5620,N_5614);
or U5728 (N_5728,N_5669,N_5685);
or U5729 (N_5729,N_5672,N_5609);
nand U5730 (N_5730,N_5642,N_5628);
nor U5731 (N_5731,N_5681,N_5665);
or U5732 (N_5732,N_5696,N_5616);
xor U5733 (N_5733,N_5633,N_5635);
and U5734 (N_5734,N_5624,N_5630);
nand U5735 (N_5735,N_5668,N_5693);
nand U5736 (N_5736,N_5636,N_5641);
or U5737 (N_5737,N_5627,N_5606);
and U5738 (N_5738,N_5661,N_5689);
nor U5739 (N_5739,N_5604,N_5621);
and U5740 (N_5740,N_5617,N_5646);
nand U5741 (N_5741,N_5654,N_5645);
nor U5742 (N_5742,N_5694,N_5697);
or U5743 (N_5743,N_5655,N_5659);
and U5744 (N_5744,N_5603,N_5698);
or U5745 (N_5745,N_5690,N_5649);
and U5746 (N_5746,N_5695,N_5631);
or U5747 (N_5747,N_5651,N_5674);
xor U5748 (N_5748,N_5619,N_5653);
and U5749 (N_5749,N_5648,N_5612);
or U5750 (N_5750,N_5602,N_5636);
nand U5751 (N_5751,N_5672,N_5616);
nor U5752 (N_5752,N_5633,N_5647);
nand U5753 (N_5753,N_5680,N_5665);
and U5754 (N_5754,N_5619,N_5663);
xor U5755 (N_5755,N_5695,N_5658);
nand U5756 (N_5756,N_5656,N_5637);
nand U5757 (N_5757,N_5646,N_5657);
and U5758 (N_5758,N_5666,N_5644);
xnor U5759 (N_5759,N_5625,N_5628);
nor U5760 (N_5760,N_5650,N_5657);
and U5761 (N_5761,N_5638,N_5600);
nor U5762 (N_5762,N_5613,N_5645);
or U5763 (N_5763,N_5635,N_5674);
xor U5764 (N_5764,N_5663,N_5609);
xor U5765 (N_5765,N_5642,N_5683);
xor U5766 (N_5766,N_5657,N_5687);
or U5767 (N_5767,N_5646,N_5610);
xnor U5768 (N_5768,N_5602,N_5653);
xnor U5769 (N_5769,N_5698,N_5653);
nor U5770 (N_5770,N_5625,N_5616);
xnor U5771 (N_5771,N_5657,N_5638);
nand U5772 (N_5772,N_5642,N_5641);
nand U5773 (N_5773,N_5619,N_5608);
and U5774 (N_5774,N_5698,N_5656);
nor U5775 (N_5775,N_5687,N_5664);
xnor U5776 (N_5776,N_5684,N_5639);
nand U5777 (N_5777,N_5687,N_5608);
xor U5778 (N_5778,N_5690,N_5604);
nand U5779 (N_5779,N_5618,N_5658);
and U5780 (N_5780,N_5638,N_5696);
and U5781 (N_5781,N_5661,N_5673);
nor U5782 (N_5782,N_5661,N_5608);
xor U5783 (N_5783,N_5640,N_5658);
and U5784 (N_5784,N_5644,N_5673);
and U5785 (N_5785,N_5647,N_5615);
xor U5786 (N_5786,N_5663,N_5658);
or U5787 (N_5787,N_5624,N_5658);
nor U5788 (N_5788,N_5694,N_5682);
nor U5789 (N_5789,N_5669,N_5603);
xor U5790 (N_5790,N_5647,N_5638);
nand U5791 (N_5791,N_5682,N_5613);
xnor U5792 (N_5792,N_5675,N_5681);
nand U5793 (N_5793,N_5639,N_5681);
xor U5794 (N_5794,N_5684,N_5669);
or U5795 (N_5795,N_5602,N_5692);
nor U5796 (N_5796,N_5652,N_5681);
or U5797 (N_5797,N_5680,N_5696);
nor U5798 (N_5798,N_5609,N_5647);
xnor U5799 (N_5799,N_5692,N_5608);
nand U5800 (N_5800,N_5769,N_5750);
or U5801 (N_5801,N_5727,N_5780);
and U5802 (N_5802,N_5740,N_5785);
and U5803 (N_5803,N_5734,N_5707);
and U5804 (N_5804,N_5758,N_5768);
and U5805 (N_5805,N_5773,N_5762);
nor U5806 (N_5806,N_5784,N_5726);
and U5807 (N_5807,N_5711,N_5744);
or U5808 (N_5808,N_5738,N_5781);
nand U5809 (N_5809,N_5755,N_5700);
nor U5810 (N_5810,N_5771,N_5717);
or U5811 (N_5811,N_5730,N_5779);
nand U5812 (N_5812,N_5728,N_5718);
xor U5813 (N_5813,N_5793,N_5757);
nand U5814 (N_5814,N_5701,N_5747);
or U5815 (N_5815,N_5715,N_5776);
and U5816 (N_5816,N_5742,N_5731);
xor U5817 (N_5817,N_5795,N_5788);
nand U5818 (N_5818,N_5770,N_5704);
xnor U5819 (N_5819,N_5782,N_5778);
and U5820 (N_5820,N_5732,N_5789);
xor U5821 (N_5821,N_5716,N_5767);
nand U5822 (N_5822,N_5729,N_5745);
xnor U5823 (N_5823,N_5765,N_5733);
and U5824 (N_5824,N_5760,N_5766);
and U5825 (N_5825,N_5763,N_5705);
and U5826 (N_5826,N_5721,N_5796);
and U5827 (N_5827,N_5741,N_5720);
xnor U5828 (N_5828,N_5797,N_5764);
xor U5829 (N_5829,N_5794,N_5709);
or U5830 (N_5830,N_5799,N_5759);
nand U5831 (N_5831,N_5787,N_5792);
nor U5832 (N_5832,N_5774,N_5706);
nand U5833 (N_5833,N_5708,N_5756);
nand U5834 (N_5834,N_5791,N_5739);
xnor U5835 (N_5835,N_5761,N_5748);
nor U5836 (N_5836,N_5754,N_5743);
nand U5837 (N_5837,N_5751,N_5786);
and U5838 (N_5838,N_5777,N_5737);
xnor U5839 (N_5839,N_5736,N_5723);
xor U5840 (N_5840,N_5790,N_5798);
nor U5841 (N_5841,N_5752,N_5722);
or U5842 (N_5842,N_5713,N_5735);
nand U5843 (N_5843,N_5783,N_5710);
and U5844 (N_5844,N_5725,N_5724);
xor U5845 (N_5845,N_5772,N_5775);
or U5846 (N_5846,N_5703,N_5753);
xor U5847 (N_5847,N_5714,N_5746);
nand U5848 (N_5848,N_5749,N_5719);
xor U5849 (N_5849,N_5702,N_5712);
and U5850 (N_5850,N_5733,N_5728);
nand U5851 (N_5851,N_5754,N_5776);
nor U5852 (N_5852,N_5757,N_5732);
xnor U5853 (N_5853,N_5795,N_5720);
or U5854 (N_5854,N_5714,N_5708);
xor U5855 (N_5855,N_5766,N_5738);
nand U5856 (N_5856,N_5797,N_5773);
nor U5857 (N_5857,N_5732,N_5721);
or U5858 (N_5858,N_5751,N_5793);
and U5859 (N_5859,N_5747,N_5776);
xor U5860 (N_5860,N_5701,N_5708);
and U5861 (N_5861,N_5740,N_5792);
nor U5862 (N_5862,N_5799,N_5768);
nand U5863 (N_5863,N_5773,N_5746);
or U5864 (N_5864,N_5749,N_5754);
nand U5865 (N_5865,N_5766,N_5735);
and U5866 (N_5866,N_5727,N_5737);
and U5867 (N_5867,N_5716,N_5730);
or U5868 (N_5868,N_5764,N_5732);
and U5869 (N_5869,N_5775,N_5724);
xnor U5870 (N_5870,N_5749,N_5770);
xnor U5871 (N_5871,N_5764,N_5777);
and U5872 (N_5872,N_5759,N_5772);
xnor U5873 (N_5873,N_5739,N_5771);
nand U5874 (N_5874,N_5744,N_5776);
or U5875 (N_5875,N_5711,N_5709);
or U5876 (N_5876,N_5769,N_5709);
xor U5877 (N_5877,N_5778,N_5784);
or U5878 (N_5878,N_5760,N_5724);
nand U5879 (N_5879,N_5712,N_5748);
nand U5880 (N_5880,N_5769,N_5775);
or U5881 (N_5881,N_5742,N_5752);
or U5882 (N_5882,N_5700,N_5719);
nor U5883 (N_5883,N_5700,N_5762);
xor U5884 (N_5884,N_5786,N_5709);
nand U5885 (N_5885,N_5713,N_5793);
nand U5886 (N_5886,N_5784,N_5753);
xor U5887 (N_5887,N_5744,N_5703);
nor U5888 (N_5888,N_5795,N_5701);
and U5889 (N_5889,N_5735,N_5798);
and U5890 (N_5890,N_5754,N_5709);
or U5891 (N_5891,N_5756,N_5775);
and U5892 (N_5892,N_5733,N_5727);
and U5893 (N_5893,N_5773,N_5748);
and U5894 (N_5894,N_5795,N_5752);
nand U5895 (N_5895,N_5790,N_5744);
or U5896 (N_5896,N_5718,N_5739);
xnor U5897 (N_5897,N_5757,N_5740);
nor U5898 (N_5898,N_5792,N_5704);
xnor U5899 (N_5899,N_5796,N_5719);
nand U5900 (N_5900,N_5829,N_5857);
or U5901 (N_5901,N_5833,N_5811);
nand U5902 (N_5902,N_5819,N_5841);
nor U5903 (N_5903,N_5879,N_5874);
nand U5904 (N_5904,N_5867,N_5800);
or U5905 (N_5905,N_5854,N_5802);
xor U5906 (N_5906,N_5839,N_5838);
nor U5907 (N_5907,N_5842,N_5897);
and U5908 (N_5908,N_5866,N_5852);
nor U5909 (N_5909,N_5815,N_5887);
xnor U5910 (N_5910,N_5805,N_5846);
and U5911 (N_5911,N_5865,N_5826);
or U5912 (N_5912,N_5885,N_5883);
nand U5913 (N_5913,N_5803,N_5880);
and U5914 (N_5914,N_5817,N_5896);
nor U5915 (N_5915,N_5888,N_5832);
xnor U5916 (N_5916,N_5823,N_5812);
nand U5917 (N_5917,N_5898,N_5830);
and U5918 (N_5918,N_5871,N_5816);
xor U5919 (N_5919,N_5859,N_5849);
and U5920 (N_5920,N_5870,N_5831);
nand U5921 (N_5921,N_5899,N_5890);
or U5922 (N_5922,N_5894,N_5827);
and U5923 (N_5923,N_5844,N_5860);
and U5924 (N_5924,N_5806,N_5807);
or U5925 (N_5925,N_5878,N_5851);
xor U5926 (N_5926,N_5834,N_5845);
or U5927 (N_5927,N_5889,N_5821);
and U5928 (N_5928,N_5825,N_5813);
or U5929 (N_5929,N_5835,N_5818);
and U5930 (N_5930,N_5855,N_5861);
or U5931 (N_5931,N_5892,N_5886);
and U5932 (N_5932,N_5810,N_5820);
nor U5933 (N_5933,N_5856,N_5872);
xnor U5934 (N_5934,N_5801,N_5862);
and U5935 (N_5935,N_5876,N_5869);
and U5936 (N_5936,N_5848,N_5875);
nand U5937 (N_5937,N_5824,N_5895);
xnor U5938 (N_5938,N_5804,N_5853);
and U5939 (N_5939,N_5808,N_5847);
nor U5940 (N_5940,N_5891,N_5850);
or U5941 (N_5941,N_5884,N_5828);
or U5942 (N_5942,N_5836,N_5809);
nand U5943 (N_5943,N_5822,N_5858);
nand U5944 (N_5944,N_5882,N_5873);
xor U5945 (N_5945,N_5840,N_5864);
nand U5946 (N_5946,N_5843,N_5868);
or U5947 (N_5947,N_5863,N_5837);
or U5948 (N_5948,N_5881,N_5877);
or U5949 (N_5949,N_5814,N_5893);
nand U5950 (N_5950,N_5866,N_5821);
xor U5951 (N_5951,N_5893,N_5842);
or U5952 (N_5952,N_5841,N_5812);
nor U5953 (N_5953,N_5847,N_5829);
xnor U5954 (N_5954,N_5860,N_5897);
and U5955 (N_5955,N_5871,N_5843);
or U5956 (N_5956,N_5882,N_5823);
nor U5957 (N_5957,N_5801,N_5898);
nor U5958 (N_5958,N_5841,N_5861);
or U5959 (N_5959,N_5816,N_5803);
and U5960 (N_5960,N_5850,N_5843);
and U5961 (N_5961,N_5855,N_5802);
and U5962 (N_5962,N_5870,N_5815);
nor U5963 (N_5963,N_5849,N_5874);
nor U5964 (N_5964,N_5822,N_5848);
nand U5965 (N_5965,N_5812,N_5821);
and U5966 (N_5966,N_5834,N_5821);
and U5967 (N_5967,N_5877,N_5849);
xnor U5968 (N_5968,N_5807,N_5883);
xor U5969 (N_5969,N_5841,N_5840);
and U5970 (N_5970,N_5809,N_5864);
or U5971 (N_5971,N_5887,N_5834);
and U5972 (N_5972,N_5806,N_5811);
nor U5973 (N_5973,N_5894,N_5891);
and U5974 (N_5974,N_5857,N_5810);
xnor U5975 (N_5975,N_5858,N_5852);
nor U5976 (N_5976,N_5833,N_5846);
and U5977 (N_5977,N_5878,N_5859);
xnor U5978 (N_5978,N_5819,N_5802);
and U5979 (N_5979,N_5898,N_5894);
xor U5980 (N_5980,N_5807,N_5891);
or U5981 (N_5981,N_5876,N_5877);
and U5982 (N_5982,N_5859,N_5891);
nor U5983 (N_5983,N_5806,N_5863);
or U5984 (N_5984,N_5882,N_5890);
xor U5985 (N_5985,N_5891,N_5837);
or U5986 (N_5986,N_5837,N_5856);
nand U5987 (N_5987,N_5867,N_5806);
and U5988 (N_5988,N_5812,N_5831);
nor U5989 (N_5989,N_5867,N_5849);
and U5990 (N_5990,N_5886,N_5835);
or U5991 (N_5991,N_5885,N_5842);
nand U5992 (N_5992,N_5884,N_5843);
nor U5993 (N_5993,N_5855,N_5837);
xnor U5994 (N_5994,N_5877,N_5892);
and U5995 (N_5995,N_5883,N_5810);
nor U5996 (N_5996,N_5843,N_5882);
nor U5997 (N_5997,N_5832,N_5868);
and U5998 (N_5998,N_5888,N_5811);
nor U5999 (N_5999,N_5877,N_5810);
or U6000 (N_6000,N_5962,N_5942);
or U6001 (N_6001,N_5989,N_5961);
and U6002 (N_6002,N_5974,N_5999);
or U6003 (N_6003,N_5978,N_5946);
and U6004 (N_6004,N_5902,N_5915);
nor U6005 (N_6005,N_5949,N_5900);
or U6006 (N_6006,N_5943,N_5924);
xor U6007 (N_6007,N_5919,N_5923);
xnor U6008 (N_6008,N_5939,N_5972);
nand U6009 (N_6009,N_5965,N_5967);
xnor U6010 (N_6010,N_5968,N_5983);
or U6011 (N_6011,N_5953,N_5971);
nand U6012 (N_6012,N_5980,N_5938);
nand U6013 (N_6013,N_5912,N_5907);
xor U6014 (N_6014,N_5950,N_5935);
xor U6015 (N_6015,N_5990,N_5913);
nor U6016 (N_6016,N_5917,N_5987);
nand U6017 (N_6017,N_5994,N_5914);
and U6018 (N_6018,N_5958,N_5925);
and U6019 (N_6019,N_5906,N_5916);
or U6020 (N_6020,N_5908,N_5922);
xor U6021 (N_6021,N_5970,N_5984);
xor U6022 (N_6022,N_5985,N_5944);
nor U6023 (N_6023,N_5920,N_5973);
nor U6024 (N_6024,N_5948,N_5954);
and U6025 (N_6025,N_5941,N_5991);
or U6026 (N_6026,N_5910,N_5926);
and U6027 (N_6027,N_5918,N_5937);
or U6028 (N_6028,N_5982,N_5969);
and U6029 (N_6029,N_5927,N_5963);
and U6030 (N_6030,N_5997,N_5921);
or U6031 (N_6031,N_5928,N_5905);
or U6032 (N_6032,N_5909,N_5931);
or U6033 (N_6033,N_5955,N_5956);
xnor U6034 (N_6034,N_5903,N_5995);
nor U6035 (N_6035,N_5981,N_5998);
nand U6036 (N_6036,N_5957,N_5959);
and U6037 (N_6037,N_5933,N_5932);
nor U6038 (N_6038,N_5979,N_5929);
xnor U6039 (N_6039,N_5940,N_5934);
nand U6040 (N_6040,N_5975,N_5911);
and U6041 (N_6041,N_5986,N_5977);
nor U6042 (N_6042,N_5996,N_5960);
and U6043 (N_6043,N_5988,N_5966);
and U6044 (N_6044,N_5901,N_5993);
nor U6045 (N_6045,N_5992,N_5976);
xor U6046 (N_6046,N_5945,N_5964);
nor U6047 (N_6047,N_5947,N_5952);
or U6048 (N_6048,N_5951,N_5936);
nor U6049 (N_6049,N_5904,N_5930);
or U6050 (N_6050,N_5988,N_5977);
and U6051 (N_6051,N_5900,N_5932);
nor U6052 (N_6052,N_5934,N_5993);
nor U6053 (N_6053,N_5946,N_5980);
nor U6054 (N_6054,N_5919,N_5977);
and U6055 (N_6055,N_5951,N_5926);
nand U6056 (N_6056,N_5994,N_5908);
xnor U6057 (N_6057,N_5949,N_5943);
nand U6058 (N_6058,N_5949,N_5992);
or U6059 (N_6059,N_5969,N_5957);
or U6060 (N_6060,N_5932,N_5961);
and U6061 (N_6061,N_5987,N_5963);
nand U6062 (N_6062,N_5998,N_5969);
or U6063 (N_6063,N_5904,N_5907);
nor U6064 (N_6064,N_5969,N_5991);
xnor U6065 (N_6065,N_5943,N_5956);
or U6066 (N_6066,N_5900,N_5916);
nand U6067 (N_6067,N_5975,N_5933);
or U6068 (N_6068,N_5949,N_5904);
xor U6069 (N_6069,N_5927,N_5925);
or U6070 (N_6070,N_5905,N_5990);
nand U6071 (N_6071,N_5950,N_5966);
nand U6072 (N_6072,N_5957,N_5943);
and U6073 (N_6073,N_5929,N_5915);
nand U6074 (N_6074,N_5959,N_5967);
xor U6075 (N_6075,N_5900,N_5931);
xnor U6076 (N_6076,N_5990,N_5994);
nand U6077 (N_6077,N_5974,N_5983);
or U6078 (N_6078,N_5904,N_5953);
nand U6079 (N_6079,N_5999,N_5906);
or U6080 (N_6080,N_5964,N_5965);
and U6081 (N_6081,N_5951,N_5919);
nand U6082 (N_6082,N_5940,N_5955);
and U6083 (N_6083,N_5994,N_5937);
nand U6084 (N_6084,N_5992,N_5937);
or U6085 (N_6085,N_5965,N_5918);
nand U6086 (N_6086,N_5916,N_5964);
nor U6087 (N_6087,N_5909,N_5977);
xnor U6088 (N_6088,N_5940,N_5918);
and U6089 (N_6089,N_5943,N_5990);
nor U6090 (N_6090,N_5987,N_5982);
nand U6091 (N_6091,N_5919,N_5903);
xnor U6092 (N_6092,N_5910,N_5931);
nor U6093 (N_6093,N_5901,N_5906);
xnor U6094 (N_6094,N_5923,N_5912);
nor U6095 (N_6095,N_5922,N_5903);
or U6096 (N_6096,N_5902,N_5904);
or U6097 (N_6097,N_5960,N_5971);
or U6098 (N_6098,N_5904,N_5936);
nor U6099 (N_6099,N_5958,N_5961);
nand U6100 (N_6100,N_6054,N_6011);
nand U6101 (N_6101,N_6050,N_6094);
nand U6102 (N_6102,N_6009,N_6067);
nor U6103 (N_6103,N_6042,N_6013);
and U6104 (N_6104,N_6056,N_6037);
xor U6105 (N_6105,N_6022,N_6052);
or U6106 (N_6106,N_6051,N_6058);
xor U6107 (N_6107,N_6080,N_6039);
nor U6108 (N_6108,N_6083,N_6096);
nand U6109 (N_6109,N_6076,N_6073);
and U6110 (N_6110,N_6033,N_6007);
and U6111 (N_6111,N_6085,N_6020);
xnor U6112 (N_6112,N_6008,N_6026);
nor U6113 (N_6113,N_6040,N_6074);
nand U6114 (N_6114,N_6046,N_6065);
xor U6115 (N_6115,N_6098,N_6014);
xnor U6116 (N_6116,N_6018,N_6075);
nor U6117 (N_6117,N_6077,N_6035);
and U6118 (N_6118,N_6063,N_6064);
and U6119 (N_6119,N_6068,N_6082);
nor U6120 (N_6120,N_6071,N_6048);
xnor U6121 (N_6121,N_6004,N_6034);
and U6122 (N_6122,N_6055,N_6024);
nor U6123 (N_6123,N_6093,N_6006);
nor U6124 (N_6124,N_6081,N_6069);
xor U6125 (N_6125,N_6043,N_6057);
and U6126 (N_6126,N_6062,N_6044);
nor U6127 (N_6127,N_6012,N_6002);
nor U6128 (N_6128,N_6047,N_6001);
and U6129 (N_6129,N_6028,N_6097);
nand U6130 (N_6130,N_6059,N_6015);
nand U6131 (N_6131,N_6019,N_6023);
and U6132 (N_6132,N_6032,N_6029);
nand U6133 (N_6133,N_6045,N_6090);
and U6134 (N_6134,N_6010,N_6088);
nand U6135 (N_6135,N_6031,N_6000);
or U6136 (N_6136,N_6095,N_6078);
or U6137 (N_6137,N_6017,N_6053);
and U6138 (N_6138,N_6066,N_6092);
nand U6139 (N_6139,N_6027,N_6021);
and U6140 (N_6140,N_6005,N_6061);
nor U6141 (N_6141,N_6038,N_6091);
or U6142 (N_6142,N_6087,N_6025);
nor U6143 (N_6143,N_6041,N_6072);
xnor U6144 (N_6144,N_6016,N_6030);
nor U6145 (N_6145,N_6070,N_6079);
and U6146 (N_6146,N_6049,N_6089);
and U6147 (N_6147,N_6086,N_6036);
or U6148 (N_6148,N_6099,N_6060);
xor U6149 (N_6149,N_6084,N_6003);
xor U6150 (N_6150,N_6017,N_6094);
or U6151 (N_6151,N_6075,N_6043);
xor U6152 (N_6152,N_6047,N_6092);
nand U6153 (N_6153,N_6055,N_6071);
nor U6154 (N_6154,N_6045,N_6024);
nand U6155 (N_6155,N_6067,N_6015);
nor U6156 (N_6156,N_6054,N_6027);
nand U6157 (N_6157,N_6030,N_6026);
xor U6158 (N_6158,N_6012,N_6090);
nor U6159 (N_6159,N_6031,N_6033);
nand U6160 (N_6160,N_6094,N_6059);
nor U6161 (N_6161,N_6016,N_6052);
nor U6162 (N_6162,N_6051,N_6077);
and U6163 (N_6163,N_6081,N_6078);
xor U6164 (N_6164,N_6009,N_6020);
or U6165 (N_6165,N_6094,N_6058);
nand U6166 (N_6166,N_6010,N_6007);
and U6167 (N_6167,N_6088,N_6082);
nor U6168 (N_6168,N_6003,N_6083);
and U6169 (N_6169,N_6037,N_6039);
and U6170 (N_6170,N_6046,N_6088);
nand U6171 (N_6171,N_6090,N_6058);
xor U6172 (N_6172,N_6058,N_6046);
nor U6173 (N_6173,N_6024,N_6032);
xor U6174 (N_6174,N_6038,N_6098);
and U6175 (N_6175,N_6023,N_6024);
xor U6176 (N_6176,N_6070,N_6012);
and U6177 (N_6177,N_6095,N_6030);
nand U6178 (N_6178,N_6072,N_6054);
nor U6179 (N_6179,N_6021,N_6037);
and U6180 (N_6180,N_6098,N_6054);
and U6181 (N_6181,N_6024,N_6016);
xnor U6182 (N_6182,N_6096,N_6033);
nor U6183 (N_6183,N_6023,N_6025);
xnor U6184 (N_6184,N_6024,N_6000);
or U6185 (N_6185,N_6070,N_6040);
xnor U6186 (N_6186,N_6003,N_6019);
nor U6187 (N_6187,N_6026,N_6048);
and U6188 (N_6188,N_6029,N_6084);
and U6189 (N_6189,N_6006,N_6065);
nor U6190 (N_6190,N_6071,N_6095);
xnor U6191 (N_6191,N_6031,N_6029);
and U6192 (N_6192,N_6093,N_6074);
xnor U6193 (N_6193,N_6040,N_6097);
nand U6194 (N_6194,N_6051,N_6039);
or U6195 (N_6195,N_6028,N_6022);
xor U6196 (N_6196,N_6039,N_6005);
nand U6197 (N_6197,N_6013,N_6031);
nor U6198 (N_6198,N_6011,N_6017);
nor U6199 (N_6199,N_6097,N_6076);
and U6200 (N_6200,N_6159,N_6136);
nand U6201 (N_6201,N_6192,N_6121);
nor U6202 (N_6202,N_6115,N_6158);
xnor U6203 (N_6203,N_6165,N_6146);
nand U6204 (N_6204,N_6176,N_6174);
nand U6205 (N_6205,N_6139,N_6172);
and U6206 (N_6206,N_6168,N_6106);
and U6207 (N_6207,N_6117,N_6156);
nor U6208 (N_6208,N_6114,N_6179);
nand U6209 (N_6209,N_6113,N_6128);
nand U6210 (N_6210,N_6185,N_6101);
nand U6211 (N_6211,N_6148,N_6180);
or U6212 (N_6212,N_6191,N_6197);
nor U6213 (N_6213,N_6122,N_6190);
and U6214 (N_6214,N_6182,N_6162);
or U6215 (N_6215,N_6131,N_6195);
nor U6216 (N_6216,N_6107,N_6102);
and U6217 (N_6217,N_6100,N_6187);
and U6218 (N_6218,N_6132,N_6175);
nand U6219 (N_6219,N_6183,N_6164);
nand U6220 (N_6220,N_6140,N_6130);
or U6221 (N_6221,N_6134,N_6119);
or U6222 (N_6222,N_6103,N_6189);
or U6223 (N_6223,N_6111,N_6184);
xor U6224 (N_6224,N_6124,N_6170);
or U6225 (N_6225,N_6150,N_6177);
nand U6226 (N_6226,N_6104,N_6196);
nand U6227 (N_6227,N_6152,N_6147);
nand U6228 (N_6228,N_6105,N_6178);
xnor U6229 (N_6229,N_6123,N_6149);
xnor U6230 (N_6230,N_6194,N_6181);
nor U6231 (N_6231,N_6198,N_6157);
or U6232 (N_6232,N_6125,N_6151);
nand U6233 (N_6233,N_6167,N_6186);
nor U6234 (N_6234,N_6137,N_6154);
and U6235 (N_6235,N_6116,N_6138);
or U6236 (N_6236,N_6120,N_6171);
nand U6237 (N_6237,N_6112,N_6145);
and U6238 (N_6238,N_6199,N_6129);
nor U6239 (N_6239,N_6193,N_6141);
nand U6240 (N_6240,N_6160,N_6169);
nor U6241 (N_6241,N_6143,N_6133);
nand U6242 (N_6242,N_6135,N_6163);
and U6243 (N_6243,N_6109,N_6118);
nor U6244 (N_6244,N_6110,N_6108);
and U6245 (N_6245,N_6188,N_6173);
or U6246 (N_6246,N_6153,N_6127);
nand U6247 (N_6247,N_6166,N_6144);
nor U6248 (N_6248,N_6161,N_6142);
or U6249 (N_6249,N_6155,N_6126);
or U6250 (N_6250,N_6199,N_6145);
nor U6251 (N_6251,N_6167,N_6192);
nand U6252 (N_6252,N_6176,N_6175);
xnor U6253 (N_6253,N_6126,N_6123);
xor U6254 (N_6254,N_6132,N_6100);
nand U6255 (N_6255,N_6106,N_6181);
nor U6256 (N_6256,N_6175,N_6196);
and U6257 (N_6257,N_6172,N_6198);
nand U6258 (N_6258,N_6184,N_6193);
and U6259 (N_6259,N_6123,N_6110);
nor U6260 (N_6260,N_6154,N_6197);
xnor U6261 (N_6261,N_6169,N_6159);
nand U6262 (N_6262,N_6146,N_6105);
xnor U6263 (N_6263,N_6145,N_6111);
nand U6264 (N_6264,N_6178,N_6154);
and U6265 (N_6265,N_6188,N_6103);
nor U6266 (N_6266,N_6116,N_6196);
nand U6267 (N_6267,N_6110,N_6146);
or U6268 (N_6268,N_6111,N_6166);
and U6269 (N_6269,N_6162,N_6118);
and U6270 (N_6270,N_6199,N_6138);
or U6271 (N_6271,N_6136,N_6198);
and U6272 (N_6272,N_6124,N_6159);
or U6273 (N_6273,N_6175,N_6126);
or U6274 (N_6274,N_6176,N_6124);
nand U6275 (N_6275,N_6148,N_6113);
xnor U6276 (N_6276,N_6163,N_6124);
nor U6277 (N_6277,N_6110,N_6102);
or U6278 (N_6278,N_6118,N_6107);
and U6279 (N_6279,N_6185,N_6175);
nand U6280 (N_6280,N_6152,N_6165);
nand U6281 (N_6281,N_6163,N_6174);
nand U6282 (N_6282,N_6169,N_6119);
or U6283 (N_6283,N_6149,N_6180);
xnor U6284 (N_6284,N_6122,N_6182);
nand U6285 (N_6285,N_6104,N_6190);
or U6286 (N_6286,N_6159,N_6116);
nand U6287 (N_6287,N_6113,N_6185);
and U6288 (N_6288,N_6100,N_6103);
nand U6289 (N_6289,N_6116,N_6193);
nand U6290 (N_6290,N_6144,N_6159);
and U6291 (N_6291,N_6181,N_6136);
nand U6292 (N_6292,N_6175,N_6162);
xnor U6293 (N_6293,N_6105,N_6153);
and U6294 (N_6294,N_6177,N_6158);
or U6295 (N_6295,N_6152,N_6185);
and U6296 (N_6296,N_6177,N_6115);
and U6297 (N_6297,N_6125,N_6144);
nor U6298 (N_6298,N_6150,N_6144);
xnor U6299 (N_6299,N_6135,N_6123);
nor U6300 (N_6300,N_6239,N_6281);
nand U6301 (N_6301,N_6242,N_6271);
nor U6302 (N_6302,N_6269,N_6227);
and U6303 (N_6303,N_6266,N_6249);
nand U6304 (N_6304,N_6257,N_6237);
or U6305 (N_6305,N_6220,N_6245);
and U6306 (N_6306,N_6289,N_6259);
and U6307 (N_6307,N_6284,N_6268);
xnor U6308 (N_6308,N_6246,N_6263);
nand U6309 (N_6309,N_6288,N_6294);
and U6310 (N_6310,N_6272,N_6273);
and U6311 (N_6311,N_6292,N_6206);
xor U6312 (N_6312,N_6258,N_6255);
xor U6313 (N_6313,N_6247,N_6250);
nand U6314 (N_6314,N_6279,N_6204);
and U6315 (N_6315,N_6275,N_6261);
or U6316 (N_6316,N_6248,N_6212);
or U6317 (N_6317,N_6213,N_6277);
nor U6318 (N_6318,N_6210,N_6207);
xnor U6319 (N_6319,N_6236,N_6291);
nor U6320 (N_6320,N_6270,N_6208);
xnor U6321 (N_6321,N_6202,N_6282);
nand U6322 (N_6322,N_6235,N_6278);
or U6323 (N_6323,N_6203,N_6293);
or U6324 (N_6324,N_6240,N_6286);
xor U6325 (N_6325,N_6228,N_6298);
xnor U6326 (N_6326,N_6226,N_6295);
or U6327 (N_6327,N_6296,N_6243);
nor U6328 (N_6328,N_6200,N_6265);
and U6329 (N_6329,N_6254,N_6224);
nor U6330 (N_6330,N_6215,N_6297);
nor U6331 (N_6331,N_6260,N_6211);
and U6332 (N_6332,N_6217,N_6214);
nand U6333 (N_6333,N_6244,N_6219);
nand U6334 (N_6334,N_6222,N_6267);
or U6335 (N_6335,N_6231,N_6232);
xor U6336 (N_6336,N_6274,N_6230);
nand U6337 (N_6337,N_6299,N_6285);
and U6338 (N_6338,N_6287,N_6280);
or U6339 (N_6339,N_6201,N_6218);
and U6340 (N_6340,N_6234,N_6276);
nor U6341 (N_6341,N_6256,N_6264);
and U6342 (N_6342,N_6241,N_6229);
and U6343 (N_6343,N_6209,N_6253);
and U6344 (N_6344,N_6223,N_6225);
nand U6345 (N_6345,N_6252,N_6233);
nor U6346 (N_6346,N_6216,N_6283);
xnor U6347 (N_6347,N_6221,N_6262);
xnor U6348 (N_6348,N_6238,N_6205);
nor U6349 (N_6349,N_6251,N_6290);
nor U6350 (N_6350,N_6200,N_6256);
and U6351 (N_6351,N_6235,N_6208);
and U6352 (N_6352,N_6220,N_6268);
nor U6353 (N_6353,N_6272,N_6222);
nand U6354 (N_6354,N_6265,N_6246);
and U6355 (N_6355,N_6233,N_6222);
nand U6356 (N_6356,N_6240,N_6250);
or U6357 (N_6357,N_6263,N_6295);
or U6358 (N_6358,N_6248,N_6208);
nand U6359 (N_6359,N_6268,N_6226);
nor U6360 (N_6360,N_6298,N_6261);
and U6361 (N_6361,N_6209,N_6264);
nand U6362 (N_6362,N_6278,N_6283);
nand U6363 (N_6363,N_6282,N_6240);
or U6364 (N_6364,N_6276,N_6208);
or U6365 (N_6365,N_6256,N_6292);
and U6366 (N_6366,N_6211,N_6205);
xnor U6367 (N_6367,N_6239,N_6286);
xor U6368 (N_6368,N_6229,N_6236);
nand U6369 (N_6369,N_6285,N_6224);
xnor U6370 (N_6370,N_6230,N_6293);
nand U6371 (N_6371,N_6220,N_6285);
nor U6372 (N_6372,N_6202,N_6293);
nand U6373 (N_6373,N_6243,N_6225);
and U6374 (N_6374,N_6246,N_6268);
or U6375 (N_6375,N_6297,N_6214);
nand U6376 (N_6376,N_6218,N_6247);
xor U6377 (N_6377,N_6213,N_6238);
and U6378 (N_6378,N_6214,N_6237);
nor U6379 (N_6379,N_6223,N_6230);
nor U6380 (N_6380,N_6201,N_6232);
and U6381 (N_6381,N_6261,N_6274);
and U6382 (N_6382,N_6295,N_6222);
and U6383 (N_6383,N_6227,N_6298);
and U6384 (N_6384,N_6210,N_6228);
xor U6385 (N_6385,N_6248,N_6250);
xor U6386 (N_6386,N_6267,N_6235);
nor U6387 (N_6387,N_6214,N_6292);
nand U6388 (N_6388,N_6260,N_6232);
nor U6389 (N_6389,N_6260,N_6225);
nor U6390 (N_6390,N_6293,N_6242);
nor U6391 (N_6391,N_6230,N_6260);
nor U6392 (N_6392,N_6248,N_6294);
xnor U6393 (N_6393,N_6299,N_6220);
and U6394 (N_6394,N_6280,N_6202);
nand U6395 (N_6395,N_6202,N_6250);
and U6396 (N_6396,N_6210,N_6241);
or U6397 (N_6397,N_6259,N_6204);
or U6398 (N_6398,N_6277,N_6268);
nand U6399 (N_6399,N_6242,N_6223);
nand U6400 (N_6400,N_6392,N_6341);
nand U6401 (N_6401,N_6315,N_6311);
and U6402 (N_6402,N_6380,N_6360);
nand U6403 (N_6403,N_6367,N_6373);
or U6404 (N_6404,N_6366,N_6348);
nand U6405 (N_6405,N_6330,N_6362);
xor U6406 (N_6406,N_6356,N_6314);
nor U6407 (N_6407,N_6316,N_6300);
or U6408 (N_6408,N_6381,N_6399);
nor U6409 (N_6409,N_6361,N_6393);
nand U6410 (N_6410,N_6390,N_6397);
nand U6411 (N_6411,N_6370,N_6365);
or U6412 (N_6412,N_6309,N_6351);
nor U6413 (N_6413,N_6306,N_6343);
and U6414 (N_6414,N_6308,N_6327);
and U6415 (N_6415,N_6322,N_6387);
or U6416 (N_6416,N_6323,N_6302);
nand U6417 (N_6417,N_6369,N_6346);
and U6418 (N_6418,N_6391,N_6350);
nor U6419 (N_6419,N_6318,N_6342);
or U6420 (N_6420,N_6304,N_6368);
xor U6421 (N_6421,N_6319,N_6332);
xnor U6422 (N_6422,N_6374,N_6301);
and U6423 (N_6423,N_6310,N_6386);
xor U6424 (N_6424,N_6345,N_6320);
and U6425 (N_6425,N_6324,N_6347);
or U6426 (N_6426,N_6364,N_6388);
xor U6427 (N_6427,N_6335,N_6398);
nand U6428 (N_6428,N_6337,N_6305);
xor U6429 (N_6429,N_6313,N_6375);
nor U6430 (N_6430,N_6371,N_6329);
xnor U6431 (N_6431,N_6331,N_6378);
xor U6432 (N_6432,N_6372,N_6396);
and U6433 (N_6433,N_6303,N_6355);
and U6434 (N_6434,N_6389,N_6340);
and U6435 (N_6435,N_6385,N_6384);
or U6436 (N_6436,N_6336,N_6377);
nand U6437 (N_6437,N_6312,N_6317);
xnor U6438 (N_6438,N_6333,N_6353);
and U6439 (N_6439,N_6358,N_6326);
nand U6440 (N_6440,N_6395,N_6383);
nand U6441 (N_6441,N_6359,N_6394);
and U6442 (N_6442,N_6325,N_6328);
xor U6443 (N_6443,N_6321,N_6334);
xor U6444 (N_6444,N_6344,N_6339);
or U6445 (N_6445,N_6307,N_6357);
nand U6446 (N_6446,N_6338,N_6349);
or U6447 (N_6447,N_6382,N_6363);
nand U6448 (N_6448,N_6379,N_6376);
nand U6449 (N_6449,N_6354,N_6352);
or U6450 (N_6450,N_6386,N_6378);
or U6451 (N_6451,N_6381,N_6343);
and U6452 (N_6452,N_6372,N_6347);
and U6453 (N_6453,N_6342,N_6335);
xor U6454 (N_6454,N_6350,N_6346);
or U6455 (N_6455,N_6325,N_6311);
xor U6456 (N_6456,N_6347,N_6337);
nand U6457 (N_6457,N_6398,N_6358);
or U6458 (N_6458,N_6340,N_6374);
or U6459 (N_6459,N_6376,N_6302);
and U6460 (N_6460,N_6389,N_6399);
nor U6461 (N_6461,N_6323,N_6346);
or U6462 (N_6462,N_6311,N_6326);
or U6463 (N_6463,N_6345,N_6307);
nand U6464 (N_6464,N_6387,N_6363);
xnor U6465 (N_6465,N_6324,N_6335);
or U6466 (N_6466,N_6319,N_6337);
or U6467 (N_6467,N_6326,N_6382);
nor U6468 (N_6468,N_6336,N_6314);
and U6469 (N_6469,N_6380,N_6310);
xor U6470 (N_6470,N_6324,N_6393);
nor U6471 (N_6471,N_6390,N_6326);
and U6472 (N_6472,N_6374,N_6357);
nor U6473 (N_6473,N_6393,N_6358);
nor U6474 (N_6474,N_6333,N_6363);
and U6475 (N_6475,N_6396,N_6311);
xnor U6476 (N_6476,N_6352,N_6377);
and U6477 (N_6477,N_6392,N_6358);
or U6478 (N_6478,N_6302,N_6392);
nor U6479 (N_6479,N_6347,N_6377);
nand U6480 (N_6480,N_6346,N_6353);
nor U6481 (N_6481,N_6334,N_6319);
nor U6482 (N_6482,N_6335,N_6392);
xor U6483 (N_6483,N_6323,N_6318);
nor U6484 (N_6484,N_6316,N_6318);
nor U6485 (N_6485,N_6315,N_6349);
and U6486 (N_6486,N_6330,N_6335);
nor U6487 (N_6487,N_6340,N_6361);
nand U6488 (N_6488,N_6353,N_6342);
nor U6489 (N_6489,N_6357,N_6371);
nand U6490 (N_6490,N_6306,N_6327);
nand U6491 (N_6491,N_6365,N_6331);
or U6492 (N_6492,N_6396,N_6357);
nand U6493 (N_6493,N_6306,N_6355);
or U6494 (N_6494,N_6388,N_6310);
nor U6495 (N_6495,N_6367,N_6392);
xnor U6496 (N_6496,N_6379,N_6393);
nor U6497 (N_6497,N_6367,N_6372);
or U6498 (N_6498,N_6314,N_6398);
and U6499 (N_6499,N_6339,N_6361);
or U6500 (N_6500,N_6459,N_6479);
xor U6501 (N_6501,N_6488,N_6444);
or U6502 (N_6502,N_6422,N_6456);
xnor U6503 (N_6503,N_6427,N_6471);
or U6504 (N_6504,N_6436,N_6421);
nand U6505 (N_6505,N_6498,N_6496);
nor U6506 (N_6506,N_6424,N_6438);
and U6507 (N_6507,N_6454,N_6484);
or U6508 (N_6508,N_6453,N_6475);
or U6509 (N_6509,N_6435,N_6426);
xor U6510 (N_6510,N_6463,N_6461);
xnor U6511 (N_6511,N_6474,N_6442);
xor U6512 (N_6512,N_6400,N_6465);
and U6513 (N_6513,N_6440,N_6443);
xnor U6514 (N_6514,N_6493,N_6486);
or U6515 (N_6515,N_6416,N_6457);
xor U6516 (N_6516,N_6429,N_6450);
or U6517 (N_6517,N_6476,N_6412);
nor U6518 (N_6518,N_6495,N_6418);
xnor U6519 (N_6519,N_6439,N_6462);
or U6520 (N_6520,N_6428,N_6409);
or U6521 (N_6521,N_6464,N_6452);
or U6522 (N_6522,N_6490,N_6455);
nor U6523 (N_6523,N_6437,N_6472);
nor U6524 (N_6524,N_6415,N_6413);
nor U6525 (N_6525,N_6478,N_6404);
xnor U6526 (N_6526,N_6410,N_6485);
and U6527 (N_6527,N_6467,N_6403);
and U6528 (N_6528,N_6497,N_6458);
nor U6529 (N_6529,N_6477,N_6447);
xnor U6530 (N_6530,N_6420,N_6492);
nand U6531 (N_6531,N_6417,N_6448);
or U6532 (N_6532,N_6430,N_6460);
xor U6533 (N_6533,N_6433,N_6431);
and U6534 (N_6534,N_6470,N_6408);
xnor U6535 (N_6535,N_6407,N_6499);
and U6536 (N_6536,N_6451,N_6466);
nand U6537 (N_6537,N_6449,N_6445);
and U6538 (N_6538,N_6468,N_6482);
and U6539 (N_6539,N_6441,N_6483);
and U6540 (N_6540,N_6423,N_6401);
and U6541 (N_6541,N_6405,N_6425);
xnor U6542 (N_6542,N_6480,N_6491);
nor U6543 (N_6543,N_6406,N_6481);
and U6544 (N_6544,N_6494,N_6414);
and U6545 (N_6545,N_6469,N_6446);
and U6546 (N_6546,N_6432,N_6434);
and U6547 (N_6547,N_6489,N_6402);
nand U6548 (N_6548,N_6419,N_6487);
nor U6549 (N_6549,N_6411,N_6473);
xor U6550 (N_6550,N_6416,N_6430);
and U6551 (N_6551,N_6487,N_6421);
and U6552 (N_6552,N_6492,N_6494);
and U6553 (N_6553,N_6479,N_6422);
nand U6554 (N_6554,N_6437,N_6462);
or U6555 (N_6555,N_6435,N_6434);
xor U6556 (N_6556,N_6457,N_6497);
nand U6557 (N_6557,N_6473,N_6418);
nand U6558 (N_6558,N_6422,N_6464);
or U6559 (N_6559,N_6403,N_6410);
or U6560 (N_6560,N_6403,N_6491);
and U6561 (N_6561,N_6463,N_6487);
or U6562 (N_6562,N_6431,N_6404);
or U6563 (N_6563,N_6476,N_6478);
or U6564 (N_6564,N_6430,N_6422);
or U6565 (N_6565,N_6447,N_6457);
nand U6566 (N_6566,N_6471,N_6472);
or U6567 (N_6567,N_6489,N_6471);
nor U6568 (N_6568,N_6447,N_6463);
or U6569 (N_6569,N_6473,N_6440);
nor U6570 (N_6570,N_6408,N_6455);
nor U6571 (N_6571,N_6483,N_6479);
and U6572 (N_6572,N_6482,N_6428);
nor U6573 (N_6573,N_6486,N_6432);
xnor U6574 (N_6574,N_6417,N_6440);
or U6575 (N_6575,N_6482,N_6457);
xor U6576 (N_6576,N_6438,N_6469);
and U6577 (N_6577,N_6445,N_6415);
nand U6578 (N_6578,N_6477,N_6444);
nor U6579 (N_6579,N_6474,N_6413);
nor U6580 (N_6580,N_6498,N_6474);
nand U6581 (N_6581,N_6409,N_6440);
or U6582 (N_6582,N_6450,N_6412);
and U6583 (N_6583,N_6471,N_6434);
nor U6584 (N_6584,N_6496,N_6432);
nand U6585 (N_6585,N_6461,N_6493);
or U6586 (N_6586,N_6479,N_6402);
nand U6587 (N_6587,N_6440,N_6464);
and U6588 (N_6588,N_6499,N_6473);
xnor U6589 (N_6589,N_6494,N_6473);
and U6590 (N_6590,N_6415,N_6417);
xnor U6591 (N_6591,N_6431,N_6443);
nor U6592 (N_6592,N_6418,N_6409);
and U6593 (N_6593,N_6455,N_6481);
or U6594 (N_6594,N_6409,N_6408);
xor U6595 (N_6595,N_6428,N_6405);
and U6596 (N_6596,N_6499,N_6409);
nor U6597 (N_6597,N_6494,N_6412);
nor U6598 (N_6598,N_6452,N_6405);
nor U6599 (N_6599,N_6420,N_6445);
xnor U6600 (N_6600,N_6524,N_6541);
and U6601 (N_6601,N_6554,N_6561);
xor U6602 (N_6602,N_6560,N_6574);
xnor U6603 (N_6603,N_6505,N_6550);
and U6604 (N_6604,N_6523,N_6581);
nand U6605 (N_6605,N_6519,N_6573);
xnor U6606 (N_6606,N_6528,N_6544);
nand U6607 (N_6607,N_6587,N_6527);
or U6608 (N_6608,N_6545,N_6580);
nor U6609 (N_6609,N_6534,N_6584);
nor U6610 (N_6610,N_6552,N_6532);
and U6611 (N_6611,N_6563,N_6502);
and U6612 (N_6612,N_6586,N_6595);
and U6613 (N_6613,N_6509,N_6510);
or U6614 (N_6614,N_6596,N_6521);
xnor U6615 (N_6615,N_6514,N_6522);
nand U6616 (N_6616,N_6533,N_6513);
nand U6617 (N_6617,N_6537,N_6501);
nor U6618 (N_6618,N_6559,N_6568);
or U6619 (N_6619,N_6548,N_6593);
and U6620 (N_6620,N_6531,N_6577);
xor U6621 (N_6621,N_6578,N_6590);
nor U6622 (N_6622,N_6536,N_6538);
xnor U6623 (N_6623,N_6557,N_6582);
nand U6624 (N_6624,N_6535,N_6506);
and U6625 (N_6625,N_6575,N_6551);
and U6626 (N_6626,N_6504,N_6585);
or U6627 (N_6627,N_6549,N_6576);
or U6628 (N_6628,N_6529,N_6567);
nand U6629 (N_6629,N_6571,N_6597);
nor U6630 (N_6630,N_6598,N_6555);
nand U6631 (N_6631,N_6547,N_6583);
nor U6632 (N_6632,N_6507,N_6539);
xor U6633 (N_6633,N_6518,N_6594);
xor U6634 (N_6634,N_6540,N_6520);
nand U6635 (N_6635,N_6525,N_6565);
xnor U6636 (N_6636,N_6566,N_6508);
xnor U6637 (N_6637,N_6579,N_6543);
nor U6638 (N_6638,N_6564,N_6542);
nand U6639 (N_6639,N_6503,N_6589);
nor U6640 (N_6640,N_6588,N_6530);
and U6641 (N_6641,N_6562,N_6553);
or U6642 (N_6642,N_6515,N_6570);
and U6643 (N_6643,N_6592,N_6599);
or U6644 (N_6644,N_6558,N_6516);
and U6645 (N_6645,N_6517,N_6512);
and U6646 (N_6646,N_6591,N_6569);
xnor U6647 (N_6647,N_6526,N_6546);
xnor U6648 (N_6648,N_6572,N_6556);
nand U6649 (N_6649,N_6500,N_6511);
xnor U6650 (N_6650,N_6513,N_6572);
xor U6651 (N_6651,N_6585,N_6501);
nand U6652 (N_6652,N_6503,N_6532);
nor U6653 (N_6653,N_6570,N_6517);
xor U6654 (N_6654,N_6500,N_6591);
or U6655 (N_6655,N_6537,N_6520);
and U6656 (N_6656,N_6582,N_6546);
nor U6657 (N_6657,N_6588,N_6551);
nor U6658 (N_6658,N_6506,N_6551);
nand U6659 (N_6659,N_6590,N_6573);
xor U6660 (N_6660,N_6547,N_6549);
nand U6661 (N_6661,N_6589,N_6569);
xnor U6662 (N_6662,N_6509,N_6562);
and U6663 (N_6663,N_6539,N_6581);
nor U6664 (N_6664,N_6524,N_6506);
nor U6665 (N_6665,N_6593,N_6570);
xor U6666 (N_6666,N_6576,N_6571);
nor U6667 (N_6667,N_6531,N_6515);
nand U6668 (N_6668,N_6570,N_6506);
nand U6669 (N_6669,N_6540,N_6538);
or U6670 (N_6670,N_6543,N_6504);
and U6671 (N_6671,N_6571,N_6585);
and U6672 (N_6672,N_6590,N_6529);
nand U6673 (N_6673,N_6588,N_6589);
nor U6674 (N_6674,N_6570,N_6559);
and U6675 (N_6675,N_6511,N_6580);
nand U6676 (N_6676,N_6550,N_6527);
or U6677 (N_6677,N_6568,N_6579);
nor U6678 (N_6678,N_6571,N_6543);
or U6679 (N_6679,N_6513,N_6537);
nand U6680 (N_6680,N_6594,N_6564);
and U6681 (N_6681,N_6538,N_6532);
nand U6682 (N_6682,N_6544,N_6565);
nand U6683 (N_6683,N_6510,N_6556);
xor U6684 (N_6684,N_6576,N_6557);
nor U6685 (N_6685,N_6538,N_6570);
and U6686 (N_6686,N_6548,N_6509);
or U6687 (N_6687,N_6513,N_6589);
nand U6688 (N_6688,N_6546,N_6503);
xor U6689 (N_6689,N_6585,N_6578);
and U6690 (N_6690,N_6540,N_6544);
xor U6691 (N_6691,N_6561,N_6599);
and U6692 (N_6692,N_6580,N_6575);
xor U6693 (N_6693,N_6574,N_6572);
nand U6694 (N_6694,N_6523,N_6583);
nand U6695 (N_6695,N_6525,N_6522);
nor U6696 (N_6696,N_6578,N_6549);
nand U6697 (N_6697,N_6597,N_6529);
nor U6698 (N_6698,N_6595,N_6594);
xor U6699 (N_6699,N_6554,N_6562);
nand U6700 (N_6700,N_6610,N_6655);
nand U6701 (N_6701,N_6654,N_6641);
or U6702 (N_6702,N_6609,N_6639);
nor U6703 (N_6703,N_6624,N_6640);
and U6704 (N_6704,N_6684,N_6662);
or U6705 (N_6705,N_6633,N_6607);
or U6706 (N_6706,N_6623,N_6658);
nor U6707 (N_6707,N_6629,N_6645);
nor U6708 (N_6708,N_6697,N_6665);
nand U6709 (N_6709,N_6614,N_6671);
and U6710 (N_6710,N_6634,N_6668);
and U6711 (N_6711,N_6657,N_6622);
and U6712 (N_6712,N_6601,N_6648);
or U6713 (N_6713,N_6660,N_6667);
nand U6714 (N_6714,N_6625,N_6600);
nor U6715 (N_6715,N_6675,N_6682);
nand U6716 (N_6716,N_6687,N_6694);
nor U6717 (N_6717,N_6652,N_6632);
or U6718 (N_6718,N_6683,N_6613);
nor U6719 (N_6719,N_6647,N_6678);
nor U6720 (N_6720,N_6685,N_6619);
and U6721 (N_6721,N_6664,N_6692);
and U6722 (N_6722,N_6656,N_6650);
nand U6723 (N_6723,N_6602,N_6680);
and U6724 (N_6724,N_6626,N_6611);
and U6725 (N_6725,N_6688,N_6676);
or U6726 (N_6726,N_6666,N_6642);
xnor U6727 (N_6727,N_6698,N_6679);
or U6728 (N_6728,N_6699,N_6603);
nand U6729 (N_6729,N_6627,N_6659);
xnor U6730 (N_6730,N_6643,N_6612);
or U6731 (N_6731,N_6628,N_6661);
nor U6732 (N_6732,N_6673,N_6638);
nor U6733 (N_6733,N_6606,N_6631);
nand U6734 (N_6734,N_6674,N_6690);
xnor U6735 (N_6735,N_6691,N_6646);
nand U6736 (N_6736,N_6637,N_6681);
or U6737 (N_6737,N_6630,N_6621);
or U6738 (N_6738,N_6644,N_6649);
nand U6739 (N_6739,N_6669,N_6672);
or U6740 (N_6740,N_6651,N_6604);
nor U6741 (N_6741,N_6616,N_6615);
or U6742 (N_6742,N_6605,N_6686);
nor U6743 (N_6743,N_6635,N_6618);
nand U6744 (N_6744,N_6689,N_6608);
nand U6745 (N_6745,N_6693,N_6653);
xnor U6746 (N_6746,N_6677,N_6663);
and U6747 (N_6747,N_6695,N_6670);
and U6748 (N_6748,N_6696,N_6636);
nor U6749 (N_6749,N_6620,N_6617);
xnor U6750 (N_6750,N_6621,N_6666);
nand U6751 (N_6751,N_6654,N_6622);
xor U6752 (N_6752,N_6639,N_6659);
xnor U6753 (N_6753,N_6679,N_6690);
nor U6754 (N_6754,N_6659,N_6633);
and U6755 (N_6755,N_6682,N_6672);
nand U6756 (N_6756,N_6669,N_6613);
nand U6757 (N_6757,N_6614,N_6634);
nor U6758 (N_6758,N_6624,N_6681);
xor U6759 (N_6759,N_6678,N_6641);
nor U6760 (N_6760,N_6637,N_6624);
or U6761 (N_6761,N_6652,N_6607);
or U6762 (N_6762,N_6673,N_6620);
nor U6763 (N_6763,N_6614,N_6677);
xnor U6764 (N_6764,N_6678,N_6673);
nor U6765 (N_6765,N_6680,N_6660);
xor U6766 (N_6766,N_6647,N_6668);
and U6767 (N_6767,N_6609,N_6644);
or U6768 (N_6768,N_6677,N_6637);
or U6769 (N_6769,N_6612,N_6631);
or U6770 (N_6770,N_6675,N_6695);
nand U6771 (N_6771,N_6635,N_6615);
nor U6772 (N_6772,N_6640,N_6634);
nand U6773 (N_6773,N_6672,N_6649);
xor U6774 (N_6774,N_6650,N_6604);
or U6775 (N_6775,N_6660,N_6600);
and U6776 (N_6776,N_6662,N_6639);
xnor U6777 (N_6777,N_6689,N_6606);
nand U6778 (N_6778,N_6608,N_6686);
or U6779 (N_6779,N_6686,N_6690);
or U6780 (N_6780,N_6630,N_6637);
or U6781 (N_6781,N_6687,N_6602);
and U6782 (N_6782,N_6614,N_6685);
nand U6783 (N_6783,N_6635,N_6662);
nand U6784 (N_6784,N_6607,N_6663);
nor U6785 (N_6785,N_6663,N_6661);
and U6786 (N_6786,N_6675,N_6652);
nand U6787 (N_6787,N_6606,N_6637);
or U6788 (N_6788,N_6607,N_6619);
xor U6789 (N_6789,N_6638,N_6625);
and U6790 (N_6790,N_6634,N_6696);
nand U6791 (N_6791,N_6693,N_6610);
nand U6792 (N_6792,N_6601,N_6609);
or U6793 (N_6793,N_6641,N_6614);
xor U6794 (N_6794,N_6654,N_6694);
nand U6795 (N_6795,N_6630,N_6697);
and U6796 (N_6796,N_6631,N_6673);
nand U6797 (N_6797,N_6644,N_6672);
nand U6798 (N_6798,N_6602,N_6612);
xnor U6799 (N_6799,N_6636,N_6614);
nand U6800 (N_6800,N_6739,N_6722);
nor U6801 (N_6801,N_6703,N_6700);
or U6802 (N_6802,N_6759,N_6701);
nor U6803 (N_6803,N_6758,N_6719);
or U6804 (N_6804,N_6786,N_6751);
and U6805 (N_6805,N_6709,N_6710);
nor U6806 (N_6806,N_6728,N_6782);
nor U6807 (N_6807,N_6732,N_6793);
nand U6808 (N_6808,N_6725,N_6715);
nand U6809 (N_6809,N_6778,N_6717);
nor U6810 (N_6810,N_6761,N_6738);
and U6811 (N_6811,N_6727,N_6757);
nand U6812 (N_6812,N_6718,N_6784);
nand U6813 (N_6813,N_6705,N_6762);
and U6814 (N_6814,N_6796,N_6797);
xnor U6815 (N_6815,N_6737,N_6733);
or U6816 (N_6816,N_6744,N_6734);
xnor U6817 (N_6817,N_6724,N_6736);
or U6818 (N_6818,N_6706,N_6772);
or U6819 (N_6819,N_6735,N_6794);
and U6820 (N_6820,N_6765,N_6798);
nand U6821 (N_6821,N_6752,N_6767);
nand U6822 (N_6822,N_6774,N_6766);
or U6823 (N_6823,N_6750,N_6747);
and U6824 (N_6824,N_6776,N_6771);
nor U6825 (N_6825,N_6729,N_6777);
and U6826 (N_6826,N_6783,N_6779);
nand U6827 (N_6827,N_6788,N_6742);
or U6828 (N_6828,N_6769,N_6712);
nor U6829 (N_6829,N_6799,N_6789);
nor U6830 (N_6830,N_6763,N_6708);
nor U6831 (N_6831,N_6768,N_6731);
xor U6832 (N_6832,N_6780,N_6764);
and U6833 (N_6833,N_6730,N_6723);
xnor U6834 (N_6834,N_6721,N_6745);
nand U6835 (N_6835,N_6741,N_6773);
nand U6836 (N_6836,N_6726,N_6702);
xor U6837 (N_6837,N_6748,N_6756);
xnor U6838 (N_6838,N_6791,N_6740);
nand U6839 (N_6839,N_6746,N_6720);
xnor U6840 (N_6840,N_6753,N_6743);
nor U6841 (N_6841,N_6787,N_6790);
nand U6842 (N_6842,N_6714,N_6704);
xor U6843 (N_6843,N_6775,N_6754);
xnor U6844 (N_6844,N_6770,N_6785);
nor U6845 (N_6845,N_6795,N_6713);
or U6846 (N_6846,N_6792,N_6707);
nor U6847 (N_6847,N_6749,N_6755);
and U6848 (N_6848,N_6716,N_6781);
nor U6849 (N_6849,N_6711,N_6760);
or U6850 (N_6850,N_6741,N_6783);
nor U6851 (N_6851,N_6704,N_6734);
nor U6852 (N_6852,N_6708,N_6740);
or U6853 (N_6853,N_6728,N_6761);
nand U6854 (N_6854,N_6752,N_6748);
xnor U6855 (N_6855,N_6734,N_6770);
xnor U6856 (N_6856,N_6735,N_6770);
or U6857 (N_6857,N_6739,N_6735);
nand U6858 (N_6858,N_6750,N_6772);
and U6859 (N_6859,N_6718,N_6739);
xnor U6860 (N_6860,N_6759,N_6732);
nand U6861 (N_6861,N_6726,N_6705);
xor U6862 (N_6862,N_6796,N_6769);
or U6863 (N_6863,N_6790,N_6796);
or U6864 (N_6864,N_6787,N_6797);
nand U6865 (N_6865,N_6773,N_6747);
or U6866 (N_6866,N_6758,N_6779);
xnor U6867 (N_6867,N_6768,N_6700);
nand U6868 (N_6868,N_6796,N_6723);
nand U6869 (N_6869,N_6786,N_6716);
or U6870 (N_6870,N_6719,N_6706);
or U6871 (N_6871,N_6704,N_6702);
nor U6872 (N_6872,N_6714,N_6756);
xnor U6873 (N_6873,N_6704,N_6725);
and U6874 (N_6874,N_6752,N_6782);
and U6875 (N_6875,N_6757,N_6737);
or U6876 (N_6876,N_6703,N_6713);
and U6877 (N_6877,N_6768,N_6726);
and U6878 (N_6878,N_6730,N_6720);
nor U6879 (N_6879,N_6706,N_6745);
nor U6880 (N_6880,N_6740,N_6741);
or U6881 (N_6881,N_6758,N_6723);
nand U6882 (N_6882,N_6720,N_6761);
nand U6883 (N_6883,N_6775,N_6730);
nor U6884 (N_6884,N_6774,N_6779);
and U6885 (N_6885,N_6784,N_6728);
and U6886 (N_6886,N_6763,N_6718);
xor U6887 (N_6887,N_6780,N_6797);
or U6888 (N_6888,N_6701,N_6735);
nor U6889 (N_6889,N_6780,N_6755);
and U6890 (N_6890,N_6793,N_6725);
nand U6891 (N_6891,N_6781,N_6715);
nor U6892 (N_6892,N_6744,N_6710);
nor U6893 (N_6893,N_6799,N_6763);
xnor U6894 (N_6894,N_6727,N_6782);
and U6895 (N_6895,N_6772,N_6713);
nand U6896 (N_6896,N_6749,N_6798);
or U6897 (N_6897,N_6702,N_6732);
nor U6898 (N_6898,N_6764,N_6709);
xor U6899 (N_6899,N_6735,N_6752);
nand U6900 (N_6900,N_6856,N_6843);
and U6901 (N_6901,N_6861,N_6830);
xor U6902 (N_6902,N_6823,N_6842);
xnor U6903 (N_6903,N_6837,N_6857);
xnor U6904 (N_6904,N_6893,N_6800);
or U6905 (N_6905,N_6824,N_6812);
and U6906 (N_6906,N_6895,N_6816);
nand U6907 (N_6907,N_6880,N_6885);
nor U6908 (N_6908,N_6834,N_6873);
nand U6909 (N_6909,N_6896,N_6858);
and U6910 (N_6910,N_6839,N_6831);
nand U6911 (N_6911,N_6818,N_6892);
nand U6912 (N_6912,N_6815,N_6869);
or U6913 (N_6913,N_6810,N_6864);
xnor U6914 (N_6914,N_6886,N_6868);
nand U6915 (N_6915,N_6891,N_6820);
nor U6916 (N_6916,N_6840,N_6870);
or U6917 (N_6917,N_6887,N_6883);
or U6918 (N_6918,N_6898,N_6803);
xnor U6919 (N_6919,N_6836,N_6855);
nand U6920 (N_6920,N_6809,N_6849);
nand U6921 (N_6921,N_6850,N_6890);
nor U6922 (N_6922,N_6827,N_6806);
xnor U6923 (N_6923,N_6835,N_6841);
and U6924 (N_6924,N_6872,N_6814);
nor U6925 (N_6925,N_6807,N_6882);
xnor U6926 (N_6926,N_6899,N_6860);
and U6927 (N_6927,N_6889,N_6833);
nand U6928 (N_6928,N_6829,N_6862);
and U6929 (N_6929,N_6875,N_6813);
nand U6930 (N_6930,N_6838,N_6876);
xnor U6931 (N_6931,N_6867,N_6863);
xor U6932 (N_6932,N_6846,N_6804);
nor U6933 (N_6933,N_6805,N_6811);
nor U6934 (N_6934,N_6865,N_6821);
and U6935 (N_6935,N_6874,N_6844);
nor U6936 (N_6936,N_6884,N_6847);
or U6937 (N_6937,N_6866,N_6879);
xor U6938 (N_6938,N_6881,N_6828);
nand U6939 (N_6939,N_6852,N_6854);
xnor U6940 (N_6940,N_6802,N_6825);
nand U6941 (N_6941,N_6832,N_6897);
xor U6942 (N_6942,N_6845,N_6859);
and U6943 (N_6943,N_6871,N_6808);
xnor U6944 (N_6944,N_6878,N_6817);
and U6945 (N_6945,N_6822,N_6877);
or U6946 (N_6946,N_6894,N_6888);
xnor U6947 (N_6947,N_6826,N_6853);
nor U6948 (N_6948,N_6819,N_6848);
nand U6949 (N_6949,N_6851,N_6801);
nor U6950 (N_6950,N_6832,N_6818);
and U6951 (N_6951,N_6849,N_6854);
xor U6952 (N_6952,N_6815,N_6854);
xnor U6953 (N_6953,N_6896,N_6869);
or U6954 (N_6954,N_6891,N_6869);
or U6955 (N_6955,N_6815,N_6857);
and U6956 (N_6956,N_6876,N_6820);
or U6957 (N_6957,N_6872,N_6850);
nand U6958 (N_6958,N_6811,N_6817);
nand U6959 (N_6959,N_6889,N_6804);
and U6960 (N_6960,N_6886,N_6897);
nand U6961 (N_6961,N_6859,N_6876);
nand U6962 (N_6962,N_6881,N_6807);
and U6963 (N_6963,N_6838,N_6833);
and U6964 (N_6964,N_6872,N_6861);
nand U6965 (N_6965,N_6823,N_6851);
and U6966 (N_6966,N_6847,N_6889);
and U6967 (N_6967,N_6896,N_6823);
and U6968 (N_6968,N_6832,N_6831);
nor U6969 (N_6969,N_6869,N_6833);
and U6970 (N_6970,N_6846,N_6837);
or U6971 (N_6971,N_6860,N_6897);
nand U6972 (N_6972,N_6858,N_6838);
nand U6973 (N_6973,N_6893,N_6806);
and U6974 (N_6974,N_6806,N_6839);
xnor U6975 (N_6975,N_6854,N_6872);
nand U6976 (N_6976,N_6863,N_6890);
nand U6977 (N_6977,N_6828,N_6886);
nand U6978 (N_6978,N_6849,N_6873);
xor U6979 (N_6979,N_6890,N_6844);
nor U6980 (N_6980,N_6839,N_6812);
and U6981 (N_6981,N_6828,N_6896);
or U6982 (N_6982,N_6801,N_6815);
and U6983 (N_6983,N_6831,N_6801);
nand U6984 (N_6984,N_6857,N_6875);
nand U6985 (N_6985,N_6815,N_6891);
nor U6986 (N_6986,N_6835,N_6898);
or U6987 (N_6987,N_6859,N_6870);
xor U6988 (N_6988,N_6865,N_6892);
nand U6989 (N_6989,N_6873,N_6828);
or U6990 (N_6990,N_6816,N_6829);
xor U6991 (N_6991,N_6846,N_6849);
nor U6992 (N_6992,N_6888,N_6843);
xor U6993 (N_6993,N_6896,N_6829);
and U6994 (N_6994,N_6876,N_6888);
or U6995 (N_6995,N_6880,N_6888);
nor U6996 (N_6996,N_6894,N_6824);
xor U6997 (N_6997,N_6872,N_6822);
or U6998 (N_6998,N_6834,N_6868);
nand U6999 (N_6999,N_6867,N_6864);
nand U7000 (N_7000,N_6999,N_6983);
and U7001 (N_7001,N_6903,N_6922);
nand U7002 (N_7002,N_6908,N_6995);
nor U7003 (N_7003,N_6915,N_6941);
or U7004 (N_7004,N_6998,N_6986);
and U7005 (N_7005,N_6947,N_6921);
nor U7006 (N_7006,N_6914,N_6967);
or U7007 (N_7007,N_6969,N_6926);
nor U7008 (N_7008,N_6989,N_6976);
and U7009 (N_7009,N_6979,N_6959);
and U7010 (N_7010,N_6997,N_6945);
or U7011 (N_7011,N_6980,N_6900);
nor U7012 (N_7012,N_6933,N_6958);
nor U7013 (N_7013,N_6906,N_6990);
and U7014 (N_7014,N_6910,N_6974);
nor U7015 (N_7015,N_6975,N_6918);
xnor U7016 (N_7016,N_6988,N_6909);
xor U7017 (N_7017,N_6902,N_6984);
and U7018 (N_7018,N_6951,N_6964);
nor U7019 (N_7019,N_6977,N_6911);
xnor U7020 (N_7020,N_6907,N_6928);
xor U7021 (N_7021,N_6935,N_6973);
nand U7022 (N_7022,N_6904,N_6923);
or U7023 (N_7023,N_6913,N_6978);
or U7024 (N_7024,N_6962,N_6938);
nand U7025 (N_7025,N_6960,N_6929);
xnor U7026 (N_7026,N_6931,N_6965);
nor U7027 (N_7027,N_6963,N_6919);
xnor U7028 (N_7028,N_6982,N_6985);
or U7029 (N_7029,N_6981,N_6992);
nor U7030 (N_7030,N_6942,N_6944);
or U7031 (N_7031,N_6936,N_6972);
and U7032 (N_7032,N_6952,N_6956);
or U7033 (N_7033,N_6920,N_6993);
xnor U7034 (N_7034,N_6991,N_6954);
xnor U7035 (N_7035,N_6994,N_6939);
and U7036 (N_7036,N_6940,N_6955);
xnor U7037 (N_7037,N_6901,N_6971);
and U7038 (N_7038,N_6966,N_6905);
nor U7039 (N_7039,N_6930,N_6948);
and U7040 (N_7040,N_6937,N_6949);
xor U7041 (N_7041,N_6927,N_6925);
nor U7042 (N_7042,N_6917,N_6961);
nand U7043 (N_7043,N_6912,N_6957);
and U7044 (N_7044,N_6968,N_6953);
xor U7045 (N_7045,N_6932,N_6924);
nor U7046 (N_7046,N_6934,N_6996);
and U7047 (N_7047,N_6950,N_6987);
nand U7048 (N_7048,N_6943,N_6970);
nor U7049 (N_7049,N_6916,N_6946);
nand U7050 (N_7050,N_6969,N_6948);
nand U7051 (N_7051,N_6982,N_6988);
and U7052 (N_7052,N_6965,N_6949);
xor U7053 (N_7053,N_6918,N_6969);
or U7054 (N_7054,N_6945,N_6957);
and U7055 (N_7055,N_6943,N_6945);
and U7056 (N_7056,N_6958,N_6964);
nor U7057 (N_7057,N_6942,N_6956);
nor U7058 (N_7058,N_6985,N_6906);
nand U7059 (N_7059,N_6946,N_6984);
nand U7060 (N_7060,N_6977,N_6995);
xor U7061 (N_7061,N_6997,N_6979);
or U7062 (N_7062,N_6963,N_6905);
or U7063 (N_7063,N_6997,N_6960);
nor U7064 (N_7064,N_6946,N_6985);
or U7065 (N_7065,N_6947,N_6901);
and U7066 (N_7066,N_6913,N_6966);
nor U7067 (N_7067,N_6952,N_6997);
xnor U7068 (N_7068,N_6978,N_6988);
and U7069 (N_7069,N_6916,N_6957);
or U7070 (N_7070,N_6968,N_6908);
or U7071 (N_7071,N_6943,N_6988);
xnor U7072 (N_7072,N_6971,N_6932);
nor U7073 (N_7073,N_6918,N_6931);
xor U7074 (N_7074,N_6978,N_6919);
nand U7075 (N_7075,N_6938,N_6934);
nor U7076 (N_7076,N_6934,N_6943);
nand U7077 (N_7077,N_6956,N_6938);
and U7078 (N_7078,N_6908,N_6925);
nor U7079 (N_7079,N_6962,N_6984);
xor U7080 (N_7080,N_6957,N_6994);
nand U7081 (N_7081,N_6981,N_6954);
and U7082 (N_7082,N_6965,N_6925);
nor U7083 (N_7083,N_6997,N_6992);
xnor U7084 (N_7084,N_6905,N_6914);
nand U7085 (N_7085,N_6990,N_6907);
or U7086 (N_7086,N_6970,N_6986);
or U7087 (N_7087,N_6926,N_6959);
xnor U7088 (N_7088,N_6971,N_6998);
xor U7089 (N_7089,N_6904,N_6981);
nor U7090 (N_7090,N_6955,N_6975);
and U7091 (N_7091,N_6935,N_6914);
nor U7092 (N_7092,N_6961,N_6963);
xor U7093 (N_7093,N_6992,N_6998);
nor U7094 (N_7094,N_6918,N_6977);
xor U7095 (N_7095,N_6946,N_6908);
nor U7096 (N_7096,N_6919,N_6959);
xnor U7097 (N_7097,N_6941,N_6926);
and U7098 (N_7098,N_6910,N_6993);
and U7099 (N_7099,N_6990,N_6916);
or U7100 (N_7100,N_7039,N_7049);
nor U7101 (N_7101,N_7069,N_7021);
nor U7102 (N_7102,N_7057,N_7001);
xnor U7103 (N_7103,N_7036,N_7009);
nor U7104 (N_7104,N_7077,N_7025);
or U7105 (N_7105,N_7080,N_7048);
xor U7106 (N_7106,N_7033,N_7086);
nand U7107 (N_7107,N_7040,N_7059);
nor U7108 (N_7108,N_7089,N_7075);
nand U7109 (N_7109,N_7004,N_7045);
nor U7110 (N_7110,N_7019,N_7041);
and U7111 (N_7111,N_7097,N_7098);
and U7112 (N_7112,N_7003,N_7081);
nand U7113 (N_7113,N_7034,N_7068);
and U7114 (N_7114,N_7099,N_7029);
xor U7115 (N_7115,N_7007,N_7060);
or U7116 (N_7116,N_7066,N_7076);
or U7117 (N_7117,N_7042,N_7010);
and U7118 (N_7118,N_7022,N_7017);
nand U7119 (N_7119,N_7074,N_7043);
nor U7120 (N_7120,N_7064,N_7037);
xor U7121 (N_7121,N_7054,N_7024);
xor U7122 (N_7122,N_7005,N_7084);
and U7123 (N_7123,N_7056,N_7093);
nor U7124 (N_7124,N_7061,N_7006);
and U7125 (N_7125,N_7065,N_7027);
xor U7126 (N_7126,N_7031,N_7008);
xnor U7127 (N_7127,N_7002,N_7011);
nand U7128 (N_7128,N_7058,N_7015);
nand U7129 (N_7129,N_7090,N_7083);
nor U7130 (N_7130,N_7073,N_7053);
xor U7131 (N_7131,N_7062,N_7088);
nand U7132 (N_7132,N_7091,N_7085);
xnor U7133 (N_7133,N_7020,N_7072);
nand U7134 (N_7134,N_7030,N_7050);
nor U7135 (N_7135,N_7023,N_7087);
or U7136 (N_7136,N_7044,N_7018);
xnor U7137 (N_7137,N_7000,N_7035);
and U7138 (N_7138,N_7047,N_7013);
and U7139 (N_7139,N_7026,N_7051);
nand U7140 (N_7140,N_7055,N_7063);
nand U7141 (N_7141,N_7095,N_7038);
nor U7142 (N_7142,N_7082,N_7046);
and U7143 (N_7143,N_7028,N_7092);
and U7144 (N_7144,N_7096,N_7070);
xnor U7145 (N_7145,N_7014,N_7071);
or U7146 (N_7146,N_7078,N_7094);
or U7147 (N_7147,N_7052,N_7032);
and U7148 (N_7148,N_7016,N_7067);
and U7149 (N_7149,N_7012,N_7079);
or U7150 (N_7150,N_7083,N_7059);
xor U7151 (N_7151,N_7037,N_7048);
or U7152 (N_7152,N_7066,N_7079);
or U7153 (N_7153,N_7053,N_7052);
nand U7154 (N_7154,N_7042,N_7009);
and U7155 (N_7155,N_7089,N_7018);
nor U7156 (N_7156,N_7047,N_7051);
and U7157 (N_7157,N_7082,N_7074);
and U7158 (N_7158,N_7051,N_7030);
or U7159 (N_7159,N_7036,N_7026);
nand U7160 (N_7160,N_7087,N_7054);
and U7161 (N_7161,N_7090,N_7061);
nand U7162 (N_7162,N_7045,N_7030);
nand U7163 (N_7163,N_7048,N_7040);
and U7164 (N_7164,N_7067,N_7018);
xnor U7165 (N_7165,N_7026,N_7050);
or U7166 (N_7166,N_7002,N_7056);
or U7167 (N_7167,N_7067,N_7023);
or U7168 (N_7168,N_7048,N_7058);
xnor U7169 (N_7169,N_7038,N_7015);
or U7170 (N_7170,N_7084,N_7067);
xor U7171 (N_7171,N_7094,N_7033);
nor U7172 (N_7172,N_7024,N_7077);
and U7173 (N_7173,N_7072,N_7005);
nand U7174 (N_7174,N_7032,N_7069);
nand U7175 (N_7175,N_7034,N_7027);
and U7176 (N_7176,N_7082,N_7004);
nand U7177 (N_7177,N_7026,N_7002);
nor U7178 (N_7178,N_7072,N_7066);
or U7179 (N_7179,N_7010,N_7006);
and U7180 (N_7180,N_7028,N_7002);
and U7181 (N_7181,N_7026,N_7065);
nor U7182 (N_7182,N_7037,N_7005);
nor U7183 (N_7183,N_7080,N_7011);
nand U7184 (N_7184,N_7002,N_7075);
nand U7185 (N_7185,N_7021,N_7064);
or U7186 (N_7186,N_7019,N_7026);
or U7187 (N_7187,N_7016,N_7069);
nor U7188 (N_7188,N_7038,N_7065);
xor U7189 (N_7189,N_7017,N_7099);
nand U7190 (N_7190,N_7043,N_7024);
and U7191 (N_7191,N_7037,N_7055);
and U7192 (N_7192,N_7074,N_7045);
and U7193 (N_7193,N_7017,N_7041);
and U7194 (N_7194,N_7008,N_7017);
nand U7195 (N_7195,N_7056,N_7005);
nor U7196 (N_7196,N_7002,N_7067);
xor U7197 (N_7197,N_7098,N_7089);
and U7198 (N_7198,N_7068,N_7072);
or U7199 (N_7199,N_7009,N_7073);
nor U7200 (N_7200,N_7164,N_7125);
nor U7201 (N_7201,N_7143,N_7152);
nand U7202 (N_7202,N_7139,N_7169);
nor U7203 (N_7203,N_7153,N_7172);
nor U7204 (N_7204,N_7106,N_7171);
and U7205 (N_7205,N_7199,N_7145);
nor U7206 (N_7206,N_7188,N_7194);
nand U7207 (N_7207,N_7185,N_7110);
nor U7208 (N_7208,N_7168,N_7177);
and U7209 (N_7209,N_7138,N_7118);
or U7210 (N_7210,N_7119,N_7173);
nor U7211 (N_7211,N_7197,N_7140);
or U7212 (N_7212,N_7127,N_7189);
xor U7213 (N_7213,N_7151,N_7186);
or U7214 (N_7214,N_7128,N_7192);
nand U7215 (N_7215,N_7112,N_7178);
nor U7216 (N_7216,N_7144,N_7108);
and U7217 (N_7217,N_7176,N_7123);
xor U7218 (N_7218,N_7102,N_7161);
nor U7219 (N_7219,N_7148,N_7103);
or U7220 (N_7220,N_7100,N_7154);
or U7221 (N_7221,N_7157,N_7158);
xnor U7222 (N_7222,N_7136,N_7124);
or U7223 (N_7223,N_7142,N_7162);
nor U7224 (N_7224,N_7149,N_7141);
and U7225 (N_7225,N_7134,N_7156);
nor U7226 (N_7226,N_7129,N_7196);
and U7227 (N_7227,N_7181,N_7160);
or U7228 (N_7228,N_7146,N_7126);
xnor U7229 (N_7229,N_7183,N_7150);
or U7230 (N_7230,N_7195,N_7120);
and U7231 (N_7231,N_7147,N_7105);
xnor U7232 (N_7232,N_7101,N_7184);
nand U7233 (N_7233,N_7165,N_7131);
or U7234 (N_7234,N_7111,N_7132);
nor U7235 (N_7235,N_7174,N_7115);
xor U7236 (N_7236,N_7130,N_7193);
nand U7237 (N_7237,N_7180,N_7182);
or U7238 (N_7238,N_7179,N_7109);
nand U7239 (N_7239,N_7122,N_7114);
xor U7240 (N_7240,N_7116,N_7170);
and U7241 (N_7241,N_7191,N_7104);
xnor U7242 (N_7242,N_7107,N_7163);
or U7243 (N_7243,N_7121,N_7167);
nand U7244 (N_7244,N_7113,N_7133);
xnor U7245 (N_7245,N_7198,N_7135);
nor U7246 (N_7246,N_7159,N_7166);
nor U7247 (N_7247,N_7137,N_7187);
or U7248 (N_7248,N_7175,N_7117);
nand U7249 (N_7249,N_7190,N_7155);
nor U7250 (N_7250,N_7186,N_7149);
nand U7251 (N_7251,N_7190,N_7180);
xor U7252 (N_7252,N_7165,N_7116);
and U7253 (N_7253,N_7171,N_7109);
nand U7254 (N_7254,N_7121,N_7125);
xnor U7255 (N_7255,N_7174,N_7109);
or U7256 (N_7256,N_7198,N_7103);
nand U7257 (N_7257,N_7182,N_7132);
or U7258 (N_7258,N_7157,N_7146);
xor U7259 (N_7259,N_7153,N_7155);
nand U7260 (N_7260,N_7116,N_7113);
or U7261 (N_7261,N_7125,N_7102);
xor U7262 (N_7262,N_7148,N_7119);
xnor U7263 (N_7263,N_7130,N_7170);
or U7264 (N_7264,N_7155,N_7129);
xnor U7265 (N_7265,N_7115,N_7170);
xor U7266 (N_7266,N_7182,N_7118);
and U7267 (N_7267,N_7149,N_7123);
or U7268 (N_7268,N_7142,N_7157);
or U7269 (N_7269,N_7130,N_7197);
xor U7270 (N_7270,N_7149,N_7104);
xor U7271 (N_7271,N_7160,N_7182);
nor U7272 (N_7272,N_7106,N_7130);
or U7273 (N_7273,N_7122,N_7157);
nor U7274 (N_7274,N_7178,N_7158);
and U7275 (N_7275,N_7156,N_7182);
or U7276 (N_7276,N_7151,N_7142);
nand U7277 (N_7277,N_7127,N_7128);
nor U7278 (N_7278,N_7138,N_7133);
xor U7279 (N_7279,N_7147,N_7176);
xor U7280 (N_7280,N_7102,N_7168);
nor U7281 (N_7281,N_7165,N_7112);
or U7282 (N_7282,N_7114,N_7176);
nor U7283 (N_7283,N_7130,N_7188);
nand U7284 (N_7284,N_7169,N_7168);
nand U7285 (N_7285,N_7194,N_7173);
and U7286 (N_7286,N_7141,N_7112);
nand U7287 (N_7287,N_7130,N_7149);
nand U7288 (N_7288,N_7159,N_7156);
xnor U7289 (N_7289,N_7129,N_7179);
or U7290 (N_7290,N_7125,N_7135);
nand U7291 (N_7291,N_7116,N_7127);
and U7292 (N_7292,N_7189,N_7185);
or U7293 (N_7293,N_7103,N_7150);
and U7294 (N_7294,N_7142,N_7198);
nand U7295 (N_7295,N_7116,N_7114);
and U7296 (N_7296,N_7158,N_7184);
nor U7297 (N_7297,N_7119,N_7123);
nand U7298 (N_7298,N_7173,N_7177);
and U7299 (N_7299,N_7141,N_7165);
xor U7300 (N_7300,N_7201,N_7294);
nand U7301 (N_7301,N_7210,N_7269);
and U7302 (N_7302,N_7263,N_7273);
and U7303 (N_7303,N_7249,N_7232);
nand U7304 (N_7304,N_7220,N_7254);
xor U7305 (N_7305,N_7258,N_7245);
nand U7306 (N_7306,N_7285,N_7222);
xnor U7307 (N_7307,N_7224,N_7225);
nand U7308 (N_7308,N_7290,N_7274);
nand U7309 (N_7309,N_7253,N_7241);
xor U7310 (N_7310,N_7239,N_7227);
xnor U7311 (N_7311,N_7287,N_7275);
xnor U7312 (N_7312,N_7212,N_7234);
and U7313 (N_7313,N_7236,N_7219);
xnor U7314 (N_7314,N_7215,N_7237);
nor U7315 (N_7315,N_7291,N_7268);
nand U7316 (N_7316,N_7250,N_7209);
nand U7317 (N_7317,N_7213,N_7233);
nand U7318 (N_7318,N_7217,N_7208);
and U7319 (N_7319,N_7299,N_7270);
xnor U7320 (N_7320,N_7296,N_7280);
xor U7321 (N_7321,N_7262,N_7211);
and U7322 (N_7322,N_7255,N_7251);
or U7323 (N_7323,N_7205,N_7228);
xnor U7324 (N_7324,N_7293,N_7284);
and U7325 (N_7325,N_7247,N_7216);
xnor U7326 (N_7326,N_7243,N_7257);
or U7327 (N_7327,N_7278,N_7229);
nand U7328 (N_7328,N_7202,N_7230);
nand U7329 (N_7329,N_7286,N_7277);
xor U7330 (N_7330,N_7289,N_7261);
xor U7331 (N_7331,N_7200,N_7226);
and U7332 (N_7332,N_7264,N_7248);
nand U7333 (N_7333,N_7246,N_7282);
or U7334 (N_7334,N_7203,N_7204);
nand U7335 (N_7335,N_7288,N_7218);
nor U7336 (N_7336,N_7206,N_7279);
or U7337 (N_7337,N_7244,N_7276);
nor U7338 (N_7338,N_7221,N_7238);
xor U7339 (N_7339,N_7259,N_7235);
or U7340 (N_7340,N_7223,N_7252);
or U7341 (N_7341,N_7297,N_7295);
and U7342 (N_7342,N_7260,N_7240);
or U7343 (N_7343,N_7298,N_7256);
nand U7344 (N_7344,N_7266,N_7265);
nor U7345 (N_7345,N_7267,N_7231);
nand U7346 (N_7346,N_7292,N_7207);
and U7347 (N_7347,N_7242,N_7214);
and U7348 (N_7348,N_7283,N_7281);
and U7349 (N_7349,N_7272,N_7271);
xor U7350 (N_7350,N_7214,N_7251);
and U7351 (N_7351,N_7262,N_7201);
or U7352 (N_7352,N_7216,N_7221);
and U7353 (N_7353,N_7272,N_7246);
nor U7354 (N_7354,N_7252,N_7291);
or U7355 (N_7355,N_7274,N_7260);
xor U7356 (N_7356,N_7255,N_7297);
xnor U7357 (N_7357,N_7239,N_7206);
nand U7358 (N_7358,N_7283,N_7289);
nor U7359 (N_7359,N_7224,N_7243);
nand U7360 (N_7360,N_7254,N_7264);
nand U7361 (N_7361,N_7270,N_7227);
nor U7362 (N_7362,N_7261,N_7215);
and U7363 (N_7363,N_7251,N_7299);
nand U7364 (N_7364,N_7239,N_7225);
xnor U7365 (N_7365,N_7240,N_7277);
nand U7366 (N_7366,N_7255,N_7227);
xnor U7367 (N_7367,N_7269,N_7238);
or U7368 (N_7368,N_7263,N_7262);
or U7369 (N_7369,N_7210,N_7203);
nand U7370 (N_7370,N_7263,N_7277);
nand U7371 (N_7371,N_7245,N_7232);
nand U7372 (N_7372,N_7259,N_7213);
and U7373 (N_7373,N_7238,N_7217);
or U7374 (N_7374,N_7292,N_7232);
nand U7375 (N_7375,N_7224,N_7268);
nor U7376 (N_7376,N_7222,N_7237);
xor U7377 (N_7377,N_7268,N_7275);
or U7378 (N_7378,N_7275,N_7213);
and U7379 (N_7379,N_7290,N_7253);
nor U7380 (N_7380,N_7252,N_7262);
or U7381 (N_7381,N_7249,N_7222);
xnor U7382 (N_7382,N_7295,N_7296);
and U7383 (N_7383,N_7213,N_7205);
or U7384 (N_7384,N_7247,N_7251);
or U7385 (N_7385,N_7222,N_7208);
or U7386 (N_7386,N_7292,N_7252);
xnor U7387 (N_7387,N_7292,N_7276);
xor U7388 (N_7388,N_7200,N_7275);
xor U7389 (N_7389,N_7251,N_7260);
or U7390 (N_7390,N_7269,N_7216);
xor U7391 (N_7391,N_7249,N_7245);
xor U7392 (N_7392,N_7231,N_7243);
or U7393 (N_7393,N_7279,N_7222);
nor U7394 (N_7394,N_7254,N_7249);
nand U7395 (N_7395,N_7266,N_7275);
or U7396 (N_7396,N_7203,N_7202);
xnor U7397 (N_7397,N_7235,N_7239);
or U7398 (N_7398,N_7241,N_7288);
or U7399 (N_7399,N_7296,N_7230);
nor U7400 (N_7400,N_7312,N_7331);
or U7401 (N_7401,N_7352,N_7346);
or U7402 (N_7402,N_7327,N_7348);
nor U7403 (N_7403,N_7387,N_7313);
xor U7404 (N_7404,N_7391,N_7340);
nor U7405 (N_7405,N_7334,N_7320);
xnor U7406 (N_7406,N_7370,N_7372);
nand U7407 (N_7407,N_7399,N_7323);
nand U7408 (N_7408,N_7300,N_7381);
and U7409 (N_7409,N_7341,N_7395);
and U7410 (N_7410,N_7339,N_7394);
and U7411 (N_7411,N_7365,N_7371);
nand U7412 (N_7412,N_7347,N_7393);
nand U7413 (N_7413,N_7353,N_7378);
xnor U7414 (N_7414,N_7373,N_7383);
nand U7415 (N_7415,N_7310,N_7359);
nand U7416 (N_7416,N_7330,N_7389);
nor U7417 (N_7417,N_7345,N_7349);
or U7418 (N_7418,N_7380,N_7369);
and U7419 (N_7419,N_7385,N_7360);
nor U7420 (N_7420,N_7333,N_7398);
or U7421 (N_7421,N_7319,N_7311);
or U7422 (N_7422,N_7304,N_7354);
nand U7423 (N_7423,N_7350,N_7325);
nor U7424 (N_7424,N_7361,N_7375);
nand U7425 (N_7425,N_7338,N_7306);
nand U7426 (N_7426,N_7362,N_7384);
or U7427 (N_7427,N_7366,N_7329);
and U7428 (N_7428,N_7303,N_7337);
and U7429 (N_7429,N_7382,N_7332);
nor U7430 (N_7430,N_7322,N_7321);
or U7431 (N_7431,N_7326,N_7342);
or U7432 (N_7432,N_7301,N_7305);
nor U7433 (N_7433,N_7351,N_7379);
nor U7434 (N_7434,N_7358,N_7302);
or U7435 (N_7435,N_7392,N_7355);
nand U7436 (N_7436,N_7374,N_7363);
nor U7437 (N_7437,N_7328,N_7317);
or U7438 (N_7438,N_7397,N_7308);
and U7439 (N_7439,N_7388,N_7335);
xnor U7440 (N_7440,N_7318,N_7314);
nor U7441 (N_7441,N_7357,N_7336);
and U7442 (N_7442,N_7386,N_7316);
and U7443 (N_7443,N_7344,N_7315);
nor U7444 (N_7444,N_7376,N_7396);
xor U7445 (N_7445,N_7364,N_7309);
nor U7446 (N_7446,N_7356,N_7367);
xor U7447 (N_7447,N_7343,N_7368);
and U7448 (N_7448,N_7390,N_7377);
or U7449 (N_7449,N_7324,N_7307);
nand U7450 (N_7450,N_7396,N_7370);
or U7451 (N_7451,N_7336,N_7374);
or U7452 (N_7452,N_7361,N_7383);
xnor U7453 (N_7453,N_7347,N_7349);
and U7454 (N_7454,N_7389,N_7397);
xor U7455 (N_7455,N_7377,N_7323);
xor U7456 (N_7456,N_7380,N_7306);
nor U7457 (N_7457,N_7365,N_7339);
xor U7458 (N_7458,N_7359,N_7362);
nand U7459 (N_7459,N_7390,N_7388);
xnor U7460 (N_7460,N_7332,N_7383);
xor U7461 (N_7461,N_7363,N_7313);
xnor U7462 (N_7462,N_7392,N_7348);
or U7463 (N_7463,N_7378,N_7321);
nand U7464 (N_7464,N_7390,N_7328);
and U7465 (N_7465,N_7351,N_7323);
or U7466 (N_7466,N_7313,N_7386);
nand U7467 (N_7467,N_7363,N_7307);
or U7468 (N_7468,N_7371,N_7386);
nand U7469 (N_7469,N_7349,N_7372);
nor U7470 (N_7470,N_7359,N_7323);
or U7471 (N_7471,N_7389,N_7392);
and U7472 (N_7472,N_7308,N_7382);
nor U7473 (N_7473,N_7346,N_7369);
and U7474 (N_7474,N_7342,N_7349);
and U7475 (N_7475,N_7359,N_7333);
nand U7476 (N_7476,N_7392,N_7367);
or U7477 (N_7477,N_7333,N_7368);
and U7478 (N_7478,N_7385,N_7324);
nand U7479 (N_7479,N_7340,N_7379);
and U7480 (N_7480,N_7334,N_7329);
or U7481 (N_7481,N_7316,N_7326);
nand U7482 (N_7482,N_7348,N_7366);
nor U7483 (N_7483,N_7371,N_7377);
or U7484 (N_7484,N_7372,N_7317);
xor U7485 (N_7485,N_7352,N_7395);
or U7486 (N_7486,N_7354,N_7340);
nand U7487 (N_7487,N_7385,N_7336);
or U7488 (N_7488,N_7360,N_7382);
nand U7489 (N_7489,N_7389,N_7362);
xor U7490 (N_7490,N_7378,N_7320);
nor U7491 (N_7491,N_7316,N_7314);
nor U7492 (N_7492,N_7307,N_7355);
and U7493 (N_7493,N_7329,N_7308);
or U7494 (N_7494,N_7348,N_7345);
nand U7495 (N_7495,N_7399,N_7329);
nor U7496 (N_7496,N_7355,N_7335);
xor U7497 (N_7497,N_7337,N_7359);
nand U7498 (N_7498,N_7356,N_7353);
xnor U7499 (N_7499,N_7390,N_7389);
xnor U7500 (N_7500,N_7484,N_7441);
or U7501 (N_7501,N_7487,N_7466);
or U7502 (N_7502,N_7405,N_7479);
or U7503 (N_7503,N_7435,N_7434);
nor U7504 (N_7504,N_7414,N_7433);
nand U7505 (N_7505,N_7493,N_7492);
and U7506 (N_7506,N_7418,N_7453);
nor U7507 (N_7507,N_7498,N_7440);
nor U7508 (N_7508,N_7469,N_7421);
nor U7509 (N_7509,N_7409,N_7422);
or U7510 (N_7510,N_7449,N_7432);
nand U7511 (N_7511,N_7404,N_7459);
nor U7512 (N_7512,N_7465,N_7442);
or U7513 (N_7513,N_7430,N_7473);
nor U7514 (N_7514,N_7447,N_7420);
or U7515 (N_7515,N_7490,N_7486);
xnor U7516 (N_7516,N_7454,N_7452);
or U7517 (N_7517,N_7411,N_7445);
nand U7518 (N_7518,N_7419,N_7410);
nor U7519 (N_7519,N_7450,N_7496);
or U7520 (N_7520,N_7403,N_7437);
xnor U7521 (N_7521,N_7491,N_7423);
nor U7522 (N_7522,N_7474,N_7489);
or U7523 (N_7523,N_7436,N_7464);
or U7524 (N_7524,N_7448,N_7415);
and U7525 (N_7525,N_7475,N_7451);
xnor U7526 (N_7526,N_7416,N_7478);
and U7527 (N_7527,N_7456,N_7417);
or U7528 (N_7528,N_7408,N_7495);
and U7529 (N_7529,N_7461,N_7413);
nor U7530 (N_7530,N_7406,N_7467);
and U7531 (N_7531,N_7426,N_7427);
nand U7532 (N_7532,N_7407,N_7457);
or U7533 (N_7533,N_7431,N_7497);
nand U7534 (N_7534,N_7402,N_7477);
or U7535 (N_7535,N_7481,N_7400);
nor U7536 (N_7536,N_7499,N_7480);
nand U7537 (N_7537,N_7429,N_7458);
nand U7538 (N_7538,N_7468,N_7460);
xor U7539 (N_7539,N_7482,N_7463);
xor U7540 (N_7540,N_7438,N_7439);
nor U7541 (N_7541,N_7485,N_7476);
nor U7542 (N_7542,N_7412,N_7443);
nand U7543 (N_7543,N_7455,N_7470);
or U7544 (N_7544,N_7462,N_7494);
nor U7545 (N_7545,N_7444,N_7471);
and U7546 (N_7546,N_7472,N_7401);
nor U7547 (N_7547,N_7488,N_7428);
and U7548 (N_7548,N_7424,N_7446);
xor U7549 (N_7549,N_7483,N_7425);
xnor U7550 (N_7550,N_7406,N_7430);
and U7551 (N_7551,N_7471,N_7434);
and U7552 (N_7552,N_7471,N_7422);
xnor U7553 (N_7553,N_7434,N_7429);
nand U7554 (N_7554,N_7438,N_7430);
xor U7555 (N_7555,N_7451,N_7455);
or U7556 (N_7556,N_7400,N_7429);
nor U7557 (N_7557,N_7433,N_7407);
xnor U7558 (N_7558,N_7491,N_7459);
and U7559 (N_7559,N_7447,N_7487);
or U7560 (N_7560,N_7410,N_7424);
or U7561 (N_7561,N_7490,N_7474);
and U7562 (N_7562,N_7434,N_7473);
nand U7563 (N_7563,N_7429,N_7468);
nor U7564 (N_7564,N_7417,N_7485);
nor U7565 (N_7565,N_7410,N_7461);
nand U7566 (N_7566,N_7411,N_7459);
nor U7567 (N_7567,N_7499,N_7466);
nand U7568 (N_7568,N_7456,N_7472);
nor U7569 (N_7569,N_7443,N_7465);
nor U7570 (N_7570,N_7479,N_7465);
and U7571 (N_7571,N_7455,N_7483);
or U7572 (N_7572,N_7419,N_7431);
or U7573 (N_7573,N_7435,N_7403);
and U7574 (N_7574,N_7435,N_7429);
or U7575 (N_7575,N_7473,N_7429);
and U7576 (N_7576,N_7423,N_7467);
xor U7577 (N_7577,N_7470,N_7400);
nor U7578 (N_7578,N_7484,N_7480);
nor U7579 (N_7579,N_7440,N_7462);
nor U7580 (N_7580,N_7415,N_7463);
nor U7581 (N_7581,N_7465,N_7466);
nand U7582 (N_7582,N_7429,N_7443);
or U7583 (N_7583,N_7428,N_7451);
nand U7584 (N_7584,N_7469,N_7487);
or U7585 (N_7585,N_7400,N_7450);
nand U7586 (N_7586,N_7414,N_7481);
nor U7587 (N_7587,N_7463,N_7481);
and U7588 (N_7588,N_7426,N_7429);
xor U7589 (N_7589,N_7454,N_7432);
nand U7590 (N_7590,N_7449,N_7428);
or U7591 (N_7591,N_7435,N_7450);
xnor U7592 (N_7592,N_7420,N_7435);
and U7593 (N_7593,N_7458,N_7479);
nand U7594 (N_7594,N_7417,N_7438);
nand U7595 (N_7595,N_7426,N_7458);
nor U7596 (N_7596,N_7449,N_7405);
and U7597 (N_7597,N_7441,N_7409);
or U7598 (N_7598,N_7452,N_7433);
nand U7599 (N_7599,N_7478,N_7428);
xor U7600 (N_7600,N_7543,N_7574);
nand U7601 (N_7601,N_7581,N_7532);
nor U7602 (N_7602,N_7565,N_7503);
nor U7603 (N_7603,N_7544,N_7540);
and U7604 (N_7604,N_7566,N_7546);
xor U7605 (N_7605,N_7545,N_7528);
or U7606 (N_7606,N_7576,N_7580);
nand U7607 (N_7607,N_7522,N_7567);
or U7608 (N_7608,N_7510,N_7598);
and U7609 (N_7609,N_7537,N_7518);
nor U7610 (N_7610,N_7534,N_7551);
nor U7611 (N_7611,N_7595,N_7559);
or U7612 (N_7612,N_7570,N_7526);
and U7613 (N_7613,N_7578,N_7516);
nand U7614 (N_7614,N_7501,N_7575);
nor U7615 (N_7615,N_7505,N_7594);
xnor U7616 (N_7616,N_7539,N_7564);
nor U7617 (N_7617,N_7558,N_7583);
nand U7618 (N_7618,N_7563,N_7555);
xnor U7619 (N_7619,N_7509,N_7589);
xor U7620 (N_7620,N_7552,N_7584);
nor U7621 (N_7621,N_7529,N_7550);
nor U7622 (N_7622,N_7582,N_7536);
nand U7623 (N_7623,N_7512,N_7535);
nor U7624 (N_7624,N_7547,N_7511);
and U7625 (N_7625,N_7521,N_7524);
or U7626 (N_7626,N_7586,N_7591);
xnor U7627 (N_7627,N_7560,N_7548);
nand U7628 (N_7628,N_7568,N_7587);
nand U7629 (N_7629,N_7530,N_7531);
and U7630 (N_7630,N_7538,N_7579);
nand U7631 (N_7631,N_7599,N_7541);
nor U7632 (N_7632,N_7549,N_7500);
xnor U7633 (N_7633,N_7557,N_7527);
nand U7634 (N_7634,N_7592,N_7542);
nor U7635 (N_7635,N_7590,N_7513);
nor U7636 (N_7636,N_7556,N_7507);
and U7637 (N_7637,N_7585,N_7553);
nor U7638 (N_7638,N_7569,N_7554);
and U7639 (N_7639,N_7504,N_7506);
xnor U7640 (N_7640,N_7533,N_7573);
and U7641 (N_7641,N_7572,N_7525);
nand U7642 (N_7642,N_7515,N_7519);
xor U7643 (N_7643,N_7596,N_7561);
or U7644 (N_7644,N_7508,N_7588);
and U7645 (N_7645,N_7577,N_7571);
xor U7646 (N_7646,N_7520,N_7517);
and U7647 (N_7647,N_7597,N_7562);
nand U7648 (N_7648,N_7593,N_7502);
or U7649 (N_7649,N_7514,N_7523);
nand U7650 (N_7650,N_7536,N_7557);
or U7651 (N_7651,N_7554,N_7520);
xor U7652 (N_7652,N_7578,N_7545);
nand U7653 (N_7653,N_7575,N_7513);
nand U7654 (N_7654,N_7567,N_7570);
nor U7655 (N_7655,N_7599,N_7545);
nor U7656 (N_7656,N_7508,N_7538);
nor U7657 (N_7657,N_7577,N_7537);
nand U7658 (N_7658,N_7596,N_7510);
nor U7659 (N_7659,N_7522,N_7589);
nand U7660 (N_7660,N_7574,N_7540);
and U7661 (N_7661,N_7545,N_7574);
nor U7662 (N_7662,N_7574,N_7594);
or U7663 (N_7663,N_7563,N_7599);
xor U7664 (N_7664,N_7518,N_7587);
and U7665 (N_7665,N_7523,N_7574);
nand U7666 (N_7666,N_7515,N_7562);
or U7667 (N_7667,N_7534,N_7535);
and U7668 (N_7668,N_7509,N_7534);
nor U7669 (N_7669,N_7577,N_7504);
nor U7670 (N_7670,N_7524,N_7500);
and U7671 (N_7671,N_7597,N_7564);
nand U7672 (N_7672,N_7537,N_7540);
and U7673 (N_7673,N_7567,N_7542);
nand U7674 (N_7674,N_7535,N_7523);
or U7675 (N_7675,N_7514,N_7521);
nor U7676 (N_7676,N_7548,N_7505);
nor U7677 (N_7677,N_7522,N_7559);
xnor U7678 (N_7678,N_7533,N_7595);
nand U7679 (N_7679,N_7524,N_7532);
nor U7680 (N_7680,N_7510,N_7589);
or U7681 (N_7681,N_7515,N_7596);
nand U7682 (N_7682,N_7520,N_7598);
nor U7683 (N_7683,N_7507,N_7560);
nor U7684 (N_7684,N_7569,N_7562);
nand U7685 (N_7685,N_7577,N_7586);
xnor U7686 (N_7686,N_7559,N_7581);
xor U7687 (N_7687,N_7500,N_7543);
nand U7688 (N_7688,N_7564,N_7535);
nand U7689 (N_7689,N_7501,N_7574);
and U7690 (N_7690,N_7578,N_7561);
or U7691 (N_7691,N_7515,N_7563);
or U7692 (N_7692,N_7509,N_7502);
or U7693 (N_7693,N_7532,N_7544);
or U7694 (N_7694,N_7511,N_7519);
nor U7695 (N_7695,N_7532,N_7563);
nor U7696 (N_7696,N_7572,N_7504);
xnor U7697 (N_7697,N_7524,N_7589);
nand U7698 (N_7698,N_7534,N_7538);
xor U7699 (N_7699,N_7599,N_7549);
nand U7700 (N_7700,N_7691,N_7605);
and U7701 (N_7701,N_7662,N_7654);
and U7702 (N_7702,N_7677,N_7629);
nand U7703 (N_7703,N_7621,N_7699);
xnor U7704 (N_7704,N_7604,N_7660);
xnor U7705 (N_7705,N_7695,N_7664);
and U7706 (N_7706,N_7618,N_7686);
and U7707 (N_7707,N_7667,N_7638);
and U7708 (N_7708,N_7649,N_7607);
or U7709 (N_7709,N_7606,N_7684);
and U7710 (N_7710,N_7678,N_7601);
and U7711 (N_7711,N_7685,N_7692);
or U7712 (N_7712,N_7647,N_7679);
or U7713 (N_7713,N_7603,N_7682);
and U7714 (N_7714,N_7693,N_7617);
and U7715 (N_7715,N_7602,N_7611);
xnor U7716 (N_7716,N_7633,N_7675);
and U7717 (N_7717,N_7600,N_7652);
or U7718 (N_7718,N_7614,N_7661);
and U7719 (N_7719,N_7613,N_7625);
or U7720 (N_7720,N_7612,N_7640);
nor U7721 (N_7721,N_7676,N_7656);
nand U7722 (N_7722,N_7637,N_7626);
or U7723 (N_7723,N_7620,N_7622);
xnor U7724 (N_7724,N_7624,N_7610);
nand U7725 (N_7725,N_7651,N_7641);
nor U7726 (N_7726,N_7646,N_7632);
nand U7727 (N_7727,N_7680,N_7609);
and U7728 (N_7728,N_7630,N_7683);
nand U7729 (N_7729,N_7619,N_7615);
nand U7730 (N_7730,N_7694,N_7671);
xor U7731 (N_7731,N_7689,N_7653);
or U7732 (N_7732,N_7628,N_7666);
nand U7733 (N_7733,N_7608,N_7698);
nor U7734 (N_7734,N_7616,N_7642);
and U7735 (N_7735,N_7673,N_7635);
nand U7736 (N_7736,N_7655,N_7634);
and U7737 (N_7737,N_7657,N_7623);
or U7738 (N_7738,N_7690,N_7670);
nand U7739 (N_7739,N_7674,N_7681);
or U7740 (N_7740,N_7669,N_7639);
nor U7741 (N_7741,N_7696,N_7631);
nor U7742 (N_7742,N_7687,N_7648);
nor U7743 (N_7743,N_7659,N_7697);
and U7744 (N_7744,N_7627,N_7688);
xor U7745 (N_7745,N_7650,N_7644);
or U7746 (N_7746,N_7636,N_7672);
or U7747 (N_7747,N_7643,N_7665);
or U7748 (N_7748,N_7658,N_7668);
nor U7749 (N_7749,N_7663,N_7645);
and U7750 (N_7750,N_7699,N_7667);
and U7751 (N_7751,N_7640,N_7661);
nor U7752 (N_7752,N_7671,N_7610);
xnor U7753 (N_7753,N_7610,N_7640);
xor U7754 (N_7754,N_7603,N_7676);
or U7755 (N_7755,N_7625,N_7624);
and U7756 (N_7756,N_7663,N_7672);
or U7757 (N_7757,N_7649,N_7638);
and U7758 (N_7758,N_7624,N_7660);
xnor U7759 (N_7759,N_7612,N_7643);
xnor U7760 (N_7760,N_7682,N_7640);
and U7761 (N_7761,N_7651,N_7606);
or U7762 (N_7762,N_7662,N_7681);
or U7763 (N_7763,N_7603,N_7660);
and U7764 (N_7764,N_7690,N_7655);
nor U7765 (N_7765,N_7635,N_7663);
xor U7766 (N_7766,N_7624,N_7613);
xor U7767 (N_7767,N_7631,N_7671);
xnor U7768 (N_7768,N_7684,N_7690);
and U7769 (N_7769,N_7637,N_7693);
and U7770 (N_7770,N_7631,N_7693);
nor U7771 (N_7771,N_7648,N_7664);
or U7772 (N_7772,N_7644,N_7687);
nand U7773 (N_7773,N_7627,N_7692);
xor U7774 (N_7774,N_7691,N_7687);
xor U7775 (N_7775,N_7634,N_7652);
nand U7776 (N_7776,N_7676,N_7680);
or U7777 (N_7777,N_7612,N_7667);
and U7778 (N_7778,N_7677,N_7609);
and U7779 (N_7779,N_7618,N_7692);
nor U7780 (N_7780,N_7603,N_7619);
nor U7781 (N_7781,N_7630,N_7694);
and U7782 (N_7782,N_7673,N_7650);
or U7783 (N_7783,N_7657,N_7671);
or U7784 (N_7784,N_7641,N_7691);
nor U7785 (N_7785,N_7648,N_7690);
nor U7786 (N_7786,N_7641,N_7643);
xor U7787 (N_7787,N_7697,N_7691);
nand U7788 (N_7788,N_7696,N_7612);
or U7789 (N_7789,N_7680,N_7651);
nor U7790 (N_7790,N_7639,N_7644);
or U7791 (N_7791,N_7622,N_7659);
nand U7792 (N_7792,N_7668,N_7694);
or U7793 (N_7793,N_7652,N_7639);
and U7794 (N_7794,N_7682,N_7632);
nor U7795 (N_7795,N_7627,N_7631);
and U7796 (N_7796,N_7614,N_7678);
or U7797 (N_7797,N_7659,N_7658);
xor U7798 (N_7798,N_7692,N_7676);
and U7799 (N_7799,N_7668,N_7640);
or U7800 (N_7800,N_7765,N_7746);
nor U7801 (N_7801,N_7768,N_7762);
xnor U7802 (N_7802,N_7730,N_7717);
or U7803 (N_7803,N_7703,N_7780);
nand U7804 (N_7804,N_7735,N_7713);
and U7805 (N_7805,N_7740,N_7786);
nor U7806 (N_7806,N_7720,N_7727);
or U7807 (N_7807,N_7724,N_7733);
xor U7808 (N_7808,N_7721,N_7756);
nand U7809 (N_7809,N_7704,N_7745);
nor U7810 (N_7810,N_7785,N_7788);
nand U7811 (N_7811,N_7761,N_7783);
and U7812 (N_7812,N_7750,N_7728);
nand U7813 (N_7813,N_7719,N_7779);
or U7814 (N_7814,N_7706,N_7771);
or U7815 (N_7815,N_7742,N_7725);
xnor U7816 (N_7816,N_7794,N_7715);
nand U7817 (N_7817,N_7793,N_7753);
nor U7818 (N_7818,N_7743,N_7770);
or U7819 (N_7819,N_7782,N_7723);
nand U7820 (N_7820,N_7755,N_7792);
and U7821 (N_7821,N_7726,N_7766);
or U7822 (N_7822,N_7732,N_7716);
and U7823 (N_7823,N_7777,N_7778);
or U7824 (N_7824,N_7749,N_7747);
nand U7825 (N_7825,N_7701,N_7700);
xnor U7826 (N_7826,N_7711,N_7739);
xnor U7827 (N_7827,N_7705,N_7772);
and U7828 (N_7828,N_7712,N_7707);
nor U7829 (N_7829,N_7789,N_7752);
or U7830 (N_7830,N_7751,N_7797);
or U7831 (N_7831,N_7763,N_7799);
nand U7832 (N_7832,N_7790,N_7781);
and U7833 (N_7833,N_7760,N_7795);
nor U7834 (N_7834,N_7787,N_7748);
nor U7835 (N_7835,N_7757,N_7709);
and U7836 (N_7836,N_7798,N_7769);
or U7837 (N_7837,N_7776,N_7744);
and U7838 (N_7838,N_7791,N_7702);
xnor U7839 (N_7839,N_7718,N_7708);
and U7840 (N_7840,N_7773,N_7759);
and U7841 (N_7841,N_7737,N_7796);
nand U7842 (N_7842,N_7722,N_7784);
xnor U7843 (N_7843,N_7774,N_7764);
xor U7844 (N_7844,N_7775,N_7741);
and U7845 (N_7845,N_7758,N_7729);
and U7846 (N_7846,N_7738,N_7714);
or U7847 (N_7847,N_7710,N_7754);
and U7848 (N_7848,N_7736,N_7731);
nor U7849 (N_7849,N_7734,N_7767);
and U7850 (N_7850,N_7766,N_7716);
and U7851 (N_7851,N_7723,N_7705);
and U7852 (N_7852,N_7715,N_7786);
or U7853 (N_7853,N_7799,N_7757);
nor U7854 (N_7854,N_7733,N_7743);
nand U7855 (N_7855,N_7770,N_7752);
or U7856 (N_7856,N_7747,N_7774);
xnor U7857 (N_7857,N_7785,N_7730);
and U7858 (N_7858,N_7722,N_7786);
nand U7859 (N_7859,N_7706,N_7756);
xor U7860 (N_7860,N_7798,N_7762);
or U7861 (N_7861,N_7715,N_7754);
xor U7862 (N_7862,N_7789,N_7796);
nor U7863 (N_7863,N_7736,N_7769);
nand U7864 (N_7864,N_7771,N_7729);
xor U7865 (N_7865,N_7704,N_7719);
xor U7866 (N_7866,N_7759,N_7720);
xor U7867 (N_7867,N_7732,N_7775);
nand U7868 (N_7868,N_7739,N_7789);
or U7869 (N_7869,N_7736,N_7761);
or U7870 (N_7870,N_7761,N_7737);
nor U7871 (N_7871,N_7763,N_7796);
xnor U7872 (N_7872,N_7705,N_7700);
xor U7873 (N_7873,N_7740,N_7710);
nor U7874 (N_7874,N_7779,N_7706);
xnor U7875 (N_7875,N_7794,N_7741);
xnor U7876 (N_7876,N_7721,N_7755);
or U7877 (N_7877,N_7769,N_7725);
or U7878 (N_7878,N_7763,N_7731);
and U7879 (N_7879,N_7765,N_7763);
nor U7880 (N_7880,N_7737,N_7734);
nor U7881 (N_7881,N_7732,N_7780);
and U7882 (N_7882,N_7799,N_7706);
xor U7883 (N_7883,N_7775,N_7709);
nand U7884 (N_7884,N_7717,N_7754);
or U7885 (N_7885,N_7741,N_7772);
or U7886 (N_7886,N_7757,N_7734);
nand U7887 (N_7887,N_7728,N_7714);
or U7888 (N_7888,N_7747,N_7734);
or U7889 (N_7889,N_7706,N_7753);
nor U7890 (N_7890,N_7749,N_7765);
nand U7891 (N_7891,N_7741,N_7715);
xor U7892 (N_7892,N_7739,N_7769);
nor U7893 (N_7893,N_7774,N_7738);
xnor U7894 (N_7894,N_7763,N_7708);
nand U7895 (N_7895,N_7757,N_7743);
or U7896 (N_7896,N_7701,N_7729);
nor U7897 (N_7897,N_7792,N_7796);
nor U7898 (N_7898,N_7771,N_7753);
nand U7899 (N_7899,N_7726,N_7737);
and U7900 (N_7900,N_7813,N_7843);
nand U7901 (N_7901,N_7835,N_7846);
nand U7902 (N_7902,N_7831,N_7873);
or U7903 (N_7903,N_7869,N_7841);
xnor U7904 (N_7904,N_7817,N_7883);
or U7905 (N_7905,N_7888,N_7876);
nand U7906 (N_7906,N_7855,N_7893);
nor U7907 (N_7907,N_7806,N_7829);
xnor U7908 (N_7908,N_7834,N_7825);
or U7909 (N_7909,N_7810,N_7818);
and U7910 (N_7910,N_7830,N_7858);
nor U7911 (N_7911,N_7836,N_7821);
nand U7912 (N_7912,N_7851,N_7804);
xor U7913 (N_7913,N_7837,N_7899);
or U7914 (N_7914,N_7856,N_7853);
xor U7915 (N_7915,N_7838,N_7819);
nand U7916 (N_7916,N_7826,N_7879);
and U7917 (N_7917,N_7811,N_7815);
or U7918 (N_7918,N_7866,N_7845);
nand U7919 (N_7919,N_7822,N_7849);
or U7920 (N_7920,N_7802,N_7823);
or U7921 (N_7921,N_7800,N_7898);
or U7922 (N_7922,N_7875,N_7882);
and U7923 (N_7923,N_7816,N_7824);
nand U7924 (N_7924,N_7812,N_7891);
nand U7925 (N_7925,N_7895,N_7870);
nor U7926 (N_7926,N_7886,N_7878);
nor U7927 (N_7927,N_7827,N_7894);
nand U7928 (N_7928,N_7896,N_7848);
and U7929 (N_7929,N_7874,N_7860);
xnor U7930 (N_7930,N_7857,N_7852);
xor U7931 (N_7931,N_7807,N_7805);
or U7932 (N_7932,N_7862,N_7832);
or U7933 (N_7933,N_7833,N_7864);
nor U7934 (N_7934,N_7859,N_7828);
or U7935 (N_7935,N_7887,N_7897);
nor U7936 (N_7936,N_7865,N_7850);
nand U7937 (N_7937,N_7814,N_7871);
nor U7938 (N_7938,N_7861,N_7885);
and U7939 (N_7939,N_7890,N_7803);
and U7940 (N_7940,N_7884,N_7839);
xor U7941 (N_7941,N_7892,N_7844);
and U7942 (N_7942,N_7881,N_7809);
xor U7943 (N_7943,N_7872,N_7847);
nor U7944 (N_7944,N_7877,N_7854);
nand U7945 (N_7945,N_7868,N_7867);
xor U7946 (N_7946,N_7820,N_7801);
nor U7947 (N_7947,N_7880,N_7863);
or U7948 (N_7948,N_7808,N_7842);
or U7949 (N_7949,N_7889,N_7840);
and U7950 (N_7950,N_7829,N_7833);
or U7951 (N_7951,N_7800,N_7899);
nor U7952 (N_7952,N_7873,N_7818);
and U7953 (N_7953,N_7895,N_7891);
xor U7954 (N_7954,N_7844,N_7808);
and U7955 (N_7955,N_7861,N_7853);
nor U7956 (N_7956,N_7804,N_7841);
nand U7957 (N_7957,N_7829,N_7859);
nand U7958 (N_7958,N_7847,N_7874);
xnor U7959 (N_7959,N_7878,N_7854);
nand U7960 (N_7960,N_7809,N_7868);
or U7961 (N_7961,N_7837,N_7881);
and U7962 (N_7962,N_7812,N_7878);
xnor U7963 (N_7963,N_7894,N_7807);
and U7964 (N_7964,N_7882,N_7828);
and U7965 (N_7965,N_7822,N_7860);
or U7966 (N_7966,N_7891,N_7832);
nand U7967 (N_7967,N_7890,N_7833);
and U7968 (N_7968,N_7889,N_7872);
nor U7969 (N_7969,N_7837,N_7839);
nor U7970 (N_7970,N_7858,N_7874);
nand U7971 (N_7971,N_7818,N_7811);
nor U7972 (N_7972,N_7869,N_7836);
xnor U7973 (N_7973,N_7856,N_7888);
nor U7974 (N_7974,N_7848,N_7800);
nor U7975 (N_7975,N_7843,N_7890);
and U7976 (N_7976,N_7860,N_7881);
nand U7977 (N_7977,N_7815,N_7887);
or U7978 (N_7978,N_7892,N_7871);
xnor U7979 (N_7979,N_7866,N_7804);
or U7980 (N_7980,N_7895,N_7880);
nand U7981 (N_7981,N_7811,N_7852);
or U7982 (N_7982,N_7820,N_7842);
or U7983 (N_7983,N_7808,N_7854);
nand U7984 (N_7984,N_7821,N_7881);
and U7985 (N_7985,N_7818,N_7832);
nor U7986 (N_7986,N_7848,N_7872);
nand U7987 (N_7987,N_7871,N_7802);
or U7988 (N_7988,N_7863,N_7876);
nand U7989 (N_7989,N_7839,N_7866);
xnor U7990 (N_7990,N_7883,N_7814);
nor U7991 (N_7991,N_7804,N_7847);
nand U7992 (N_7992,N_7893,N_7891);
and U7993 (N_7993,N_7827,N_7820);
and U7994 (N_7994,N_7808,N_7868);
nand U7995 (N_7995,N_7865,N_7820);
and U7996 (N_7996,N_7868,N_7833);
and U7997 (N_7997,N_7816,N_7806);
nor U7998 (N_7998,N_7829,N_7890);
nor U7999 (N_7999,N_7895,N_7837);
and U8000 (N_8000,N_7975,N_7935);
and U8001 (N_8001,N_7995,N_7932);
or U8002 (N_8002,N_7970,N_7922);
and U8003 (N_8003,N_7910,N_7950);
nand U8004 (N_8004,N_7959,N_7973);
or U8005 (N_8005,N_7976,N_7944);
or U8006 (N_8006,N_7974,N_7938);
xnor U8007 (N_8007,N_7926,N_7906);
xnor U8008 (N_8008,N_7940,N_7996);
nor U8009 (N_8009,N_7981,N_7955);
xor U8010 (N_8010,N_7966,N_7998);
xor U8011 (N_8011,N_7991,N_7931);
nor U8012 (N_8012,N_7901,N_7917);
xor U8013 (N_8013,N_7915,N_7952);
nand U8014 (N_8014,N_7983,N_7960);
and U8015 (N_8015,N_7999,N_7972);
nor U8016 (N_8016,N_7925,N_7918);
and U8017 (N_8017,N_7900,N_7963);
and U8018 (N_8018,N_7968,N_7929);
and U8019 (N_8019,N_7954,N_7951);
xnor U8020 (N_8020,N_7993,N_7934);
nor U8021 (N_8021,N_7957,N_7921);
nor U8022 (N_8022,N_7942,N_7989);
xor U8023 (N_8023,N_7903,N_7978);
or U8024 (N_8024,N_7911,N_7985);
and U8025 (N_8025,N_7984,N_7927);
nand U8026 (N_8026,N_7956,N_7953);
xnor U8027 (N_8027,N_7964,N_7986);
or U8028 (N_8028,N_7937,N_7971);
nor U8029 (N_8029,N_7958,N_7902);
nand U8030 (N_8030,N_7943,N_7920);
or U8031 (N_8031,N_7965,N_7933);
or U8032 (N_8032,N_7962,N_7923);
nand U8033 (N_8033,N_7904,N_7928);
nand U8034 (N_8034,N_7969,N_7945);
nor U8035 (N_8035,N_7992,N_7946);
or U8036 (N_8036,N_7949,N_7947);
nand U8037 (N_8037,N_7913,N_7961);
or U8038 (N_8038,N_7967,N_7997);
xor U8039 (N_8039,N_7987,N_7930);
xnor U8040 (N_8040,N_7982,N_7909);
xnor U8041 (N_8041,N_7941,N_7977);
or U8042 (N_8042,N_7939,N_7988);
xor U8043 (N_8043,N_7919,N_7924);
nor U8044 (N_8044,N_7948,N_7936);
nor U8045 (N_8045,N_7905,N_7990);
xnor U8046 (N_8046,N_7914,N_7907);
and U8047 (N_8047,N_7979,N_7912);
and U8048 (N_8048,N_7916,N_7980);
or U8049 (N_8049,N_7908,N_7994);
or U8050 (N_8050,N_7920,N_7913);
or U8051 (N_8051,N_7960,N_7959);
nand U8052 (N_8052,N_7988,N_7909);
nor U8053 (N_8053,N_7900,N_7908);
nand U8054 (N_8054,N_7967,N_7986);
xnor U8055 (N_8055,N_7997,N_7960);
or U8056 (N_8056,N_7929,N_7901);
and U8057 (N_8057,N_7928,N_7989);
nand U8058 (N_8058,N_7960,N_7920);
xnor U8059 (N_8059,N_7981,N_7900);
nand U8060 (N_8060,N_7989,N_7943);
and U8061 (N_8061,N_7927,N_7948);
or U8062 (N_8062,N_7991,N_7907);
nand U8063 (N_8063,N_7992,N_7901);
xnor U8064 (N_8064,N_7937,N_7933);
or U8065 (N_8065,N_7997,N_7968);
xnor U8066 (N_8066,N_7970,N_7992);
nand U8067 (N_8067,N_7916,N_7974);
nand U8068 (N_8068,N_7924,N_7935);
or U8069 (N_8069,N_7992,N_7932);
or U8070 (N_8070,N_7984,N_7900);
and U8071 (N_8071,N_7943,N_7905);
or U8072 (N_8072,N_7930,N_7983);
nand U8073 (N_8073,N_7999,N_7966);
xnor U8074 (N_8074,N_7957,N_7964);
and U8075 (N_8075,N_7942,N_7900);
nand U8076 (N_8076,N_7937,N_7963);
nor U8077 (N_8077,N_7938,N_7905);
or U8078 (N_8078,N_7906,N_7929);
nand U8079 (N_8079,N_7990,N_7929);
nor U8080 (N_8080,N_7968,N_7946);
or U8081 (N_8081,N_7990,N_7970);
nand U8082 (N_8082,N_7981,N_7978);
nor U8083 (N_8083,N_7900,N_7987);
nor U8084 (N_8084,N_7989,N_7918);
xor U8085 (N_8085,N_7935,N_7911);
or U8086 (N_8086,N_7973,N_7905);
and U8087 (N_8087,N_7974,N_7901);
nor U8088 (N_8088,N_7920,N_7944);
and U8089 (N_8089,N_7900,N_7936);
xor U8090 (N_8090,N_7965,N_7925);
and U8091 (N_8091,N_7956,N_7986);
and U8092 (N_8092,N_7946,N_7915);
nor U8093 (N_8093,N_7909,N_7989);
nand U8094 (N_8094,N_7917,N_7910);
nand U8095 (N_8095,N_7988,N_7949);
or U8096 (N_8096,N_7943,N_7928);
nor U8097 (N_8097,N_7908,N_7980);
nand U8098 (N_8098,N_7993,N_7913);
and U8099 (N_8099,N_7995,N_7990);
and U8100 (N_8100,N_8061,N_8009);
or U8101 (N_8101,N_8067,N_8021);
xnor U8102 (N_8102,N_8008,N_8074);
xor U8103 (N_8103,N_8004,N_8097);
or U8104 (N_8104,N_8019,N_8010);
nor U8105 (N_8105,N_8023,N_8048);
xor U8106 (N_8106,N_8047,N_8003);
nor U8107 (N_8107,N_8057,N_8062);
and U8108 (N_8108,N_8056,N_8092);
nand U8109 (N_8109,N_8050,N_8011);
xnor U8110 (N_8110,N_8006,N_8018);
nor U8111 (N_8111,N_8033,N_8083);
or U8112 (N_8112,N_8060,N_8082);
nand U8113 (N_8113,N_8015,N_8093);
xnor U8114 (N_8114,N_8066,N_8080);
xnor U8115 (N_8115,N_8070,N_8090);
and U8116 (N_8116,N_8096,N_8002);
and U8117 (N_8117,N_8052,N_8063);
xor U8118 (N_8118,N_8030,N_8017);
nand U8119 (N_8119,N_8020,N_8028);
xnor U8120 (N_8120,N_8024,N_8037);
nor U8121 (N_8121,N_8016,N_8064);
and U8122 (N_8122,N_8039,N_8073);
or U8123 (N_8123,N_8086,N_8095);
or U8124 (N_8124,N_8071,N_8029);
nand U8125 (N_8125,N_8035,N_8059);
xor U8126 (N_8126,N_8091,N_8001);
nand U8127 (N_8127,N_8055,N_8078);
nand U8128 (N_8128,N_8072,N_8022);
or U8129 (N_8129,N_8046,N_8041);
xnor U8130 (N_8130,N_8077,N_8084);
or U8131 (N_8131,N_8013,N_8068);
nand U8132 (N_8132,N_8045,N_8075);
xor U8133 (N_8133,N_8085,N_8027);
nand U8134 (N_8134,N_8005,N_8044);
nor U8135 (N_8135,N_8053,N_8025);
and U8136 (N_8136,N_8076,N_8036);
nor U8137 (N_8137,N_8049,N_8032);
and U8138 (N_8138,N_8031,N_8089);
xor U8139 (N_8139,N_8065,N_8079);
and U8140 (N_8140,N_8081,N_8098);
nor U8141 (N_8141,N_8051,N_8007);
nand U8142 (N_8142,N_8054,N_8087);
or U8143 (N_8143,N_8094,N_8058);
or U8144 (N_8144,N_8000,N_8026);
or U8145 (N_8145,N_8014,N_8069);
and U8146 (N_8146,N_8043,N_8099);
nor U8147 (N_8147,N_8040,N_8042);
xor U8148 (N_8148,N_8038,N_8088);
nor U8149 (N_8149,N_8012,N_8034);
nand U8150 (N_8150,N_8074,N_8032);
nor U8151 (N_8151,N_8098,N_8072);
nor U8152 (N_8152,N_8053,N_8031);
and U8153 (N_8153,N_8029,N_8093);
nor U8154 (N_8154,N_8030,N_8021);
and U8155 (N_8155,N_8024,N_8031);
nor U8156 (N_8156,N_8050,N_8007);
xnor U8157 (N_8157,N_8004,N_8014);
nor U8158 (N_8158,N_8022,N_8099);
and U8159 (N_8159,N_8038,N_8084);
xor U8160 (N_8160,N_8062,N_8071);
and U8161 (N_8161,N_8050,N_8099);
xnor U8162 (N_8162,N_8030,N_8082);
xnor U8163 (N_8163,N_8054,N_8055);
xnor U8164 (N_8164,N_8041,N_8085);
and U8165 (N_8165,N_8089,N_8067);
and U8166 (N_8166,N_8027,N_8013);
nor U8167 (N_8167,N_8081,N_8027);
nand U8168 (N_8168,N_8036,N_8040);
nand U8169 (N_8169,N_8086,N_8010);
or U8170 (N_8170,N_8085,N_8084);
or U8171 (N_8171,N_8076,N_8031);
xor U8172 (N_8172,N_8092,N_8059);
nand U8173 (N_8173,N_8082,N_8093);
xnor U8174 (N_8174,N_8092,N_8026);
and U8175 (N_8175,N_8053,N_8065);
or U8176 (N_8176,N_8082,N_8025);
or U8177 (N_8177,N_8002,N_8026);
or U8178 (N_8178,N_8094,N_8014);
and U8179 (N_8179,N_8050,N_8008);
xnor U8180 (N_8180,N_8018,N_8085);
nor U8181 (N_8181,N_8038,N_8052);
or U8182 (N_8182,N_8018,N_8068);
xnor U8183 (N_8183,N_8051,N_8094);
nand U8184 (N_8184,N_8097,N_8085);
or U8185 (N_8185,N_8074,N_8021);
nand U8186 (N_8186,N_8061,N_8021);
nor U8187 (N_8187,N_8053,N_8085);
or U8188 (N_8188,N_8043,N_8098);
or U8189 (N_8189,N_8049,N_8087);
xnor U8190 (N_8190,N_8078,N_8017);
and U8191 (N_8191,N_8010,N_8072);
or U8192 (N_8192,N_8035,N_8095);
and U8193 (N_8193,N_8081,N_8089);
nor U8194 (N_8194,N_8027,N_8040);
nor U8195 (N_8195,N_8080,N_8093);
nor U8196 (N_8196,N_8029,N_8096);
nor U8197 (N_8197,N_8024,N_8073);
and U8198 (N_8198,N_8060,N_8006);
nand U8199 (N_8199,N_8007,N_8009);
and U8200 (N_8200,N_8172,N_8149);
or U8201 (N_8201,N_8159,N_8137);
nor U8202 (N_8202,N_8179,N_8108);
and U8203 (N_8203,N_8168,N_8173);
xor U8204 (N_8204,N_8130,N_8185);
nand U8205 (N_8205,N_8125,N_8184);
or U8206 (N_8206,N_8115,N_8187);
and U8207 (N_8207,N_8160,N_8190);
or U8208 (N_8208,N_8101,N_8171);
xnor U8209 (N_8209,N_8122,N_8110);
nor U8210 (N_8210,N_8140,N_8128);
nor U8211 (N_8211,N_8141,N_8155);
nor U8212 (N_8212,N_8151,N_8152);
or U8213 (N_8213,N_8177,N_8129);
nand U8214 (N_8214,N_8143,N_8135);
xor U8215 (N_8215,N_8181,N_8156);
nor U8216 (N_8216,N_8132,N_8175);
xnor U8217 (N_8217,N_8126,N_8180);
or U8218 (N_8218,N_8139,N_8105);
and U8219 (N_8219,N_8124,N_8142);
and U8220 (N_8220,N_8182,N_8199);
nand U8221 (N_8221,N_8102,N_8121);
and U8222 (N_8222,N_8113,N_8104);
nand U8223 (N_8223,N_8154,N_8118);
xnor U8224 (N_8224,N_8106,N_8144);
xnor U8225 (N_8225,N_8193,N_8186);
nor U8226 (N_8226,N_8100,N_8145);
and U8227 (N_8227,N_8169,N_8195);
or U8228 (N_8228,N_8117,N_8191);
and U8229 (N_8229,N_8198,N_8164);
nor U8230 (N_8230,N_8192,N_8158);
or U8231 (N_8231,N_8107,N_8119);
nand U8232 (N_8232,N_8178,N_8157);
nand U8233 (N_8233,N_8197,N_8166);
nand U8234 (N_8234,N_8147,N_8196);
nand U8235 (N_8235,N_8116,N_8161);
or U8236 (N_8236,N_8134,N_8114);
or U8237 (N_8237,N_8123,N_8162);
nand U8238 (N_8238,N_8189,N_8103);
or U8239 (N_8239,N_8150,N_8183);
nand U8240 (N_8240,N_8153,N_8120);
and U8241 (N_8241,N_8163,N_8148);
nor U8242 (N_8242,N_8194,N_8176);
or U8243 (N_8243,N_8174,N_8136);
or U8244 (N_8244,N_8170,N_8165);
and U8245 (N_8245,N_8109,N_8133);
and U8246 (N_8246,N_8188,N_8111);
and U8247 (N_8247,N_8146,N_8127);
nand U8248 (N_8248,N_8167,N_8138);
and U8249 (N_8249,N_8112,N_8131);
nand U8250 (N_8250,N_8163,N_8153);
nor U8251 (N_8251,N_8106,N_8128);
nor U8252 (N_8252,N_8104,N_8155);
xnor U8253 (N_8253,N_8177,N_8174);
xnor U8254 (N_8254,N_8107,N_8166);
or U8255 (N_8255,N_8135,N_8107);
nor U8256 (N_8256,N_8140,N_8131);
nand U8257 (N_8257,N_8140,N_8153);
or U8258 (N_8258,N_8159,N_8172);
nor U8259 (N_8259,N_8148,N_8113);
xor U8260 (N_8260,N_8178,N_8124);
nor U8261 (N_8261,N_8109,N_8197);
nand U8262 (N_8262,N_8142,N_8162);
and U8263 (N_8263,N_8107,N_8112);
and U8264 (N_8264,N_8163,N_8125);
nor U8265 (N_8265,N_8104,N_8118);
xnor U8266 (N_8266,N_8134,N_8144);
and U8267 (N_8267,N_8143,N_8118);
nand U8268 (N_8268,N_8124,N_8181);
xnor U8269 (N_8269,N_8189,N_8146);
nand U8270 (N_8270,N_8102,N_8197);
nand U8271 (N_8271,N_8172,N_8134);
and U8272 (N_8272,N_8163,N_8116);
and U8273 (N_8273,N_8195,N_8129);
nand U8274 (N_8274,N_8108,N_8154);
nor U8275 (N_8275,N_8108,N_8181);
nor U8276 (N_8276,N_8155,N_8109);
xor U8277 (N_8277,N_8146,N_8123);
xnor U8278 (N_8278,N_8173,N_8180);
nand U8279 (N_8279,N_8129,N_8148);
xnor U8280 (N_8280,N_8153,N_8121);
and U8281 (N_8281,N_8166,N_8187);
xnor U8282 (N_8282,N_8180,N_8155);
xor U8283 (N_8283,N_8144,N_8117);
nor U8284 (N_8284,N_8105,N_8117);
or U8285 (N_8285,N_8149,N_8181);
and U8286 (N_8286,N_8164,N_8155);
nand U8287 (N_8287,N_8177,N_8102);
xnor U8288 (N_8288,N_8178,N_8159);
nand U8289 (N_8289,N_8168,N_8166);
nor U8290 (N_8290,N_8179,N_8130);
and U8291 (N_8291,N_8195,N_8163);
xor U8292 (N_8292,N_8181,N_8160);
nor U8293 (N_8293,N_8198,N_8131);
nand U8294 (N_8294,N_8185,N_8144);
nor U8295 (N_8295,N_8170,N_8110);
nand U8296 (N_8296,N_8156,N_8112);
and U8297 (N_8297,N_8164,N_8131);
nor U8298 (N_8298,N_8181,N_8112);
and U8299 (N_8299,N_8148,N_8167);
or U8300 (N_8300,N_8281,N_8221);
or U8301 (N_8301,N_8233,N_8205);
nor U8302 (N_8302,N_8285,N_8292);
xnor U8303 (N_8303,N_8235,N_8241);
nor U8304 (N_8304,N_8251,N_8254);
or U8305 (N_8305,N_8200,N_8249);
nor U8306 (N_8306,N_8206,N_8259);
nor U8307 (N_8307,N_8216,N_8211);
xor U8308 (N_8308,N_8217,N_8260);
nor U8309 (N_8309,N_8296,N_8290);
and U8310 (N_8310,N_8262,N_8276);
and U8311 (N_8311,N_8252,N_8257);
nor U8312 (N_8312,N_8210,N_8250);
or U8313 (N_8313,N_8264,N_8240);
or U8314 (N_8314,N_8242,N_8212);
nand U8315 (N_8315,N_8286,N_8293);
or U8316 (N_8316,N_8223,N_8255);
nor U8317 (N_8317,N_8287,N_8204);
xor U8318 (N_8318,N_8289,N_8298);
and U8319 (N_8319,N_8297,N_8218);
or U8320 (N_8320,N_8214,N_8294);
nor U8321 (N_8321,N_8295,N_8269);
xor U8322 (N_8322,N_8220,N_8291);
xor U8323 (N_8323,N_8275,N_8279);
or U8324 (N_8324,N_8228,N_8225);
or U8325 (N_8325,N_8203,N_8288);
and U8326 (N_8326,N_8245,N_8222);
xnor U8327 (N_8327,N_8208,N_8258);
nand U8328 (N_8328,N_8256,N_8284);
xor U8329 (N_8329,N_8272,N_8266);
nor U8330 (N_8330,N_8230,N_8274);
and U8331 (N_8331,N_8244,N_8268);
nor U8332 (N_8332,N_8238,N_8267);
or U8333 (N_8333,N_8277,N_8224);
xnor U8334 (N_8334,N_8261,N_8280);
xor U8335 (N_8335,N_8270,N_8283);
and U8336 (N_8336,N_8219,N_8282);
and U8337 (N_8337,N_8237,N_8232);
xnor U8338 (N_8338,N_8207,N_8243);
xor U8339 (N_8339,N_8253,N_8246);
xor U8340 (N_8340,N_8247,N_8299);
and U8341 (N_8341,N_8248,N_8215);
and U8342 (N_8342,N_8271,N_8201);
or U8343 (N_8343,N_8213,N_8278);
nand U8344 (N_8344,N_8234,N_8229);
xor U8345 (N_8345,N_8231,N_8209);
or U8346 (N_8346,N_8202,N_8273);
nor U8347 (N_8347,N_8239,N_8227);
nor U8348 (N_8348,N_8226,N_8265);
and U8349 (N_8349,N_8263,N_8236);
and U8350 (N_8350,N_8261,N_8242);
nand U8351 (N_8351,N_8228,N_8281);
nor U8352 (N_8352,N_8287,N_8257);
xnor U8353 (N_8353,N_8254,N_8210);
or U8354 (N_8354,N_8211,N_8250);
and U8355 (N_8355,N_8267,N_8282);
or U8356 (N_8356,N_8277,N_8209);
or U8357 (N_8357,N_8289,N_8252);
nand U8358 (N_8358,N_8235,N_8206);
xnor U8359 (N_8359,N_8253,N_8221);
nand U8360 (N_8360,N_8242,N_8215);
nand U8361 (N_8361,N_8268,N_8205);
and U8362 (N_8362,N_8234,N_8228);
or U8363 (N_8363,N_8214,N_8206);
and U8364 (N_8364,N_8202,N_8282);
and U8365 (N_8365,N_8213,N_8258);
xnor U8366 (N_8366,N_8275,N_8244);
nand U8367 (N_8367,N_8265,N_8219);
xor U8368 (N_8368,N_8276,N_8218);
xnor U8369 (N_8369,N_8249,N_8218);
or U8370 (N_8370,N_8272,N_8277);
nor U8371 (N_8371,N_8254,N_8215);
nor U8372 (N_8372,N_8208,N_8242);
nor U8373 (N_8373,N_8271,N_8292);
nor U8374 (N_8374,N_8229,N_8216);
nor U8375 (N_8375,N_8230,N_8245);
nand U8376 (N_8376,N_8281,N_8258);
or U8377 (N_8377,N_8232,N_8246);
or U8378 (N_8378,N_8234,N_8232);
nor U8379 (N_8379,N_8269,N_8266);
and U8380 (N_8380,N_8215,N_8221);
or U8381 (N_8381,N_8287,N_8293);
nor U8382 (N_8382,N_8215,N_8293);
or U8383 (N_8383,N_8279,N_8220);
nand U8384 (N_8384,N_8233,N_8208);
or U8385 (N_8385,N_8221,N_8290);
nor U8386 (N_8386,N_8270,N_8236);
nand U8387 (N_8387,N_8240,N_8237);
or U8388 (N_8388,N_8226,N_8262);
or U8389 (N_8389,N_8219,N_8236);
nor U8390 (N_8390,N_8296,N_8245);
nor U8391 (N_8391,N_8236,N_8295);
nor U8392 (N_8392,N_8263,N_8249);
nor U8393 (N_8393,N_8236,N_8298);
or U8394 (N_8394,N_8290,N_8258);
or U8395 (N_8395,N_8296,N_8287);
or U8396 (N_8396,N_8278,N_8232);
nand U8397 (N_8397,N_8216,N_8204);
nand U8398 (N_8398,N_8248,N_8273);
xor U8399 (N_8399,N_8270,N_8239);
nand U8400 (N_8400,N_8348,N_8373);
and U8401 (N_8401,N_8310,N_8383);
xor U8402 (N_8402,N_8368,N_8316);
nor U8403 (N_8403,N_8333,N_8387);
and U8404 (N_8404,N_8370,N_8336);
xor U8405 (N_8405,N_8397,N_8317);
xnor U8406 (N_8406,N_8327,N_8326);
or U8407 (N_8407,N_8365,N_8330);
xnor U8408 (N_8408,N_8388,N_8301);
or U8409 (N_8409,N_8311,N_8369);
or U8410 (N_8410,N_8323,N_8334);
xor U8411 (N_8411,N_8303,N_8338);
nor U8412 (N_8412,N_8314,N_8391);
nand U8413 (N_8413,N_8312,N_8328);
or U8414 (N_8414,N_8350,N_8351);
nand U8415 (N_8415,N_8389,N_8325);
nor U8416 (N_8416,N_8331,N_8340);
and U8417 (N_8417,N_8304,N_8347);
nand U8418 (N_8418,N_8359,N_8364);
nand U8419 (N_8419,N_8362,N_8378);
or U8420 (N_8420,N_8366,N_8386);
xor U8421 (N_8421,N_8390,N_8385);
nor U8422 (N_8422,N_8376,N_8345);
nor U8423 (N_8423,N_8352,N_8354);
xor U8424 (N_8424,N_8377,N_8398);
nor U8425 (N_8425,N_8357,N_8318);
xnor U8426 (N_8426,N_8363,N_8315);
xor U8427 (N_8427,N_8356,N_8360);
or U8428 (N_8428,N_8379,N_8332);
xnor U8429 (N_8429,N_8337,N_8342);
xor U8430 (N_8430,N_8349,N_8394);
nand U8431 (N_8431,N_8355,N_8300);
and U8432 (N_8432,N_8367,N_8353);
nand U8433 (N_8433,N_8382,N_8372);
nor U8434 (N_8434,N_8375,N_8306);
and U8435 (N_8435,N_8396,N_8335);
nor U8436 (N_8436,N_8384,N_8302);
and U8437 (N_8437,N_8341,N_8380);
or U8438 (N_8438,N_8371,N_8313);
or U8439 (N_8439,N_8361,N_8343);
nor U8440 (N_8440,N_8392,N_8321);
nor U8441 (N_8441,N_8395,N_8305);
and U8442 (N_8442,N_8309,N_8308);
or U8443 (N_8443,N_8320,N_8344);
nand U8444 (N_8444,N_8319,N_8346);
xnor U8445 (N_8445,N_8374,N_8381);
nand U8446 (N_8446,N_8399,N_8307);
nor U8447 (N_8447,N_8329,N_8393);
xnor U8448 (N_8448,N_8339,N_8322);
xnor U8449 (N_8449,N_8358,N_8324);
and U8450 (N_8450,N_8343,N_8362);
and U8451 (N_8451,N_8307,N_8369);
xor U8452 (N_8452,N_8393,N_8326);
nor U8453 (N_8453,N_8372,N_8347);
nand U8454 (N_8454,N_8322,N_8360);
nand U8455 (N_8455,N_8342,N_8393);
or U8456 (N_8456,N_8397,N_8378);
xnor U8457 (N_8457,N_8371,N_8353);
nor U8458 (N_8458,N_8344,N_8356);
nor U8459 (N_8459,N_8329,N_8382);
or U8460 (N_8460,N_8357,N_8339);
nand U8461 (N_8461,N_8352,N_8370);
xnor U8462 (N_8462,N_8378,N_8391);
nand U8463 (N_8463,N_8356,N_8342);
nand U8464 (N_8464,N_8387,N_8398);
xnor U8465 (N_8465,N_8392,N_8359);
nor U8466 (N_8466,N_8331,N_8324);
nand U8467 (N_8467,N_8377,N_8375);
nand U8468 (N_8468,N_8330,N_8309);
or U8469 (N_8469,N_8314,N_8360);
and U8470 (N_8470,N_8328,N_8399);
and U8471 (N_8471,N_8323,N_8356);
or U8472 (N_8472,N_8350,N_8397);
and U8473 (N_8473,N_8328,N_8320);
and U8474 (N_8474,N_8393,N_8395);
and U8475 (N_8475,N_8350,N_8362);
or U8476 (N_8476,N_8397,N_8346);
and U8477 (N_8477,N_8325,N_8329);
and U8478 (N_8478,N_8305,N_8367);
or U8479 (N_8479,N_8377,N_8399);
or U8480 (N_8480,N_8388,N_8362);
xor U8481 (N_8481,N_8315,N_8398);
nor U8482 (N_8482,N_8387,N_8308);
and U8483 (N_8483,N_8393,N_8386);
nand U8484 (N_8484,N_8385,N_8357);
xnor U8485 (N_8485,N_8346,N_8333);
and U8486 (N_8486,N_8374,N_8386);
or U8487 (N_8487,N_8386,N_8334);
xor U8488 (N_8488,N_8368,N_8301);
or U8489 (N_8489,N_8375,N_8344);
and U8490 (N_8490,N_8381,N_8339);
or U8491 (N_8491,N_8321,N_8342);
or U8492 (N_8492,N_8374,N_8328);
nor U8493 (N_8493,N_8331,N_8323);
or U8494 (N_8494,N_8342,N_8391);
xor U8495 (N_8495,N_8348,N_8392);
and U8496 (N_8496,N_8357,N_8383);
xnor U8497 (N_8497,N_8368,N_8308);
or U8498 (N_8498,N_8305,N_8349);
and U8499 (N_8499,N_8317,N_8343);
and U8500 (N_8500,N_8474,N_8458);
nand U8501 (N_8501,N_8447,N_8407);
xnor U8502 (N_8502,N_8466,N_8424);
nand U8503 (N_8503,N_8443,N_8486);
or U8504 (N_8504,N_8448,N_8459);
or U8505 (N_8505,N_8436,N_8465);
or U8506 (N_8506,N_8472,N_8419);
nand U8507 (N_8507,N_8430,N_8422);
nand U8508 (N_8508,N_8435,N_8439);
nor U8509 (N_8509,N_8417,N_8445);
nand U8510 (N_8510,N_8434,N_8483);
xnor U8511 (N_8511,N_8457,N_8451);
nand U8512 (N_8512,N_8441,N_8491);
nor U8513 (N_8513,N_8489,N_8495);
and U8514 (N_8514,N_8473,N_8452);
and U8515 (N_8515,N_8454,N_8453);
nor U8516 (N_8516,N_8410,N_8493);
and U8517 (N_8517,N_8403,N_8461);
nor U8518 (N_8518,N_8478,N_8433);
nor U8519 (N_8519,N_8450,N_8428);
nand U8520 (N_8520,N_8449,N_8400);
nand U8521 (N_8521,N_8405,N_8496);
xor U8522 (N_8522,N_8494,N_8477);
nor U8523 (N_8523,N_8423,N_8411);
and U8524 (N_8524,N_8416,N_8426);
or U8525 (N_8525,N_8427,N_8498);
nor U8526 (N_8526,N_8404,N_8485);
and U8527 (N_8527,N_8431,N_8415);
xor U8528 (N_8528,N_8421,N_8464);
or U8529 (N_8529,N_8438,N_8409);
and U8530 (N_8530,N_8475,N_8455);
nor U8531 (N_8531,N_8440,N_8490);
and U8532 (N_8532,N_8460,N_8492);
nand U8533 (N_8533,N_8414,N_8462);
or U8534 (N_8534,N_8412,N_8484);
nor U8535 (N_8535,N_8401,N_8480);
and U8536 (N_8536,N_8463,N_8476);
nand U8537 (N_8537,N_8408,N_8470);
and U8538 (N_8538,N_8442,N_8482);
nor U8539 (N_8539,N_8481,N_8479);
nand U8540 (N_8540,N_8499,N_8402);
and U8541 (N_8541,N_8425,N_8418);
nand U8542 (N_8542,N_8469,N_8437);
nand U8543 (N_8543,N_8456,N_8406);
or U8544 (N_8544,N_8471,N_8487);
nor U8545 (N_8545,N_8488,N_8497);
and U8546 (N_8546,N_8467,N_8420);
nand U8547 (N_8547,N_8446,N_8468);
nand U8548 (N_8548,N_8444,N_8432);
nor U8549 (N_8549,N_8413,N_8429);
nor U8550 (N_8550,N_8439,N_8484);
or U8551 (N_8551,N_8488,N_8408);
xor U8552 (N_8552,N_8444,N_8409);
nand U8553 (N_8553,N_8488,N_8483);
and U8554 (N_8554,N_8415,N_8463);
and U8555 (N_8555,N_8426,N_8412);
xor U8556 (N_8556,N_8419,N_8462);
xnor U8557 (N_8557,N_8407,N_8437);
nand U8558 (N_8558,N_8485,N_8492);
xnor U8559 (N_8559,N_8439,N_8468);
xnor U8560 (N_8560,N_8451,N_8493);
or U8561 (N_8561,N_8448,N_8425);
nand U8562 (N_8562,N_8466,N_8475);
nand U8563 (N_8563,N_8423,N_8493);
xor U8564 (N_8564,N_8473,N_8405);
and U8565 (N_8565,N_8448,N_8497);
nand U8566 (N_8566,N_8459,N_8499);
nand U8567 (N_8567,N_8476,N_8418);
or U8568 (N_8568,N_8411,N_8464);
or U8569 (N_8569,N_8425,N_8467);
and U8570 (N_8570,N_8467,N_8419);
and U8571 (N_8571,N_8431,N_8403);
or U8572 (N_8572,N_8436,N_8432);
nor U8573 (N_8573,N_8440,N_8455);
or U8574 (N_8574,N_8409,N_8479);
or U8575 (N_8575,N_8459,N_8473);
nand U8576 (N_8576,N_8461,N_8427);
and U8577 (N_8577,N_8480,N_8475);
nand U8578 (N_8578,N_8465,N_8486);
and U8579 (N_8579,N_8454,N_8417);
xor U8580 (N_8580,N_8440,N_8405);
and U8581 (N_8581,N_8426,N_8453);
nand U8582 (N_8582,N_8409,N_8424);
and U8583 (N_8583,N_8468,N_8421);
xnor U8584 (N_8584,N_8476,N_8458);
nor U8585 (N_8585,N_8425,N_8452);
and U8586 (N_8586,N_8431,N_8401);
and U8587 (N_8587,N_8434,N_8415);
nand U8588 (N_8588,N_8480,N_8474);
and U8589 (N_8589,N_8470,N_8448);
xnor U8590 (N_8590,N_8489,N_8496);
nand U8591 (N_8591,N_8419,N_8421);
or U8592 (N_8592,N_8484,N_8414);
xnor U8593 (N_8593,N_8482,N_8437);
xnor U8594 (N_8594,N_8433,N_8477);
or U8595 (N_8595,N_8447,N_8401);
nand U8596 (N_8596,N_8487,N_8481);
or U8597 (N_8597,N_8408,N_8468);
or U8598 (N_8598,N_8485,N_8450);
or U8599 (N_8599,N_8485,N_8446);
nor U8600 (N_8600,N_8547,N_8546);
and U8601 (N_8601,N_8510,N_8524);
xnor U8602 (N_8602,N_8521,N_8571);
or U8603 (N_8603,N_8552,N_8563);
or U8604 (N_8604,N_8588,N_8525);
nand U8605 (N_8605,N_8504,N_8584);
nor U8606 (N_8606,N_8508,N_8570);
xor U8607 (N_8607,N_8505,N_8590);
nand U8608 (N_8608,N_8578,N_8512);
or U8609 (N_8609,N_8561,N_8581);
xnor U8610 (N_8610,N_8589,N_8577);
nor U8611 (N_8611,N_8591,N_8513);
or U8612 (N_8612,N_8569,N_8520);
or U8613 (N_8613,N_8553,N_8593);
xnor U8614 (N_8614,N_8592,N_8599);
and U8615 (N_8615,N_8507,N_8534);
or U8616 (N_8616,N_8511,N_8559);
or U8617 (N_8617,N_8551,N_8537);
nor U8618 (N_8618,N_8536,N_8500);
xor U8619 (N_8619,N_8564,N_8539);
nand U8620 (N_8620,N_8556,N_8575);
xor U8621 (N_8621,N_8568,N_8567);
or U8622 (N_8622,N_8574,N_8554);
or U8623 (N_8623,N_8565,N_8557);
or U8624 (N_8624,N_8541,N_8526);
and U8625 (N_8625,N_8515,N_8533);
nand U8626 (N_8626,N_8519,N_8550);
or U8627 (N_8627,N_8517,N_8558);
and U8628 (N_8628,N_8573,N_8518);
nor U8629 (N_8629,N_8580,N_8597);
nor U8630 (N_8630,N_8595,N_8582);
nand U8631 (N_8631,N_8528,N_8501);
xor U8632 (N_8632,N_8598,N_8543);
and U8633 (N_8633,N_8585,N_8545);
nand U8634 (N_8634,N_8540,N_8502);
and U8635 (N_8635,N_8522,N_8560);
nand U8636 (N_8636,N_8586,N_8503);
and U8637 (N_8637,N_8566,N_8538);
or U8638 (N_8638,N_8555,N_8596);
nand U8639 (N_8639,N_8583,N_8548);
nor U8640 (N_8640,N_8562,N_8509);
xor U8641 (N_8641,N_8506,N_8579);
and U8642 (N_8642,N_8572,N_8516);
or U8643 (N_8643,N_8594,N_8544);
xnor U8644 (N_8644,N_8531,N_8527);
xnor U8645 (N_8645,N_8587,N_8530);
nor U8646 (N_8646,N_8549,N_8529);
nor U8647 (N_8647,N_8514,N_8532);
nor U8648 (N_8648,N_8576,N_8523);
and U8649 (N_8649,N_8535,N_8542);
nor U8650 (N_8650,N_8559,N_8545);
xnor U8651 (N_8651,N_8554,N_8521);
nor U8652 (N_8652,N_8562,N_8529);
xnor U8653 (N_8653,N_8541,N_8537);
and U8654 (N_8654,N_8597,N_8560);
nor U8655 (N_8655,N_8595,N_8589);
xnor U8656 (N_8656,N_8519,N_8503);
nand U8657 (N_8657,N_8503,N_8557);
nand U8658 (N_8658,N_8554,N_8583);
xor U8659 (N_8659,N_8588,N_8538);
nor U8660 (N_8660,N_8571,N_8541);
and U8661 (N_8661,N_8530,N_8571);
and U8662 (N_8662,N_8534,N_8558);
nand U8663 (N_8663,N_8566,N_8534);
and U8664 (N_8664,N_8560,N_8541);
and U8665 (N_8665,N_8591,N_8597);
xor U8666 (N_8666,N_8561,N_8591);
nand U8667 (N_8667,N_8593,N_8536);
xor U8668 (N_8668,N_8505,N_8512);
xor U8669 (N_8669,N_8528,N_8568);
nor U8670 (N_8670,N_8593,N_8506);
and U8671 (N_8671,N_8564,N_8536);
or U8672 (N_8672,N_8503,N_8535);
and U8673 (N_8673,N_8521,N_8558);
nor U8674 (N_8674,N_8529,N_8582);
or U8675 (N_8675,N_8562,N_8591);
nand U8676 (N_8676,N_8570,N_8595);
nand U8677 (N_8677,N_8530,N_8585);
and U8678 (N_8678,N_8542,N_8584);
and U8679 (N_8679,N_8550,N_8588);
nand U8680 (N_8680,N_8524,N_8523);
xnor U8681 (N_8681,N_8595,N_8536);
nor U8682 (N_8682,N_8522,N_8536);
xor U8683 (N_8683,N_8507,N_8566);
or U8684 (N_8684,N_8511,N_8553);
nor U8685 (N_8685,N_8566,N_8562);
xnor U8686 (N_8686,N_8521,N_8569);
nor U8687 (N_8687,N_8530,N_8575);
and U8688 (N_8688,N_8585,N_8509);
or U8689 (N_8689,N_8543,N_8549);
or U8690 (N_8690,N_8585,N_8514);
and U8691 (N_8691,N_8561,N_8515);
nor U8692 (N_8692,N_8586,N_8501);
nand U8693 (N_8693,N_8569,N_8560);
and U8694 (N_8694,N_8597,N_8550);
or U8695 (N_8695,N_8549,N_8592);
xor U8696 (N_8696,N_8515,N_8505);
or U8697 (N_8697,N_8544,N_8506);
or U8698 (N_8698,N_8558,N_8543);
and U8699 (N_8699,N_8555,N_8563);
or U8700 (N_8700,N_8682,N_8685);
and U8701 (N_8701,N_8627,N_8650);
xor U8702 (N_8702,N_8673,N_8640);
and U8703 (N_8703,N_8602,N_8616);
xnor U8704 (N_8704,N_8658,N_8660);
or U8705 (N_8705,N_8646,N_8600);
nand U8706 (N_8706,N_8611,N_8678);
nand U8707 (N_8707,N_8648,N_8626);
nor U8708 (N_8708,N_8609,N_8676);
nor U8709 (N_8709,N_8649,N_8659);
nor U8710 (N_8710,N_8645,N_8657);
nor U8711 (N_8711,N_8621,N_8656);
or U8712 (N_8712,N_8653,N_8624);
and U8713 (N_8713,N_8647,N_8641);
or U8714 (N_8714,N_8684,N_8638);
xor U8715 (N_8715,N_8628,N_8692);
nand U8716 (N_8716,N_8669,N_8622);
or U8717 (N_8717,N_8671,N_8619);
xor U8718 (N_8718,N_8630,N_8661);
nor U8719 (N_8719,N_8634,N_8698);
nor U8720 (N_8720,N_8618,N_8690);
or U8721 (N_8721,N_8620,N_8691);
nand U8722 (N_8722,N_8695,N_8686);
or U8723 (N_8723,N_8694,N_8606);
or U8724 (N_8724,N_8625,N_8636);
nor U8725 (N_8725,N_8674,N_8672);
nand U8726 (N_8726,N_8605,N_8629);
or U8727 (N_8727,N_8668,N_8681);
nand U8728 (N_8728,N_8631,N_8607);
nor U8729 (N_8729,N_8655,N_8652);
nand U8730 (N_8730,N_8683,N_8603);
and U8731 (N_8731,N_8635,N_8617);
and U8732 (N_8732,N_8675,N_8637);
nor U8733 (N_8733,N_8664,N_8687);
nand U8734 (N_8734,N_8693,N_8665);
or U8735 (N_8735,N_8614,N_8612);
xor U8736 (N_8736,N_8639,N_8677);
and U8737 (N_8737,N_8642,N_8601);
nor U8738 (N_8738,N_8604,N_8696);
and U8739 (N_8739,N_8654,N_8651);
xor U8740 (N_8740,N_8689,N_8670);
nand U8741 (N_8741,N_8644,N_8697);
and U8742 (N_8742,N_8643,N_8699);
and U8743 (N_8743,N_8623,N_8613);
xor U8744 (N_8744,N_8679,N_8663);
or U8745 (N_8745,N_8666,N_8662);
nand U8746 (N_8746,N_8667,N_8632);
xnor U8747 (N_8747,N_8633,N_8608);
xor U8748 (N_8748,N_8680,N_8610);
nand U8749 (N_8749,N_8688,N_8615);
nand U8750 (N_8750,N_8685,N_8668);
and U8751 (N_8751,N_8698,N_8656);
xnor U8752 (N_8752,N_8604,N_8693);
xnor U8753 (N_8753,N_8695,N_8611);
xor U8754 (N_8754,N_8652,N_8624);
nand U8755 (N_8755,N_8684,N_8649);
or U8756 (N_8756,N_8686,N_8685);
nor U8757 (N_8757,N_8665,N_8644);
xor U8758 (N_8758,N_8623,N_8682);
nand U8759 (N_8759,N_8689,N_8695);
and U8760 (N_8760,N_8696,N_8605);
or U8761 (N_8761,N_8679,N_8684);
nand U8762 (N_8762,N_8662,N_8612);
or U8763 (N_8763,N_8631,N_8698);
nand U8764 (N_8764,N_8607,N_8653);
nor U8765 (N_8765,N_8685,N_8687);
nor U8766 (N_8766,N_8665,N_8603);
and U8767 (N_8767,N_8620,N_8680);
and U8768 (N_8768,N_8610,N_8645);
xnor U8769 (N_8769,N_8604,N_8690);
xnor U8770 (N_8770,N_8634,N_8690);
nand U8771 (N_8771,N_8601,N_8683);
or U8772 (N_8772,N_8670,N_8620);
or U8773 (N_8773,N_8671,N_8613);
xnor U8774 (N_8774,N_8624,N_8610);
or U8775 (N_8775,N_8639,N_8616);
nor U8776 (N_8776,N_8645,N_8611);
xnor U8777 (N_8777,N_8659,N_8620);
or U8778 (N_8778,N_8668,N_8607);
nand U8779 (N_8779,N_8671,N_8621);
nand U8780 (N_8780,N_8643,N_8634);
and U8781 (N_8781,N_8648,N_8681);
and U8782 (N_8782,N_8658,N_8604);
nand U8783 (N_8783,N_8682,N_8666);
nor U8784 (N_8784,N_8634,N_8665);
nand U8785 (N_8785,N_8696,N_8661);
xor U8786 (N_8786,N_8647,N_8686);
nor U8787 (N_8787,N_8664,N_8606);
nor U8788 (N_8788,N_8603,N_8617);
nand U8789 (N_8789,N_8613,N_8684);
or U8790 (N_8790,N_8680,N_8632);
nand U8791 (N_8791,N_8655,N_8618);
and U8792 (N_8792,N_8670,N_8674);
and U8793 (N_8793,N_8691,N_8667);
nor U8794 (N_8794,N_8649,N_8635);
xnor U8795 (N_8795,N_8672,N_8625);
nand U8796 (N_8796,N_8693,N_8690);
or U8797 (N_8797,N_8685,N_8693);
nor U8798 (N_8798,N_8684,N_8651);
nand U8799 (N_8799,N_8610,N_8657);
and U8800 (N_8800,N_8737,N_8731);
or U8801 (N_8801,N_8714,N_8722);
or U8802 (N_8802,N_8774,N_8759);
and U8803 (N_8803,N_8794,N_8718);
nand U8804 (N_8804,N_8781,N_8777);
nor U8805 (N_8805,N_8790,N_8705);
and U8806 (N_8806,N_8709,N_8746);
or U8807 (N_8807,N_8711,N_8796);
nand U8808 (N_8808,N_8784,N_8701);
xnor U8809 (N_8809,N_8773,N_8767);
nor U8810 (N_8810,N_8761,N_8712);
nor U8811 (N_8811,N_8729,N_8721);
or U8812 (N_8812,N_8710,N_8719);
and U8813 (N_8813,N_8752,N_8788);
or U8814 (N_8814,N_8785,N_8734);
xor U8815 (N_8815,N_8726,N_8708);
or U8816 (N_8816,N_8793,N_8716);
nand U8817 (N_8817,N_8736,N_8727);
or U8818 (N_8818,N_8769,N_8743);
nand U8819 (N_8819,N_8754,N_8782);
and U8820 (N_8820,N_8786,N_8768);
xor U8821 (N_8821,N_8740,N_8762);
nand U8822 (N_8822,N_8750,N_8792);
nor U8823 (N_8823,N_8733,N_8749);
nand U8824 (N_8824,N_8715,N_8730);
nor U8825 (N_8825,N_8779,N_8707);
nand U8826 (N_8826,N_8778,N_8798);
and U8827 (N_8827,N_8756,N_8775);
xnor U8828 (N_8828,N_8706,N_8765);
nor U8829 (N_8829,N_8787,N_8772);
or U8830 (N_8830,N_8735,N_8745);
nor U8831 (N_8831,N_8702,N_8725);
and U8832 (N_8832,N_8732,N_8744);
nor U8833 (N_8833,N_8783,N_8713);
xor U8834 (N_8834,N_8728,N_8724);
or U8835 (N_8835,N_8789,N_8766);
and U8836 (N_8836,N_8720,N_8753);
or U8837 (N_8837,N_8797,N_8776);
xnor U8838 (N_8838,N_8791,N_8780);
nor U8839 (N_8839,N_8704,N_8723);
nand U8840 (N_8840,N_8741,N_8748);
nand U8841 (N_8841,N_8795,N_8703);
nor U8842 (N_8842,N_8755,N_8771);
xnor U8843 (N_8843,N_8739,N_8738);
or U8844 (N_8844,N_8717,N_8763);
xor U8845 (N_8845,N_8764,N_8751);
nor U8846 (N_8846,N_8742,N_8770);
nand U8847 (N_8847,N_8747,N_8760);
and U8848 (N_8848,N_8757,N_8700);
or U8849 (N_8849,N_8758,N_8799);
and U8850 (N_8850,N_8782,N_8770);
nor U8851 (N_8851,N_8743,N_8732);
and U8852 (N_8852,N_8787,N_8788);
and U8853 (N_8853,N_8780,N_8760);
nor U8854 (N_8854,N_8751,N_8742);
or U8855 (N_8855,N_8775,N_8774);
nand U8856 (N_8856,N_8702,N_8727);
or U8857 (N_8857,N_8759,N_8770);
nand U8858 (N_8858,N_8717,N_8711);
or U8859 (N_8859,N_8706,N_8713);
nand U8860 (N_8860,N_8751,N_8795);
nand U8861 (N_8861,N_8789,N_8779);
nor U8862 (N_8862,N_8762,N_8706);
or U8863 (N_8863,N_8796,N_8742);
nor U8864 (N_8864,N_8701,N_8775);
or U8865 (N_8865,N_8764,N_8741);
nor U8866 (N_8866,N_8790,N_8761);
or U8867 (N_8867,N_8772,N_8789);
xnor U8868 (N_8868,N_8768,N_8739);
xor U8869 (N_8869,N_8747,N_8709);
nor U8870 (N_8870,N_8722,N_8771);
xnor U8871 (N_8871,N_8703,N_8747);
and U8872 (N_8872,N_8756,N_8751);
and U8873 (N_8873,N_8762,N_8797);
and U8874 (N_8874,N_8735,N_8720);
nand U8875 (N_8875,N_8713,N_8765);
or U8876 (N_8876,N_8753,N_8796);
xor U8877 (N_8877,N_8703,N_8749);
xor U8878 (N_8878,N_8757,N_8794);
nor U8879 (N_8879,N_8728,N_8753);
nor U8880 (N_8880,N_8716,N_8757);
nor U8881 (N_8881,N_8791,N_8742);
nand U8882 (N_8882,N_8795,N_8735);
xnor U8883 (N_8883,N_8752,N_8798);
or U8884 (N_8884,N_8773,N_8740);
or U8885 (N_8885,N_8775,N_8742);
nand U8886 (N_8886,N_8711,N_8763);
nor U8887 (N_8887,N_8700,N_8704);
or U8888 (N_8888,N_8741,N_8731);
nand U8889 (N_8889,N_8795,N_8706);
xnor U8890 (N_8890,N_8757,N_8768);
nor U8891 (N_8891,N_8798,N_8729);
or U8892 (N_8892,N_8799,N_8736);
xnor U8893 (N_8893,N_8722,N_8710);
xnor U8894 (N_8894,N_8794,N_8785);
or U8895 (N_8895,N_8790,N_8755);
nand U8896 (N_8896,N_8715,N_8775);
and U8897 (N_8897,N_8793,N_8747);
nor U8898 (N_8898,N_8703,N_8792);
nand U8899 (N_8899,N_8729,N_8774);
and U8900 (N_8900,N_8811,N_8803);
or U8901 (N_8901,N_8892,N_8879);
nand U8902 (N_8902,N_8802,N_8804);
nor U8903 (N_8903,N_8812,N_8881);
nor U8904 (N_8904,N_8841,N_8815);
and U8905 (N_8905,N_8859,N_8860);
xnor U8906 (N_8906,N_8864,N_8883);
or U8907 (N_8907,N_8897,N_8844);
nor U8908 (N_8908,N_8895,N_8828);
nor U8909 (N_8909,N_8869,N_8855);
xor U8910 (N_8910,N_8850,N_8849);
or U8911 (N_8911,N_8848,N_8831);
and U8912 (N_8912,N_8874,N_8805);
nor U8913 (N_8913,N_8870,N_8889);
or U8914 (N_8914,N_8851,N_8830);
nand U8915 (N_8915,N_8840,N_8878);
or U8916 (N_8916,N_8833,N_8838);
and U8917 (N_8917,N_8886,N_8842);
nand U8918 (N_8918,N_8807,N_8884);
and U8919 (N_8919,N_8827,N_8819);
xnor U8920 (N_8920,N_8877,N_8865);
and U8921 (N_8921,N_8809,N_8836);
or U8922 (N_8922,N_8834,N_8832);
xnor U8923 (N_8923,N_8888,N_8854);
xor U8924 (N_8924,N_8891,N_8867);
nand U8925 (N_8925,N_8835,N_8861);
xnor U8926 (N_8926,N_8856,N_8818);
and U8927 (N_8927,N_8837,N_8885);
or U8928 (N_8928,N_8847,N_8871);
nand U8929 (N_8929,N_8813,N_8800);
and U8930 (N_8930,N_8887,N_8825);
and U8931 (N_8931,N_8823,N_8820);
xor U8932 (N_8932,N_8882,N_8817);
xnor U8933 (N_8933,N_8829,N_8898);
or U8934 (N_8934,N_8866,N_8808);
nand U8935 (N_8935,N_8857,N_8826);
nand U8936 (N_8936,N_8806,N_8868);
or U8937 (N_8937,N_8846,N_8858);
and U8938 (N_8938,N_8872,N_8824);
nand U8939 (N_8939,N_8899,N_8875);
nand U8940 (N_8940,N_8894,N_8839);
nand U8941 (N_8941,N_8880,N_8893);
nand U8942 (N_8942,N_8873,N_8801);
xnor U8943 (N_8943,N_8896,N_8853);
nor U8944 (N_8944,N_8845,N_8822);
xnor U8945 (N_8945,N_8814,N_8890);
or U8946 (N_8946,N_8821,N_8852);
nand U8947 (N_8947,N_8816,N_8863);
nor U8948 (N_8948,N_8876,N_8810);
and U8949 (N_8949,N_8843,N_8862);
xor U8950 (N_8950,N_8844,N_8801);
xor U8951 (N_8951,N_8851,N_8896);
and U8952 (N_8952,N_8888,N_8837);
nand U8953 (N_8953,N_8803,N_8852);
nand U8954 (N_8954,N_8804,N_8895);
nor U8955 (N_8955,N_8801,N_8867);
nand U8956 (N_8956,N_8851,N_8852);
and U8957 (N_8957,N_8804,N_8821);
and U8958 (N_8958,N_8811,N_8834);
nand U8959 (N_8959,N_8862,N_8848);
nor U8960 (N_8960,N_8809,N_8874);
xnor U8961 (N_8961,N_8824,N_8893);
nand U8962 (N_8962,N_8850,N_8893);
nand U8963 (N_8963,N_8808,N_8855);
nor U8964 (N_8964,N_8850,N_8853);
or U8965 (N_8965,N_8856,N_8896);
nor U8966 (N_8966,N_8885,N_8842);
xnor U8967 (N_8967,N_8825,N_8883);
or U8968 (N_8968,N_8815,N_8833);
and U8969 (N_8969,N_8806,N_8829);
nor U8970 (N_8970,N_8800,N_8893);
nor U8971 (N_8971,N_8823,N_8821);
nor U8972 (N_8972,N_8832,N_8824);
or U8973 (N_8973,N_8855,N_8879);
or U8974 (N_8974,N_8859,N_8886);
nand U8975 (N_8975,N_8853,N_8871);
and U8976 (N_8976,N_8869,N_8848);
or U8977 (N_8977,N_8814,N_8869);
xnor U8978 (N_8978,N_8840,N_8846);
or U8979 (N_8979,N_8882,N_8849);
and U8980 (N_8980,N_8802,N_8816);
nand U8981 (N_8981,N_8850,N_8828);
nor U8982 (N_8982,N_8809,N_8817);
xor U8983 (N_8983,N_8885,N_8819);
or U8984 (N_8984,N_8877,N_8891);
or U8985 (N_8985,N_8858,N_8898);
xnor U8986 (N_8986,N_8875,N_8866);
and U8987 (N_8987,N_8853,N_8820);
or U8988 (N_8988,N_8863,N_8800);
nand U8989 (N_8989,N_8815,N_8831);
nand U8990 (N_8990,N_8856,N_8881);
nor U8991 (N_8991,N_8823,N_8846);
nand U8992 (N_8992,N_8809,N_8855);
and U8993 (N_8993,N_8897,N_8801);
nand U8994 (N_8994,N_8829,N_8864);
and U8995 (N_8995,N_8825,N_8878);
xor U8996 (N_8996,N_8821,N_8814);
or U8997 (N_8997,N_8853,N_8858);
nand U8998 (N_8998,N_8890,N_8839);
nor U8999 (N_8999,N_8893,N_8869);
and U9000 (N_9000,N_8934,N_8984);
nand U9001 (N_9001,N_8906,N_8926);
and U9002 (N_9002,N_8933,N_8917);
and U9003 (N_9003,N_8967,N_8935);
xor U9004 (N_9004,N_8937,N_8980);
or U9005 (N_9005,N_8914,N_8954);
nor U9006 (N_9006,N_8998,N_8989);
or U9007 (N_9007,N_8952,N_8949);
or U9008 (N_9008,N_8997,N_8901);
or U9009 (N_9009,N_8922,N_8921);
and U9010 (N_9010,N_8902,N_8929);
or U9011 (N_9011,N_8981,N_8945);
or U9012 (N_9012,N_8968,N_8931);
nor U9013 (N_9013,N_8900,N_8932);
nor U9014 (N_9014,N_8969,N_8919);
or U9015 (N_9015,N_8973,N_8999);
and U9016 (N_9016,N_8985,N_8951);
and U9017 (N_9017,N_8909,N_8944);
or U9018 (N_9018,N_8913,N_8971);
and U9019 (N_9019,N_8930,N_8943);
and U9020 (N_9020,N_8965,N_8963);
nor U9021 (N_9021,N_8987,N_8941);
and U9022 (N_9022,N_8915,N_8918);
nand U9023 (N_9023,N_8908,N_8978);
xor U9024 (N_9024,N_8962,N_8972);
nor U9025 (N_9025,N_8916,N_8912);
and U9026 (N_9026,N_8955,N_8996);
or U9027 (N_9027,N_8920,N_8975);
xnor U9028 (N_9028,N_8905,N_8961);
nor U9029 (N_9029,N_8979,N_8947);
nor U9030 (N_9030,N_8924,N_8904);
xor U9031 (N_9031,N_8942,N_8957);
xnor U9032 (N_9032,N_8946,N_8960);
or U9033 (N_9033,N_8976,N_8990);
nor U9034 (N_9034,N_8948,N_8910);
nor U9035 (N_9035,N_8982,N_8995);
and U9036 (N_9036,N_8994,N_8992);
or U9037 (N_9037,N_8966,N_8938);
nor U9038 (N_9038,N_8940,N_8956);
nand U9039 (N_9039,N_8964,N_8923);
nand U9040 (N_9040,N_8983,N_8939);
xor U9041 (N_9041,N_8950,N_8927);
or U9042 (N_9042,N_8959,N_8958);
and U9043 (N_9043,N_8903,N_8936);
nand U9044 (N_9044,N_8988,N_8970);
nand U9045 (N_9045,N_8953,N_8986);
nor U9046 (N_9046,N_8911,N_8993);
or U9047 (N_9047,N_8925,N_8977);
and U9048 (N_9048,N_8974,N_8928);
nand U9049 (N_9049,N_8907,N_8991);
xor U9050 (N_9050,N_8996,N_8932);
xor U9051 (N_9051,N_8970,N_8980);
or U9052 (N_9052,N_8979,N_8977);
nor U9053 (N_9053,N_8901,N_8956);
or U9054 (N_9054,N_8952,N_8929);
nor U9055 (N_9055,N_8911,N_8929);
xnor U9056 (N_9056,N_8979,N_8922);
xnor U9057 (N_9057,N_8926,N_8909);
or U9058 (N_9058,N_8988,N_8937);
and U9059 (N_9059,N_8947,N_8918);
nand U9060 (N_9060,N_8942,N_8974);
nor U9061 (N_9061,N_8997,N_8922);
nand U9062 (N_9062,N_8912,N_8917);
and U9063 (N_9063,N_8903,N_8983);
xnor U9064 (N_9064,N_8950,N_8908);
and U9065 (N_9065,N_8997,N_8985);
and U9066 (N_9066,N_8912,N_8973);
xor U9067 (N_9067,N_8995,N_8926);
and U9068 (N_9068,N_8938,N_8970);
xor U9069 (N_9069,N_8913,N_8942);
and U9070 (N_9070,N_8999,N_8949);
or U9071 (N_9071,N_8932,N_8947);
xnor U9072 (N_9072,N_8934,N_8971);
and U9073 (N_9073,N_8911,N_8907);
nand U9074 (N_9074,N_8997,N_8912);
and U9075 (N_9075,N_8996,N_8988);
nand U9076 (N_9076,N_8992,N_8956);
xor U9077 (N_9077,N_8968,N_8998);
and U9078 (N_9078,N_8978,N_8926);
and U9079 (N_9079,N_8992,N_8909);
or U9080 (N_9080,N_8994,N_8950);
or U9081 (N_9081,N_8917,N_8944);
nand U9082 (N_9082,N_8955,N_8950);
and U9083 (N_9083,N_8947,N_8923);
xnor U9084 (N_9084,N_8955,N_8918);
or U9085 (N_9085,N_8909,N_8907);
and U9086 (N_9086,N_8929,N_8998);
nor U9087 (N_9087,N_8969,N_8943);
or U9088 (N_9088,N_8945,N_8987);
nand U9089 (N_9089,N_8927,N_8981);
nor U9090 (N_9090,N_8932,N_8978);
nand U9091 (N_9091,N_8999,N_8954);
nand U9092 (N_9092,N_8948,N_8998);
nand U9093 (N_9093,N_8965,N_8920);
xnor U9094 (N_9094,N_8942,N_8960);
and U9095 (N_9095,N_8964,N_8938);
nor U9096 (N_9096,N_8995,N_8976);
nand U9097 (N_9097,N_8960,N_8970);
xnor U9098 (N_9098,N_8943,N_8923);
xnor U9099 (N_9099,N_8971,N_8939);
and U9100 (N_9100,N_9017,N_9063);
or U9101 (N_9101,N_9083,N_9073);
nor U9102 (N_9102,N_9009,N_9027);
xnor U9103 (N_9103,N_9053,N_9041);
or U9104 (N_9104,N_9067,N_9085);
and U9105 (N_9105,N_9005,N_9084);
and U9106 (N_9106,N_9064,N_9087);
and U9107 (N_9107,N_9056,N_9057);
and U9108 (N_9108,N_9000,N_9079);
or U9109 (N_9109,N_9062,N_9013);
nor U9110 (N_9110,N_9030,N_9043);
nand U9111 (N_9111,N_9035,N_9022);
nor U9112 (N_9112,N_9003,N_9093);
nor U9113 (N_9113,N_9065,N_9008);
xor U9114 (N_9114,N_9042,N_9066);
nand U9115 (N_9115,N_9026,N_9058);
nor U9116 (N_9116,N_9034,N_9089);
nand U9117 (N_9117,N_9045,N_9007);
or U9118 (N_9118,N_9049,N_9018);
nor U9119 (N_9119,N_9046,N_9016);
or U9120 (N_9120,N_9069,N_9038);
xnor U9121 (N_9121,N_9047,N_9012);
nand U9122 (N_9122,N_9094,N_9052);
or U9123 (N_9123,N_9075,N_9039);
nand U9124 (N_9124,N_9004,N_9070);
nand U9125 (N_9125,N_9074,N_9082);
and U9126 (N_9126,N_9081,N_9090);
nand U9127 (N_9127,N_9061,N_9023);
xnor U9128 (N_9128,N_9068,N_9099);
nand U9129 (N_9129,N_9037,N_9051);
and U9130 (N_9130,N_9060,N_9033);
nand U9131 (N_9131,N_9072,N_9015);
xnor U9132 (N_9132,N_9019,N_9029);
or U9133 (N_9133,N_9076,N_9097);
nor U9134 (N_9134,N_9011,N_9086);
or U9135 (N_9135,N_9088,N_9092);
xnor U9136 (N_9136,N_9031,N_9077);
and U9137 (N_9137,N_9048,N_9040);
xor U9138 (N_9138,N_9006,N_9096);
and U9139 (N_9139,N_9050,N_9024);
or U9140 (N_9140,N_9071,N_9021);
and U9141 (N_9141,N_9014,N_9080);
xor U9142 (N_9142,N_9036,N_9059);
nor U9143 (N_9143,N_9032,N_9078);
xnor U9144 (N_9144,N_9055,N_9028);
or U9145 (N_9145,N_9054,N_9095);
nand U9146 (N_9146,N_9010,N_9044);
or U9147 (N_9147,N_9025,N_9001);
and U9148 (N_9148,N_9091,N_9098);
and U9149 (N_9149,N_9020,N_9002);
nand U9150 (N_9150,N_9095,N_9005);
nor U9151 (N_9151,N_9015,N_9009);
xor U9152 (N_9152,N_9050,N_9059);
nor U9153 (N_9153,N_9037,N_9065);
xnor U9154 (N_9154,N_9080,N_9096);
and U9155 (N_9155,N_9084,N_9094);
nand U9156 (N_9156,N_9075,N_9081);
or U9157 (N_9157,N_9077,N_9014);
nor U9158 (N_9158,N_9046,N_9058);
nor U9159 (N_9159,N_9029,N_9060);
nand U9160 (N_9160,N_9077,N_9006);
nor U9161 (N_9161,N_9093,N_9074);
xor U9162 (N_9162,N_9082,N_9018);
nor U9163 (N_9163,N_9024,N_9033);
xnor U9164 (N_9164,N_9034,N_9044);
or U9165 (N_9165,N_9019,N_9077);
xnor U9166 (N_9166,N_9072,N_9090);
xor U9167 (N_9167,N_9089,N_9015);
nand U9168 (N_9168,N_9080,N_9020);
or U9169 (N_9169,N_9090,N_9088);
and U9170 (N_9170,N_9046,N_9076);
nand U9171 (N_9171,N_9018,N_9003);
and U9172 (N_9172,N_9091,N_9089);
xor U9173 (N_9173,N_9082,N_9027);
or U9174 (N_9174,N_9047,N_9069);
nor U9175 (N_9175,N_9055,N_9080);
nor U9176 (N_9176,N_9078,N_9017);
nand U9177 (N_9177,N_9093,N_9031);
or U9178 (N_9178,N_9030,N_9032);
xor U9179 (N_9179,N_9030,N_9040);
xnor U9180 (N_9180,N_9042,N_9096);
nand U9181 (N_9181,N_9063,N_9050);
nor U9182 (N_9182,N_9050,N_9011);
nand U9183 (N_9183,N_9088,N_9036);
nand U9184 (N_9184,N_9037,N_9014);
and U9185 (N_9185,N_9025,N_9062);
nand U9186 (N_9186,N_9096,N_9001);
nor U9187 (N_9187,N_9052,N_9077);
and U9188 (N_9188,N_9088,N_9035);
nor U9189 (N_9189,N_9031,N_9060);
and U9190 (N_9190,N_9058,N_9060);
nand U9191 (N_9191,N_9025,N_9040);
xor U9192 (N_9192,N_9001,N_9038);
xor U9193 (N_9193,N_9099,N_9095);
and U9194 (N_9194,N_9022,N_9074);
nor U9195 (N_9195,N_9092,N_9032);
nor U9196 (N_9196,N_9071,N_9068);
or U9197 (N_9197,N_9033,N_9058);
and U9198 (N_9198,N_9076,N_9037);
nor U9199 (N_9199,N_9063,N_9008);
or U9200 (N_9200,N_9166,N_9163);
nand U9201 (N_9201,N_9179,N_9183);
nor U9202 (N_9202,N_9191,N_9196);
xnor U9203 (N_9203,N_9198,N_9195);
and U9204 (N_9204,N_9103,N_9128);
xnor U9205 (N_9205,N_9168,N_9169);
nand U9206 (N_9206,N_9123,N_9127);
nand U9207 (N_9207,N_9100,N_9124);
nand U9208 (N_9208,N_9162,N_9199);
xnor U9209 (N_9209,N_9176,N_9170);
xnor U9210 (N_9210,N_9133,N_9137);
nor U9211 (N_9211,N_9154,N_9151);
nand U9212 (N_9212,N_9145,N_9165);
or U9213 (N_9213,N_9104,N_9114);
or U9214 (N_9214,N_9186,N_9140);
or U9215 (N_9215,N_9105,N_9129);
nor U9216 (N_9216,N_9190,N_9184);
and U9217 (N_9217,N_9138,N_9119);
or U9218 (N_9218,N_9153,N_9171);
and U9219 (N_9219,N_9141,N_9150);
nand U9220 (N_9220,N_9108,N_9106);
xnor U9221 (N_9221,N_9120,N_9117);
nand U9222 (N_9222,N_9110,N_9102);
or U9223 (N_9223,N_9172,N_9155);
nor U9224 (N_9224,N_9136,N_9160);
nor U9225 (N_9225,N_9157,N_9126);
and U9226 (N_9226,N_9132,N_9152);
xnor U9227 (N_9227,N_9115,N_9156);
nand U9228 (N_9228,N_9142,N_9146);
and U9229 (N_9229,N_9118,N_9122);
and U9230 (N_9230,N_9148,N_9107);
or U9231 (N_9231,N_9144,N_9193);
xor U9232 (N_9232,N_9139,N_9164);
xor U9233 (N_9233,N_9113,N_9189);
and U9234 (N_9234,N_9161,N_9109);
nand U9235 (N_9235,N_9130,N_9147);
nor U9236 (N_9236,N_9159,N_9111);
or U9237 (N_9237,N_9116,N_9180);
nand U9238 (N_9238,N_9178,N_9182);
xnor U9239 (N_9239,N_9134,N_9158);
and U9240 (N_9240,N_9121,N_9173);
or U9241 (N_9241,N_9101,N_9112);
or U9242 (N_9242,N_9194,N_9125);
or U9243 (N_9243,N_9197,N_9177);
nand U9244 (N_9244,N_9174,N_9167);
nand U9245 (N_9245,N_9192,N_9188);
nor U9246 (N_9246,N_9143,N_9131);
nor U9247 (N_9247,N_9185,N_9175);
nor U9248 (N_9248,N_9149,N_9135);
or U9249 (N_9249,N_9187,N_9181);
and U9250 (N_9250,N_9149,N_9178);
nand U9251 (N_9251,N_9178,N_9123);
nand U9252 (N_9252,N_9192,N_9153);
xor U9253 (N_9253,N_9137,N_9116);
nand U9254 (N_9254,N_9197,N_9110);
nor U9255 (N_9255,N_9158,N_9173);
nand U9256 (N_9256,N_9169,N_9192);
nand U9257 (N_9257,N_9105,N_9161);
nor U9258 (N_9258,N_9109,N_9183);
nor U9259 (N_9259,N_9156,N_9160);
and U9260 (N_9260,N_9162,N_9150);
xor U9261 (N_9261,N_9121,N_9109);
nand U9262 (N_9262,N_9182,N_9119);
xnor U9263 (N_9263,N_9122,N_9129);
or U9264 (N_9264,N_9193,N_9131);
nand U9265 (N_9265,N_9194,N_9148);
or U9266 (N_9266,N_9175,N_9123);
nor U9267 (N_9267,N_9177,N_9151);
nor U9268 (N_9268,N_9166,N_9109);
nor U9269 (N_9269,N_9116,N_9100);
or U9270 (N_9270,N_9176,N_9190);
nor U9271 (N_9271,N_9136,N_9131);
nor U9272 (N_9272,N_9169,N_9152);
xor U9273 (N_9273,N_9189,N_9170);
and U9274 (N_9274,N_9147,N_9101);
nand U9275 (N_9275,N_9137,N_9140);
or U9276 (N_9276,N_9151,N_9199);
nor U9277 (N_9277,N_9179,N_9128);
or U9278 (N_9278,N_9116,N_9171);
nand U9279 (N_9279,N_9152,N_9165);
nand U9280 (N_9280,N_9186,N_9134);
nand U9281 (N_9281,N_9169,N_9181);
and U9282 (N_9282,N_9153,N_9127);
xor U9283 (N_9283,N_9130,N_9178);
or U9284 (N_9284,N_9157,N_9138);
xnor U9285 (N_9285,N_9192,N_9149);
xnor U9286 (N_9286,N_9114,N_9130);
xor U9287 (N_9287,N_9100,N_9134);
nor U9288 (N_9288,N_9185,N_9146);
nor U9289 (N_9289,N_9157,N_9102);
and U9290 (N_9290,N_9146,N_9104);
nand U9291 (N_9291,N_9148,N_9104);
or U9292 (N_9292,N_9100,N_9125);
xnor U9293 (N_9293,N_9184,N_9192);
nand U9294 (N_9294,N_9193,N_9142);
nand U9295 (N_9295,N_9164,N_9193);
and U9296 (N_9296,N_9137,N_9154);
and U9297 (N_9297,N_9187,N_9145);
or U9298 (N_9298,N_9104,N_9195);
or U9299 (N_9299,N_9179,N_9139);
and U9300 (N_9300,N_9219,N_9285);
xor U9301 (N_9301,N_9273,N_9266);
nor U9302 (N_9302,N_9242,N_9256);
and U9303 (N_9303,N_9252,N_9289);
nor U9304 (N_9304,N_9265,N_9294);
xor U9305 (N_9305,N_9278,N_9282);
xnor U9306 (N_9306,N_9248,N_9232);
xor U9307 (N_9307,N_9209,N_9241);
or U9308 (N_9308,N_9286,N_9246);
nand U9309 (N_9309,N_9261,N_9220);
nand U9310 (N_9310,N_9217,N_9203);
or U9311 (N_9311,N_9269,N_9293);
or U9312 (N_9312,N_9243,N_9283);
nor U9313 (N_9313,N_9224,N_9277);
nor U9314 (N_9314,N_9250,N_9247);
nand U9315 (N_9315,N_9244,N_9234);
nand U9316 (N_9316,N_9267,N_9264);
and U9317 (N_9317,N_9279,N_9290);
and U9318 (N_9318,N_9254,N_9226);
or U9319 (N_9319,N_9238,N_9263);
or U9320 (N_9320,N_9214,N_9211);
or U9321 (N_9321,N_9258,N_9291);
and U9322 (N_9322,N_9213,N_9288);
nor U9323 (N_9323,N_9268,N_9245);
nor U9324 (N_9324,N_9299,N_9201);
and U9325 (N_9325,N_9249,N_9270);
xor U9326 (N_9326,N_9284,N_9271);
nor U9327 (N_9327,N_9276,N_9210);
nor U9328 (N_9328,N_9223,N_9230);
and U9329 (N_9329,N_9235,N_9253);
xnor U9330 (N_9330,N_9233,N_9208);
nor U9331 (N_9331,N_9274,N_9292);
nand U9332 (N_9332,N_9218,N_9260);
xor U9333 (N_9333,N_9212,N_9257);
xor U9334 (N_9334,N_9296,N_9222);
and U9335 (N_9335,N_9259,N_9240);
and U9336 (N_9336,N_9295,N_9216);
nor U9337 (N_9337,N_9272,N_9215);
nor U9338 (N_9338,N_9229,N_9227);
and U9339 (N_9339,N_9206,N_9236);
nor U9340 (N_9340,N_9281,N_9205);
nand U9341 (N_9341,N_9297,N_9280);
and U9342 (N_9342,N_9239,N_9255);
nor U9343 (N_9343,N_9275,N_9204);
xnor U9344 (N_9344,N_9231,N_9237);
nor U9345 (N_9345,N_9228,N_9298);
xnor U9346 (N_9346,N_9287,N_9225);
xor U9347 (N_9347,N_9251,N_9221);
xor U9348 (N_9348,N_9202,N_9207);
nand U9349 (N_9349,N_9200,N_9262);
or U9350 (N_9350,N_9287,N_9282);
or U9351 (N_9351,N_9235,N_9292);
nor U9352 (N_9352,N_9201,N_9238);
xor U9353 (N_9353,N_9202,N_9232);
and U9354 (N_9354,N_9298,N_9292);
and U9355 (N_9355,N_9229,N_9223);
or U9356 (N_9356,N_9237,N_9201);
and U9357 (N_9357,N_9292,N_9277);
xnor U9358 (N_9358,N_9220,N_9249);
nand U9359 (N_9359,N_9242,N_9210);
nor U9360 (N_9360,N_9260,N_9264);
nand U9361 (N_9361,N_9240,N_9282);
nor U9362 (N_9362,N_9247,N_9248);
xnor U9363 (N_9363,N_9283,N_9297);
or U9364 (N_9364,N_9275,N_9246);
nor U9365 (N_9365,N_9242,N_9204);
nand U9366 (N_9366,N_9226,N_9251);
or U9367 (N_9367,N_9205,N_9268);
xor U9368 (N_9368,N_9260,N_9283);
xnor U9369 (N_9369,N_9265,N_9269);
and U9370 (N_9370,N_9220,N_9228);
nand U9371 (N_9371,N_9221,N_9215);
nand U9372 (N_9372,N_9235,N_9217);
nor U9373 (N_9373,N_9271,N_9269);
and U9374 (N_9374,N_9277,N_9220);
and U9375 (N_9375,N_9252,N_9238);
nor U9376 (N_9376,N_9258,N_9218);
nor U9377 (N_9377,N_9207,N_9249);
or U9378 (N_9378,N_9288,N_9259);
nor U9379 (N_9379,N_9211,N_9224);
nor U9380 (N_9380,N_9263,N_9266);
and U9381 (N_9381,N_9254,N_9296);
nand U9382 (N_9382,N_9206,N_9274);
xor U9383 (N_9383,N_9297,N_9282);
nand U9384 (N_9384,N_9265,N_9214);
or U9385 (N_9385,N_9209,N_9230);
xor U9386 (N_9386,N_9213,N_9221);
xnor U9387 (N_9387,N_9202,N_9209);
nand U9388 (N_9388,N_9299,N_9273);
or U9389 (N_9389,N_9206,N_9286);
or U9390 (N_9390,N_9260,N_9256);
or U9391 (N_9391,N_9283,N_9204);
and U9392 (N_9392,N_9275,N_9251);
or U9393 (N_9393,N_9245,N_9252);
xnor U9394 (N_9394,N_9273,N_9279);
nand U9395 (N_9395,N_9299,N_9211);
nand U9396 (N_9396,N_9215,N_9284);
nand U9397 (N_9397,N_9241,N_9238);
xnor U9398 (N_9398,N_9239,N_9261);
or U9399 (N_9399,N_9282,N_9238);
or U9400 (N_9400,N_9338,N_9343);
nand U9401 (N_9401,N_9378,N_9388);
nand U9402 (N_9402,N_9311,N_9353);
xor U9403 (N_9403,N_9323,N_9382);
and U9404 (N_9404,N_9384,N_9394);
and U9405 (N_9405,N_9308,N_9340);
or U9406 (N_9406,N_9328,N_9393);
nand U9407 (N_9407,N_9321,N_9330);
or U9408 (N_9408,N_9309,N_9376);
nand U9409 (N_9409,N_9359,N_9365);
nand U9410 (N_9410,N_9341,N_9305);
or U9411 (N_9411,N_9337,N_9395);
nand U9412 (N_9412,N_9366,N_9354);
nand U9413 (N_9413,N_9377,N_9368);
xor U9414 (N_9414,N_9398,N_9332);
nand U9415 (N_9415,N_9381,N_9371);
or U9416 (N_9416,N_9344,N_9303);
and U9417 (N_9417,N_9300,N_9333);
nor U9418 (N_9418,N_9383,N_9396);
nand U9419 (N_9419,N_9369,N_9346);
or U9420 (N_9420,N_9315,N_9319);
and U9421 (N_9421,N_9373,N_9392);
xor U9422 (N_9422,N_9345,N_9389);
nor U9423 (N_9423,N_9301,N_9397);
nand U9424 (N_9424,N_9314,N_9307);
or U9425 (N_9425,N_9327,N_9310);
and U9426 (N_9426,N_9342,N_9390);
nor U9427 (N_9427,N_9313,N_9357);
xnor U9428 (N_9428,N_9336,N_9326);
nor U9429 (N_9429,N_9302,N_9374);
nand U9430 (N_9430,N_9386,N_9348);
nor U9431 (N_9431,N_9351,N_9347);
nand U9432 (N_9432,N_9379,N_9391);
nand U9433 (N_9433,N_9329,N_9349);
or U9434 (N_9434,N_9352,N_9339);
xor U9435 (N_9435,N_9316,N_9350);
nand U9436 (N_9436,N_9375,N_9358);
or U9437 (N_9437,N_9362,N_9399);
xor U9438 (N_9438,N_9370,N_9312);
or U9439 (N_9439,N_9331,N_9320);
nand U9440 (N_9440,N_9364,N_9318);
nor U9441 (N_9441,N_9361,N_9385);
xor U9442 (N_9442,N_9363,N_9334);
nand U9443 (N_9443,N_9372,N_9380);
nand U9444 (N_9444,N_9317,N_9325);
nor U9445 (N_9445,N_9306,N_9367);
or U9446 (N_9446,N_9322,N_9356);
or U9447 (N_9447,N_9360,N_9387);
nand U9448 (N_9448,N_9324,N_9304);
nor U9449 (N_9449,N_9355,N_9335);
and U9450 (N_9450,N_9303,N_9399);
nor U9451 (N_9451,N_9391,N_9348);
nor U9452 (N_9452,N_9348,N_9372);
and U9453 (N_9453,N_9363,N_9307);
or U9454 (N_9454,N_9382,N_9380);
xor U9455 (N_9455,N_9380,N_9367);
nor U9456 (N_9456,N_9365,N_9381);
nor U9457 (N_9457,N_9351,N_9307);
and U9458 (N_9458,N_9363,N_9376);
nand U9459 (N_9459,N_9361,N_9362);
nor U9460 (N_9460,N_9320,N_9360);
or U9461 (N_9461,N_9336,N_9341);
xnor U9462 (N_9462,N_9339,N_9396);
xor U9463 (N_9463,N_9360,N_9352);
or U9464 (N_9464,N_9305,N_9397);
or U9465 (N_9465,N_9367,N_9358);
and U9466 (N_9466,N_9391,N_9319);
nand U9467 (N_9467,N_9333,N_9311);
nand U9468 (N_9468,N_9302,N_9300);
nor U9469 (N_9469,N_9315,N_9387);
and U9470 (N_9470,N_9339,N_9328);
or U9471 (N_9471,N_9348,N_9310);
or U9472 (N_9472,N_9346,N_9309);
or U9473 (N_9473,N_9392,N_9364);
and U9474 (N_9474,N_9319,N_9395);
xnor U9475 (N_9475,N_9391,N_9356);
and U9476 (N_9476,N_9386,N_9359);
nor U9477 (N_9477,N_9313,N_9385);
xor U9478 (N_9478,N_9338,N_9363);
nand U9479 (N_9479,N_9363,N_9317);
nand U9480 (N_9480,N_9311,N_9372);
nand U9481 (N_9481,N_9347,N_9307);
and U9482 (N_9482,N_9333,N_9382);
and U9483 (N_9483,N_9326,N_9323);
nor U9484 (N_9484,N_9349,N_9341);
xnor U9485 (N_9485,N_9382,N_9389);
and U9486 (N_9486,N_9376,N_9373);
nand U9487 (N_9487,N_9371,N_9344);
and U9488 (N_9488,N_9334,N_9371);
nand U9489 (N_9489,N_9357,N_9347);
and U9490 (N_9490,N_9345,N_9313);
or U9491 (N_9491,N_9311,N_9391);
nand U9492 (N_9492,N_9364,N_9366);
and U9493 (N_9493,N_9376,N_9365);
or U9494 (N_9494,N_9395,N_9336);
and U9495 (N_9495,N_9376,N_9359);
xnor U9496 (N_9496,N_9372,N_9329);
nor U9497 (N_9497,N_9391,N_9355);
or U9498 (N_9498,N_9323,N_9393);
xnor U9499 (N_9499,N_9371,N_9325);
nand U9500 (N_9500,N_9475,N_9491);
nor U9501 (N_9501,N_9436,N_9468);
nor U9502 (N_9502,N_9490,N_9403);
nand U9503 (N_9503,N_9412,N_9481);
or U9504 (N_9504,N_9414,N_9427);
and U9505 (N_9505,N_9429,N_9477);
and U9506 (N_9506,N_9463,N_9415);
nand U9507 (N_9507,N_9497,N_9401);
or U9508 (N_9508,N_9434,N_9409);
nand U9509 (N_9509,N_9410,N_9443);
and U9510 (N_9510,N_9456,N_9492);
nand U9511 (N_9511,N_9474,N_9454);
or U9512 (N_9512,N_9405,N_9479);
nand U9513 (N_9513,N_9451,N_9417);
or U9514 (N_9514,N_9483,N_9421);
and U9515 (N_9515,N_9440,N_9448);
or U9516 (N_9516,N_9478,N_9420);
nor U9517 (N_9517,N_9496,N_9487);
and U9518 (N_9518,N_9488,N_9430);
and U9519 (N_9519,N_9452,N_9489);
or U9520 (N_9520,N_9499,N_9418);
and U9521 (N_9521,N_9462,N_9447);
nor U9522 (N_9522,N_9466,N_9404);
nor U9523 (N_9523,N_9407,N_9480);
and U9524 (N_9524,N_9449,N_9484);
nand U9525 (N_9525,N_9444,N_9457);
or U9526 (N_9526,N_9485,N_9467);
xor U9527 (N_9527,N_9445,N_9446);
and U9528 (N_9528,N_9433,N_9413);
nor U9529 (N_9529,N_9419,N_9432);
nand U9530 (N_9530,N_9423,N_9460);
and U9531 (N_9531,N_9470,N_9455);
or U9532 (N_9532,N_9476,N_9473);
nand U9533 (N_9533,N_9424,N_9472);
and U9534 (N_9534,N_9425,N_9486);
and U9535 (N_9535,N_9435,N_9422);
xnor U9536 (N_9536,N_9437,N_9453);
nand U9537 (N_9537,N_9469,N_9498);
nand U9538 (N_9538,N_9402,N_9465);
and U9539 (N_9539,N_9442,N_9408);
nor U9540 (N_9540,N_9493,N_9458);
and U9541 (N_9541,N_9464,N_9459);
nand U9542 (N_9542,N_9406,N_9431);
or U9543 (N_9543,N_9439,N_9428);
and U9544 (N_9544,N_9482,N_9441);
and U9545 (N_9545,N_9494,N_9411);
and U9546 (N_9546,N_9495,N_9416);
and U9547 (N_9547,N_9400,N_9471);
or U9548 (N_9548,N_9450,N_9461);
xor U9549 (N_9549,N_9426,N_9438);
and U9550 (N_9550,N_9402,N_9453);
xor U9551 (N_9551,N_9481,N_9444);
nor U9552 (N_9552,N_9437,N_9461);
and U9553 (N_9553,N_9410,N_9468);
nand U9554 (N_9554,N_9465,N_9490);
nor U9555 (N_9555,N_9440,N_9446);
xnor U9556 (N_9556,N_9451,N_9464);
and U9557 (N_9557,N_9435,N_9444);
xor U9558 (N_9558,N_9495,N_9441);
and U9559 (N_9559,N_9491,N_9415);
nor U9560 (N_9560,N_9436,N_9443);
nor U9561 (N_9561,N_9418,N_9420);
xnor U9562 (N_9562,N_9454,N_9480);
xor U9563 (N_9563,N_9454,N_9434);
nand U9564 (N_9564,N_9418,N_9472);
and U9565 (N_9565,N_9455,N_9466);
nand U9566 (N_9566,N_9458,N_9401);
nor U9567 (N_9567,N_9419,N_9489);
xnor U9568 (N_9568,N_9482,N_9424);
nand U9569 (N_9569,N_9452,N_9474);
nor U9570 (N_9570,N_9462,N_9434);
or U9571 (N_9571,N_9449,N_9402);
or U9572 (N_9572,N_9471,N_9481);
xnor U9573 (N_9573,N_9494,N_9461);
and U9574 (N_9574,N_9445,N_9406);
or U9575 (N_9575,N_9425,N_9485);
nand U9576 (N_9576,N_9472,N_9459);
nor U9577 (N_9577,N_9429,N_9421);
nand U9578 (N_9578,N_9467,N_9438);
nand U9579 (N_9579,N_9470,N_9438);
and U9580 (N_9580,N_9420,N_9434);
nand U9581 (N_9581,N_9498,N_9487);
nand U9582 (N_9582,N_9403,N_9462);
or U9583 (N_9583,N_9428,N_9450);
xor U9584 (N_9584,N_9430,N_9462);
or U9585 (N_9585,N_9448,N_9435);
nand U9586 (N_9586,N_9404,N_9463);
or U9587 (N_9587,N_9499,N_9417);
nand U9588 (N_9588,N_9404,N_9413);
nand U9589 (N_9589,N_9427,N_9493);
nor U9590 (N_9590,N_9421,N_9444);
nor U9591 (N_9591,N_9436,N_9461);
nand U9592 (N_9592,N_9485,N_9435);
xor U9593 (N_9593,N_9402,N_9451);
nand U9594 (N_9594,N_9451,N_9449);
and U9595 (N_9595,N_9498,N_9471);
nor U9596 (N_9596,N_9476,N_9458);
nand U9597 (N_9597,N_9408,N_9461);
xnor U9598 (N_9598,N_9419,N_9417);
xnor U9599 (N_9599,N_9479,N_9432);
nor U9600 (N_9600,N_9552,N_9549);
nand U9601 (N_9601,N_9528,N_9564);
or U9602 (N_9602,N_9550,N_9517);
nand U9603 (N_9603,N_9587,N_9567);
nor U9604 (N_9604,N_9503,N_9506);
nor U9605 (N_9605,N_9575,N_9592);
or U9606 (N_9606,N_9509,N_9535);
or U9607 (N_9607,N_9598,N_9581);
or U9608 (N_9608,N_9584,N_9594);
or U9609 (N_9609,N_9515,N_9537);
nand U9610 (N_9610,N_9530,N_9514);
and U9611 (N_9611,N_9541,N_9526);
nor U9612 (N_9612,N_9512,N_9556);
nor U9613 (N_9613,N_9500,N_9570);
and U9614 (N_9614,N_9543,N_9545);
or U9615 (N_9615,N_9501,N_9518);
nor U9616 (N_9616,N_9533,N_9523);
nand U9617 (N_9617,N_9586,N_9544);
nor U9618 (N_9618,N_9516,N_9519);
or U9619 (N_9619,N_9559,N_9572);
nor U9620 (N_9620,N_9502,N_9511);
nand U9621 (N_9621,N_9571,N_9563);
and U9622 (N_9622,N_9580,N_9591);
and U9623 (N_9623,N_9573,N_9577);
xor U9624 (N_9624,N_9558,N_9555);
nor U9625 (N_9625,N_9582,N_9585);
xnor U9626 (N_9626,N_9527,N_9554);
or U9627 (N_9627,N_9561,N_9557);
nor U9628 (N_9628,N_9569,N_9599);
nand U9629 (N_9629,N_9551,N_9505);
xnor U9630 (N_9630,N_9560,N_9529);
nand U9631 (N_9631,N_9588,N_9524);
and U9632 (N_9632,N_9525,N_9520);
nor U9633 (N_9633,N_9548,N_9595);
nand U9634 (N_9634,N_9540,N_9596);
nor U9635 (N_9635,N_9568,N_9583);
xnor U9636 (N_9636,N_9553,N_9576);
or U9637 (N_9637,N_9532,N_9566);
and U9638 (N_9638,N_9531,N_9547);
xor U9639 (N_9639,N_9590,N_9539);
xor U9640 (N_9640,N_9597,N_9508);
nand U9641 (N_9641,N_9565,N_9579);
or U9642 (N_9642,N_9546,N_9589);
or U9643 (N_9643,N_9574,N_9578);
nor U9644 (N_9644,N_9534,N_9507);
or U9645 (N_9645,N_9521,N_9510);
nor U9646 (N_9646,N_9504,N_9522);
or U9647 (N_9647,N_9513,N_9538);
nand U9648 (N_9648,N_9536,N_9593);
or U9649 (N_9649,N_9562,N_9542);
or U9650 (N_9650,N_9522,N_9581);
xnor U9651 (N_9651,N_9555,N_9562);
nand U9652 (N_9652,N_9566,N_9547);
or U9653 (N_9653,N_9585,N_9566);
or U9654 (N_9654,N_9598,N_9516);
or U9655 (N_9655,N_9506,N_9530);
and U9656 (N_9656,N_9538,N_9576);
nand U9657 (N_9657,N_9548,N_9566);
nor U9658 (N_9658,N_9589,N_9578);
xor U9659 (N_9659,N_9535,N_9502);
nor U9660 (N_9660,N_9567,N_9554);
nand U9661 (N_9661,N_9583,N_9553);
or U9662 (N_9662,N_9501,N_9581);
nand U9663 (N_9663,N_9573,N_9558);
xnor U9664 (N_9664,N_9562,N_9578);
or U9665 (N_9665,N_9518,N_9522);
nand U9666 (N_9666,N_9588,N_9536);
or U9667 (N_9667,N_9519,N_9538);
nor U9668 (N_9668,N_9545,N_9583);
nand U9669 (N_9669,N_9512,N_9587);
nand U9670 (N_9670,N_9584,N_9589);
xor U9671 (N_9671,N_9567,N_9543);
and U9672 (N_9672,N_9573,N_9549);
nand U9673 (N_9673,N_9540,N_9595);
nor U9674 (N_9674,N_9598,N_9565);
nand U9675 (N_9675,N_9502,N_9591);
nand U9676 (N_9676,N_9504,N_9511);
and U9677 (N_9677,N_9518,N_9507);
and U9678 (N_9678,N_9548,N_9525);
and U9679 (N_9679,N_9509,N_9543);
nor U9680 (N_9680,N_9546,N_9569);
nor U9681 (N_9681,N_9523,N_9598);
xor U9682 (N_9682,N_9586,N_9532);
or U9683 (N_9683,N_9520,N_9582);
and U9684 (N_9684,N_9530,N_9531);
or U9685 (N_9685,N_9598,N_9564);
and U9686 (N_9686,N_9589,N_9516);
and U9687 (N_9687,N_9591,N_9557);
xor U9688 (N_9688,N_9509,N_9525);
xnor U9689 (N_9689,N_9518,N_9588);
and U9690 (N_9690,N_9526,N_9593);
xnor U9691 (N_9691,N_9531,N_9579);
and U9692 (N_9692,N_9521,N_9518);
nand U9693 (N_9693,N_9508,N_9561);
xnor U9694 (N_9694,N_9554,N_9556);
or U9695 (N_9695,N_9550,N_9501);
or U9696 (N_9696,N_9562,N_9588);
xnor U9697 (N_9697,N_9504,N_9565);
xor U9698 (N_9698,N_9596,N_9517);
xor U9699 (N_9699,N_9564,N_9584);
xor U9700 (N_9700,N_9613,N_9623);
xnor U9701 (N_9701,N_9674,N_9669);
nand U9702 (N_9702,N_9670,N_9663);
nand U9703 (N_9703,N_9671,N_9626);
nor U9704 (N_9704,N_9644,N_9682);
nor U9705 (N_9705,N_9685,N_9680);
nand U9706 (N_9706,N_9611,N_9637);
and U9707 (N_9707,N_9692,N_9625);
or U9708 (N_9708,N_9636,N_9668);
and U9709 (N_9709,N_9694,N_9699);
and U9710 (N_9710,N_9686,N_9624);
or U9711 (N_9711,N_9643,N_9654);
or U9712 (N_9712,N_9675,N_9631);
or U9713 (N_9713,N_9696,N_9657);
nand U9714 (N_9714,N_9653,N_9608);
xor U9715 (N_9715,N_9642,N_9627);
nor U9716 (N_9716,N_9618,N_9677);
xor U9717 (N_9717,N_9603,N_9635);
or U9718 (N_9718,N_9662,N_9672);
xnor U9719 (N_9719,N_9676,N_9681);
and U9720 (N_9720,N_9678,N_9610);
nand U9721 (N_9721,N_9684,N_9665);
or U9722 (N_9722,N_9695,N_9649);
nor U9723 (N_9723,N_9691,N_9673);
or U9724 (N_9724,N_9698,N_9658);
xor U9725 (N_9725,N_9688,N_9619);
nand U9726 (N_9726,N_9606,N_9632);
nand U9727 (N_9727,N_9607,N_9652);
or U9728 (N_9728,N_9634,N_9655);
or U9729 (N_9729,N_9612,N_9664);
or U9730 (N_9730,N_9689,N_9604);
xnor U9731 (N_9731,N_9640,N_9617);
and U9732 (N_9732,N_9600,N_9647);
nor U9733 (N_9733,N_9621,N_9622);
and U9734 (N_9734,N_9667,N_9620);
or U9735 (N_9735,N_9650,N_9629);
or U9736 (N_9736,N_9697,N_9648);
or U9737 (N_9737,N_9616,N_9638);
nand U9738 (N_9738,N_9630,N_9614);
xor U9739 (N_9739,N_9639,N_9633);
xnor U9740 (N_9740,N_9646,N_9659);
and U9741 (N_9741,N_9628,N_9690);
and U9742 (N_9742,N_9601,N_9602);
and U9743 (N_9743,N_9693,N_9660);
or U9744 (N_9744,N_9687,N_9656);
or U9745 (N_9745,N_9651,N_9641);
or U9746 (N_9746,N_9683,N_9605);
xor U9747 (N_9747,N_9661,N_9615);
or U9748 (N_9748,N_9609,N_9645);
or U9749 (N_9749,N_9666,N_9679);
or U9750 (N_9750,N_9638,N_9664);
xnor U9751 (N_9751,N_9632,N_9687);
nand U9752 (N_9752,N_9611,N_9679);
nor U9753 (N_9753,N_9687,N_9616);
nand U9754 (N_9754,N_9698,N_9610);
xor U9755 (N_9755,N_9670,N_9628);
nor U9756 (N_9756,N_9614,N_9692);
or U9757 (N_9757,N_9648,N_9663);
nor U9758 (N_9758,N_9647,N_9639);
and U9759 (N_9759,N_9669,N_9611);
or U9760 (N_9760,N_9666,N_9663);
or U9761 (N_9761,N_9674,N_9686);
nand U9762 (N_9762,N_9678,N_9605);
nand U9763 (N_9763,N_9687,N_9603);
nor U9764 (N_9764,N_9677,N_9608);
or U9765 (N_9765,N_9693,N_9612);
nor U9766 (N_9766,N_9681,N_9641);
and U9767 (N_9767,N_9615,N_9664);
xnor U9768 (N_9768,N_9600,N_9641);
nand U9769 (N_9769,N_9620,N_9648);
xor U9770 (N_9770,N_9691,N_9648);
and U9771 (N_9771,N_9630,N_9682);
or U9772 (N_9772,N_9676,N_9680);
nand U9773 (N_9773,N_9607,N_9699);
nor U9774 (N_9774,N_9631,N_9669);
nand U9775 (N_9775,N_9693,N_9602);
nor U9776 (N_9776,N_9600,N_9608);
or U9777 (N_9777,N_9602,N_9657);
nand U9778 (N_9778,N_9608,N_9695);
nor U9779 (N_9779,N_9651,N_9674);
and U9780 (N_9780,N_9667,N_9674);
or U9781 (N_9781,N_9666,N_9635);
and U9782 (N_9782,N_9627,N_9658);
xnor U9783 (N_9783,N_9670,N_9679);
xor U9784 (N_9784,N_9622,N_9692);
nand U9785 (N_9785,N_9658,N_9654);
nor U9786 (N_9786,N_9636,N_9631);
nand U9787 (N_9787,N_9649,N_9622);
or U9788 (N_9788,N_9654,N_9681);
or U9789 (N_9789,N_9681,N_9629);
nor U9790 (N_9790,N_9640,N_9695);
and U9791 (N_9791,N_9632,N_9613);
nor U9792 (N_9792,N_9665,N_9612);
or U9793 (N_9793,N_9648,N_9684);
xnor U9794 (N_9794,N_9649,N_9672);
or U9795 (N_9795,N_9687,N_9679);
and U9796 (N_9796,N_9681,N_9696);
xor U9797 (N_9797,N_9631,N_9630);
or U9798 (N_9798,N_9634,N_9624);
and U9799 (N_9799,N_9646,N_9650);
or U9800 (N_9800,N_9717,N_9798);
xor U9801 (N_9801,N_9782,N_9710);
and U9802 (N_9802,N_9759,N_9788);
or U9803 (N_9803,N_9775,N_9704);
or U9804 (N_9804,N_9757,N_9713);
and U9805 (N_9805,N_9737,N_9747);
nand U9806 (N_9806,N_9744,N_9745);
xnor U9807 (N_9807,N_9738,N_9700);
nand U9808 (N_9808,N_9731,N_9705);
nand U9809 (N_9809,N_9766,N_9721);
nand U9810 (N_9810,N_9702,N_9791);
and U9811 (N_9811,N_9781,N_9784);
or U9812 (N_9812,N_9715,N_9786);
xnor U9813 (N_9813,N_9720,N_9701);
nand U9814 (N_9814,N_9750,N_9742);
or U9815 (N_9815,N_9796,N_9764);
and U9816 (N_9816,N_9780,N_9792);
xor U9817 (N_9817,N_9754,N_9778);
nand U9818 (N_9818,N_9730,N_9707);
nor U9819 (N_9819,N_9740,N_9732);
nand U9820 (N_9820,N_9746,N_9712);
nor U9821 (N_9821,N_9714,N_9739);
or U9822 (N_9822,N_9777,N_9709);
and U9823 (N_9823,N_9785,N_9733);
nand U9824 (N_9824,N_9793,N_9765);
and U9825 (N_9825,N_9756,N_9752);
nand U9826 (N_9826,N_9751,N_9728);
nor U9827 (N_9827,N_9723,N_9735);
or U9828 (N_9828,N_9755,N_9767);
nor U9829 (N_9829,N_9789,N_9724);
and U9830 (N_9830,N_9726,N_9719);
xnor U9831 (N_9831,N_9795,N_9774);
nor U9832 (N_9832,N_9768,N_9736);
xnor U9833 (N_9833,N_9779,N_9727);
xor U9834 (N_9834,N_9771,N_9776);
or U9835 (N_9835,N_9769,N_9770);
nor U9836 (N_9836,N_9753,N_9773);
nor U9837 (N_9837,N_9787,N_9783);
and U9838 (N_9838,N_9790,N_9743);
nor U9839 (N_9839,N_9741,N_9729);
or U9840 (N_9840,N_9722,N_9760);
nor U9841 (N_9841,N_9762,N_9772);
nor U9842 (N_9842,N_9797,N_9708);
xor U9843 (N_9843,N_9794,N_9799);
nor U9844 (N_9844,N_9716,N_9763);
xor U9845 (N_9845,N_9718,N_9748);
or U9846 (N_9846,N_9703,N_9758);
nor U9847 (N_9847,N_9761,N_9749);
nor U9848 (N_9848,N_9711,N_9725);
nor U9849 (N_9849,N_9734,N_9706);
xor U9850 (N_9850,N_9714,N_9722);
xor U9851 (N_9851,N_9712,N_9763);
nand U9852 (N_9852,N_9717,N_9780);
and U9853 (N_9853,N_9788,N_9799);
xor U9854 (N_9854,N_9765,N_9701);
xnor U9855 (N_9855,N_9709,N_9768);
nor U9856 (N_9856,N_9746,N_9733);
and U9857 (N_9857,N_9724,N_9790);
xnor U9858 (N_9858,N_9770,N_9754);
nand U9859 (N_9859,N_9759,N_9783);
nor U9860 (N_9860,N_9795,N_9765);
nand U9861 (N_9861,N_9781,N_9794);
nand U9862 (N_9862,N_9757,N_9752);
nor U9863 (N_9863,N_9774,N_9779);
or U9864 (N_9864,N_9737,N_9766);
and U9865 (N_9865,N_9774,N_9750);
nand U9866 (N_9866,N_9789,N_9765);
nor U9867 (N_9867,N_9792,N_9747);
and U9868 (N_9868,N_9793,N_9731);
xor U9869 (N_9869,N_9788,N_9746);
nand U9870 (N_9870,N_9742,N_9727);
or U9871 (N_9871,N_9737,N_9792);
nand U9872 (N_9872,N_9719,N_9767);
nor U9873 (N_9873,N_9706,N_9745);
xor U9874 (N_9874,N_9729,N_9778);
or U9875 (N_9875,N_9716,N_9728);
or U9876 (N_9876,N_9792,N_9736);
nand U9877 (N_9877,N_9744,N_9739);
and U9878 (N_9878,N_9701,N_9741);
nand U9879 (N_9879,N_9746,N_9729);
xnor U9880 (N_9880,N_9724,N_9738);
nand U9881 (N_9881,N_9712,N_9731);
and U9882 (N_9882,N_9712,N_9792);
and U9883 (N_9883,N_9780,N_9740);
nor U9884 (N_9884,N_9755,N_9746);
or U9885 (N_9885,N_9796,N_9759);
nand U9886 (N_9886,N_9721,N_9790);
xor U9887 (N_9887,N_9775,N_9768);
nand U9888 (N_9888,N_9775,N_9777);
and U9889 (N_9889,N_9761,N_9726);
or U9890 (N_9890,N_9756,N_9702);
and U9891 (N_9891,N_9748,N_9762);
xnor U9892 (N_9892,N_9729,N_9771);
nor U9893 (N_9893,N_9765,N_9703);
nand U9894 (N_9894,N_9738,N_9718);
xnor U9895 (N_9895,N_9722,N_9710);
or U9896 (N_9896,N_9747,N_9715);
nand U9897 (N_9897,N_9730,N_9737);
or U9898 (N_9898,N_9792,N_9796);
nand U9899 (N_9899,N_9796,N_9747);
nor U9900 (N_9900,N_9833,N_9817);
and U9901 (N_9901,N_9802,N_9842);
or U9902 (N_9902,N_9857,N_9886);
nand U9903 (N_9903,N_9828,N_9847);
and U9904 (N_9904,N_9804,N_9830);
and U9905 (N_9905,N_9848,N_9890);
or U9906 (N_9906,N_9803,N_9839);
nor U9907 (N_9907,N_9815,N_9859);
xnor U9908 (N_9908,N_9888,N_9891);
xnor U9909 (N_9909,N_9852,N_9869);
nand U9910 (N_9910,N_9867,N_9827);
nand U9911 (N_9911,N_9816,N_9898);
nor U9912 (N_9912,N_9810,N_9863);
and U9913 (N_9913,N_9820,N_9872);
and U9914 (N_9914,N_9861,N_9811);
or U9915 (N_9915,N_9885,N_9894);
or U9916 (N_9916,N_9892,N_9813);
or U9917 (N_9917,N_9812,N_9870);
nand U9918 (N_9918,N_9821,N_9868);
nand U9919 (N_9919,N_9807,N_9809);
nor U9920 (N_9920,N_9831,N_9873);
nor U9921 (N_9921,N_9855,N_9871);
or U9922 (N_9922,N_9805,N_9823);
xnor U9923 (N_9923,N_9806,N_9824);
and U9924 (N_9924,N_9856,N_9858);
and U9925 (N_9925,N_9834,N_9838);
or U9926 (N_9926,N_9829,N_9846);
and U9927 (N_9927,N_9879,N_9819);
or U9928 (N_9928,N_9878,N_9866);
and U9929 (N_9929,N_9808,N_9880);
nand U9930 (N_9930,N_9832,N_9893);
and U9931 (N_9931,N_9825,N_9889);
or U9932 (N_9932,N_9818,N_9895);
and U9933 (N_9933,N_9853,N_9874);
nor U9934 (N_9934,N_9884,N_9841);
and U9935 (N_9935,N_9896,N_9840);
or U9936 (N_9936,N_9883,N_9887);
and U9937 (N_9937,N_9822,N_9865);
nand U9938 (N_9938,N_9835,N_9875);
xnor U9939 (N_9939,N_9897,N_9843);
nand U9940 (N_9940,N_9862,N_9854);
or U9941 (N_9941,N_9851,N_9881);
xor U9942 (N_9942,N_9800,N_9836);
nor U9943 (N_9943,N_9882,N_9850);
nand U9944 (N_9944,N_9864,N_9845);
nand U9945 (N_9945,N_9801,N_9899);
or U9946 (N_9946,N_9877,N_9860);
nor U9947 (N_9947,N_9844,N_9849);
nor U9948 (N_9948,N_9876,N_9814);
nand U9949 (N_9949,N_9826,N_9837);
and U9950 (N_9950,N_9873,N_9805);
xnor U9951 (N_9951,N_9833,N_9829);
nor U9952 (N_9952,N_9882,N_9886);
xor U9953 (N_9953,N_9807,N_9816);
or U9954 (N_9954,N_9861,N_9802);
nor U9955 (N_9955,N_9824,N_9848);
nand U9956 (N_9956,N_9856,N_9881);
xor U9957 (N_9957,N_9843,N_9842);
and U9958 (N_9958,N_9855,N_9887);
xnor U9959 (N_9959,N_9831,N_9828);
xnor U9960 (N_9960,N_9866,N_9846);
nor U9961 (N_9961,N_9841,N_9827);
and U9962 (N_9962,N_9878,N_9827);
and U9963 (N_9963,N_9855,N_9853);
xor U9964 (N_9964,N_9858,N_9860);
xnor U9965 (N_9965,N_9858,N_9850);
xor U9966 (N_9966,N_9835,N_9800);
and U9967 (N_9967,N_9849,N_9848);
xnor U9968 (N_9968,N_9853,N_9835);
nand U9969 (N_9969,N_9846,N_9817);
nor U9970 (N_9970,N_9820,N_9849);
nand U9971 (N_9971,N_9894,N_9820);
nand U9972 (N_9972,N_9803,N_9809);
nor U9973 (N_9973,N_9831,N_9849);
and U9974 (N_9974,N_9846,N_9850);
and U9975 (N_9975,N_9898,N_9815);
and U9976 (N_9976,N_9825,N_9897);
nor U9977 (N_9977,N_9895,N_9880);
nor U9978 (N_9978,N_9896,N_9845);
and U9979 (N_9979,N_9882,N_9884);
xnor U9980 (N_9980,N_9856,N_9885);
and U9981 (N_9981,N_9892,N_9826);
or U9982 (N_9982,N_9861,N_9847);
nand U9983 (N_9983,N_9853,N_9895);
nand U9984 (N_9984,N_9802,N_9845);
xor U9985 (N_9985,N_9821,N_9851);
xor U9986 (N_9986,N_9850,N_9809);
nand U9987 (N_9987,N_9892,N_9881);
nor U9988 (N_9988,N_9892,N_9873);
nor U9989 (N_9989,N_9811,N_9857);
and U9990 (N_9990,N_9862,N_9875);
nand U9991 (N_9991,N_9813,N_9893);
or U9992 (N_9992,N_9874,N_9823);
xor U9993 (N_9993,N_9831,N_9800);
xor U9994 (N_9994,N_9866,N_9816);
xnor U9995 (N_9995,N_9815,N_9855);
nor U9996 (N_9996,N_9859,N_9820);
and U9997 (N_9997,N_9860,N_9897);
xnor U9998 (N_9998,N_9868,N_9891);
and U9999 (N_9999,N_9865,N_9869);
nor UO_0 (O_0,N_9991,N_9923);
xor UO_1 (O_1,N_9927,N_9929);
or UO_2 (O_2,N_9986,N_9901);
nor UO_3 (O_3,N_9950,N_9914);
nor UO_4 (O_4,N_9984,N_9946);
or UO_5 (O_5,N_9900,N_9919);
xnor UO_6 (O_6,N_9953,N_9939);
or UO_7 (O_7,N_9990,N_9962);
xor UO_8 (O_8,N_9957,N_9998);
and UO_9 (O_9,N_9935,N_9949);
xor UO_10 (O_10,N_9997,N_9976);
and UO_11 (O_11,N_9910,N_9954);
nand UO_12 (O_12,N_9928,N_9941);
and UO_13 (O_13,N_9909,N_9952);
xnor UO_14 (O_14,N_9934,N_9922);
and UO_15 (O_15,N_9958,N_9959);
nand UO_16 (O_16,N_9982,N_9972);
nor UO_17 (O_17,N_9921,N_9996);
xnor UO_18 (O_18,N_9993,N_9969);
or UO_19 (O_19,N_9947,N_9999);
nor UO_20 (O_20,N_9963,N_9912);
or UO_21 (O_21,N_9924,N_9979);
and UO_22 (O_22,N_9989,N_9964);
and UO_23 (O_23,N_9978,N_9992);
xnor UO_24 (O_24,N_9933,N_9937);
xor UO_25 (O_25,N_9907,N_9971);
nand UO_26 (O_26,N_9983,N_9913);
and UO_27 (O_27,N_9938,N_9926);
or UO_28 (O_28,N_9966,N_9987);
or UO_29 (O_29,N_9968,N_9915);
nand UO_30 (O_30,N_9905,N_9961);
and UO_31 (O_31,N_9951,N_9940);
and UO_32 (O_32,N_9931,N_9918);
and UO_33 (O_33,N_9973,N_9904);
or UO_34 (O_34,N_9960,N_9988);
nor UO_35 (O_35,N_9943,N_9902);
xnor UO_36 (O_36,N_9977,N_9967);
and UO_37 (O_37,N_9911,N_9916);
and UO_38 (O_38,N_9980,N_9936);
xor UO_39 (O_39,N_9925,N_9948);
xnor UO_40 (O_40,N_9903,N_9995);
xor UO_41 (O_41,N_9906,N_9975);
and UO_42 (O_42,N_9945,N_9994);
or UO_43 (O_43,N_9956,N_9955);
nand UO_44 (O_44,N_9985,N_9917);
nor UO_45 (O_45,N_9908,N_9965);
nor UO_46 (O_46,N_9970,N_9920);
xnor UO_47 (O_47,N_9932,N_9930);
nand UO_48 (O_48,N_9974,N_9942);
nor UO_49 (O_49,N_9944,N_9981);
and UO_50 (O_50,N_9939,N_9969);
and UO_51 (O_51,N_9939,N_9951);
or UO_52 (O_52,N_9940,N_9931);
or UO_53 (O_53,N_9940,N_9977);
or UO_54 (O_54,N_9957,N_9944);
nor UO_55 (O_55,N_9991,N_9992);
xor UO_56 (O_56,N_9992,N_9997);
xnor UO_57 (O_57,N_9948,N_9937);
xnor UO_58 (O_58,N_9934,N_9907);
xor UO_59 (O_59,N_9937,N_9913);
nor UO_60 (O_60,N_9905,N_9984);
or UO_61 (O_61,N_9968,N_9964);
nand UO_62 (O_62,N_9916,N_9941);
nor UO_63 (O_63,N_9949,N_9954);
nor UO_64 (O_64,N_9928,N_9943);
nor UO_65 (O_65,N_9936,N_9949);
nand UO_66 (O_66,N_9900,N_9967);
and UO_67 (O_67,N_9955,N_9962);
xor UO_68 (O_68,N_9965,N_9938);
nand UO_69 (O_69,N_9909,N_9939);
nor UO_70 (O_70,N_9957,N_9901);
nand UO_71 (O_71,N_9967,N_9972);
and UO_72 (O_72,N_9953,N_9964);
or UO_73 (O_73,N_9916,N_9963);
xnor UO_74 (O_74,N_9904,N_9960);
nand UO_75 (O_75,N_9975,N_9944);
nand UO_76 (O_76,N_9932,N_9928);
and UO_77 (O_77,N_9948,N_9904);
and UO_78 (O_78,N_9998,N_9937);
nand UO_79 (O_79,N_9962,N_9984);
xor UO_80 (O_80,N_9940,N_9923);
nand UO_81 (O_81,N_9973,N_9967);
xor UO_82 (O_82,N_9939,N_9972);
nand UO_83 (O_83,N_9947,N_9960);
nor UO_84 (O_84,N_9977,N_9987);
xor UO_85 (O_85,N_9940,N_9970);
or UO_86 (O_86,N_9924,N_9965);
nand UO_87 (O_87,N_9924,N_9962);
and UO_88 (O_88,N_9925,N_9961);
xor UO_89 (O_89,N_9934,N_9944);
and UO_90 (O_90,N_9995,N_9939);
nand UO_91 (O_91,N_9958,N_9976);
xnor UO_92 (O_92,N_9990,N_9995);
or UO_93 (O_93,N_9957,N_9913);
nor UO_94 (O_94,N_9925,N_9926);
nand UO_95 (O_95,N_9991,N_9983);
xnor UO_96 (O_96,N_9959,N_9989);
or UO_97 (O_97,N_9927,N_9925);
or UO_98 (O_98,N_9986,N_9979);
or UO_99 (O_99,N_9954,N_9952);
and UO_100 (O_100,N_9958,N_9987);
nor UO_101 (O_101,N_9961,N_9986);
xor UO_102 (O_102,N_9935,N_9962);
nand UO_103 (O_103,N_9961,N_9940);
and UO_104 (O_104,N_9933,N_9999);
nor UO_105 (O_105,N_9953,N_9947);
nand UO_106 (O_106,N_9904,N_9949);
and UO_107 (O_107,N_9905,N_9950);
xnor UO_108 (O_108,N_9911,N_9910);
nor UO_109 (O_109,N_9973,N_9970);
nor UO_110 (O_110,N_9932,N_9913);
nor UO_111 (O_111,N_9974,N_9941);
nand UO_112 (O_112,N_9996,N_9936);
nand UO_113 (O_113,N_9938,N_9909);
nor UO_114 (O_114,N_9986,N_9910);
and UO_115 (O_115,N_9991,N_9942);
nand UO_116 (O_116,N_9993,N_9926);
xor UO_117 (O_117,N_9990,N_9982);
nor UO_118 (O_118,N_9997,N_9963);
nand UO_119 (O_119,N_9983,N_9953);
nor UO_120 (O_120,N_9900,N_9944);
nor UO_121 (O_121,N_9955,N_9977);
xor UO_122 (O_122,N_9970,N_9994);
and UO_123 (O_123,N_9957,N_9911);
nand UO_124 (O_124,N_9985,N_9993);
and UO_125 (O_125,N_9935,N_9938);
nand UO_126 (O_126,N_9994,N_9941);
xnor UO_127 (O_127,N_9939,N_9992);
and UO_128 (O_128,N_9978,N_9962);
and UO_129 (O_129,N_9933,N_9974);
xnor UO_130 (O_130,N_9948,N_9934);
nor UO_131 (O_131,N_9935,N_9901);
xor UO_132 (O_132,N_9997,N_9964);
xor UO_133 (O_133,N_9905,N_9978);
and UO_134 (O_134,N_9980,N_9934);
xor UO_135 (O_135,N_9989,N_9970);
and UO_136 (O_136,N_9993,N_9923);
xor UO_137 (O_137,N_9940,N_9929);
nand UO_138 (O_138,N_9955,N_9912);
or UO_139 (O_139,N_9982,N_9959);
or UO_140 (O_140,N_9934,N_9988);
and UO_141 (O_141,N_9973,N_9964);
nor UO_142 (O_142,N_9945,N_9934);
xor UO_143 (O_143,N_9952,N_9985);
xnor UO_144 (O_144,N_9996,N_9984);
nor UO_145 (O_145,N_9966,N_9968);
and UO_146 (O_146,N_9980,N_9923);
or UO_147 (O_147,N_9944,N_9903);
nor UO_148 (O_148,N_9927,N_9975);
nand UO_149 (O_149,N_9951,N_9932);
or UO_150 (O_150,N_9999,N_9907);
xnor UO_151 (O_151,N_9926,N_9952);
nand UO_152 (O_152,N_9945,N_9959);
nor UO_153 (O_153,N_9996,N_9978);
or UO_154 (O_154,N_9926,N_9931);
and UO_155 (O_155,N_9944,N_9987);
and UO_156 (O_156,N_9983,N_9924);
or UO_157 (O_157,N_9994,N_9906);
and UO_158 (O_158,N_9975,N_9952);
or UO_159 (O_159,N_9996,N_9927);
and UO_160 (O_160,N_9970,N_9969);
nand UO_161 (O_161,N_9913,N_9904);
and UO_162 (O_162,N_9957,N_9993);
nand UO_163 (O_163,N_9986,N_9903);
or UO_164 (O_164,N_9984,N_9916);
nand UO_165 (O_165,N_9922,N_9903);
and UO_166 (O_166,N_9998,N_9972);
and UO_167 (O_167,N_9984,N_9951);
nor UO_168 (O_168,N_9919,N_9932);
and UO_169 (O_169,N_9918,N_9906);
nand UO_170 (O_170,N_9999,N_9910);
nor UO_171 (O_171,N_9925,N_9933);
and UO_172 (O_172,N_9928,N_9955);
xnor UO_173 (O_173,N_9926,N_9964);
nor UO_174 (O_174,N_9936,N_9937);
xnor UO_175 (O_175,N_9971,N_9942);
nand UO_176 (O_176,N_9995,N_9919);
and UO_177 (O_177,N_9937,N_9906);
and UO_178 (O_178,N_9927,N_9918);
and UO_179 (O_179,N_9957,N_9966);
or UO_180 (O_180,N_9941,N_9981);
nand UO_181 (O_181,N_9918,N_9954);
nand UO_182 (O_182,N_9936,N_9919);
and UO_183 (O_183,N_9994,N_9976);
xor UO_184 (O_184,N_9911,N_9931);
nor UO_185 (O_185,N_9936,N_9931);
nand UO_186 (O_186,N_9936,N_9933);
nand UO_187 (O_187,N_9946,N_9973);
and UO_188 (O_188,N_9931,N_9903);
or UO_189 (O_189,N_9936,N_9942);
nand UO_190 (O_190,N_9944,N_9995);
and UO_191 (O_191,N_9955,N_9999);
or UO_192 (O_192,N_9952,N_9905);
xor UO_193 (O_193,N_9906,N_9976);
xnor UO_194 (O_194,N_9936,N_9911);
nand UO_195 (O_195,N_9961,N_9976);
nand UO_196 (O_196,N_9921,N_9934);
nand UO_197 (O_197,N_9986,N_9926);
or UO_198 (O_198,N_9953,N_9913);
nor UO_199 (O_199,N_9938,N_9902);
nand UO_200 (O_200,N_9969,N_9935);
nor UO_201 (O_201,N_9960,N_9967);
xnor UO_202 (O_202,N_9994,N_9986);
nor UO_203 (O_203,N_9927,N_9945);
and UO_204 (O_204,N_9949,N_9966);
or UO_205 (O_205,N_9983,N_9930);
xor UO_206 (O_206,N_9931,N_9965);
nor UO_207 (O_207,N_9944,N_9961);
xor UO_208 (O_208,N_9938,N_9943);
xnor UO_209 (O_209,N_9929,N_9990);
or UO_210 (O_210,N_9911,N_9986);
or UO_211 (O_211,N_9952,N_9942);
and UO_212 (O_212,N_9938,N_9951);
and UO_213 (O_213,N_9941,N_9985);
nor UO_214 (O_214,N_9952,N_9981);
and UO_215 (O_215,N_9947,N_9919);
and UO_216 (O_216,N_9991,N_9957);
nor UO_217 (O_217,N_9901,N_9996);
xnor UO_218 (O_218,N_9910,N_9964);
nand UO_219 (O_219,N_9985,N_9971);
or UO_220 (O_220,N_9958,N_9926);
nand UO_221 (O_221,N_9957,N_9987);
or UO_222 (O_222,N_9982,N_9943);
nand UO_223 (O_223,N_9994,N_9958);
or UO_224 (O_224,N_9960,N_9934);
nor UO_225 (O_225,N_9956,N_9932);
and UO_226 (O_226,N_9966,N_9974);
xnor UO_227 (O_227,N_9957,N_9917);
nor UO_228 (O_228,N_9904,N_9956);
or UO_229 (O_229,N_9948,N_9969);
nor UO_230 (O_230,N_9936,N_9916);
xnor UO_231 (O_231,N_9980,N_9948);
nor UO_232 (O_232,N_9952,N_9949);
nand UO_233 (O_233,N_9977,N_9908);
xor UO_234 (O_234,N_9965,N_9935);
or UO_235 (O_235,N_9956,N_9977);
or UO_236 (O_236,N_9944,N_9955);
xnor UO_237 (O_237,N_9991,N_9906);
and UO_238 (O_238,N_9986,N_9925);
xnor UO_239 (O_239,N_9928,N_9987);
and UO_240 (O_240,N_9963,N_9908);
nand UO_241 (O_241,N_9969,N_9958);
nand UO_242 (O_242,N_9963,N_9917);
nor UO_243 (O_243,N_9996,N_9918);
or UO_244 (O_244,N_9912,N_9932);
or UO_245 (O_245,N_9946,N_9995);
nand UO_246 (O_246,N_9969,N_9959);
nand UO_247 (O_247,N_9951,N_9952);
nor UO_248 (O_248,N_9990,N_9976);
or UO_249 (O_249,N_9944,N_9959);
nand UO_250 (O_250,N_9967,N_9992);
nand UO_251 (O_251,N_9974,N_9961);
nor UO_252 (O_252,N_9961,N_9957);
or UO_253 (O_253,N_9952,N_9919);
or UO_254 (O_254,N_9921,N_9915);
and UO_255 (O_255,N_9953,N_9928);
nor UO_256 (O_256,N_9946,N_9912);
xor UO_257 (O_257,N_9952,N_9928);
and UO_258 (O_258,N_9942,N_9988);
and UO_259 (O_259,N_9995,N_9996);
and UO_260 (O_260,N_9936,N_9966);
xnor UO_261 (O_261,N_9992,N_9945);
nor UO_262 (O_262,N_9915,N_9938);
nor UO_263 (O_263,N_9936,N_9953);
xnor UO_264 (O_264,N_9964,N_9999);
xor UO_265 (O_265,N_9946,N_9958);
and UO_266 (O_266,N_9930,N_9967);
or UO_267 (O_267,N_9970,N_9952);
and UO_268 (O_268,N_9989,N_9917);
xnor UO_269 (O_269,N_9945,N_9953);
nor UO_270 (O_270,N_9918,N_9963);
nand UO_271 (O_271,N_9912,N_9969);
and UO_272 (O_272,N_9959,N_9968);
nand UO_273 (O_273,N_9987,N_9914);
nor UO_274 (O_274,N_9938,N_9903);
nand UO_275 (O_275,N_9983,N_9962);
and UO_276 (O_276,N_9941,N_9977);
nand UO_277 (O_277,N_9922,N_9989);
or UO_278 (O_278,N_9993,N_9904);
nor UO_279 (O_279,N_9933,N_9914);
and UO_280 (O_280,N_9958,N_9942);
or UO_281 (O_281,N_9988,N_9950);
or UO_282 (O_282,N_9914,N_9964);
nand UO_283 (O_283,N_9981,N_9990);
or UO_284 (O_284,N_9966,N_9915);
or UO_285 (O_285,N_9922,N_9927);
nand UO_286 (O_286,N_9960,N_9982);
nand UO_287 (O_287,N_9996,N_9911);
and UO_288 (O_288,N_9929,N_9908);
xor UO_289 (O_289,N_9969,N_9926);
and UO_290 (O_290,N_9988,N_9998);
and UO_291 (O_291,N_9999,N_9992);
nor UO_292 (O_292,N_9926,N_9992);
or UO_293 (O_293,N_9909,N_9923);
and UO_294 (O_294,N_9938,N_9972);
xnor UO_295 (O_295,N_9927,N_9919);
or UO_296 (O_296,N_9922,N_9916);
xor UO_297 (O_297,N_9940,N_9958);
and UO_298 (O_298,N_9962,N_9941);
nor UO_299 (O_299,N_9986,N_9921);
xnor UO_300 (O_300,N_9981,N_9934);
and UO_301 (O_301,N_9935,N_9910);
and UO_302 (O_302,N_9928,N_9959);
xor UO_303 (O_303,N_9975,N_9917);
or UO_304 (O_304,N_9954,N_9947);
nand UO_305 (O_305,N_9925,N_9908);
and UO_306 (O_306,N_9904,N_9994);
nand UO_307 (O_307,N_9983,N_9969);
or UO_308 (O_308,N_9918,N_9953);
or UO_309 (O_309,N_9939,N_9990);
xnor UO_310 (O_310,N_9905,N_9934);
and UO_311 (O_311,N_9947,N_9996);
or UO_312 (O_312,N_9910,N_9952);
nand UO_313 (O_313,N_9975,N_9958);
nor UO_314 (O_314,N_9988,N_9957);
and UO_315 (O_315,N_9922,N_9919);
or UO_316 (O_316,N_9986,N_9907);
or UO_317 (O_317,N_9989,N_9925);
xnor UO_318 (O_318,N_9979,N_9912);
and UO_319 (O_319,N_9903,N_9958);
or UO_320 (O_320,N_9916,N_9909);
nand UO_321 (O_321,N_9932,N_9967);
nand UO_322 (O_322,N_9901,N_9926);
xnor UO_323 (O_323,N_9996,N_9922);
and UO_324 (O_324,N_9902,N_9963);
nor UO_325 (O_325,N_9924,N_9910);
nand UO_326 (O_326,N_9929,N_9961);
xnor UO_327 (O_327,N_9945,N_9964);
or UO_328 (O_328,N_9942,N_9993);
and UO_329 (O_329,N_9978,N_9945);
and UO_330 (O_330,N_9993,N_9938);
nand UO_331 (O_331,N_9903,N_9911);
nand UO_332 (O_332,N_9976,N_9986);
and UO_333 (O_333,N_9990,N_9925);
xnor UO_334 (O_334,N_9988,N_9945);
or UO_335 (O_335,N_9948,N_9930);
or UO_336 (O_336,N_9992,N_9919);
xor UO_337 (O_337,N_9970,N_9924);
nor UO_338 (O_338,N_9977,N_9984);
or UO_339 (O_339,N_9962,N_9982);
nor UO_340 (O_340,N_9979,N_9922);
and UO_341 (O_341,N_9900,N_9973);
nor UO_342 (O_342,N_9984,N_9974);
or UO_343 (O_343,N_9997,N_9939);
and UO_344 (O_344,N_9929,N_9949);
and UO_345 (O_345,N_9982,N_9956);
and UO_346 (O_346,N_9942,N_9946);
nand UO_347 (O_347,N_9966,N_9952);
xor UO_348 (O_348,N_9960,N_9946);
xor UO_349 (O_349,N_9923,N_9939);
nor UO_350 (O_350,N_9957,N_9952);
or UO_351 (O_351,N_9955,N_9986);
xor UO_352 (O_352,N_9994,N_9982);
and UO_353 (O_353,N_9922,N_9924);
nand UO_354 (O_354,N_9916,N_9993);
or UO_355 (O_355,N_9974,N_9959);
nand UO_356 (O_356,N_9958,N_9952);
xor UO_357 (O_357,N_9900,N_9966);
and UO_358 (O_358,N_9943,N_9986);
nor UO_359 (O_359,N_9909,N_9956);
nand UO_360 (O_360,N_9973,N_9958);
xnor UO_361 (O_361,N_9947,N_9983);
nor UO_362 (O_362,N_9924,N_9919);
nand UO_363 (O_363,N_9997,N_9974);
nor UO_364 (O_364,N_9952,N_9901);
nand UO_365 (O_365,N_9983,N_9979);
nand UO_366 (O_366,N_9971,N_9938);
nor UO_367 (O_367,N_9967,N_9937);
nor UO_368 (O_368,N_9955,N_9957);
nor UO_369 (O_369,N_9923,N_9935);
nand UO_370 (O_370,N_9920,N_9986);
nand UO_371 (O_371,N_9900,N_9935);
and UO_372 (O_372,N_9975,N_9942);
xnor UO_373 (O_373,N_9960,N_9920);
and UO_374 (O_374,N_9923,N_9966);
and UO_375 (O_375,N_9950,N_9977);
xnor UO_376 (O_376,N_9996,N_9941);
and UO_377 (O_377,N_9988,N_9962);
and UO_378 (O_378,N_9996,N_9940);
and UO_379 (O_379,N_9980,N_9991);
or UO_380 (O_380,N_9971,N_9978);
nand UO_381 (O_381,N_9977,N_9960);
xor UO_382 (O_382,N_9961,N_9903);
nand UO_383 (O_383,N_9993,N_9932);
nor UO_384 (O_384,N_9934,N_9972);
or UO_385 (O_385,N_9979,N_9993);
nand UO_386 (O_386,N_9912,N_9921);
nand UO_387 (O_387,N_9968,N_9919);
nor UO_388 (O_388,N_9993,N_9954);
or UO_389 (O_389,N_9966,N_9929);
nor UO_390 (O_390,N_9974,N_9956);
and UO_391 (O_391,N_9944,N_9914);
nor UO_392 (O_392,N_9939,N_9958);
or UO_393 (O_393,N_9988,N_9939);
nor UO_394 (O_394,N_9951,N_9960);
nor UO_395 (O_395,N_9912,N_9901);
or UO_396 (O_396,N_9942,N_9985);
and UO_397 (O_397,N_9951,N_9935);
nor UO_398 (O_398,N_9927,N_9924);
nor UO_399 (O_399,N_9910,N_9940);
xor UO_400 (O_400,N_9936,N_9998);
nor UO_401 (O_401,N_9933,N_9935);
nand UO_402 (O_402,N_9925,N_9934);
nor UO_403 (O_403,N_9956,N_9939);
and UO_404 (O_404,N_9990,N_9960);
xor UO_405 (O_405,N_9928,N_9927);
nand UO_406 (O_406,N_9964,N_9940);
nor UO_407 (O_407,N_9994,N_9940);
or UO_408 (O_408,N_9980,N_9916);
nand UO_409 (O_409,N_9983,N_9905);
and UO_410 (O_410,N_9926,N_9930);
or UO_411 (O_411,N_9918,N_9994);
xnor UO_412 (O_412,N_9978,N_9941);
nor UO_413 (O_413,N_9953,N_9952);
xor UO_414 (O_414,N_9942,N_9953);
nand UO_415 (O_415,N_9991,N_9928);
xnor UO_416 (O_416,N_9983,N_9978);
or UO_417 (O_417,N_9982,N_9926);
and UO_418 (O_418,N_9981,N_9907);
nand UO_419 (O_419,N_9903,N_9935);
xor UO_420 (O_420,N_9949,N_9978);
or UO_421 (O_421,N_9921,N_9955);
nand UO_422 (O_422,N_9900,N_9937);
or UO_423 (O_423,N_9961,N_9933);
or UO_424 (O_424,N_9972,N_9923);
and UO_425 (O_425,N_9919,N_9959);
nand UO_426 (O_426,N_9969,N_9991);
or UO_427 (O_427,N_9984,N_9910);
nand UO_428 (O_428,N_9909,N_9946);
nand UO_429 (O_429,N_9979,N_9929);
nand UO_430 (O_430,N_9939,N_9987);
xor UO_431 (O_431,N_9933,N_9948);
nand UO_432 (O_432,N_9988,N_9959);
xnor UO_433 (O_433,N_9972,N_9914);
nand UO_434 (O_434,N_9945,N_9929);
nor UO_435 (O_435,N_9945,N_9956);
or UO_436 (O_436,N_9975,N_9953);
xor UO_437 (O_437,N_9957,N_9916);
nand UO_438 (O_438,N_9935,N_9963);
nand UO_439 (O_439,N_9942,N_9963);
nor UO_440 (O_440,N_9909,N_9902);
nand UO_441 (O_441,N_9908,N_9996);
xor UO_442 (O_442,N_9915,N_9911);
and UO_443 (O_443,N_9973,N_9903);
nor UO_444 (O_444,N_9976,N_9969);
or UO_445 (O_445,N_9922,N_9972);
xnor UO_446 (O_446,N_9947,N_9902);
xor UO_447 (O_447,N_9915,N_9935);
or UO_448 (O_448,N_9901,N_9989);
nand UO_449 (O_449,N_9903,N_9999);
nand UO_450 (O_450,N_9978,N_9970);
and UO_451 (O_451,N_9980,N_9942);
xor UO_452 (O_452,N_9946,N_9957);
or UO_453 (O_453,N_9918,N_9987);
xnor UO_454 (O_454,N_9930,N_9956);
xnor UO_455 (O_455,N_9936,N_9918);
xor UO_456 (O_456,N_9978,N_9956);
nor UO_457 (O_457,N_9968,N_9925);
or UO_458 (O_458,N_9933,N_9949);
xnor UO_459 (O_459,N_9937,N_9982);
and UO_460 (O_460,N_9949,N_9941);
nor UO_461 (O_461,N_9922,N_9947);
and UO_462 (O_462,N_9904,N_9990);
xnor UO_463 (O_463,N_9956,N_9912);
nor UO_464 (O_464,N_9937,N_9976);
nor UO_465 (O_465,N_9998,N_9983);
nor UO_466 (O_466,N_9997,N_9986);
nor UO_467 (O_467,N_9983,N_9982);
xor UO_468 (O_468,N_9992,N_9953);
and UO_469 (O_469,N_9922,N_9973);
xor UO_470 (O_470,N_9909,N_9919);
nor UO_471 (O_471,N_9980,N_9996);
or UO_472 (O_472,N_9972,N_9983);
nand UO_473 (O_473,N_9909,N_9973);
nand UO_474 (O_474,N_9942,N_9926);
xnor UO_475 (O_475,N_9959,N_9952);
nand UO_476 (O_476,N_9991,N_9956);
nor UO_477 (O_477,N_9986,N_9930);
nand UO_478 (O_478,N_9937,N_9995);
nor UO_479 (O_479,N_9960,N_9986);
nand UO_480 (O_480,N_9993,N_9931);
nor UO_481 (O_481,N_9989,N_9980);
xnor UO_482 (O_482,N_9993,N_9944);
xnor UO_483 (O_483,N_9957,N_9920);
nand UO_484 (O_484,N_9929,N_9974);
nand UO_485 (O_485,N_9943,N_9955);
nor UO_486 (O_486,N_9986,N_9906);
or UO_487 (O_487,N_9991,N_9979);
xor UO_488 (O_488,N_9970,N_9929);
xor UO_489 (O_489,N_9928,N_9935);
or UO_490 (O_490,N_9977,N_9937);
xnor UO_491 (O_491,N_9943,N_9999);
nor UO_492 (O_492,N_9945,N_9981);
xor UO_493 (O_493,N_9975,N_9950);
and UO_494 (O_494,N_9906,N_9990);
or UO_495 (O_495,N_9975,N_9932);
nor UO_496 (O_496,N_9956,N_9938);
nand UO_497 (O_497,N_9925,N_9976);
or UO_498 (O_498,N_9927,N_9959);
nand UO_499 (O_499,N_9999,N_9938);
nor UO_500 (O_500,N_9931,N_9906);
nor UO_501 (O_501,N_9931,N_9995);
nand UO_502 (O_502,N_9966,N_9927);
and UO_503 (O_503,N_9999,N_9901);
nand UO_504 (O_504,N_9975,N_9915);
nor UO_505 (O_505,N_9975,N_9967);
xnor UO_506 (O_506,N_9916,N_9940);
and UO_507 (O_507,N_9944,N_9978);
or UO_508 (O_508,N_9987,N_9965);
nand UO_509 (O_509,N_9940,N_9990);
and UO_510 (O_510,N_9902,N_9996);
nor UO_511 (O_511,N_9951,N_9988);
or UO_512 (O_512,N_9917,N_9936);
and UO_513 (O_513,N_9965,N_9969);
nand UO_514 (O_514,N_9906,N_9997);
xnor UO_515 (O_515,N_9906,N_9943);
xor UO_516 (O_516,N_9988,N_9926);
nand UO_517 (O_517,N_9928,N_9947);
or UO_518 (O_518,N_9980,N_9906);
nor UO_519 (O_519,N_9958,N_9997);
or UO_520 (O_520,N_9972,N_9970);
nand UO_521 (O_521,N_9968,N_9967);
and UO_522 (O_522,N_9988,N_9976);
and UO_523 (O_523,N_9960,N_9949);
and UO_524 (O_524,N_9996,N_9952);
nor UO_525 (O_525,N_9999,N_9970);
and UO_526 (O_526,N_9929,N_9934);
nand UO_527 (O_527,N_9918,N_9921);
nand UO_528 (O_528,N_9937,N_9914);
and UO_529 (O_529,N_9999,N_9944);
or UO_530 (O_530,N_9964,N_9990);
xnor UO_531 (O_531,N_9940,N_9905);
nor UO_532 (O_532,N_9975,N_9969);
nand UO_533 (O_533,N_9979,N_9970);
or UO_534 (O_534,N_9915,N_9931);
nor UO_535 (O_535,N_9944,N_9908);
nor UO_536 (O_536,N_9999,N_9996);
xnor UO_537 (O_537,N_9974,N_9925);
xnor UO_538 (O_538,N_9928,N_9961);
xnor UO_539 (O_539,N_9922,N_9951);
or UO_540 (O_540,N_9925,N_9918);
nand UO_541 (O_541,N_9942,N_9979);
and UO_542 (O_542,N_9997,N_9967);
and UO_543 (O_543,N_9942,N_9908);
or UO_544 (O_544,N_9938,N_9978);
and UO_545 (O_545,N_9986,N_9931);
and UO_546 (O_546,N_9909,N_9953);
xnor UO_547 (O_547,N_9939,N_9955);
nand UO_548 (O_548,N_9900,N_9959);
nand UO_549 (O_549,N_9903,N_9983);
xnor UO_550 (O_550,N_9999,N_9971);
nand UO_551 (O_551,N_9943,N_9922);
nand UO_552 (O_552,N_9945,N_9930);
and UO_553 (O_553,N_9986,N_9905);
and UO_554 (O_554,N_9953,N_9934);
nor UO_555 (O_555,N_9975,N_9945);
nor UO_556 (O_556,N_9909,N_9951);
or UO_557 (O_557,N_9946,N_9901);
or UO_558 (O_558,N_9940,N_9938);
nor UO_559 (O_559,N_9977,N_9933);
xor UO_560 (O_560,N_9939,N_9934);
xnor UO_561 (O_561,N_9923,N_9905);
and UO_562 (O_562,N_9924,N_9920);
xor UO_563 (O_563,N_9928,N_9962);
and UO_564 (O_564,N_9956,N_9996);
nand UO_565 (O_565,N_9999,N_9946);
or UO_566 (O_566,N_9916,N_9944);
and UO_567 (O_567,N_9973,N_9994);
nor UO_568 (O_568,N_9913,N_9971);
nor UO_569 (O_569,N_9929,N_9942);
and UO_570 (O_570,N_9978,N_9927);
nor UO_571 (O_571,N_9918,N_9914);
nor UO_572 (O_572,N_9935,N_9902);
and UO_573 (O_573,N_9936,N_9988);
or UO_574 (O_574,N_9923,N_9984);
xor UO_575 (O_575,N_9978,N_9958);
and UO_576 (O_576,N_9999,N_9974);
nand UO_577 (O_577,N_9955,N_9978);
xnor UO_578 (O_578,N_9992,N_9968);
xor UO_579 (O_579,N_9923,N_9925);
nor UO_580 (O_580,N_9975,N_9931);
xnor UO_581 (O_581,N_9926,N_9916);
nor UO_582 (O_582,N_9955,N_9946);
xor UO_583 (O_583,N_9957,N_9984);
or UO_584 (O_584,N_9937,N_9927);
nor UO_585 (O_585,N_9919,N_9939);
and UO_586 (O_586,N_9935,N_9929);
or UO_587 (O_587,N_9913,N_9940);
or UO_588 (O_588,N_9938,N_9933);
or UO_589 (O_589,N_9938,N_9970);
and UO_590 (O_590,N_9983,N_9934);
nor UO_591 (O_591,N_9940,N_9936);
and UO_592 (O_592,N_9952,N_9944);
or UO_593 (O_593,N_9965,N_9983);
xor UO_594 (O_594,N_9906,N_9902);
nor UO_595 (O_595,N_9981,N_9970);
nand UO_596 (O_596,N_9982,N_9936);
and UO_597 (O_597,N_9980,N_9950);
nand UO_598 (O_598,N_9986,N_9998);
or UO_599 (O_599,N_9922,N_9954);
xnor UO_600 (O_600,N_9924,N_9980);
nor UO_601 (O_601,N_9905,N_9931);
nand UO_602 (O_602,N_9962,N_9931);
nor UO_603 (O_603,N_9958,N_9923);
or UO_604 (O_604,N_9949,N_9975);
and UO_605 (O_605,N_9976,N_9964);
nand UO_606 (O_606,N_9907,N_9998);
and UO_607 (O_607,N_9970,N_9930);
nor UO_608 (O_608,N_9938,N_9961);
nand UO_609 (O_609,N_9963,N_9968);
nand UO_610 (O_610,N_9911,N_9909);
or UO_611 (O_611,N_9918,N_9989);
xor UO_612 (O_612,N_9924,N_9953);
nor UO_613 (O_613,N_9963,N_9984);
and UO_614 (O_614,N_9949,N_9912);
nand UO_615 (O_615,N_9903,N_9981);
xor UO_616 (O_616,N_9974,N_9940);
nor UO_617 (O_617,N_9921,N_9992);
nor UO_618 (O_618,N_9944,N_9909);
nor UO_619 (O_619,N_9937,N_9956);
xor UO_620 (O_620,N_9935,N_9937);
nor UO_621 (O_621,N_9979,N_9999);
xnor UO_622 (O_622,N_9906,N_9957);
xor UO_623 (O_623,N_9972,N_9989);
and UO_624 (O_624,N_9971,N_9956);
and UO_625 (O_625,N_9990,N_9961);
xnor UO_626 (O_626,N_9919,N_9944);
xnor UO_627 (O_627,N_9941,N_9921);
nand UO_628 (O_628,N_9921,N_9997);
nand UO_629 (O_629,N_9973,N_9945);
nor UO_630 (O_630,N_9927,N_9998);
nand UO_631 (O_631,N_9935,N_9939);
xnor UO_632 (O_632,N_9966,N_9932);
nor UO_633 (O_633,N_9945,N_9937);
xnor UO_634 (O_634,N_9904,N_9947);
nor UO_635 (O_635,N_9964,N_9952);
xnor UO_636 (O_636,N_9987,N_9904);
and UO_637 (O_637,N_9942,N_9982);
or UO_638 (O_638,N_9983,N_9990);
and UO_639 (O_639,N_9998,N_9993);
or UO_640 (O_640,N_9955,N_9933);
nand UO_641 (O_641,N_9979,N_9963);
and UO_642 (O_642,N_9928,N_9939);
nand UO_643 (O_643,N_9900,N_9980);
nand UO_644 (O_644,N_9958,N_9962);
or UO_645 (O_645,N_9924,N_9934);
xnor UO_646 (O_646,N_9997,N_9903);
or UO_647 (O_647,N_9938,N_9964);
xor UO_648 (O_648,N_9942,N_9918);
nand UO_649 (O_649,N_9932,N_9965);
and UO_650 (O_650,N_9999,N_9957);
xor UO_651 (O_651,N_9927,N_9985);
nand UO_652 (O_652,N_9989,N_9999);
or UO_653 (O_653,N_9961,N_9936);
and UO_654 (O_654,N_9950,N_9948);
or UO_655 (O_655,N_9962,N_9977);
nand UO_656 (O_656,N_9921,N_9967);
or UO_657 (O_657,N_9979,N_9944);
nor UO_658 (O_658,N_9972,N_9992);
xor UO_659 (O_659,N_9987,N_9995);
and UO_660 (O_660,N_9981,N_9929);
xnor UO_661 (O_661,N_9973,N_9977);
xnor UO_662 (O_662,N_9904,N_9911);
xnor UO_663 (O_663,N_9915,N_9973);
xnor UO_664 (O_664,N_9965,N_9989);
nor UO_665 (O_665,N_9904,N_9943);
nor UO_666 (O_666,N_9989,N_9932);
and UO_667 (O_667,N_9915,N_9941);
nor UO_668 (O_668,N_9906,N_9909);
xor UO_669 (O_669,N_9990,N_9915);
or UO_670 (O_670,N_9957,N_9939);
or UO_671 (O_671,N_9912,N_9992);
xor UO_672 (O_672,N_9991,N_9945);
nand UO_673 (O_673,N_9990,N_9920);
xnor UO_674 (O_674,N_9985,N_9935);
or UO_675 (O_675,N_9919,N_9998);
or UO_676 (O_676,N_9983,N_9997);
xor UO_677 (O_677,N_9951,N_9967);
nand UO_678 (O_678,N_9922,N_9967);
xnor UO_679 (O_679,N_9960,N_9925);
or UO_680 (O_680,N_9924,N_9915);
nand UO_681 (O_681,N_9930,N_9904);
and UO_682 (O_682,N_9963,N_9956);
xnor UO_683 (O_683,N_9996,N_9939);
and UO_684 (O_684,N_9957,N_9922);
or UO_685 (O_685,N_9927,N_9954);
and UO_686 (O_686,N_9933,N_9990);
and UO_687 (O_687,N_9977,N_9983);
nor UO_688 (O_688,N_9943,N_9929);
and UO_689 (O_689,N_9909,N_9922);
or UO_690 (O_690,N_9933,N_9921);
or UO_691 (O_691,N_9947,N_9962);
xor UO_692 (O_692,N_9998,N_9938);
nor UO_693 (O_693,N_9985,N_9909);
nor UO_694 (O_694,N_9934,N_9998);
nor UO_695 (O_695,N_9902,N_9966);
and UO_696 (O_696,N_9900,N_9902);
xnor UO_697 (O_697,N_9936,N_9965);
nor UO_698 (O_698,N_9943,N_9900);
xor UO_699 (O_699,N_9982,N_9928);
or UO_700 (O_700,N_9988,N_9941);
or UO_701 (O_701,N_9941,N_9951);
or UO_702 (O_702,N_9901,N_9945);
and UO_703 (O_703,N_9939,N_9977);
and UO_704 (O_704,N_9940,N_9992);
and UO_705 (O_705,N_9922,N_9930);
nand UO_706 (O_706,N_9921,N_9984);
and UO_707 (O_707,N_9948,N_9945);
and UO_708 (O_708,N_9984,N_9978);
xnor UO_709 (O_709,N_9911,N_9913);
or UO_710 (O_710,N_9941,N_9993);
and UO_711 (O_711,N_9949,N_9995);
or UO_712 (O_712,N_9907,N_9962);
nand UO_713 (O_713,N_9907,N_9905);
nand UO_714 (O_714,N_9996,N_9963);
xor UO_715 (O_715,N_9975,N_9938);
or UO_716 (O_716,N_9996,N_9958);
nand UO_717 (O_717,N_9982,N_9964);
and UO_718 (O_718,N_9952,N_9925);
or UO_719 (O_719,N_9919,N_9948);
xor UO_720 (O_720,N_9952,N_9913);
and UO_721 (O_721,N_9968,N_9905);
xnor UO_722 (O_722,N_9901,N_9994);
or UO_723 (O_723,N_9924,N_9945);
nand UO_724 (O_724,N_9934,N_9984);
xor UO_725 (O_725,N_9980,N_9954);
or UO_726 (O_726,N_9971,N_9917);
and UO_727 (O_727,N_9949,N_9946);
nor UO_728 (O_728,N_9983,N_9995);
or UO_729 (O_729,N_9923,N_9956);
xor UO_730 (O_730,N_9961,N_9977);
and UO_731 (O_731,N_9960,N_9900);
and UO_732 (O_732,N_9966,N_9926);
xor UO_733 (O_733,N_9977,N_9934);
nand UO_734 (O_734,N_9909,N_9941);
or UO_735 (O_735,N_9992,N_9908);
xnor UO_736 (O_736,N_9978,N_9952);
nand UO_737 (O_737,N_9966,N_9916);
or UO_738 (O_738,N_9927,N_9946);
xor UO_739 (O_739,N_9977,N_9917);
or UO_740 (O_740,N_9970,N_9903);
xor UO_741 (O_741,N_9973,N_9939);
and UO_742 (O_742,N_9993,N_9902);
or UO_743 (O_743,N_9963,N_9998);
nor UO_744 (O_744,N_9967,N_9939);
and UO_745 (O_745,N_9959,N_9901);
xor UO_746 (O_746,N_9965,N_9985);
xor UO_747 (O_747,N_9959,N_9985);
nand UO_748 (O_748,N_9981,N_9921);
xor UO_749 (O_749,N_9984,N_9900);
and UO_750 (O_750,N_9937,N_9920);
nand UO_751 (O_751,N_9955,N_9950);
xnor UO_752 (O_752,N_9971,N_9969);
nor UO_753 (O_753,N_9991,N_9982);
nand UO_754 (O_754,N_9917,N_9950);
nor UO_755 (O_755,N_9900,N_9939);
or UO_756 (O_756,N_9935,N_9974);
nor UO_757 (O_757,N_9994,N_9988);
nand UO_758 (O_758,N_9980,N_9940);
and UO_759 (O_759,N_9971,N_9909);
or UO_760 (O_760,N_9905,N_9943);
nand UO_761 (O_761,N_9907,N_9901);
and UO_762 (O_762,N_9983,N_9929);
nand UO_763 (O_763,N_9926,N_9947);
or UO_764 (O_764,N_9970,N_9918);
nand UO_765 (O_765,N_9995,N_9917);
xnor UO_766 (O_766,N_9962,N_9912);
and UO_767 (O_767,N_9992,N_9959);
xor UO_768 (O_768,N_9964,N_9963);
and UO_769 (O_769,N_9908,N_9912);
nand UO_770 (O_770,N_9976,N_9965);
xor UO_771 (O_771,N_9959,N_9922);
nor UO_772 (O_772,N_9979,N_9928);
or UO_773 (O_773,N_9956,N_9935);
xnor UO_774 (O_774,N_9967,N_9963);
xnor UO_775 (O_775,N_9901,N_9998);
or UO_776 (O_776,N_9971,N_9962);
xor UO_777 (O_777,N_9903,N_9967);
nand UO_778 (O_778,N_9964,N_9939);
nor UO_779 (O_779,N_9994,N_9979);
nor UO_780 (O_780,N_9948,N_9960);
and UO_781 (O_781,N_9941,N_9931);
xor UO_782 (O_782,N_9975,N_9984);
nor UO_783 (O_783,N_9981,N_9900);
nor UO_784 (O_784,N_9978,N_9919);
and UO_785 (O_785,N_9911,N_9989);
xnor UO_786 (O_786,N_9989,N_9947);
nor UO_787 (O_787,N_9946,N_9969);
xor UO_788 (O_788,N_9901,N_9978);
nor UO_789 (O_789,N_9957,N_9937);
nor UO_790 (O_790,N_9949,N_9987);
and UO_791 (O_791,N_9916,N_9996);
nor UO_792 (O_792,N_9907,N_9953);
nand UO_793 (O_793,N_9965,N_9974);
nor UO_794 (O_794,N_9990,N_9916);
nand UO_795 (O_795,N_9978,N_9930);
and UO_796 (O_796,N_9904,N_9972);
nand UO_797 (O_797,N_9964,N_9969);
and UO_798 (O_798,N_9942,N_9922);
or UO_799 (O_799,N_9953,N_9968);
nand UO_800 (O_800,N_9979,N_9982);
xnor UO_801 (O_801,N_9937,N_9974);
or UO_802 (O_802,N_9967,N_9964);
nand UO_803 (O_803,N_9999,N_9930);
xnor UO_804 (O_804,N_9970,N_9941);
xnor UO_805 (O_805,N_9998,N_9965);
xnor UO_806 (O_806,N_9999,N_9942);
nand UO_807 (O_807,N_9911,N_9988);
and UO_808 (O_808,N_9952,N_9989);
or UO_809 (O_809,N_9939,N_9946);
nor UO_810 (O_810,N_9962,N_9953);
and UO_811 (O_811,N_9913,N_9930);
nand UO_812 (O_812,N_9951,N_9925);
xor UO_813 (O_813,N_9981,N_9928);
nor UO_814 (O_814,N_9918,N_9976);
nor UO_815 (O_815,N_9917,N_9982);
nand UO_816 (O_816,N_9917,N_9922);
or UO_817 (O_817,N_9910,N_9989);
xnor UO_818 (O_818,N_9907,N_9973);
nand UO_819 (O_819,N_9923,N_9929);
and UO_820 (O_820,N_9908,N_9915);
nand UO_821 (O_821,N_9908,N_9941);
nand UO_822 (O_822,N_9939,N_9985);
nor UO_823 (O_823,N_9991,N_9914);
nor UO_824 (O_824,N_9993,N_9992);
or UO_825 (O_825,N_9917,N_9949);
nor UO_826 (O_826,N_9975,N_9980);
or UO_827 (O_827,N_9977,N_9915);
nor UO_828 (O_828,N_9950,N_9996);
or UO_829 (O_829,N_9932,N_9905);
nand UO_830 (O_830,N_9999,N_9945);
and UO_831 (O_831,N_9986,N_9948);
and UO_832 (O_832,N_9955,N_9902);
and UO_833 (O_833,N_9907,N_9925);
and UO_834 (O_834,N_9939,N_9910);
nand UO_835 (O_835,N_9914,N_9901);
and UO_836 (O_836,N_9914,N_9953);
nor UO_837 (O_837,N_9922,N_9940);
and UO_838 (O_838,N_9995,N_9955);
nor UO_839 (O_839,N_9938,N_9952);
or UO_840 (O_840,N_9911,N_9960);
xnor UO_841 (O_841,N_9955,N_9951);
nor UO_842 (O_842,N_9934,N_9943);
nand UO_843 (O_843,N_9904,N_9969);
nor UO_844 (O_844,N_9954,N_9981);
nand UO_845 (O_845,N_9952,N_9939);
and UO_846 (O_846,N_9993,N_9922);
or UO_847 (O_847,N_9917,N_9900);
xnor UO_848 (O_848,N_9954,N_9911);
nand UO_849 (O_849,N_9953,N_9915);
nor UO_850 (O_850,N_9967,N_9906);
nor UO_851 (O_851,N_9985,N_9932);
nor UO_852 (O_852,N_9931,N_9923);
or UO_853 (O_853,N_9947,N_9965);
xnor UO_854 (O_854,N_9908,N_9961);
nor UO_855 (O_855,N_9930,N_9963);
nand UO_856 (O_856,N_9983,N_9921);
xnor UO_857 (O_857,N_9941,N_9966);
xnor UO_858 (O_858,N_9929,N_9959);
nor UO_859 (O_859,N_9916,N_9951);
xnor UO_860 (O_860,N_9984,N_9917);
xor UO_861 (O_861,N_9936,N_9924);
and UO_862 (O_862,N_9996,N_9989);
nand UO_863 (O_863,N_9980,N_9952);
nand UO_864 (O_864,N_9981,N_9961);
and UO_865 (O_865,N_9936,N_9900);
or UO_866 (O_866,N_9934,N_9994);
xor UO_867 (O_867,N_9953,N_9994);
and UO_868 (O_868,N_9906,N_9999);
nand UO_869 (O_869,N_9923,N_9937);
or UO_870 (O_870,N_9914,N_9935);
xnor UO_871 (O_871,N_9907,N_9937);
xnor UO_872 (O_872,N_9972,N_9978);
and UO_873 (O_873,N_9953,N_9987);
or UO_874 (O_874,N_9975,N_9986);
or UO_875 (O_875,N_9900,N_9908);
and UO_876 (O_876,N_9916,N_9929);
or UO_877 (O_877,N_9969,N_9955);
nor UO_878 (O_878,N_9936,N_9934);
nor UO_879 (O_879,N_9966,N_9960);
or UO_880 (O_880,N_9915,N_9932);
or UO_881 (O_881,N_9930,N_9920);
nand UO_882 (O_882,N_9910,N_9946);
nand UO_883 (O_883,N_9906,N_9992);
nand UO_884 (O_884,N_9917,N_9974);
or UO_885 (O_885,N_9950,N_9976);
nor UO_886 (O_886,N_9938,N_9913);
or UO_887 (O_887,N_9906,N_9921);
nor UO_888 (O_888,N_9997,N_9940);
nand UO_889 (O_889,N_9992,N_9990);
nor UO_890 (O_890,N_9925,N_9900);
xor UO_891 (O_891,N_9964,N_9932);
and UO_892 (O_892,N_9930,N_9918);
and UO_893 (O_893,N_9934,N_9915);
nor UO_894 (O_894,N_9901,N_9933);
nor UO_895 (O_895,N_9913,N_9972);
nor UO_896 (O_896,N_9989,N_9933);
nand UO_897 (O_897,N_9954,N_9932);
nand UO_898 (O_898,N_9962,N_9968);
xor UO_899 (O_899,N_9954,N_9934);
or UO_900 (O_900,N_9950,N_9985);
and UO_901 (O_901,N_9913,N_9986);
or UO_902 (O_902,N_9970,N_9912);
or UO_903 (O_903,N_9917,N_9994);
and UO_904 (O_904,N_9947,N_9966);
xor UO_905 (O_905,N_9909,N_9940);
nor UO_906 (O_906,N_9963,N_9944);
xnor UO_907 (O_907,N_9982,N_9971);
nand UO_908 (O_908,N_9940,N_9941);
and UO_909 (O_909,N_9958,N_9936);
nor UO_910 (O_910,N_9955,N_9916);
and UO_911 (O_911,N_9906,N_9932);
nor UO_912 (O_912,N_9948,N_9926);
nand UO_913 (O_913,N_9966,N_9997);
and UO_914 (O_914,N_9906,N_9929);
nor UO_915 (O_915,N_9945,N_9965);
xor UO_916 (O_916,N_9967,N_9917);
and UO_917 (O_917,N_9972,N_9929);
nor UO_918 (O_918,N_9986,N_9946);
nand UO_919 (O_919,N_9976,N_9932);
or UO_920 (O_920,N_9903,N_9910);
nor UO_921 (O_921,N_9948,N_9968);
or UO_922 (O_922,N_9957,N_9959);
xor UO_923 (O_923,N_9933,N_9982);
nand UO_924 (O_924,N_9936,N_9975);
xnor UO_925 (O_925,N_9938,N_9904);
nand UO_926 (O_926,N_9960,N_9921);
or UO_927 (O_927,N_9976,N_9916);
xor UO_928 (O_928,N_9967,N_9907);
nor UO_929 (O_929,N_9967,N_9929);
or UO_930 (O_930,N_9936,N_9957);
and UO_931 (O_931,N_9957,N_9902);
nor UO_932 (O_932,N_9966,N_9954);
xor UO_933 (O_933,N_9972,N_9988);
nor UO_934 (O_934,N_9941,N_9945);
and UO_935 (O_935,N_9921,N_9990);
xor UO_936 (O_936,N_9901,N_9921);
nor UO_937 (O_937,N_9980,N_9926);
and UO_938 (O_938,N_9965,N_9911);
nor UO_939 (O_939,N_9955,N_9998);
nand UO_940 (O_940,N_9945,N_9900);
nand UO_941 (O_941,N_9915,N_9969);
or UO_942 (O_942,N_9974,N_9991);
nor UO_943 (O_943,N_9955,N_9959);
and UO_944 (O_944,N_9929,N_9994);
nor UO_945 (O_945,N_9977,N_9988);
nand UO_946 (O_946,N_9961,N_9956);
xor UO_947 (O_947,N_9979,N_9955);
and UO_948 (O_948,N_9983,N_9939);
nand UO_949 (O_949,N_9947,N_9977);
nand UO_950 (O_950,N_9975,N_9901);
nor UO_951 (O_951,N_9990,N_9971);
or UO_952 (O_952,N_9951,N_9995);
xor UO_953 (O_953,N_9917,N_9955);
and UO_954 (O_954,N_9912,N_9919);
xnor UO_955 (O_955,N_9932,N_9992);
and UO_956 (O_956,N_9983,N_9911);
xnor UO_957 (O_957,N_9915,N_9916);
xnor UO_958 (O_958,N_9992,N_9979);
xor UO_959 (O_959,N_9972,N_9928);
and UO_960 (O_960,N_9986,N_9939);
xnor UO_961 (O_961,N_9903,N_9979);
nor UO_962 (O_962,N_9978,N_9990);
or UO_963 (O_963,N_9967,N_9985);
or UO_964 (O_964,N_9945,N_9996);
nand UO_965 (O_965,N_9957,N_9909);
xor UO_966 (O_966,N_9915,N_9963);
nand UO_967 (O_967,N_9971,N_9933);
xnor UO_968 (O_968,N_9907,N_9903);
or UO_969 (O_969,N_9996,N_9928);
or UO_970 (O_970,N_9925,N_9987);
nand UO_971 (O_971,N_9993,N_9940);
and UO_972 (O_972,N_9986,N_9942);
nand UO_973 (O_973,N_9942,N_9990);
and UO_974 (O_974,N_9993,N_9952);
nand UO_975 (O_975,N_9935,N_9905);
or UO_976 (O_976,N_9934,N_9976);
nor UO_977 (O_977,N_9926,N_9951);
nand UO_978 (O_978,N_9983,N_9992);
nor UO_979 (O_979,N_9933,N_9939);
and UO_980 (O_980,N_9922,N_9963);
xnor UO_981 (O_981,N_9994,N_9902);
nor UO_982 (O_982,N_9949,N_9997);
nor UO_983 (O_983,N_9960,N_9959);
nor UO_984 (O_984,N_9981,N_9935);
and UO_985 (O_985,N_9977,N_9982);
nand UO_986 (O_986,N_9950,N_9978);
nand UO_987 (O_987,N_9920,N_9942);
and UO_988 (O_988,N_9938,N_9945);
xor UO_989 (O_989,N_9912,N_9922);
or UO_990 (O_990,N_9953,N_9998);
xnor UO_991 (O_991,N_9960,N_9970);
xor UO_992 (O_992,N_9940,N_9904);
xor UO_993 (O_993,N_9937,N_9975);
xnor UO_994 (O_994,N_9911,N_9976);
and UO_995 (O_995,N_9978,N_9977);
nand UO_996 (O_996,N_9962,N_9923);
xnor UO_997 (O_997,N_9962,N_9986);
or UO_998 (O_998,N_9943,N_9946);
nand UO_999 (O_999,N_9902,N_9975);
or UO_1000 (O_1000,N_9973,N_9934);
xnor UO_1001 (O_1001,N_9908,N_9958);
or UO_1002 (O_1002,N_9953,N_9985);
nor UO_1003 (O_1003,N_9994,N_9900);
or UO_1004 (O_1004,N_9904,N_9955);
or UO_1005 (O_1005,N_9903,N_9900);
and UO_1006 (O_1006,N_9955,N_9981);
xor UO_1007 (O_1007,N_9978,N_9907);
nor UO_1008 (O_1008,N_9927,N_9942);
nor UO_1009 (O_1009,N_9935,N_9924);
or UO_1010 (O_1010,N_9924,N_9923);
nand UO_1011 (O_1011,N_9937,N_9988);
and UO_1012 (O_1012,N_9967,N_9901);
nand UO_1013 (O_1013,N_9902,N_9925);
and UO_1014 (O_1014,N_9915,N_9917);
nor UO_1015 (O_1015,N_9931,N_9979);
or UO_1016 (O_1016,N_9922,N_9921);
nor UO_1017 (O_1017,N_9986,N_9934);
xnor UO_1018 (O_1018,N_9943,N_9961);
xnor UO_1019 (O_1019,N_9922,N_9931);
or UO_1020 (O_1020,N_9974,N_9912);
or UO_1021 (O_1021,N_9938,N_9928);
xnor UO_1022 (O_1022,N_9943,N_9923);
and UO_1023 (O_1023,N_9917,N_9906);
and UO_1024 (O_1024,N_9937,N_9972);
nand UO_1025 (O_1025,N_9988,N_9990);
or UO_1026 (O_1026,N_9989,N_9938);
or UO_1027 (O_1027,N_9934,N_9992);
xnor UO_1028 (O_1028,N_9973,N_9957);
xnor UO_1029 (O_1029,N_9907,N_9915);
nand UO_1030 (O_1030,N_9905,N_9908);
nor UO_1031 (O_1031,N_9966,N_9984);
nor UO_1032 (O_1032,N_9908,N_9918);
nand UO_1033 (O_1033,N_9918,N_9979);
nor UO_1034 (O_1034,N_9915,N_9974);
and UO_1035 (O_1035,N_9961,N_9983);
nand UO_1036 (O_1036,N_9907,N_9922);
or UO_1037 (O_1037,N_9990,N_9993);
nor UO_1038 (O_1038,N_9971,N_9979);
nand UO_1039 (O_1039,N_9997,N_9926);
nor UO_1040 (O_1040,N_9981,N_9939);
or UO_1041 (O_1041,N_9924,N_9940);
nand UO_1042 (O_1042,N_9945,N_9902);
xnor UO_1043 (O_1043,N_9995,N_9918);
and UO_1044 (O_1044,N_9910,N_9909);
or UO_1045 (O_1045,N_9997,N_9923);
nand UO_1046 (O_1046,N_9986,N_9940);
nor UO_1047 (O_1047,N_9914,N_9934);
or UO_1048 (O_1048,N_9922,N_9999);
nor UO_1049 (O_1049,N_9969,N_9913);
or UO_1050 (O_1050,N_9918,N_9993);
and UO_1051 (O_1051,N_9953,N_9938);
and UO_1052 (O_1052,N_9928,N_9918);
and UO_1053 (O_1053,N_9921,N_9961);
and UO_1054 (O_1054,N_9932,N_9963);
xnor UO_1055 (O_1055,N_9915,N_9988);
and UO_1056 (O_1056,N_9978,N_9997);
nor UO_1057 (O_1057,N_9906,N_9969);
nor UO_1058 (O_1058,N_9900,N_9972);
nor UO_1059 (O_1059,N_9979,N_9972);
nor UO_1060 (O_1060,N_9953,N_9949);
and UO_1061 (O_1061,N_9975,N_9998);
nor UO_1062 (O_1062,N_9930,N_9917);
or UO_1063 (O_1063,N_9996,N_9967);
nand UO_1064 (O_1064,N_9900,N_9969);
nand UO_1065 (O_1065,N_9958,N_9920);
or UO_1066 (O_1066,N_9944,N_9924);
or UO_1067 (O_1067,N_9960,N_9933);
xor UO_1068 (O_1068,N_9955,N_9983);
nor UO_1069 (O_1069,N_9921,N_9965);
xor UO_1070 (O_1070,N_9911,N_9929);
nand UO_1071 (O_1071,N_9960,N_9927);
and UO_1072 (O_1072,N_9966,N_9970);
and UO_1073 (O_1073,N_9916,N_9943);
and UO_1074 (O_1074,N_9998,N_9954);
nor UO_1075 (O_1075,N_9955,N_9988);
nand UO_1076 (O_1076,N_9901,N_9991);
and UO_1077 (O_1077,N_9972,N_9944);
and UO_1078 (O_1078,N_9988,N_9961);
or UO_1079 (O_1079,N_9985,N_9969);
or UO_1080 (O_1080,N_9994,N_9983);
nor UO_1081 (O_1081,N_9949,N_9982);
and UO_1082 (O_1082,N_9923,N_9967);
or UO_1083 (O_1083,N_9960,N_9916);
or UO_1084 (O_1084,N_9964,N_9905);
and UO_1085 (O_1085,N_9960,N_9913);
nor UO_1086 (O_1086,N_9962,N_9951);
nand UO_1087 (O_1087,N_9950,N_9994);
nand UO_1088 (O_1088,N_9926,N_9967);
and UO_1089 (O_1089,N_9967,N_9990);
xor UO_1090 (O_1090,N_9923,N_9981);
and UO_1091 (O_1091,N_9932,N_9950);
xnor UO_1092 (O_1092,N_9903,N_9954);
nor UO_1093 (O_1093,N_9926,N_9922);
xnor UO_1094 (O_1094,N_9939,N_9938);
xnor UO_1095 (O_1095,N_9944,N_9960);
nand UO_1096 (O_1096,N_9944,N_9939);
nor UO_1097 (O_1097,N_9960,N_9971);
or UO_1098 (O_1098,N_9958,N_9927);
nor UO_1099 (O_1099,N_9982,N_9978);
and UO_1100 (O_1100,N_9973,N_9918);
and UO_1101 (O_1101,N_9962,N_9927);
nor UO_1102 (O_1102,N_9993,N_9939);
nand UO_1103 (O_1103,N_9910,N_9915);
and UO_1104 (O_1104,N_9935,N_9976);
and UO_1105 (O_1105,N_9954,N_9945);
or UO_1106 (O_1106,N_9997,N_9951);
nand UO_1107 (O_1107,N_9962,N_9975);
nand UO_1108 (O_1108,N_9967,N_9988);
nor UO_1109 (O_1109,N_9964,N_9985);
nand UO_1110 (O_1110,N_9961,N_9960);
nand UO_1111 (O_1111,N_9930,N_9939);
nand UO_1112 (O_1112,N_9952,N_9912);
nand UO_1113 (O_1113,N_9980,N_9922);
nor UO_1114 (O_1114,N_9939,N_9906);
xor UO_1115 (O_1115,N_9985,N_9949);
nand UO_1116 (O_1116,N_9975,N_9920);
nand UO_1117 (O_1117,N_9928,N_9974);
and UO_1118 (O_1118,N_9964,N_9908);
nand UO_1119 (O_1119,N_9929,N_9973);
nand UO_1120 (O_1120,N_9920,N_9946);
or UO_1121 (O_1121,N_9923,N_9963);
nor UO_1122 (O_1122,N_9948,N_9946);
nor UO_1123 (O_1123,N_9928,N_9963);
nor UO_1124 (O_1124,N_9989,N_9987);
xor UO_1125 (O_1125,N_9938,N_9906);
xnor UO_1126 (O_1126,N_9935,N_9980);
nor UO_1127 (O_1127,N_9904,N_9967);
and UO_1128 (O_1128,N_9907,N_9908);
or UO_1129 (O_1129,N_9918,N_9948);
nand UO_1130 (O_1130,N_9921,N_9985);
and UO_1131 (O_1131,N_9936,N_9990);
nand UO_1132 (O_1132,N_9948,N_9992);
or UO_1133 (O_1133,N_9964,N_9935);
xnor UO_1134 (O_1134,N_9921,N_9940);
or UO_1135 (O_1135,N_9907,N_9995);
nor UO_1136 (O_1136,N_9942,N_9970);
and UO_1137 (O_1137,N_9953,N_9993);
nor UO_1138 (O_1138,N_9927,N_9988);
xor UO_1139 (O_1139,N_9990,N_9966);
xor UO_1140 (O_1140,N_9989,N_9978);
nor UO_1141 (O_1141,N_9971,N_9903);
xnor UO_1142 (O_1142,N_9954,N_9942);
xor UO_1143 (O_1143,N_9944,N_9923);
nand UO_1144 (O_1144,N_9998,N_9913);
xor UO_1145 (O_1145,N_9937,N_9947);
xnor UO_1146 (O_1146,N_9919,N_9943);
or UO_1147 (O_1147,N_9915,N_9978);
nor UO_1148 (O_1148,N_9995,N_9906);
nand UO_1149 (O_1149,N_9914,N_9909);
nand UO_1150 (O_1150,N_9995,N_9925);
nor UO_1151 (O_1151,N_9967,N_9961);
or UO_1152 (O_1152,N_9920,N_9953);
nor UO_1153 (O_1153,N_9991,N_9977);
xnor UO_1154 (O_1154,N_9930,N_9949);
or UO_1155 (O_1155,N_9977,N_9952);
and UO_1156 (O_1156,N_9981,N_9914);
xnor UO_1157 (O_1157,N_9990,N_9943);
nor UO_1158 (O_1158,N_9926,N_9981);
or UO_1159 (O_1159,N_9945,N_9940);
nand UO_1160 (O_1160,N_9927,N_9916);
and UO_1161 (O_1161,N_9993,N_9943);
nand UO_1162 (O_1162,N_9928,N_9946);
nor UO_1163 (O_1163,N_9981,N_9987);
and UO_1164 (O_1164,N_9912,N_9984);
or UO_1165 (O_1165,N_9974,N_9983);
and UO_1166 (O_1166,N_9977,N_9998);
nor UO_1167 (O_1167,N_9989,N_9957);
xnor UO_1168 (O_1168,N_9992,N_9985);
xor UO_1169 (O_1169,N_9959,N_9994);
xor UO_1170 (O_1170,N_9991,N_9964);
nand UO_1171 (O_1171,N_9998,N_9920);
xnor UO_1172 (O_1172,N_9907,N_9940);
nand UO_1173 (O_1173,N_9959,N_9991);
and UO_1174 (O_1174,N_9929,N_9991);
or UO_1175 (O_1175,N_9915,N_9971);
nor UO_1176 (O_1176,N_9950,N_9936);
or UO_1177 (O_1177,N_9922,N_9932);
nor UO_1178 (O_1178,N_9951,N_9973);
or UO_1179 (O_1179,N_9922,N_9918);
xor UO_1180 (O_1180,N_9999,N_9937);
nand UO_1181 (O_1181,N_9968,N_9971);
nor UO_1182 (O_1182,N_9973,N_9906);
or UO_1183 (O_1183,N_9996,N_9998);
or UO_1184 (O_1184,N_9990,N_9941);
nor UO_1185 (O_1185,N_9912,N_9991);
nor UO_1186 (O_1186,N_9971,N_9941);
xor UO_1187 (O_1187,N_9962,N_9976);
nor UO_1188 (O_1188,N_9938,N_9929);
or UO_1189 (O_1189,N_9969,N_9921);
or UO_1190 (O_1190,N_9936,N_9955);
xnor UO_1191 (O_1191,N_9932,N_9918);
xnor UO_1192 (O_1192,N_9914,N_9962);
and UO_1193 (O_1193,N_9969,N_9930);
nand UO_1194 (O_1194,N_9900,N_9911);
nor UO_1195 (O_1195,N_9923,N_9986);
or UO_1196 (O_1196,N_9986,N_9958);
or UO_1197 (O_1197,N_9987,N_9906);
xor UO_1198 (O_1198,N_9918,N_9974);
and UO_1199 (O_1199,N_9990,N_9908);
nand UO_1200 (O_1200,N_9974,N_9978);
nand UO_1201 (O_1201,N_9930,N_9950);
and UO_1202 (O_1202,N_9958,N_9933);
nor UO_1203 (O_1203,N_9967,N_9984);
or UO_1204 (O_1204,N_9966,N_9935);
nand UO_1205 (O_1205,N_9922,N_9944);
nand UO_1206 (O_1206,N_9994,N_9914);
or UO_1207 (O_1207,N_9962,N_9957);
nor UO_1208 (O_1208,N_9956,N_9942);
nand UO_1209 (O_1209,N_9910,N_9995);
and UO_1210 (O_1210,N_9987,N_9967);
xnor UO_1211 (O_1211,N_9981,N_9967);
xnor UO_1212 (O_1212,N_9921,N_9923);
nor UO_1213 (O_1213,N_9991,N_9949);
nand UO_1214 (O_1214,N_9937,N_9978);
nand UO_1215 (O_1215,N_9956,N_9944);
nor UO_1216 (O_1216,N_9956,N_9948);
nand UO_1217 (O_1217,N_9999,N_9932);
nor UO_1218 (O_1218,N_9994,N_9907);
nor UO_1219 (O_1219,N_9913,N_9924);
or UO_1220 (O_1220,N_9918,N_9903);
nor UO_1221 (O_1221,N_9937,N_9951);
and UO_1222 (O_1222,N_9968,N_9999);
or UO_1223 (O_1223,N_9987,N_9937);
or UO_1224 (O_1224,N_9986,N_9995);
xnor UO_1225 (O_1225,N_9907,N_9913);
nand UO_1226 (O_1226,N_9909,N_9912);
and UO_1227 (O_1227,N_9908,N_9954);
xnor UO_1228 (O_1228,N_9998,N_9964);
xor UO_1229 (O_1229,N_9935,N_9908);
nand UO_1230 (O_1230,N_9946,N_9922);
or UO_1231 (O_1231,N_9976,N_9966);
and UO_1232 (O_1232,N_9971,N_9994);
and UO_1233 (O_1233,N_9915,N_9987);
xor UO_1234 (O_1234,N_9986,N_9952);
or UO_1235 (O_1235,N_9951,N_9947);
nand UO_1236 (O_1236,N_9965,N_9954);
or UO_1237 (O_1237,N_9949,N_9948);
xor UO_1238 (O_1238,N_9944,N_9921);
and UO_1239 (O_1239,N_9990,N_9938);
xnor UO_1240 (O_1240,N_9990,N_9949);
or UO_1241 (O_1241,N_9982,N_9950);
nand UO_1242 (O_1242,N_9985,N_9946);
nor UO_1243 (O_1243,N_9952,N_9904);
nand UO_1244 (O_1244,N_9965,N_9920);
or UO_1245 (O_1245,N_9980,N_9990);
xor UO_1246 (O_1246,N_9998,N_9939);
nor UO_1247 (O_1247,N_9921,N_9979);
xor UO_1248 (O_1248,N_9939,N_9947);
xnor UO_1249 (O_1249,N_9911,N_9999);
or UO_1250 (O_1250,N_9922,N_9985);
xor UO_1251 (O_1251,N_9927,N_9992);
nand UO_1252 (O_1252,N_9978,N_9931);
nand UO_1253 (O_1253,N_9986,N_9936);
xor UO_1254 (O_1254,N_9930,N_9989);
and UO_1255 (O_1255,N_9944,N_9927);
xor UO_1256 (O_1256,N_9994,N_9923);
nand UO_1257 (O_1257,N_9907,N_9996);
nand UO_1258 (O_1258,N_9922,N_9937);
xnor UO_1259 (O_1259,N_9983,N_9938);
xnor UO_1260 (O_1260,N_9973,N_9993);
nor UO_1261 (O_1261,N_9936,N_9952);
xnor UO_1262 (O_1262,N_9913,N_9959);
nor UO_1263 (O_1263,N_9979,N_9989);
nand UO_1264 (O_1264,N_9949,N_9962);
or UO_1265 (O_1265,N_9904,N_9984);
nand UO_1266 (O_1266,N_9925,N_9909);
nor UO_1267 (O_1267,N_9929,N_9985);
nand UO_1268 (O_1268,N_9983,N_9966);
and UO_1269 (O_1269,N_9975,N_9995);
nor UO_1270 (O_1270,N_9904,N_9933);
nor UO_1271 (O_1271,N_9996,N_9900);
and UO_1272 (O_1272,N_9902,N_9921);
nor UO_1273 (O_1273,N_9982,N_9954);
or UO_1274 (O_1274,N_9918,N_9934);
and UO_1275 (O_1275,N_9967,N_9920);
and UO_1276 (O_1276,N_9941,N_9907);
xor UO_1277 (O_1277,N_9999,N_9949);
nand UO_1278 (O_1278,N_9976,N_9905);
nand UO_1279 (O_1279,N_9932,N_9900);
xnor UO_1280 (O_1280,N_9988,N_9987);
or UO_1281 (O_1281,N_9964,N_9983);
and UO_1282 (O_1282,N_9927,N_9973);
xnor UO_1283 (O_1283,N_9958,N_9909);
and UO_1284 (O_1284,N_9990,N_9909);
nand UO_1285 (O_1285,N_9945,N_9912);
or UO_1286 (O_1286,N_9942,N_9902);
nor UO_1287 (O_1287,N_9945,N_9931);
nand UO_1288 (O_1288,N_9980,N_9974);
nor UO_1289 (O_1289,N_9976,N_9907);
nand UO_1290 (O_1290,N_9907,N_9932);
or UO_1291 (O_1291,N_9997,N_9913);
or UO_1292 (O_1292,N_9913,N_9968);
xor UO_1293 (O_1293,N_9908,N_9952);
or UO_1294 (O_1294,N_9974,N_9960);
nand UO_1295 (O_1295,N_9901,N_9954);
nor UO_1296 (O_1296,N_9974,N_9923);
and UO_1297 (O_1297,N_9902,N_9926);
nand UO_1298 (O_1298,N_9973,N_9998);
nor UO_1299 (O_1299,N_9981,N_9948);
nor UO_1300 (O_1300,N_9931,N_9934);
and UO_1301 (O_1301,N_9935,N_9917);
and UO_1302 (O_1302,N_9910,N_9966);
or UO_1303 (O_1303,N_9982,N_9975);
nor UO_1304 (O_1304,N_9933,N_9953);
xnor UO_1305 (O_1305,N_9939,N_9942);
nand UO_1306 (O_1306,N_9968,N_9936);
and UO_1307 (O_1307,N_9927,N_9908);
nand UO_1308 (O_1308,N_9978,N_9957);
nor UO_1309 (O_1309,N_9953,N_9955);
nor UO_1310 (O_1310,N_9958,N_9955);
nand UO_1311 (O_1311,N_9973,N_9940);
nor UO_1312 (O_1312,N_9932,N_9939);
or UO_1313 (O_1313,N_9977,N_9901);
and UO_1314 (O_1314,N_9903,N_9951);
or UO_1315 (O_1315,N_9924,N_9981);
xnor UO_1316 (O_1316,N_9979,N_9916);
or UO_1317 (O_1317,N_9971,N_9966);
or UO_1318 (O_1318,N_9952,N_9972);
xor UO_1319 (O_1319,N_9987,N_9938);
nor UO_1320 (O_1320,N_9904,N_9996);
nand UO_1321 (O_1321,N_9987,N_9993);
xor UO_1322 (O_1322,N_9993,N_9978);
nor UO_1323 (O_1323,N_9968,N_9941);
nor UO_1324 (O_1324,N_9997,N_9907);
nor UO_1325 (O_1325,N_9994,N_9915);
nand UO_1326 (O_1326,N_9984,N_9968);
nor UO_1327 (O_1327,N_9961,N_9969);
nor UO_1328 (O_1328,N_9973,N_9937);
and UO_1329 (O_1329,N_9938,N_9992);
and UO_1330 (O_1330,N_9960,N_9939);
nand UO_1331 (O_1331,N_9970,N_9959);
nand UO_1332 (O_1332,N_9911,N_9973);
nand UO_1333 (O_1333,N_9957,N_9903);
and UO_1334 (O_1334,N_9903,N_9963);
nor UO_1335 (O_1335,N_9984,N_9972);
and UO_1336 (O_1336,N_9914,N_9969);
nand UO_1337 (O_1337,N_9953,N_9978);
nor UO_1338 (O_1338,N_9920,N_9907);
nand UO_1339 (O_1339,N_9971,N_9925);
and UO_1340 (O_1340,N_9905,N_9999);
and UO_1341 (O_1341,N_9978,N_9979);
nand UO_1342 (O_1342,N_9922,N_9976);
nor UO_1343 (O_1343,N_9962,N_9921);
nand UO_1344 (O_1344,N_9910,N_9982);
and UO_1345 (O_1345,N_9929,N_9965);
nor UO_1346 (O_1346,N_9912,N_9943);
or UO_1347 (O_1347,N_9947,N_9900);
and UO_1348 (O_1348,N_9963,N_9925);
xnor UO_1349 (O_1349,N_9929,N_9904);
and UO_1350 (O_1350,N_9983,N_9902);
and UO_1351 (O_1351,N_9968,N_9985);
or UO_1352 (O_1352,N_9926,N_9946);
nor UO_1353 (O_1353,N_9902,N_9971);
xor UO_1354 (O_1354,N_9936,N_9945);
or UO_1355 (O_1355,N_9953,N_9977);
nand UO_1356 (O_1356,N_9920,N_9940);
nor UO_1357 (O_1357,N_9952,N_9902);
nor UO_1358 (O_1358,N_9992,N_9986);
xnor UO_1359 (O_1359,N_9993,N_9970);
xor UO_1360 (O_1360,N_9911,N_9905);
or UO_1361 (O_1361,N_9970,N_9934);
nor UO_1362 (O_1362,N_9953,N_9961);
nand UO_1363 (O_1363,N_9992,N_9933);
nor UO_1364 (O_1364,N_9979,N_9926);
xnor UO_1365 (O_1365,N_9992,N_9984);
or UO_1366 (O_1366,N_9938,N_9944);
nor UO_1367 (O_1367,N_9995,N_9900);
xnor UO_1368 (O_1368,N_9999,N_9993);
nor UO_1369 (O_1369,N_9908,N_9943);
and UO_1370 (O_1370,N_9994,N_9942);
or UO_1371 (O_1371,N_9949,N_9939);
or UO_1372 (O_1372,N_9971,N_9989);
nor UO_1373 (O_1373,N_9969,N_9951);
nor UO_1374 (O_1374,N_9986,N_9944);
nand UO_1375 (O_1375,N_9920,N_9996);
and UO_1376 (O_1376,N_9974,N_9943);
nand UO_1377 (O_1377,N_9932,N_9994);
nand UO_1378 (O_1378,N_9940,N_9928);
nand UO_1379 (O_1379,N_9901,N_9992);
or UO_1380 (O_1380,N_9933,N_9946);
nand UO_1381 (O_1381,N_9954,N_9976);
or UO_1382 (O_1382,N_9939,N_9984);
nand UO_1383 (O_1383,N_9901,N_9979);
or UO_1384 (O_1384,N_9918,N_9978);
or UO_1385 (O_1385,N_9907,N_9954);
nand UO_1386 (O_1386,N_9927,N_9900);
nor UO_1387 (O_1387,N_9967,N_9940);
nor UO_1388 (O_1388,N_9977,N_9996);
nand UO_1389 (O_1389,N_9931,N_9984);
nand UO_1390 (O_1390,N_9990,N_9979);
nor UO_1391 (O_1391,N_9964,N_9917);
or UO_1392 (O_1392,N_9976,N_9991);
xor UO_1393 (O_1393,N_9923,N_9920);
and UO_1394 (O_1394,N_9920,N_9949);
or UO_1395 (O_1395,N_9960,N_9923);
and UO_1396 (O_1396,N_9969,N_9957);
nand UO_1397 (O_1397,N_9934,N_9950);
or UO_1398 (O_1398,N_9977,N_9990);
nor UO_1399 (O_1399,N_9952,N_9920);
or UO_1400 (O_1400,N_9979,N_9981);
and UO_1401 (O_1401,N_9985,N_9915);
nand UO_1402 (O_1402,N_9976,N_9921);
xnor UO_1403 (O_1403,N_9964,N_9996);
nor UO_1404 (O_1404,N_9960,N_9919);
or UO_1405 (O_1405,N_9965,N_9995);
nor UO_1406 (O_1406,N_9908,N_9989);
xor UO_1407 (O_1407,N_9968,N_9922);
nor UO_1408 (O_1408,N_9992,N_9952);
nand UO_1409 (O_1409,N_9910,N_9934);
nor UO_1410 (O_1410,N_9990,N_9901);
nand UO_1411 (O_1411,N_9977,N_9921);
or UO_1412 (O_1412,N_9928,N_9931);
and UO_1413 (O_1413,N_9961,N_9919);
nand UO_1414 (O_1414,N_9921,N_9905);
and UO_1415 (O_1415,N_9968,N_9917);
and UO_1416 (O_1416,N_9928,N_9970);
xnor UO_1417 (O_1417,N_9901,N_9924);
nand UO_1418 (O_1418,N_9946,N_9983);
and UO_1419 (O_1419,N_9948,N_9959);
nand UO_1420 (O_1420,N_9969,N_9942);
nand UO_1421 (O_1421,N_9986,N_9927);
and UO_1422 (O_1422,N_9936,N_9976);
xnor UO_1423 (O_1423,N_9918,N_9915);
xor UO_1424 (O_1424,N_9959,N_9973);
nand UO_1425 (O_1425,N_9917,N_9938);
and UO_1426 (O_1426,N_9969,N_9902);
nand UO_1427 (O_1427,N_9954,N_9913);
nand UO_1428 (O_1428,N_9946,N_9915);
nand UO_1429 (O_1429,N_9951,N_9943);
or UO_1430 (O_1430,N_9904,N_9971);
or UO_1431 (O_1431,N_9994,N_9968);
and UO_1432 (O_1432,N_9950,N_9940);
or UO_1433 (O_1433,N_9939,N_9965);
xnor UO_1434 (O_1434,N_9966,N_9945);
nand UO_1435 (O_1435,N_9925,N_9953);
and UO_1436 (O_1436,N_9998,N_9930);
nor UO_1437 (O_1437,N_9945,N_9990);
nor UO_1438 (O_1438,N_9935,N_9918);
xnor UO_1439 (O_1439,N_9920,N_9921);
nand UO_1440 (O_1440,N_9962,N_9926);
nor UO_1441 (O_1441,N_9941,N_9989);
or UO_1442 (O_1442,N_9900,N_9985);
xnor UO_1443 (O_1443,N_9946,N_9997);
nor UO_1444 (O_1444,N_9926,N_9987);
and UO_1445 (O_1445,N_9959,N_9966);
or UO_1446 (O_1446,N_9997,N_9968);
xor UO_1447 (O_1447,N_9919,N_9951);
or UO_1448 (O_1448,N_9909,N_9955);
nand UO_1449 (O_1449,N_9982,N_9930);
nor UO_1450 (O_1450,N_9996,N_9932);
xor UO_1451 (O_1451,N_9921,N_9999);
nand UO_1452 (O_1452,N_9976,N_9917);
nand UO_1453 (O_1453,N_9950,N_9970);
nand UO_1454 (O_1454,N_9929,N_9919);
xor UO_1455 (O_1455,N_9959,N_9918);
and UO_1456 (O_1456,N_9942,N_9966);
nor UO_1457 (O_1457,N_9995,N_9967);
and UO_1458 (O_1458,N_9981,N_9999);
xor UO_1459 (O_1459,N_9960,N_9980);
nand UO_1460 (O_1460,N_9976,N_9968);
xnor UO_1461 (O_1461,N_9980,N_9914);
nor UO_1462 (O_1462,N_9945,N_9961);
xnor UO_1463 (O_1463,N_9983,N_9980);
nor UO_1464 (O_1464,N_9901,N_9960);
or UO_1465 (O_1465,N_9900,N_9931);
and UO_1466 (O_1466,N_9910,N_9978);
xnor UO_1467 (O_1467,N_9987,N_9916);
or UO_1468 (O_1468,N_9967,N_9911);
and UO_1469 (O_1469,N_9977,N_9963);
or UO_1470 (O_1470,N_9910,N_9928);
or UO_1471 (O_1471,N_9933,N_9919);
xor UO_1472 (O_1472,N_9921,N_9924);
nand UO_1473 (O_1473,N_9932,N_9909);
or UO_1474 (O_1474,N_9925,N_9935);
nand UO_1475 (O_1475,N_9991,N_9919);
and UO_1476 (O_1476,N_9960,N_9985);
or UO_1477 (O_1477,N_9958,N_9913);
and UO_1478 (O_1478,N_9989,N_9966);
and UO_1479 (O_1479,N_9910,N_9988);
or UO_1480 (O_1480,N_9956,N_9917);
nand UO_1481 (O_1481,N_9994,N_9955);
xnor UO_1482 (O_1482,N_9967,N_9976);
nand UO_1483 (O_1483,N_9927,N_9997);
and UO_1484 (O_1484,N_9955,N_9923);
xor UO_1485 (O_1485,N_9963,N_9904);
or UO_1486 (O_1486,N_9914,N_9983);
xor UO_1487 (O_1487,N_9904,N_9902);
nand UO_1488 (O_1488,N_9974,N_9905);
xnor UO_1489 (O_1489,N_9937,N_9917);
and UO_1490 (O_1490,N_9992,N_9917);
nor UO_1491 (O_1491,N_9920,N_9978);
or UO_1492 (O_1492,N_9970,N_9949);
nand UO_1493 (O_1493,N_9914,N_9977);
and UO_1494 (O_1494,N_9905,N_9996);
and UO_1495 (O_1495,N_9995,N_9940);
nor UO_1496 (O_1496,N_9979,N_9909);
nor UO_1497 (O_1497,N_9931,N_9930);
xnor UO_1498 (O_1498,N_9986,N_9904);
xnor UO_1499 (O_1499,N_9963,N_9994);
endmodule