module basic_1500_15000_2000_10_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_1301,In_820);
or U1 (N_1,In_628,In_1222);
or U2 (N_2,In_1152,In_9);
xor U3 (N_3,In_1199,In_1292);
nor U4 (N_4,In_239,In_1440);
and U5 (N_5,In_616,In_482);
xnor U6 (N_6,In_362,In_1089);
nand U7 (N_7,In_739,In_161);
and U8 (N_8,In_1155,In_887);
xnor U9 (N_9,In_311,In_941);
nor U10 (N_10,In_1165,In_1285);
nand U11 (N_11,In_814,In_1101);
nand U12 (N_12,In_1184,In_1499);
or U13 (N_13,In_1493,In_1200);
or U14 (N_14,In_787,In_590);
and U15 (N_15,In_1486,In_1489);
and U16 (N_16,In_782,In_217);
nor U17 (N_17,In_699,In_1314);
xor U18 (N_18,In_421,In_519);
nor U19 (N_19,In_532,In_1176);
nand U20 (N_20,In_1462,In_1298);
nand U21 (N_21,In_642,In_911);
and U22 (N_22,In_412,In_526);
xor U23 (N_23,In_1013,In_181);
or U24 (N_24,In_818,In_1276);
nand U25 (N_25,In_821,In_729);
nor U26 (N_26,In_1198,In_811);
and U27 (N_27,In_1123,In_518);
nand U28 (N_28,In_543,In_1179);
nor U29 (N_29,In_393,In_1208);
or U30 (N_30,In_120,In_149);
and U31 (N_31,In_1379,In_358);
or U32 (N_32,In_7,In_1187);
nor U33 (N_33,In_115,In_420);
nor U34 (N_34,In_755,In_446);
or U35 (N_35,In_418,In_512);
nor U36 (N_36,In_1017,In_551);
xnor U37 (N_37,In_1269,In_944);
or U38 (N_38,In_1359,In_364);
nand U39 (N_39,In_1289,In_647);
nor U40 (N_40,In_1307,In_277);
or U41 (N_41,In_188,In_14);
and U42 (N_42,In_688,In_1175);
nor U43 (N_43,In_874,In_1043);
and U44 (N_44,In_338,In_1401);
nor U45 (N_45,In_506,In_803);
nand U46 (N_46,In_806,In_654);
nor U47 (N_47,In_243,In_389);
nand U48 (N_48,In_842,In_67);
nand U49 (N_49,In_17,In_232);
nor U50 (N_50,In_223,In_841);
nand U51 (N_51,In_1044,In_305);
and U52 (N_52,In_744,In_658);
or U53 (N_53,In_1052,In_1386);
nand U54 (N_54,In_1480,In_585);
nor U55 (N_55,In_676,In_1116);
nand U56 (N_56,In_423,In_308);
and U57 (N_57,In_839,In_1069);
nor U58 (N_58,In_296,In_269);
or U59 (N_59,In_380,In_948);
and U60 (N_60,In_1470,In_1164);
or U61 (N_61,In_1231,In_973);
nand U62 (N_62,In_465,In_721);
or U63 (N_63,In_1374,In_934);
xnor U64 (N_64,In_21,In_609);
nand U65 (N_65,In_582,In_703);
and U66 (N_66,In_187,In_580);
nor U67 (N_67,In_52,In_772);
and U68 (N_68,In_660,In_317);
nor U69 (N_69,In_480,In_1243);
or U70 (N_70,In_817,In_1111);
or U71 (N_71,In_1346,In_13);
or U72 (N_72,In_159,In_606);
or U73 (N_73,In_1084,In_527);
nand U74 (N_74,In_1079,In_765);
or U75 (N_75,In_1065,In_35);
or U76 (N_76,In_1206,In_6);
nor U77 (N_77,In_1425,In_1355);
nand U78 (N_78,In_1191,In_978);
or U79 (N_79,In_1186,In_1154);
nand U80 (N_80,In_597,In_466);
or U81 (N_81,In_348,In_877);
nor U82 (N_82,In_1118,In_865);
nor U83 (N_83,In_1254,In_454);
xor U84 (N_84,In_1145,In_1059);
or U85 (N_85,In_139,In_1410);
nand U86 (N_86,In_1082,In_1037);
nor U87 (N_87,In_185,In_1136);
nand U88 (N_88,In_1189,In_176);
or U89 (N_89,In_146,In_416);
nand U90 (N_90,In_241,In_1467);
nand U91 (N_91,In_550,In_411);
xnor U92 (N_92,In_426,In_233);
or U93 (N_93,In_205,In_212);
nand U94 (N_94,In_991,In_1125);
nor U95 (N_95,In_867,In_838);
or U96 (N_96,In_124,In_754);
and U97 (N_97,In_1441,In_180);
nand U98 (N_98,In_912,In_963);
or U99 (N_99,In_1146,In_1034);
or U100 (N_100,In_1324,In_1361);
nor U101 (N_101,In_468,In_975);
and U102 (N_102,In_336,In_1005);
or U103 (N_103,In_1063,In_123);
and U104 (N_104,In_538,In_516);
or U105 (N_105,In_164,In_409);
and U106 (N_106,In_278,In_1287);
nor U107 (N_107,In_1453,In_1102);
nor U108 (N_108,In_780,In_1469);
xnor U109 (N_109,In_671,In_1029);
nor U110 (N_110,In_113,In_1259);
xnor U111 (N_111,In_273,In_111);
xnor U112 (N_112,In_990,In_1099);
nand U113 (N_113,In_249,In_96);
or U114 (N_114,In_1087,In_491);
nand U115 (N_115,In_881,In_1150);
nand U116 (N_116,In_927,In_75);
nand U117 (N_117,In_715,In_899);
nand U118 (N_118,In_318,In_596);
and U119 (N_119,In_1336,In_783);
or U120 (N_120,In_982,In_352);
or U121 (N_121,In_496,In_1422);
and U122 (N_122,In_425,In_1140);
or U123 (N_123,In_987,In_165);
nand U124 (N_124,In_1246,In_464);
and U125 (N_125,In_28,In_622);
nand U126 (N_126,In_377,In_697);
or U127 (N_127,In_835,In_327);
nand U128 (N_128,In_663,In_222);
nor U129 (N_129,In_1487,In_826);
nor U130 (N_130,In_434,In_1076);
xnor U131 (N_131,In_231,In_404);
or U132 (N_132,In_333,In_186);
nor U133 (N_133,In_369,In_134);
nor U134 (N_134,In_1394,In_225);
xnor U135 (N_135,In_873,In_1390);
or U136 (N_136,In_895,In_1098);
or U137 (N_137,In_350,In_335);
and U138 (N_138,In_1117,In_695);
and U139 (N_139,In_626,In_353);
nand U140 (N_140,In_769,In_1383);
and U141 (N_141,In_70,In_716);
and U142 (N_142,In_966,In_1448);
xor U143 (N_143,In_455,In_1442);
nand U144 (N_144,In_923,In_145);
nor U145 (N_145,In_11,In_786);
nor U146 (N_146,In_177,In_756);
nand U147 (N_147,In_1053,In_1077);
and U148 (N_148,In_796,In_447);
nor U149 (N_149,In_1270,In_1153);
or U150 (N_150,In_85,In_517);
xnor U151 (N_151,In_275,In_50);
and U152 (N_152,In_1400,In_90);
and U153 (N_153,In_727,In_552);
and U154 (N_154,In_690,In_1284);
and U155 (N_155,In_984,In_725);
nor U156 (N_156,In_375,In_1419);
nand U157 (N_157,In_515,In_1327);
or U158 (N_158,In_40,In_629);
xnor U159 (N_159,In_649,In_809);
nand U160 (N_160,In_386,In_199);
or U161 (N_161,In_789,In_299);
nor U162 (N_162,In_732,In_957);
and U163 (N_163,In_1347,In_870);
or U164 (N_164,In_23,In_1466);
nor U165 (N_165,In_940,In_121);
nor U166 (N_166,In_1315,In_1388);
and U167 (N_167,In_371,In_861);
and U168 (N_168,In_497,In_1064);
and U169 (N_169,In_652,In_36);
and U170 (N_170,In_1478,In_80);
nor U171 (N_171,In_977,In_160);
and U172 (N_172,In_1423,In_972);
nand U173 (N_173,In_356,In_1332);
nor U174 (N_174,In_900,In_1134);
nand U175 (N_175,In_200,In_326);
and U176 (N_176,In_288,In_860);
nor U177 (N_177,In_938,In_1039);
or U178 (N_178,In_508,In_791);
nor U179 (N_179,In_1326,In_8);
and U180 (N_180,In_397,In_960);
xor U181 (N_181,In_1148,In_1119);
or U182 (N_182,In_875,In_445);
xnor U183 (N_183,In_1011,In_1003);
xnor U184 (N_184,In_757,In_933);
or U185 (N_185,In_565,In_1278);
and U186 (N_186,In_1072,In_1429);
or U187 (N_187,In_293,In_1216);
or U188 (N_188,In_41,In_469);
and U189 (N_189,In_129,In_1433);
or U190 (N_190,In_687,In_436);
or U191 (N_191,In_829,In_1370);
xor U192 (N_192,In_993,In_15);
and U193 (N_193,In_728,In_584);
nand U194 (N_194,In_66,In_254);
nand U195 (N_195,In_1248,In_1245);
or U196 (N_196,In_1019,In_1348);
xnor U197 (N_197,In_1073,In_1086);
nand U198 (N_198,In_31,In_560);
or U199 (N_199,In_827,In_1190);
or U200 (N_200,In_674,In_534);
xnor U201 (N_201,In_73,In_19);
or U202 (N_202,In_184,In_471);
nand U203 (N_203,In_605,In_578);
nor U204 (N_204,In_1350,In_271);
nor U205 (N_205,In_921,In_89);
xnor U206 (N_206,In_1445,In_1223);
or U207 (N_207,In_1295,In_272);
or U208 (N_208,In_1294,In_481);
or U209 (N_209,In_167,In_1311);
nor U210 (N_210,In_905,In_183);
xor U211 (N_211,In_1300,In_1413);
nor U212 (N_212,In_300,In_234);
or U213 (N_213,In_825,In_410);
or U214 (N_214,In_935,In_1051);
nand U215 (N_215,In_888,In_920);
nor U216 (N_216,In_156,In_1396);
nor U217 (N_217,In_850,In_1282);
or U218 (N_218,In_1364,In_1468);
and U219 (N_219,In_1058,In_268);
nor U220 (N_220,In_286,In_1427);
xor U221 (N_221,In_78,In_1337);
nor U222 (N_222,In_1219,In_673);
or U223 (N_223,In_717,In_1021);
and U224 (N_224,In_1430,In_114);
or U225 (N_225,In_1320,In_1022);
nor U226 (N_226,In_489,In_545);
or U227 (N_227,In_1497,In_1351);
or U228 (N_228,In_880,In_1060);
and U229 (N_229,In_214,In_325);
nand U230 (N_230,In_1121,In_747);
nand U231 (N_231,In_637,In_132);
or U232 (N_232,In_857,In_1461);
or U233 (N_233,In_346,In_202);
and U234 (N_234,In_247,In_97);
or U235 (N_235,In_492,In_633);
nor U236 (N_236,In_315,In_262);
and U237 (N_237,In_967,In_235);
and U238 (N_238,In_292,In_986);
nor U239 (N_239,In_1014,In_166);
nor U240 (N_240,In_1403,In_1023);
and U241 (N_241,In_953,In_979);
nor U242 (N_242,In_730,In_112);
nand U243 (N_243,In_60,In_504);
and U244 (N_244,In_891,In_1109);
nand U245 (N_245,In_619,In_567);
xor U246 (N_246,In_1090,In_102);
xor U247 (N_247,In_1103,In_258);
nor U248 (N_248,In_854,In_558);
nor U249 (N_249,In_540,In_44);
and U250 (N_250,In_1291,In_1047);
nor U251 (N_251,In_890,In_54);
and U252 (N_252,In_1180,In_1074);
or U253 (N_253,In_639,In_12);
and U254 (N_254,In_726,In_408);
and U255 (N_255,In_896,In_163);
and U256 (N_256,In_705,In_86);
nand U257 (N_257,In_1001,In_1352);
xnor U258 (N_258,In_301,In_1450);
and U259 (N_259,In_1368,In_270);
nor U260 (N_260,In_204,In_1197);
or U261 (N_261,In_949,In_1166);
nor U262 (N_262,In_995,In_541);
nand U263 (N_263,In_926,In_1476);
or U264 (N_264,In_255,In_1473);
or U265 (N_265,In_678,In_141);
nand U266 (N_266,In_1272,In_1159);
nand U267 (N_267,In_903,In_1369);
nor U268 (N_268,In_345,In_707);
nor U269 (N_269,In_1345,In_10);
and U270 (N_270,In_1033,In_1308);
nor U271 (N_271,In_475,In_1066);
nand U272 (N_272,In_250,In_452);
and U273 (N_273,In_670,In_98);
and U274 (N_274,In_367,In_1397);
and U275 (N_275,In_844,In_368);
and U276 (N_276,In_65,In_1096);
nor U277 (N_277,In_1088,In_1215);
nor U278 (N_278,In_474,In_513);
and U279 (N_279,In_1083,In_287);
nor U280 (N_280,In_897,In_357);
nor U281 (N_281,In_1411,In_1085);
nor U282 (N_282,In_1274,In_980);
and U283 (N_283,In_81,In_441);
xor U284 (N_284,In_1267,In_523);
xnor U285 (N_285,In_1207,In_958);
and U286 (N_286,In_55,In_61);
and U287 (N_287,In_974,In_1229);
or U288 (N_288,In_321,In_470);
or U289 (N_289,In_1490,In_555);
nor U290 (N_290,In_804,In_1457);
nand U291 (N_291,In_1151,In_38);
nor U292 (N_292,In_240,In_1233);
nand U293 (N_293,In_63,In_313);
and U294 (N_294,In_1218,In_383);
nor U295 (N_295,In_463,In_1035);
or U296 (N_296,In_432,In_1363);
nor U297 (N_297,In_443,In_1196);
xnor U298 (N_298,In_88,In_599);
nand U299 (N_299,In_686,In_1234);
nand U300 (N_300,In_1256,In_947);
and U301 (N_301,In_1168,In_856);
or U302 (N_302,In_908,In_117);
nor U303 (N_303,In_1288,In_810);
xnor U304 (N_304,In_939,In_328);
nand U305 (N_305,In_1177,In_151);
or U306 (N_306,In_1050,In_193);
nor U307 (N_307,In_1237,In_125);
or U308 (N_308,In_442,In_433);
nand U309 (N_309,In_749,In_138);
xnor U310 (N_310,In_562,In_531);
nand U311 (N_311,In_266,In_501);
nor U312 (N_312,In_689,In_407);
nand U313 (N_313,In_1142,In_467);
nor U314 (N_314,In_1031,In_107);
nor U315 (N_315,In_901,In_487);
nor U316 (N_316,In_1,In_713);
or U317 (N_317,In_220,In_698);
nor U318 (N_318,In_849,In_430);
nor U319 (N_319,In_1451,In_680);
nor U320 (N_320,In_1230,In_219);
nand U321 (N_321,In_359,In_221);
or U322 (N_322,In_595,In_1178);
xor U323 (N_323,In_57,In_1008);
nand U324 (N_324,In_909,In_274);
or U325 (N_325,In_962,In_158);
nand U326 (N_326,In_51,In_1439);
nor U327 (N_327,In_365,In_1204);
nor U328 (N_328,In_312,In_1431);
nor U329 (N_329,In_495,In_845);
nor U330 (N_330,In_290,In_691);
or U331 (N_331,In_770,In_675);
nand U332 (N_332,In_319,In_1414);
or U333 (N_333,In_795,In_1316);
and U334 (N_334,In_1376,In_1362);
or U335 (N_335,In_1263,In_602);
and U336 (N_336,In_655,In_440);
or U337 (N_337,In_1126,In_510);
nand U338 (N_338,In_363,In_737);
nor U339 (N_339,In_893,In_322);
and U340 (N_340,In_1262,In_238);
and U341 (N_341,In_871,In_946);
and U342 (N_342,In_704,In_591);
nor U343 (N_343,In_307,In_1193);
xor U344 (N_344,In_1062,In_417);
nand U345 (N_345,In_280,In_405);
and U346 (N_346,In_1036,In_1471);
nor U347 (N_347,In_265,In_1238);
or U348 (N_348,In_1139,In_1106);
and U349 (N_349,In_836,In_1436);
and U350 (N_350,In_916,In_997);
or U351 (N_351,In_521,In_583);
and U352 (N_352,In_625,In_477);
nor U353 (N_353,In_1054,In_195);
and U354 (N_354,In_1426,In_323);
nor U355 (N_355,In_1365,In_910);
nor U356 (N_356,In_883,In_1214);
or U357 (N_357,In_714,In_24);
nand U358 (N_358,In_734,In_776);
nand U359 (N_359,In_959,In_969);
or U360 (N_360,In_1286,In_279);
and U361 (N_361,In_1349,In_589);
and U362 (N_362,In_812,In_906);
nand U363 (N_363,In_1172,In_1041);
xnor U364 (N_364,In_1163,In_1183);
nand U365 (N_365,In_104,In_840);
xor U366 (N_366,In_485,In_372);
nand U367 (N_367,In_556,In_1016);
and U368 (N_368,In_502,In_246);
or U369 (N_369,In_33,In_257);
and U370 (N_370,In_396,In_788);
and U371 (N_371,In_415,In_1241);
nand U372 (N_372,In_878,In_473);
nand U373 (N_373,In_722,In_1167);
nor U374 (N_374,In_1402,In_1078);
or U375 (N_375,In_331,In_53);
xnor U376 (N_376,In_661,In_864);
nand U377 (N_377,In_168,In_1158);
nand U378 (N_378,In_1244,In_520);
nand U379 (N_379,In_1143,In_101);
nor U380 (N_380,In_1202,In_344);
or U381 (N_381,In_1484,In_267);
or U382 (N_382,In_42,In_402);
or U383 (N_383,In_641,In_1275);
nor U384 (N_384,In_931,In_922);
nor U385 (N_385,In_1201,In_347);
or U386 (N_386,In_656,In_1366);
nand U387 (N_387,In_914,In_745);
or U388 (N_388,In_354,In_1339);
and U389 (N_389,In_1104,In_1306);
and U390 (N_390,In_612,In_457);
xnor U391 (N_391,In_1344,In_1067);
or U392 (N_392,In_621,In_581);
nor U393 (N_393,In_529,In_610);
or U394 (N_394,In_808,In_572);
xor U395 (N_395,In_259,In_179);
and U396 (N_396,In_95,In_724);
nand U397 (N_397,In_1325,In_741);
nand U398 (N_398,In_1299,In_1107);
nand U399 (N_399,In_1080,In_700);
nor U400 (N_400,In_965,In_1387);
nor U401 (N_401,In_828,In_570);
nor U402 (N_402,In_1373,In_1252);
nor U403 (N_403,In_1113,In_69);
and U404 (N_404,In_453,In_892);
or U405 (N_405,In_968,In_1004);
and U406 (N_406,In_1195,In_669);
nand U407 (N_407,In_1182,In_182);
and U408 (N_408,In_197,In_1482);
and U409 (N_409,In_1416,In_767);
or U410 (N_410,In_952,In_150);
and U411 (N_411,In_82,In_108);
nand U412 (N_412,In_711,In_1156);
xor U413 (N_413,In_623,In_1334);
nor U414 (N_414,In_1494,In_1211);
nor U415 (N_415,In_25,In_133);
and U416 (N_416,In_748,In_919);
nand U417 (N_417,In_395,In_1412);
nor U418 (N_418,In_553,In_542);
and U419 (N_419,In_252,In_955);
and U420 (N_420,In_1097,In_566);
and U421 (N_421,In_964,In_1105);
nor U422 (N_422,In_937,In_384);
or U423 (N_423,In_731,In_792);
nor U424 (N_424,In_302,In_932);
and U425 (N_425,In_740,In_1112);
nand U426 (N_426,In_1046,In_1188);
or U427 (N_427,In_1372,In_1110);
nand U428 (N_428,In_1015,In_406);
nor U429 (N_429,In_831,In_450);
nand U430 (N_430,In_760,In_853);
nor U431 (N_431,In_904,In_889);
nor U432 (N_432,In_1277,In_46);
nand U433 (N_433,In_500,In_785);
nand U434 (N_434,In_136,In_1273);
and U435 (N_435,In_1405,In_1000);
and U436 (N_436,In_2,In_45);
nand U437 (N_437,In_1319,In_1446);
nor U438 (N_438,In_1157,In_175);
and U439 (N_439,In_1049,In_43);
and U440 (N_440,In_449,In_1173);
or U441 (N_441,In_484,In_366);
or U442 (N_442,In_1463,In_653);
nor U443 (N_443,In_999,In_1456);
nor U444 (N_444,In_1265,In_1389);
nor U445 (N_445,In_340,In_989);
nand U446 (N_446,In_1428,In_1240);
or U447 (N_447,In_458,In_1225);
and U448 (N_448,In_805,In_1024);
and U449 (N_449,In_1149,In_644);
or U450 (N_450,In_832,In_99);
nor U451 (N_451,In_793,In_1266);
nor U452 (N_452,In_208,In_1305);
and U453 (N_453,In_603,In_303);
nand U454 (N_454,In_848,In_781);
or U455 (N_455,In_951,In_211);
or U456 (N_456,In_373,In_846);
and U457 (N_457,In_1010,In_1492);
nand U458 (N_458,In_646,In_1382);
nor U459 (N_459,In_683,In_524);
or U460 (N_460,In_1120,In_1385);
xor U461 (N_461,In_1475,In_1045);
nand U462 (N_462,In_390,In_777);
nor U463 (N_463,In_29,In_1406);
xnor U464 (N_464,In_260,In_563);
nand U465 (N_465,In_68,In_1335);
or U466 (N_466,In_548,In_438);
nand U467 (N_467,In_665,In_169);
and U468 (N_468,In_1253,In_1424);
nand U469 (N_469,In_994,In_1384);
and U470 (N_470,In_1209,In_694);
nor U471 (N_471,In_385,In_74);
or U472 (N_472,In_439,In_284);
nand U473 (N_473,In_456,In_667);
xor U474 (N_474,In_627,In_242);
or U475 (N_475,In_723,In_1210);
nor U476 (N_476,In_224,In_886);
or U477 (N_477,In_763,In_1340);
nor U478 (N_478,In_207,In_378);
nand U479 (N_479,In_925,In_918);
nor U480 (N_480,In_1081,In_588);
xnor U481 (N_481,In_659,In_657);
nand U482 (N_482,In_613,In_666);
and U483 (N_483,In_218,In_110);
nor U484 (N_484,In_882,In_1460);
nand U485 (N_485,In_309,In_636);
and U486 (N_486,In_76,In_720);
nor U487 (N_487,In_64,In_643);
nand U488 (N_488,In_1483,In_264);
and U489 (N_489,In_422,In_1444);
nor U490 (N_490,In_237,In_1393);
or U491 (N_491,In_1212,In_708);
or U492 (N_492,In_775,In_961);
or U493 (N_493,In_762,In_630);
nor U494 (N_494,In_190,In_189);
nor U495 (N_495,In_601,In_798);
nand U496 (N_496,In_894,In_546);
nor U497 (N_497,In_39,In_930);
nand U498 (N_498,In_511,In_1458);
or U499 (N_499,In_928,In_256);
or U500 (N_500,In_876,In_561);
nor U501 (N_501,In_576,In_1459);
or U502 (N_502,In_800,In_1130);
and U503 (N_503,In_30,In_1061);
nor U504 (N_504,In_483,In_1213);
or U505 (N_505,In_823,In_87);
nor U506 (N_506,In_537,In_1114);
and U507 (N_507,In_281,In_607);
xnor U508 (N_508,In_1357,In_761);
xor U509 (N_509,In_1137,In_1268);
nor U510 (N_510,In_153,In_1338);
and U511 (N_511,In_568,In_130);
nor U512 (N_512,In_1122,In_635);
nor U513 (N_513,In_1115,In_598);
nor U514 (N_514,In_1264,In_718);
or U515 (N_515,In_1169,In_1343);
nand U516 (N_516,In_1093,In_650);
and U517 (N_517,In_1464,In_651);
nor U518 (N_518,In_1310,In_843);
xnor U519 (N_519,In_915,In_790);
or U520 (N_520,In_1479,In_261);
or U521 (N_521,In_1092,In_672);
or U522 (N_522,In_1485,In_394);
xnor U523 (N_523,In_381,In_1474);
nor U524 (N_524,In_733,In_929);
or U525 (N_525,In_1496,In_1100);
nor U526 (N_526,In_1071,In_735);
and U527 (N_527,In_126,In_172);
nand U528 (N_528,In_1415,In_1472);
and U529 (N_529,In_985,In_822);
and U530 (N_530,In_196,In_815);
or U531 (N_531,In_866,In_575);
or U532 (N_532,In_324,In_924);
nand U533 (N_533,In_47,In_1048);
nor U534 (N_534,In_1302,In_355);
nor U535 (N_535,In_801,In_631);
nor U536 (N_536,In_574,In_62);
or U537 (N_537,In_1452,In_1391);
xor U538 (N_538,In_298,In_48);
nor U539 (N_539,In_1174,In_334);
nand U540 (N_540,In_600,In_1331);
or U541 (N_541,In_799,In_1007);
and U542 (N_542,In_170,In_210);
and U543 (N_543,In_1296,In_1407);
nand U544 (N_544,In_528,In_1356);
nand U545 (N_545,In_742,In_1129);
nor U546 (N_546,In_998,In_1028);
nor U547 (N_547,In_1283,In_119);
nand U548 (N_548,In_316,In_1070);
nand U549 (N_549,In_1185,In_1009);
and U550 (N_550,In_648,In_618);
and U551 (N_551,In_569,In_374);
nor U552 (N_552,In_1006,In_847);
or U553 (N_553,In_229,In_824);
nor U554 (N_554,In_662,In_1258);
or U555 (N_555,In_1192,In_379);
and U556 (N_556,In_992,In_1360);
and U557 (N_557,In_1477,In_1377);
xor U558 (N_558,In_476,In_1260);
and U559 (N_559,In_295,In_209);
nor U560 (N_560,In_1418,In_898);
or U561 (N_561,In_105,In_736);
xnor U562 (N_562,In_152,In_1147);
and U563 (N_563,In_913,In_339);
or U564 (N_564,In_403,In_615);
and U565 (N_565,In_632,In_862);
or U566 (N_566,In_1018,In_611);
nand U567 (N_567,In_1025,In_685);
nor U568 (N_568,In_1221,In_382);
and U569 (N_569,In_245,In_451);
or U570 (N_570,In_461,In_1438);
and U571 (N_571,In_1220,In_797);
nand U572 (N_572,In_4,In_306);
and U573 (N_573,In_1133,In_709);
nand U574 (N_574,In_830,In_1321);
nand U575 (N_575,In_174,In_1236);
and U576 (N_576,In_1075,In_1495);
nor U577 (N_577,In_206,In_1141);
and U578 (N_578,In_1434,In_140);
or U579 (N_579,In_976,In_1279);
nand U580 (N_580,In_640,In_1417);
nand U581 (N_581,In_1271,In_858);
and U582 (N_582,In_549,In_448);
nor U583 (N_583,In_162,In_342);
and U584 (N_584,In_1395,In_1068);
or U585 (N_585,In_16,In_429);
nand U586 (N_586,In_1227,In_539);
and U587 (N_587,In_1303,In_614);
and U588 (N_588,In_213,In_498);
nor U589 (N_589,In_594,In_431);
nor U590 (N_590,In_32,In_1341);
xnor U591 (N_591,In_83,In_337);
xnor U592 (N_592,In_1498,In_773);
or U593 (N_593,In_802,In_547);
or U594 (N_594,In_1318,In_855);
and U595 (N_595,In_198,In_807);
nand U596 (N_596,In_863,In_1309);
or U597 (N_597,In_1057,In_131);
xor U598 (N_598,In_283,In_1247);
and U599 (N_599,In_522,In_1378);
or U600 (N_600,In_349,In_681);
and U601 (N_601,In_1371,In_1012);
nand U602 (N_602,In_719,In_950);
xor U603 (N_603,In_1181,In_758);
and U604 (N_604,In_92,In_593);
and U605 (N_605,In_509,In_116);
or U606 (N_606,In_872,In_936);
nand U607 (N_607,In_1404,In_1255);
xor U608 (N_608,In_361,In_236);
nor U609 (N_609,In_1437,In_970);
and U610 (N_610,In_1409,In_1313);
nand U611 (N_611,In_388,In_320);
nand U612 (N_612,In_341,In_943);
nand U613 (N_613,In_20,In_392);
nand U614 (N_614,In_263,In_1398);
or U615 (N_615,In_1353,In_1095);
or U616 (N_616,In_462,In_696);
nor U617 (N_617,In_155,In_859);
nor U618 (N_618,In_1257,In_1027);
and U619 (N_619,In_1261,In_1251);
or U620 (N_620,In_285,In_251);
and U621 (N_621,In_1399,In_77);
nand U622 (N_622,In_3,In_1449);
and U623 (N_623,In_1091,In_1026);
and U624 (N_624,In_706,In_343);
or U625 (N_625,In_778,In_437);
xnor U626 (N_626,In_22,In_868);
nor U627 (N_627,In_1358,In_507);
or U628 (N_628,In_215,In_620);
xnor U629 (N_629,In_27,In_203);
nand U630 (N_630,In_759,In_59);
or U631 (N_631,In_248,In_276);
nor U632 (N_632,In_100,In_178);
or U633 (N_633,In_56,In_329);
nand U634 (N_634,In_1354,In_351);
xor U635 (N_635,In_137,In_535);
xor U636 (N_636,In_1138,In_869);
nor U637 (N_637,In_228,In_460);
nor U638 (N_638,In_634,In_1392);
xnor U639 (N_639,In_1228,In_1144);
and U640 (N_640,In_988,In_577);
or U641 (N_641,In_1030,In_459);
nand U642 (N_642,In_1297,In_1454);
and U643 (N_643,In_1132,In_26);
and U644 (N_644,In_1304,In_191);
nor U645 (N_645,In_693,In_1131);
and U646 (N_646,In_154,In_1330);
nor U647 (N_647,In_784,In_608);
or U648 (N_648,In_1242,In_103);
nand U649 (N_649,In_677,In_488);
nor U650 (N_650,In_834,In_664);
or U651 (N_651,In_503,In_573);
and U652 (N_652,In_360,In_297);
and U653 (N_653,In_1421,In_230);
xor U654 (N_654,In_557,In_682);
or U655 (N_655,In_544,In_692);
and U656 (N_656,In_533,In_751);
or U657 (N_657,In_514,In_1161);
and U658 (N_658,In_194,In_907);
and U659 (N_659,In_122,In_428);
nor U660 (N_660,In_884,In_127);
nand U661 (N_661,In_1465,In_314);
or U662 (N_662,In_1160,In_490);
nand U663 (N_663,In_766,In_1312);
nor U664 (N_664,In_71,In_413);
nor U665 (N_665,In_1203,In_1170);
xor U666 (N_666,In_435,In_479);
nand U667 (N_667,In_109,In_401);
nor U668 (N_668,In_813,In_833);
nor U669 (N_669,In_1367,In_954);
nand U670 (N_670,In_370,In_118);
nor U671 (N_671,In_942,In_1226);
nor U672 (N_672,In_144,In_701);
nand U673 (N_673,In_1002,In_427);
nor U674 (N_674,In_486,In_1124);
and U675 (N_675,In_391,In_106);
and U676 (N_676,In_472,In_244);
or U677 (N_677,In_226,In_94);
and U678 (N_678,In_376,In_1205);
or U679 (N_679,In_1056,In_996);
nand U680 (N_680,In_1224,In_505);
nand U681 (N_681,In_617,In_282);
or U682 (N_682,In_1217,In_1108);
nand U683 (N_683,In_478,In_253);
nor U684 (N_684,In_171,In_837);
nand U685 (N_685,In_289,In_624);
nor U686 (N_686,In_586,In_5);
nor U687 (N_687,In_1455,In_1329);
and U688 (N_688,In_1281,In_917);
and U689 (N_689,In_1235,In_304);
xor U690 (N_690,In_668,In_1171);
or U691 (N_691,In_1481,In_604);
xnor U692 (N_692,In_493,In_983);
nor U693 (N_693,In_1162,In_743);
and U694 (N_694,In_291,In_956);
and U695 (N_695,In_1135,In_419);
and U696 (N_696,In_37,In_157);
nor U697 (N_697,In_1447,In_771);
or U698 (N_698,In_1042,In_764);
and U699 (N_699,In_18,In_1055);
or U700 (N_700,In_494,In_702);
nand U701 (N_701,In_750,In_147);
and U702 (N_702,In_387,In_738);
xnor U703 (N_703,In_879,In_93);
nand U704 (N_704,In_559,In_746);
or U705 (N_705,In_536,In_645);
nor U706 (N_706,In_1094,In_227);
and U707 (N_707,In_710,In_1381);
nand U708 (N_708,In_49,In_173);
nor U709 (N_709,In_902,In_1194);
or U710 (N_710,In_414,In_201);
nor U711 (N_711,In_712,In_143);
nor U712 (N_712,In_400,In_424);
or U713 (N_713,In_1491,In_525);
or U714 (N_714,In_1435,In_444);
nor U715 (N_715,In_816,In_310);
or U716 (N_716,In_399,In_1488);
xor U717 (N_717,In_1020,In_1420);
nor U718 (N_718,In_684,In_72);
nand U719 (N_719,In_294,In_852);
xor U720 (N_720,In_1127,In_1290);
nand U721 (N_721,In_58,In_579);
or U722 (N_722,In_752,In_330);
or U723 (N_723,In_84,In_679);
xor U724 (N_724,In_794,In_398);
and U725 (N_725,In_1040,In_1038);
nor U726 (N_726,In_1032,In_79);
and U727 (N_727,In_128,In_981);
nand U728 (N_728,In_564,In_530);
nand U729 (N_729,In_135,In_592);
nor U730 (N_730,In_1293,In_1250);
xnor U731 (N_731,In_1432,In_753);
nand U732 (N_732,In_768,In_851);
nand U733 (N_733,In_779,In_571);
nor U734 (N_734,In_819,In_1239);
and U735 (N_735,In_148,In_1375);
or U736 (N_736,In_1443,In_499);
nand U737 (N_737,In_774,In_1380);
nand U738 (N_738,In_192,In_91);
nand U739 (N_739,In_1317,In_216);
and U740 (N_740,In_1408,In_638);
or U741 (N_741,In_587,In_1249);
nand U742 (N_742,In_1322,In_1128);
xor U743 (N_743,In_885,In_971);
and U744 (N_744,In_1323,In_1280);
xnor U745 (N_745,In_142,In_0);
or U746 (N_746,In_1342,In_1328);
or U747 (N_747,In_332,In_554);
nor U748 (N_748,In_1232,In_945);
or U749 (N_749,In_34,In_1333);
xor U750 (N_750,In_1394,In_987);
nor U751 (N_751,In_281,In_97);
or U752 (N_752,In_835,In_1475);
xor U753 (N_753,In_124,In_1468);
or U754 (N_754,In_1429,In_624);
nor U755 (N_755,In_1458,In_787);
and U756 (N_756,In_629,In_183);
nand U757 (N_757,In_237,In_679);
or U758 (N_758,In_478,In_483);
nor U759 (N_759,In_38,In_1229);
xnor U760 (N_760,In_878,In_120);
xor U761 (N_761,In_465,In_177);
and U762 (N_762,In_457,In_446);
or U763 (N_763,In_702,In_1180);
nand U764 (N_764,In_310,In_286);
and U765 (N_765,In_76,In_1192);
nand U766 (N_766,In_1048,In_821);
or U767 (N_767,In_1267,In_6);
nand U768 (N_768,In_984,In_862);
nor U769 (N_769,In_1421,In_580);
or U770 (N_770,In_1155,In_1484);
or U771 (N_771,In_583,In_840);
nand U772 (N_772,In_1351,In_458);
nand U773 (N_773,In_1013,In_425);
or U774 (N_774,In_960,In_1185);
or U775 (N_775,In_24,In_1469);
nand U776 (N_776,In_671,In_81);
nor U777 (N_777,In_1230,In_61);
nor U778 (N_778,In_401,In_55);
and U779 (N_779,In_881,In_247);
nand U780 (N_780,In_488,In_169);
and U781 (N_781,In_58,In_588);
nand U782 (N_782,In_258,In_1297);
nand U783 (N_783,In_581,In_285);
nor U784 (N_784,In_564,In_79);
xor U785 (N_785,In_669,In_762);
or U786 (N_786,In_897,In_109);
and U787 (N_787,In_279,In_1154);
nand U788 (N_788,In_1259,In_1040);
xor U789 (N_789,In_1484,In_927);
nor U790 (N_790,In_23,In_139);
nor U791 (N_791,In_359,In_1087);
nor U792 (N_792,In_485,In_579);
or U793 (N_793,In_177,In_1181);
nand U794 (N_794,In_1152,In_1454);
xnor U795 (N_795,In_1065,In_1061);
or U796 (N_796,In_765,In_775);
nor U797 (N_797,In_208,In_1173);
nand U798 (N_798,In_541,In_608);
or U799 (N_799,In_1436,In_1438);
or U800 (N_800,In_111,In_227);
nor U801 (N_801,In_965,In_1209);
nand U802 (N_802,In_156,In_735);
and U803 (N_803,In_830,In_875);
or U804 (N_804,In_303,In_37);
or U805 (N_805,In_663,In_206);
and U806 (N_806,In_1407,In_1081);
and U807 (N_807,In_1309,In_587);
nor U808 (N_808,In_602,In_471);
nand U809 (N_809,In_1340,In_272);
and U810 (N_810,In_1350,In_309);
or U811 (N_811,In_331,In_969);
nor U812 (N_812,In_1452,In_315);
or U813 (N_813,In_419,In_1024);
nor U814 (N_814,In_1106,In_297);
and U815 (N_815,In_479,In_868);
nor U816 (N_816,In_249,In_507);
nand U817 (N_817,In_479,In_1008);
xnor U818 (N_818,In_805,In_865);
and U819 (N_819,In_1066,In_1244);
xor U820 (N_820,In_1420,In_1389);
nand U821 (N_821,In_1389,In_506);
nand U822 (N_822,In_911,In_1080);
and U823 (N_823,In_750,In_715);
xor U824 (N_824,In_331,In_269);
or U825 (N_825,In_1083,In_65);
nor U826 (N_826,In_1332,In_1298);
nand U827 (N_827,In_1299,In_793);
nand U828 (N_828,In_654,In_525);
nand U829 (N_829,In_1172,In_33);
nor U830 (N_830,In_412,In_481);
and U831 (N_831,In_1089,In_701);
nor U832 (N_832,In_926,In_1367);
or U833 (N_833,In_1122,In_173);
or U834 (N_834,In_483,In_1325);
or U835 (N_835,In_138,In_384);
and U836 (N_836,In_354,In_489);
nand U837 (N_837,In_295,In_915);
nor U838 (N_838,In_69,In_924);
nor U839 (N_839,In_918,In_1177);
and U840 (N_840,In_241,In_1334);
and U841 (N_841,In_424,In_168);
nor U842 (N_842,In_1402,In_724);
and U843 (N_843,In_1025,In_450);
nand U844 (N_844,In_625,In_583);
nand U845 (N_845,In_306,In_335);
nor U846 (N_846,In_710,In_832);
nor U847 (N_847,In_1187,In_1249);
and U848 (N_848,In_1122,In_507);
and U849 (N_849,In_425,In_330);
nor U850 (N_850,In_758,In_1114);
or U851 (N_851,In_673,In_1052);
or U852 (N_852,In_1244,In_894);
or U853 (N_853,In_986,In_1482);
nand U854 (N_854,In_133,In_867);
and U855 (N_855,In_1084,In_229);
nand U856 (N_856,In_995,In_455);
nor U857 (N_857,In_860,In_683);
and U858 (N_858,In_1149,In_260);
or U859 (N_859,In_1078,In_570);
nand U860 (N_860,In_1064,In_1424);
and U861 (N_861,In_905,In_244);
nor U862 (N_862,In_364,In_1155);
and U863 (N_863,In_1278,In_894);
nand U864 (N_864,In_1120,In_875);
nor U865 (N_865,In_607,In_1191);
nor U866 (N_866,In_962,In_211);
and U867 (N_867,In_17,In_1201);
nor U868 (N_868,In_1046,In_691);
and U869 (N_869,In_446,In_1077);
xor U870 (N_870,In_276,In_1409);
nor U871 (N_871,In_1420,In_308);
nor U872 (N_872,In_668,In_1336);
nand U873 (N_873,In_1182,In_1019);
nor U874 (N_874,In_977,In_550);
nand U875 (N_875,In_897,In_1153);
and U876 (N_876,In_458,In_1007);
nand U877 (N_877,In_110,In_571);
nand U878 (N_878,In_751,In_1383);
and U879 (N_879,In_517,In_1200);
nand U880 (N_880,In_350,In_710);
nand U881 (N_881,In_1474,In_235);
or U882 (N_882,In_1193,In_773);
nor U883 (N_883,In_438,In_1234);
and U884 (N_884,In_501,In_917);
xor U885 (N_885,In_33,In_1433);
or U886 (N_886,In_438,In_221);
and U887 (N_887,In_420,In_350);
or U888 (N_888,In_1343,In_502);
nand U889 (N_889,In_1217,In_611);
and U890 (N_890,In_1076,In_754);
nor U891 (N_891,In_1097,In_1191);
or U892 (N_892,In_1016,In_123);
nand U893 (N_893,In_1482,In_1408);
nor U894 (N_894,In_515,In_868);
nand U895 (N_895,In_1169,In_470);
and U896 (N_896,In_469,In_1381);
xnor U897 (N_897,In_1308,In_499);
xor U898 (N_898,In_927,In_128);
and U899 (N_899,In_1370,In_1402);
nand U900 (N_900,In_1301,In_1388);
xor U901 (N_901,In_959,In_1064);
nand U902 (N_902,In_970,In_691);
xor U903 (N_903,In_97,In_1297);
nor U904 (N_904,In_1116,In_158);
or U905 (N_905,In_37,In_55);
nor U906 (N_906,In_63,In_1175);
and U907 (N_907,In_1305,In_632);
or U908 (N_908,In_381,In_550);
nand U909 (N_909,In_1390,In_1031);
xor U910 (N_910,In_873,In_582);
or U911 (N_911,In_302,In_1282);
or U912 (N_912,In_362,In_418);
and U913 (N_913,In_78,In_1112);
and U914 (N_914,In_952,In_929);
xnor U915 (N_915,In_793,In_1128);
or U916 (N_916,In_1168,In_1003);
nand U917 (N_917,In_564,In_999);
or U918 (N_918,In_909,In_1029);
xor U919 (N_919,In_1313,In_217);
and U920 (N_920,In_808,In_1405);
nand U921 (N_921,In_313,In_36);
nor U922 (N_922,In_996,In_52);
nor U923 (N_923,In_855,In_1237);
nor U924 (N_924,In_633,In_1164);
or U925 (N_925,In_1405,In_1495);
and U926 (N_926,In_970,In_6);
xnor U927 (N_927,In_105,In_1315);
or U928 (N_928,In_1326,In_115);
or U929 (N_929,In_1072,In_148);
xor U930 (N_930,In_137,In_366);
xor U931 (N_931,In_61,In_1009);
or U932 (N_932,In_314,In_1015);
nand U933 (N_933,In_964,In_1167);
or U934 (N_934,In_1409,In_28);
or U935 (N_935,In_585,In_1037);
and U936 (N_936,In_450,In_796);
and U937 (N_937,In_1058,In_949);
nor U938 (N_938,In_1176,In_618);
nand U939 (N_939,In_674,In_982);
nor U940 (N_940,In_416,In_278);
nand U941 (N_941,In_246,In_224);
or U942 (N_942,In_203,In_890);
xor U943 (N_943,In_778,In_1205);
nor U944 (N_944,In_118,In_841);
and U945 (N_945,In_1273,In_994);
and U946 (N_946,In_744,In_886);
nand U947 (N_947,In_707,In_251);
xnor U948 (N_948,In_400,In_224);
nand U949 (N_949,In_238,In_453);
or U950 (N_950,In_1017,In_1213);
or U951 (N_951,In_886,In_598);
xor U952 (N_952,In_163,In_371);
and U953 (N_953,In_832,In_47);
nor U954 (N_954,In_834,In_516);
and U955 (N_955,In_1356,In_1178);
or U956 (N_956,In_159,In_1450);
or U957 (N_957,In_452,In_997);
xor U958 (N_958,In_347,In_912);
nor U959 (N_959,In_138,In_1290);
or U960 (N_960,In_319,In_814);
and U961 (N_961,In_163,In_613);
nor U962 (N_962,In_1451,In_1300);
or U963 (N_963,In_193,In_413);
nor U964 (N_964,In_1249,In_1438);
or U965 (N_965,In_1301,In_135);
and U966 (N_966,In_256,In_1290);
nor U967 (N_967,In_1222,In_308);
nor U968 (N_968,In_128,In_1241);
nor U969 (N_969,In_1167,In_414);
nor U970 (N_970,In_1020,In_875);
nand U971 (N_971,In_507,In_1434);
nor U972 (N_972,In_951,In_413);
or U973 (N_973,In_904,In_759);
nand U974 (N_974,In_689,In_786);
and U975 (N_975,In_1031,In_133);
nor U976 (N_976,In_194,In_845);
nand U977 (N_977,In_197,In_708);
xnor U978 (N_978,In_271,In_87);
xnor U979 (N_979,In_718,In_916);
nor U980 (N_980,In_739,In_693);
and U981 (N_981,In_42,In_68);
and U982 (N_982,In_1461,In_429);
nor U983 (N_983,In_281,In_1133);
nor U984 (N_984,In_819,In_366);
nand U985 (N_985,In_145,In_1303);
or U986 (N_986,In_602,In_1390);
nand U987 (N_987,In_394,In_1153);
nand U988 (N_988,In_927,In_1059);
and U989 (N_989,In_230,In_517);
nand U990 (N_990,In_1013,In_660);
or U991 (N_991,In_1418,In_132);
nand U992 (N_992,In_1195,In_1141);
nor U993 (N_993,In_1446,In_623);
nand U994 (N_994,In_80,In_247);
and U995 (N_995,In_1341,In_1106);
nor U996 (N_996,In_1258,In_830);
nand U997 (N_997,In_839,In_1450);
nor U998 (N_998,In_744,In_637);
nand U999 (N_999,In_620,In_600);
or U1000 (N_1000,In_439,In_1237);
nor U1001 (N_1001,In_323,In_932);
or U1002 (N_1002,In_968,In_682);
and U1003 (N_1003,In_230,In_1018);
or U1004 (N_1004,In_1375,In_1199);
and U1005 (N_1005,In_1009,In_1056);
and U1006 (N_1006,In_449,In_682);
nor U1007 (N_1007,In_0,In_1272);
xor U1008 (N_1008,In_928,In_67);
xnor U1009 (N_1009,In_1074,In_434);
nand U1010 (N_1010,In_1045,In_717);
and U1011 (N_1011,In_699,In_269);
nand U1012 (N_1012,In_372,In_933);
xor U1013 (N_1013,In_439,In_1481);
nor U1014 (N_1014,In_1287,In_1065);
nor U1015 (N_1015,In_859,In_341);
and U1016 (N_1016,In_228,In_433);
nand U1017 (N_1017,In_1420,In_3);
and U1018 (N_1018,In_940,In_1082);
xnor U1019 (N_1019,In_1124,In_1209);
or U1020 (N_1020,In_1053,In_357);
nand U1021 (N_1021,In_533,In_383);
or U1022 (N_1022,In_1159,In_356);
nor U1023 (N_1023,In_1493,In_1297);
xor U1024 (N_1024,In_355,In_1313);
nor U1025 (N_1025,In_1029,In_578);
or U1026 (N_1026,In_1372,In_660);
and U1027 (N_1027,In_292,In_1358);
nor U1028 (N_1028,In_222,In_801);
xnor U1029 (N_1029,In_432,In_1121);
nor U1030 (N_1030,In_152,In_407);
or U1031 (N_1031,In_418,In_1248);
and U1032 (N_1032,In_361,In_959);
and U1033 (N_1033,In_962,In_456);
or U1034 (N_1034,In_1394,In_244);
or U1035 (N_1035,In_1183,In_1135);
nor U1036 (N_1036,In_1091,In_82);
xnor U1037 (N_1037,In_423,In_1335);
or U1038 (N_1038,In_691,In_1369);
and U1039 (N_1039,In_1172,In_701);
and U1040 (N_1040,In_916,In_259);
nand U1041 (N_1041,In_583,In_1248);
and U1042 (N_1042,In_584,In_180);
and U1043 (N_1043,In_353,In_204);
or U1044 (N_1044,In_26,In_859);
and U1045 (N_1045,In_466,In_1121);
nor U1046 (N_1046,In_72,In_765);
xor U1047 (N_1047,In_1067,In_596);
nor U1048 (N_1048,In_986,In_28);
or U1049 (N_1049,In_22,In_788);
and U1050 (N_1050,In_129,In_800);
nand U1051 (N_1051,In_1499,In_1176);
and U1052 (N_1052,In_1135,In_1084);
or U1053 (N_1053,In_1173,In_133);
nor U1054 (N_1054,In_736,In_1448);
nor U1055 (N_1055,In_1330,In_267);
or U1056 (N_1056,In_269,In_198);
nor U1057 (N_1057,In_590,In_1366);
or U1058 (N_1058,In_1390,In_41);
nand U1059 (N_1059,In_60,In_832);
or U1060 (N_1060,In_988,In_1029);
nor U1061 (N_1061,In_338,In_899);
xnor U1062 (N_1062,In_1443,In_335);
nand U1063 (N_1063,In_1,In_1327);
and U1064 (N_1064,In_897,In_716);
nand U1065 (N_1065,In_1213,In_1435);
or U1066 (N_1066,In_1253,In_1420);
or U1067 (N_1067,In_1143,In_954);
nand U1068 (N_1068,In_1222,In_200);
nand U1069 (N_1069,In_1091,In_196);
or U1070 (N_1070,In_739,In_484);
nand U1071 (N_1071,In_1058,In_713);
and U1072 (N_1072,In_1359,In_13);
nand U1073 (N_1073,In_1382,In_108);
nor U1074 (N_1074,In_611,In_1348);
nor U1075 (N_1075,In_931,In_1220);
and U1076 (N_1076,In_112,In_854);
nand U1077 (N_1077,In_863,In_192);
xnor U1078 (N_1078,In_1414,In_905);
nor U1079 (N_1079,In_1262,In_272);
or U1080 (N_1080,In_307,In_1071);
and U1081 (N_1081,In_876,In_815);
or U1082 (N_1082,In_270,In_1028);
nor U1083 (N_1083,In_6,In_360);
and U1084 (N_1084,In_286,In_447);
nand U1085 (N_1085,In_485,In_218);
or U1086 (N_1086,In_475,In_387);
nor U1087 (N_1087,In_1117,In_10);
nor U1088 (N_1088,In_49,In_163);
xnor U1089 (N_1089,In_1226,In_110);
nor U1090 (N_1090,In_945,In_897);
or U1091 (N_1091,In_190,In_224);
nor U1092 (N_1092,In_1020,In_1384);
nor U1093 (N_1093,In_306,In_1219);
or U1094 (N_1094,In_75,In_1120);
and U1095 (N_1095,In_401,In_1182);
nand U1096 (N_1096,In_749,In_673);
or U1097 (N_1097,In_437,In_779);
nor U1098 (N_1098,In_1063,In_131);
nand U1099 (N_1099,In_1152,In_758);
nand U1100 (N_1100,In_1359,In_235);
nor U1101 (N_1101,In_1156,In_135);
or U1102 (N_1102,In_901,In_1183);
and U1103 (N_1103,In_209,In_1003);
and U1104 (N_1104,In_569,In_1261);
nand U1105 (N_1105,In_1066,In_1057);
nand U1106 (N_1106,In_351,In_253);
and U1107 (N_1107,In_1101,In_679);
and U1108 (N_1108,In_1384,In_1355);
nand U1109 (N_1109,In_796,In_33);
and U1110 (N_1110,In_108,In_166);
nor U1111 (N_1111,In_1260,In_47);
and U1112 (N_1112,In_175,In_1139);
nor U1113 (N_1113,In_383,In_223);
nor U1114 (N_1114,In_183,In_742);
nand U1115 (N_1115,In_1394,In_152);
and U1116 (N_1116,In_376,In_981);
or U1117 (N_1117,In_1231,In_1168);
or U1118 (N_1118,In_49,In_719);
and U1119 (N_1119,In_33,In_50);
nand U1120 (N_1120,In_961,In_602);
and U1121 (N_1121,In_450,In_536);
nor U1122 (N_1122,In_298,In_1108);
nand U1123 (N_1123,In_667,In_986);
nand U1124 (N_1124,In_153,In_755);
nor U1125 (N_1125,In_905,In_1399);
nor U1126 (N_1126,In_1213,In_1004);
nand U1127 (N_1127,In_506,In_1444);
and U1128 (N_1128,In_249,In_1137);
or U1129 (N_1129,In_1316,In_1340);
nor U1130 (N_1130,In_1372,In_600);
and U1131 (N_1131,In_672,In_103);
or U1132 (N_1132,In_67,In_68);
xnor U1133 (N_1133,In_74,In_447);
or U1134 (N_1134,In_741,In_482);
and U1135 (N_1135,In_1109,In_1399);
nor U1136 (N_1136,In_31,In_470);
or U1137 (N_1137,In_647,In_1019);
or U1138 (N_1138,In_1413,In_1186);
or U1139 (N_1139,In_1006,In_1306);
nand U1140 (N_1140,In_658,In_269);
nand U1141 (N_1141,In_148,In_519);
nor U1142 (N_1142,In_1419,In_531);
and U1143 (N_1143,In_1036,In_1448);
nor U1144 (N_1144,In_1051,In_557);
nand U1145 (N_1145,In_193,In_999);
nand U1146 (N_1146,In_1150,In_935);
and U1147 (N_1147,In_1358,In_1023);
nand U1148 (N_1148,In_530,In_614);
xor U1149 (N_1149,In_1494,In_1481);
and U1150 (N_1150,In_872,In_226);
nand U1151 (N_1151,In_577,In_672);
and U1152 (N_1152,In_509,In_523);
nand U1153 (N_1153,In_1100,In_1488);
or U1154 (N_1154,In_831,In_1151);
nor U1155 (N_1155,In_514,In_558);
or U1156 (N_1156,In_847,In_20);
or U1157 (N_1157,In_30,In_104);
nand U1158 (N_1158,In_173,In_407);
or U1159 (N_1159,In_658,In_33);
nor U1160 (N_1160,In_1273,In_1134);
or U1161 (N_1161,In_980,In_1491);
or U1162 (N_1162,In_988,In_540);
or U1163 (N_1163,In_564,In_938);
nand U1164 (N_1164,In_469,In_1287);
nor U1165 (N_1165,In_107,In_1183);
or U1166 (N_1166,In_527,In_674);
xnor U1167 (N_1167,In_762,In_443);
and U1168 (N_1168,In_1355,In_1226);
nand U1169 (N_1169,In_24,In_915);
and U1170 (N_1170,In_290,In_794);
and U1171 (N_1171,In_204,In_1038);
xnor U1172 (N_1172,In_830,In_452);
and U1173 (N_1173,In_91,In_564);
nand U1174 (N_1174,In_323,In_763);
and U1175 (N_1175,In_1375,In_361);
nor U1176 (N_1176,In_926,In_976);
and U1177 (N_1177,In_533,In_613);
or U1178 (N_1178,In_1142,In_172);
nor U1179 (N_1179,In_605,In_447);
nand U1180 (N_1180,In_935,In_291);
or U1181 (N_1181,In_1410,In_1195);
nor U1182 (N_1182,In_1258,In_473);
or U1183 (N_1183,In_915,In_1416);
nor U1184 (N_1184,In_361,In_799);
and U1185 (N_1185,In_887,In_722);
xor U1186 (N_1186,In_202,In_67);
nor U1187 (N_1187,In_1025,In_772);
or U1188 (N_1188,In_1181,In_110);
nor U1189 (N_1189,In_641,In_1241);
xor U1190 (N_1190,In_686,In_338);
nand U1191 (N_1191,In_938,In_1043);
nand U1192 (N_1192,In_188,In_891);
xnor U1193 (N_1193,In_857,In_1112);
nor U1194 (N_1194,In_738,In_820);
xnor U1195 (N_1195,In_255,In_587);
nand U1196 (N_1196,In_646,In_452);
and U1197 (N_1197,In_259,In_569);
nor U1198 (N_1198,In_669,In_63);
and U1199 (N_1199,In_862,In_950);
xor U1200 (N_1200,In_1352,In_1068);
or U1201 (N_1201,In_555,In_1067);
nand U1202 (N_1202,In_858,In_1184);
nand U1203 (N_1203,In_1266,In_302);
xor U1204 (N_1204,In_1328,In_859);
or U1205 (N_1205,In_1413,In_246);
or U1206 (N_1206,In_27,In_1067);
nand U1207 (N_1207,In_431,In_1440);
nand U1208 (N_1208,In_41,In_468);
nand U1209 (N_1209,In_254,In_817);
nor U1210 (N_1210,In_428,In_1104);
or U1211 (N_1211,In_93,In_1109);
and U1212 (N_1212,In_718,In_1155);
nand U1213 (N_1213,In_1124,In_1213);
nand U1214 (N_1214,In_584,In_342);
or U1215 (N_1215,In_1320,In_1139);
nand U1216 (N_1216,In_1293,In_1300);
and U1217 (N_1217,In_62,In_41);
nand U1218 (N_1218,In_412,In_702);
and U1219 (N_1219,In_767,In_279);
nand U1220 (N_1220,In_449,In_237);
nand U1221 (N_1221,In_106,In_918);
or U1222 (N_1222,In_791,In_1430);
and U1223 (N_1223,In_858,In_571);
nor U1224 (N_1224,In_210,In_340);
xor U1225 (N_1225,In_1,In_238);
and U1226 (N_1226,In_1080,In_171);
nor U1227 (N_1227,In_256,In_27);
nor U1228 (N_1228,In_1198,In_1042);
nand U1229 (N_1229,In_1407,In_96);
and U1230 (N_1230,In_1217,In_612);
nand U1231 (N_1231,In_531,In_946);
xnor U1232 (N_1232,In_253,In_936);
nand U1233 (N_1233,In_1042,In_218);
or U1234 (N_1234,In_992,In_942);
or U1235 (N_1235,In_1297,In_1324);
xnor U1236 (N_1236,In_1104,In_1038);
nand U1237 (N_1237,In_1354,In_1106);
nand U1238 (N_1238,In_1124,In_223);
or U1239 (N_1239,In_306,In_255);
nor U1240 (N_1240,In_707,In_931);
and U1241 (N_1241,In_401,In_77);
or U1242 (N_1242,In_586,In_1078);
xnor U1243 (N_1243,In_1363,In_36);
or U1244 (N_1244,In_1383,In_1436);
nand U1245 (N_1245,In_984,In_534);
and U1246 (N_1246,In_928,In_263);
or U1247 (N_1247,In_902,In_384);
and U1248 (N_1248,In_612,In_178);
or U1249 (N_1249,In_966,In_152);
nand U1250 (N_1250,In_516,In_607);
nor U1251 (N_1251,In_1304,In_1263);
and U1252 (N_1252,In_1049,In_1103);
or U1253 (N_1253,In_1384,In_206);
xor U1254 (N_1254,In_1408,In_648);
nand U1255 (N_1255,In_995,In_870);
nor U1256 (N_1256,In_393,In_209);
nand U1257 (N_1257,In_685,In_1491);
nor U1258 (N_1258,In_327,In_1161);
nand U1259 (N_1259,In_1262,In_674);
and U1260 (N_1260,In_369,In_599);
nand U1261 (N_1261,In_327,In_783);
xor U1262 (N_1262,In_630,In_410);
xor U1263 (N_1263,In_905,In_1193);
xnor U1264 (N_1264,In_435,In_972);
nand U1265 (N_1265,In_1183,In_746);
nor U1266 (N_1266,In_1240,In_927);
and U1267 (N_1267,In_1082,In_115);
nor U1268 (N_1268,In_1162,In_866);
or U1269 (N_1269,In_625,In_1451);
and U1270 (N_1270,In_533,In_795);
xor U1271 (N_1271,In_448,In_807);
nor U1272 (N_1272,In_447,In_497);
nand U1273 (N_1273,In_137,In_279);
nand U1274 (N_1274,In_34,In_653);
or U1275 (N_1275,In_955,In_999);
xnor U1276 (N_1276,In_1469,In_1351);
nand U1277 (N_1277,In_977,In_271);
or U1278 (N_1278,In_717,In_41);
nand U1279 (N_1279,In_305,In_416);
nand U1280 (N_1280,In_678,In_1309);
nand U1281 (N_1281,In_618,In_859);
nor U1282 (N_1282,In_1487,In_880);
nand U1283 (N_1283,In_697,In_1068);
xnor U1284 (N_1284,In_76,In_203);
nand U1285 (N_1285,In_673,In_100);
nand U1286 (N_1286,In_277,In_1187);
xnor U1287 (N_1287,In_167,In_626);
nor U1288 (N_1288,In_961,In_744);
or U1289 (N_1289,In_973,In_1241);
nor U1290 (N_1290,In_690,In_711);
nand U1291 (N_1291,In_541,In_1044);
xor U1292 (N_1292,In_1406,In_1422);
nand U1293 (N_1293,In_778,In_36);
or U1294 (N_1294,In_1268,In_277);
nor U1295 (N_1295,In_715,In_785);
or U1296 (N_1296,In_393,In_1156);
or U1297 (N_1297,In_105,In_13);
or U1298 (N_1298,In_17,In_1198);
nor U1299 (N_1299,In_941,In_631);
or U1300 (N_1300,In_442,In_111);
nand U1301 (N_1301,In_1371,In_1210);
or U1302 (N_1302,In_1093,In_463);
nand U1303 (N_1303,In_1096,In_205);
nor U1304 (N_1304,In_1115,In_1099);
and U1305 (N_1305,In_1318,In_968);
or U1306 (N_1306,In_1350,In_719);
nor U1307 (N_1307,In_221,In_106);
or U1308 (N_1308,In_232,In_1055);
nor U1309 (N_1309,In_107,In_127);
xor U1310 (N_1310,In_1440,In_834);
and U1311 (N_1311,In_406,In_458);
or U1312 (N_1312,In_675,In_364);
nor U1313 (N_1313,In_56,In_1429);
nor U1314 (N_1314,In_1230,In_861);
nor U1315 (N_1315,In_499,In_1314);
or U1316 (N_1316,In_1119,In_209);
xor U1317 (N_1317,In_563,In_1290);
and U1318 (N_1318,In_1279,In_997);
nand U1319 (N_1319,In_576,In_599);
nor U1320 (N_1320,In_1355,In_1084);
nor U1321 (N_1321,In_1031,In_1033);
nand U1322 (N_1322,In_817,In_1007);
nand U1323 (N_1323,In_261,In_87);
nor U1324 (N_1324,In_270,In_1481);
nor U1325 (N_1325,In_675,In_1236);
or U1326 (N_1326,In_1229,In_95);
nand U1327 (N_1327,In_787,In_35);
xor U1328 (N_1328,In_998,In_536);
and U1329 (N_1329,In_207,In_1289);
xnor U1330 (N_1330,In_1494,In_1129);
or U1331 (N_1331,In_148,In_877);
and U1332 (N_1332,In_1321,In_147);
and U1333 (N_1333,In_1082,In_1225);
nor U1334 (N_1334,In_633,In_1460);
or U1335 (N_1335,In_805,In_756);
nand U1336 (N_1336,In_389,In_1225);
or U1337 (N_1337,In_304,In_1141);
and U1338 (N_1338,In_22,In_620);
and U1339 (N_1339,In_962,In_589);
xnor U1340 (N_1340,In_250,In_695);
nor U1341 (N_1341,In_873,In_83);
and U1342 (N_1342,In_1192,In_387);
or U1343 (N_1343,In_527,In_895);
xor U1344 (N_1344,In_1491,In_666);
or U1345 (N_1345,In_430,In_691);
and U1346 (N_1346,In_1004,In_1260);
nand U1347 (N_1347,In_473,In_112);
xor U1348 (N_1348,In_627,In_444);
or U1349 (N_1349,In_1277,In_484);
nor U1350 (N_1350,In_1171,In_82);
xor U1351 (N_1351,In_282,In_776);
nand U1352 (N_1352,In_1138,In_623);
nand U1353 (N_1353,In_418,In_520);
and U1354 (N_1354,In_712,In_332);
nand U1355 (N_1355,In_62,In_223);
nand U1356 (N_1356,In_552,In_1238);
nand U1357 (N_1357,In_74,In_195);
nor U1358 (N_1358,In_1386,In_753);
or U1359 (N_1359,In_1324,In_878);
or U1360 (N_1360,In_54,In_1497);
nand U1361 (N_1361,In_361,In_105);
nand U1362 (N_1362,In_1361,In_1237);
xnor U1363 (N_1363,In_1220,In_457);
nand U1364 (N_1364,In_1170,In_0);
nand U1365 (N_1365,In_59,In_525);
and U1366 (N_1366,In_68,In_1268);
or U1367 (N_1367,In_998,In_54);
nor U1368 (N_1368,In_1167,In_926);
nand U1369 (N_1369,In_627,In_451);
and U1370 (N_1370,In_1411,In_1244);
nand U1371 (N_1371,In_969,In_1044);
nor U1372 (N_1372,In_1091,In_945);
or U1373 (N_1373,In_991,In_337);
xor U1374 (N_1374,In_423,In_421);
nand U1375 (N_1375,In_518,In_1330);
nand U1376 (N_1376,In_505,In_1319);
or U1377 (N_1377,In_735,In_1381);
and U1378 (N_1378,In_1233,In_393);
xnor U1379 (N_1379,In_19,In_56);
nand U1380 (N_1380,In_333,In_661);
xor U1381 (N_1381,In_859,In_330);
and U1382 (N_1382,In_101,In_793);
nand U1383 (N_1383,In_1466,In_251);
nand U1384 (N_1384,In_613,In_463);
and U1385 (N_1385,In_768,In_405);
xor U1386 (N_1386,In_546,In_403);
nand U1387 (N_1387,In_1247,In_1395);
xor U1388 (N_1388,In_929,In_889);
nor U1389 (N_1389,In_733,In_410);
nor U1390 (N_1390,In_1095,In_1143);
or U1391 (N_1391,In_237,In_557);
nor U1392 (N_1392,In_665,In_996);
nor U1393 (N_1393,In_483,In_502);
and U1394 (N_1394,In_962,In_103);
or U1395 (N_1395,In_480,In_360);
xnor U1396 (N_1396,In_588,In_1155);
nand U1397 (N_1397,In_518,In_373);
and U1398 (N_1398,In_1456,In_950);
nor U1399 (N_1399,In_113,In_752);
and U1400 (N_1400,In_172,In_1256);
nand U1401 (N_1401,In_196,In_693);
or U1402 (N_1402,In_131,In_685);
and U1403 (N_1403,In_420,In_824);
nand U1404 (N_1404,In_1445,In_774);
nand U1405 (N_1405,In_1466,In_1173);
and U1406 (N_1406,In_1020,In_269);
or U1407 (N_1407,In_1158,In_675);
nor U1408 (N_1408,In_322,In_169);
and U1409 (N_1409,In_412,In_418);
nor U1410 (N_1410,In_286,In_213);
nor U1411 (N_1411,In_1483,In_1286);
or U1412 (N_1412,In_993,In_1289);
nor U1413 (N_1413,In_662,In_1455);
and U1414 (N_1414,In_1212,In_1452);
nor U1415 (N_1415,In_1362,In_607);
nor U1416 (N_1416,In_363,In_1129);
nor U1417 (N_1417,In_15,In_927);
nor U1418 (N_1418,In_1323,In_87);
xnor U1419 (N_1419,In_1456,In_545);
or U1420 (N_1420,In_977,In_674);
or U1421 (N_1421,In_1493,In_903);
nand U1422 (N_1422,In_1372,In_1321);
and U1423 (N_1423,In_1274,In_690);
or U1424 (N_1424,In_1470,In_740);
and U1425 (N_1425,In_436,In_807);
nand U1426 (N_1426,In_444,In_490);
or U1427 (N_1427,In_481,In_326);
nand U1428 (N_1428,In_1111,In_638);
or U1429 (N_1429,In_918,In_935);
and U1430 (N_1430,In_482,In_1472);
nor U1431 (N_1431,In_734,In_1489);
nor U1432 (N_1432,In_710,In_454);
nand U1433 (N_1433,In_220,In_1436);
nor U1434 (N_1434,In_1463,In_1316);
nand U1435 (N_1435,In_1055,In_957);
and U1436 (N_1436,In_1070,In_594);
and U1437 (N_1437,In_542,In_446);
or U1438 (N_1438,In_461,In_1300);
or U1439 (N_1439,In_717,In_1222);
nand U1440 (N_1440,In_892,In_741);
nand U1441 (N_1441,In_753,In_94);
or U1442 (N_1442,In_1165,In_870);
nand U1443 (N_1443,In_804,In_451);
nor U1444 (N_1444,In_996,In_7);
or U1445 (N_1445,In_727,In_1293);
nor U1446 (N_1446,In_770,In_71);
nand U1447 (N_1447,In_1036,In_873);
nor U1448 (N_1448,In_633,In_1149);
and U1449 (N_1449,In_26,In_978);
or U1450 (N_1450,In_287,In_580);
or U1451 (N_1451,In_701,In_671);
and U1452 (N_1452,In_1097,In_525);
and U1453 (N_1453,In_1345,In_664);
nor U1454 (N_1454,In_1300,In_1080);
nor U1455 (N_1455,In_830,In_303);
nand U1456 (N_1456,In_1437,In_875);
or U1457 (N_1457,In_518,In_496);
and U1458 (N_1458,In_1324,In_251);
nor U1459 (N_1459,In_219,In_844);
nand U1460 (N_1460,In_954,In_1232);
nor U1461 (N_1461,In_787,In_914);
xnor U1462 (N_1462,In_23,In_116);
nand U1463 (N_1463,In_1106,In_729);
and U1464 (N_1464,In_27,In_1212);
nor U1465 (N_1465,In_25,In_1430);
nor U1466 (N_1466,In_1158,In_957);
nor U1467 (N_1467,In_568,In_679);
nand U1468 (N_1468,In_952,In_1385);
nand U1469 (N_1469,In_20,In_25);
or U1470 (N_1470,In_684,In_827);
and U1471 (N_1471,In_202,In_590);
nand U1472 (N_1472,In_950,In_440);
nand U1473 (N_1473,In_1110,In_139);
xnor U1474 (N_1474,In_51,In_1497);
nand U1475 (N_1475,In_1353,In_1124);
nand U1476 (N_1476,In_624,In_406);
nor U1477 (N_1477,In_649,In_1025);
xor U1478 (N_1478,In_1437,In_1295);
nor U1479 (N_1479,In_3,In_1067);
or U1480 (N_1480,In_911,In_1215);
nor U1481 (N_1481,In_1029,In_94);
and U1482 (N_1482,In_731,In_55);
or U1483 (N_1483,In_597,In_3);
nand U1484 (N_1484,In_343,In_69);
nor U1485 (N_1485,In_446,In_223);
and U1486 (N_1486,In_534,In_91);
or U1487 (N_1487,In_1409,In_1352);
nand U1488 (N_1488,In_752,In_443);
or U1489 (N_1489,In_907,In_1039);
or U1490 (N_1490,In_30,In_1011);
nand U1491 (N_1491,In_1262,In_393);
xor U1492 (N_1492,In_419,In_757);
nand U1493 (N_1493,In_654,In_1298);
and U1494 (N_1494,In_1018,In_61);
or U1495 (N_1495,In_291,In_492);
and U1496 (N_1496,In_968,In_504);
nor U1497 (N_1497,In_1338,In_31);
nor U1498 (N_1498,In_797,In_377);
and U1499 (N_1499,In_542,In_459);
nand U1500 (N_1500,N_270,N_550);
or U1501 (N_1501,N_324,N_311);
and U1502 (N_1502,N_1312,N_1219);
and U1503 (N_1503,N_204,N_726);
nor U1504 (N_1504,N_1324,N_494);
xnor U1505 (N_1505,N_166,N_594);
and U1506 (N_1506,N_146,N_736);
nand U1507 (N_1507,N_1409,N_500);
nand U1508 (N_1508,N_915,N_1028);
nor U1509 (N_1509,N_329,N_953);
nand U1510 (N_1510,N_1194,N_247);
and U1511 (N_1511,N_144,N_506);
and U1512 (N_1512,N_918,N_147);
and U1513 (N_1513,N_339,N_56);
nor U1514 (N_1514,N_1401,N_994);
nor U1515 (N_1515,N_211,N_1211);
nand U1516 (N_1516,N_1310,N_1394);
or U1517 (N_1517,N_33,N_751);
nand U1518 (N_1518,N_416,N_0);
xor U1519 (N_1519,N_1191,N_16);
or U1520 (N_1520,N_805,N_920);
nand U1521 (N_1521,N_397,N_931);
or U1522 (N_1522,N_943,N_1300);
or U1523 (N_1523,N_8,N_951);
nand U1524 (N_1524,N_648,N_1391);
and U1525 (N_1525,N_1374,N_759);
nand U1526 (N_1526,N_677,N_539);
and U1527 (N_1527,N_502,N_496);
nor U1528 (N_1528,N_767,N_120);
and U1529 (N_1529,N_349,N_407);
nor U1530 (N_1530,N_1383,N_292);
or U1531 (N_1531,N_1359,N_1499);
or U1532 (N_1532,N_1488,N_713);
nand U1533 (N_1533,N_970,N_456);
nor U1534 (N_1534,N_145,N_794);
and U1535 (N_1535,N_1197,N_1025);
and U1536 (N_1536,N_667,N_174);
or U1537 (N_1537,N_1200,N_1269);
and U1538 (N_1538,N_1048,N_1046);
nand U1539 (N_1539,N_1436,N_1356);
or U1540 (N_1540,N_914,N_873);
nor U1541 (N_1541,N_250,N_848);
nor U1542 (N_1542,N_909,N_40);
nor U1543 (N_1543,N_1388,N_954);
or U1544 (N_1544,N_1491,N_1428);
and U1545 (N_1545,N_878,N_975);
and U1546 (N_1546,N_1152,N_714);
nand U1547 (N_1547,N_352,N_393);
nand U1548 (N_1548,N_562,N_46);
nand U1549 (N_1549,N_551,N_839);
or U1550 (N_1550,N_1495,N_179);
nand U1551 (N_1551,N_428,N_336);
and U1552 (N_1552,N_774,N_348);
nor U1553 (N_1553,N_433,N_362);
nor U1554 (N_1554,N_880,N_1060);
xor U1555 (N_1555,N_729,N_1092);
and U1556 (N_1556,N_907,N_474);
nor U1557 (N_1557,N_312,N_298);
or U1558 (N_1558,N_361,N_1478);
or U1559 (N_1559,N_269,N_1119);
or U1560 (N_1560,N_50,N_1174);
nor U1561 (N_1561,N_932,N_1369);
or U1562 (N_1562,N_1001,N_162);
and U1563 (N_1563,N_897,N_1188);
nor U1564 (N_1564,N_1402,N_644);
nand U1565 (N_1565,N_1275,N_964);
nor U1566 (N_1566,N_290,N_608);
and U1567 (N_1567,N_1266,N_514);
or U1568 (N_1568,N_183,N_257);
nor U1569 (N_1569,N_1318,N_22);
or U1570 (N_1570,N_1236,N_882);
and U1571 (N_1571,N_1009,N_947);
xor U1572 (N_1572,N_401,N_1019);
nand U1573 (N_1573,N_876,N_463);
nor U1574 (N_1574,N_696,N_906);
nand U1575 (N_1575,N_578,N_1123);
nor U1576 (N_1576,N_786,N_657);
xor U1577 (N_1577,N_414,N_626);
nand U1578 (N_1578,N_689,N_1011);
and U1579 (N_1579,N_331,N_684);
or U1580 (N_1580,N_681,N_1160);
and U1581 (N_1581,N_1425,N_475);
nand U1582 (N_1582,N_619,N_1419);
nor U1583 (N_1583,N_1187,N_161);
or U1584 (N_1584,N_1427,N_1415);
and U1585 (N_1585,N_570,N_1496);
nor U1586 (N_1586,N_1375,N_912);
or U1587 (N_1587,N_295,N_719);
nor U1588 (N_1588,N_1330,N_647);
nor U1589 (N_1589,N_1452,N_662);
nand U1590 (N_1590,N_432,N_775);
nor U1591 (N_1591,N_236,N_881);
nor U1592 (N_1592,N_106,N_1389);
and U1593 (N_1593,N_1381,N_1333);
and U1594 (N_1594,N_85,N_617);
nand U1595 (N_1595,N_235,N_1444);
nor U1596 (N_1596,N_856,N_1189);
xor U1597 (N_1597,N_1075,N_1163);
nand U1598 (N_1598,N_969,N_1338);
and U1599 (N_1599,N_1424,N_1461);
or U1600 (N_1600,N_890,N_1272);
xor U1601 (N_1601,N_1130,N_653);
or U1602 (N_1602,N_1132,N_1059);
nor U1603 (N_1603,N_338,N_755);
and U1604 (N_1604,N_251,N_1249);
and U1605 (N_1605,N_272,N_522);
or U1606 (N_1606,N_492,N_410);
or U1607 (N_1607,N_581,N_418);
nor U1608 (N_1608,N_797,N_699);
nand U1609 (N_1609,N_1454,N_1061);
nand U1610 (N_1610,N_124,N_1034);
and U1611 (N_1611,N_425,N_589);
nand U1612 (N_1612,N_1110,N_977);
nand U1613 (N_1613,N_440,N_1377);
nand U1614 (N_1614,N_521,N_1006);
or U1615 (N_1615,N_989,N_182);
nand U1616 (N_1616,N_966,N_832);
nand U1617 (N_1617,N_1407,N_239);
nand U1618 (N_1618,N_1237,N_1340);
nor U1619 (N_1619,N_605,N_412);
nor U1620 (N_1620,N_804,N_592);
or U1621 (N_1621,N_462,N_900);
or U1622 (N_1622,N_937,N_107);
or U1623 (N_1623,N_152,N_520);
or U1624 (N_1624,N_974,N_795);
nand U1625 (N_1625,N_675,N_172);
or U1626 (N_1626,N_430,N_1256);
and U1627 (N_1627,N_98,N_671);
nor U1628 (N_1628,N_700,N_1018);
nor U1629 (N_1629,N_1032,N_674);
nor U1630 (N_1630,N_524,N_1031);
or U1631 (N_1631,N_673,N_1013);
nor U1632 (N_1632,N_482,N_72);
and U1633 (N_1633,N_12,N_691);
or U1634 (N_1634,N_277,N_164);
and U1635 (N_1635,N_1255,N_125);
or U1636 (N_1636,N_1385,N_1410);
or U1637 (N_1637,N_650,N_607);
and U1638 (N_1638,N_1393,N_11);
nand U1639 (N_1639,N_1204,N_582);
or U1640 (N_1640,N_1462,N_828);
nand U1641 (N_1641,N_296,N_1198);
or U1642 (N_1642,N_228,N_1420);
nor U1643 (N_1643,N_374,N_1304);
nand U1644 (N_1644,N_1103,N_1079);
or U1645 (N_1645,N_1035,N_806);
and U1646 (N_1646,N_965,N_344);
nor U1647 (N_1647,N_762,N_346);
nor U1648 (N_1648,N_1350,N_89);
and U1649 (N_1649,N_530,N_836);
nand U1650 (N_1650,N_504,N_905);
nor U1651 (N_1651,N_988,N_353);
nor U1652 (N_1652,N_71,N_28);
or U1653 (N_1653,N_999,N_728);
nand U1654 (N_1654,N_135,N_1351);
nand U1655 (N_1655,N_244,N_950);
nand U1656 (N_1656,N_1274,N_84);
and U1657 (N_1657,N_940,N_1397);
nor U1658 (N_1658,N_253,N_574);
and U1659 (N_1659,N_889,N_819);
and U1660 (N_1660,N_1073,N_869);
nand U1661 (N_1661,N_80,N_1050);
xor U1662 (N_1662,N_771,N_784);
nand U1663 (N_1663,N_61,N_655);
xnor U1664 (N_1664,N_1475,N_1089);
and U1665 (N_1665,N_710,N_101);
xnor U1666 (N_1666,N_1071,N_1127);
nand U1667 (N_1667,N_1278,N_707);
nand U1668 (N_1668,N_109,N_248);
nor U1669 (N_1669,N_275,N_24);
xor U1670 (N_1670,N_990,N_857);
or U1671 (N_1671,N_304,N_1133);
xor U1672 (N_1672,N_82,N_1024);
or U1673 (N_1673,N_1016,N_151);
nand U1674 (N_1674,N_116,N_863);
xor U1675 (N_1675,N_1386,N_796);
nor U1676 (N_1676,N_1149,N_1457);
nand U1677 (N_1677,N_165,N_321);
or U1678 (N_1678,N_1239,N_293);
xor U1679 (N_1679,N_1208,N_1292);
or U1680 (N_1680,N_213,N_1015);
nand U1681 (N_1681,N_567,N_92);
or U1682 (N_1682,N_1322,N_380);
and U1683 (N_1683,N_249,N_534);
nor U1684 (N_1684,N_712,N_229);
or U1685 (N_1685,N_489,N_309);
nand U1686 (N_1686,N_553,N_875);
or U1687 (N_1687,N_596,N_357);
nand U1688 (N_1688,N_807,N_294);
and U1689 (N_1689,N_533,N_1376);
and U1690 (N_1690,N_434,N_1069);
and U1691 (N_1691,N_10,N_67);
or U1692 (N_1692,N_1062,N_1190);
nand U1693 (N_1693,N_883,N_171);
and U1694 (N_1694,N_316,N_464);
or U1695 (N_1695,N_478,N_859);
and U1696 (N_1696,N_1311,N_579);
nor U1697 (N_1697,N_668,N_1307);
nor U1698 (N_1698,N_426,N_1373);
nand U1699 (N_1699,N_748,N_307);
and U1700 (N_1700,N_780,N_685);
or U1701 (N_1701,N_1443,N_501);
xor U1702 (N_1702,N_25,N_600);
and U1703 (N_1703,N_402,N_201);
nand U1704 (N_1704,N_575,N_765);
nand U1705 (N_1705,N_319,N_81);
and U1706 (N_1706,N_929,N_387);
and U1707 (N_1707,N_276,N_26);
nand U1708 (N_1708,N_1433,N_1235);
or U1709 (N_1709,N_1183,N_245);
and U1710 (N_1710,N_1145,N_788);
nand U1711 (N_1711,N_1192,N_636);
nor U1712 (N_1712,N_1064,N_818);
and U1713 (N_1713,N_264,N_845);
nand U1714 (N_1714,N_716,N_835);
nand U1715 (N_1715,N_158,N_1258);
or U1716 (N_1716,N_631,N_660);
nand U1717 (N_1717,N_766,N_350);
nor U1718 (N_1718,N_370,N_1482);
nand U1719 (N_1719,N_377,N_1049);
nand U1720 (N_1720,N_654,N_115);
nand U1721 (N_1721,N_864,N_527);
nor U1722 (N_1722,N_995,N_1230);
nor U1723 (N_1723,N_824,N_692);
or U1724 (N_1724,N_868,N_955);
and U1725 (N_1725,N_511,N_70);
nor U1726 (N_1726,N_1315,N_345);
or U1727 (N_1727,N_911,N_800);
nor U1728 (N_1728,N_922,N_470);
nand U1729 (N_1729,N_776,N_1063);
nand U1730 (N_1730,N_29,N_403);
or U1731 (N_1731,N_956,N_1017);
nor U1732 (N_1732,N_602,N_261);
and U1733 (N_1733,N_96,N_396);
or U1734 (N_1734,N_9,N_442);
nor U1735 (N_1735,N_758,N_232);
and U1736 (N_1736,N_1140,N_1308);
nor U1737 (N_1737,N_708,N_916);
and U1738 (N_1738,N_595,N_341);
nor U1739 (N_1739,N_559,N_243);
or U1740 (N_1740,N_935,N_1020);
nor U1741 (N_1741,N_625,N_616);
nand U1742 (N_1742,N_733,N_112);
nand U1743 (N_1743,N_833,N_1232);
or U1744 (N_1744,N_1468,N_958);
and U1745 (N_1745,N_676,N_1405);
and U1746 (N_1746,N_821,N_1321);
or U1747 (N_1747,N_505,N_557);
or U1748 (N_1748,N_448,N_702);
xor U1749 (N_1749,N_1309,N_877);
and U1750 (N_1750,N_1466,N_6);
or U1751 (N_1751,N_356,N_1413);
nor U1752 (N_1752,N_1181,N_159);
or U1753 (N_1753,N_623,N_545);
nor U1754 (N_1754,N_1207,N_1150);
and U1755 (N_1755,N_1203,N_1037);
xnor U1756 (N_1756,N_984,N_237);
or U1757 (N_1757,N_1489,N_1240);
nand U1758 (N_1758,N_238,N_141);
nor U1759 (N_1759,N_220,N_358);
nand U1760 (N_1760,N_614,N_682);
and U1761 (N_1761,N_1378,N_1184);
and U1762 (N_1762,N_980,N_1040);
or U1763 (N_1763,N_1349,N_1328);
nand U1764 (N_1764,N_778,N_1296);
and U1765 (N_1765,N_695,N_471);
nor U1766 (N_1766,N_1421,N_639);
nand U1767 (N_1767,N_129,N_862);
nand U1768 (N_1768,N_585,N_777);
nand U1769 (N_1769,N_223,N_1158);
and U1770 (N_1770,N_254,N_571);
or U1771 (N_1771,N_1380,N_720);
and U1772 (N_1772,N_611,N_703);
nand U1773 (N_1773,N_1446,N_894);
or U1774 (N_1774,N_1165,N_1345);
nand U1775 (N_1775,N_1448,N_74);
nand U1776 (N_1776,N_1023,N_395);
and U1777 (N_1777,N_1480,N_54);
or U1778 (N_1778,N_431,N_1412);
and U1779 (N_1779,N_513,N_1367);
nand U1780 (N_1780,N_991,N_556);
or U1781 (N_1781,N_1122,N_727);
nor U1782 (N_1782,N_1193,N_764);
xor U1783 (N_1783,N_564,N_435);
and U1784 (N_1784,N_925,N_785);
or U1785 (N_1785,N_523,N_306);
xnor U1786 (N_1786,N_366,N_1418);
or U1787 (N_1787,N_711,N_643);
and U1788 (N_1788,N_1291,N_1096);
and U1789 (N_1789,N_683,N_843);
nand U1790 (N_1790,N_892,N_566);
or U1791 (N_1791,N_177,N_169);
nand U1792 (N_1792,N_1329,N_73);
and U1793 (N_1793,N_355,N_1406);
or U1794 (N_1794,N_822,N_992);
nand U1795 (N_1795,N_113,N_1005);
nand U1796 (N_1796,N_466,N_1186);
nand U1797 (N_1797,N_23,N_1481);
and U1798 (N_1798,N_133,N_688);
or U1799 (N_1799,N_749,N_802);
nand U1800 (N_1800,N_20,N_267);
nor U1801 (N_1801,N_215,N_77);
and U1802 (N_1802,N_981,N_31);
nand U1803 (N_1803,N_47,N_544);
nand U1804 (N_1804,N_216,N_1295);
nor U1805 (N_1805,N_212,N_60);
nand U1806 (N_1806,N_1259,N_1108);
nand U1807 (N_1807,N_926,N_789);
xnor U1808 (N_1808,N_1353,N_1426);
nor U1809 (N_1809,N_740,N_265);
or U1810 (N_1810,N_690,N_588);
or U1811 (N_1811,N_746,N_757);
or U1812 (N_1812,N_1484,N_1464);
and U1813 (N_1813,N_903,N_770);
nand U1814 (N_1814,N_18,N_532);
and U1815 (N_1815,N_547,N_408);
or U1816 (N_1816,N_633,N_1138);
or U1817 (N_1817,N_360,N_872);
and U1818 (N_1818,N_217,N_1348);
or U1819 (N_1819,N_1033,N_168);
nor U1820 (N_1820,N_83,N_127);
nor U1821 (N_1821,N_340,N_1166);
nand U1822 (N_1822,N_1002,N_893);
or U1823 (N_1823,N_529,N_1434);
or U1824 (N_1824,N_19,N_373);
xor U1825 (N_1825,N_678,N_866);
or U1826 (N_1826,N_149,N_1494);
nor U1827 (N_1827,N_58,N_715);
or U1828 (N_1828,N_326,N_1332);
or U1829 (N_1829,N_1238,N_732);
and U1830 (N_1830,N_1341,N_1101);
xnor U1831 (N_1831,N_1445,N_150);
nand U1832 (N_1832,N_330,N_27);
nor U1833 (N_1833,N_1107,N_308);
or U1834 (N_1834,N_1042,N_1104);
nand U1835 (N_1835,N_810,N_1408);
nand U1836 (N_1836,N_1053,N_1065);
or U1837 (N_1837,N_793,N_1144);
nor U1838 (N_1838,N_103,N_1450);
and U1839 (N_1839,N_1474,N_1263);
and U1840 (N_1840,N_1455,N_1395);
or U1841 (N_1841,N_629,N_288);
nor U1842 (N_1842,N_1347,N_630);
xor U1843 (N_1843,N_601,N_569);
nand U1844 (N_1844,N_730,N_1264);
or U1845 (N_1845,N_686,N_280);
and U1846 (N_1846,N_256,N_993);
and U1847 (N_1847,N_365,N_1159);
nand U1848 (N_1848,N_52,N_1459);
nor U1849 (N_1849,N_1326,N_1126);
and U1850 (N_1850,N_1180,N_1142);
nor U1851 (N_1851,N_1273,N_1289);
nor U1852 (N_1852,N_78,N_190);
nand U1853 (N_1853,N_901,N_525);
and U1854 (N_1854,N_450,N_772);
nand U1855 (N_1855,N_148,N_389);
nand U1856 (N_1856,N_747,N_369);
nand U1857 (N_1857,N_946,N_830);
nor U1858 (N_1858,N_1414,N_143);
or U1859 (N_1859,N_1366,N_260);
nor U1860 (N_1860,N_1319,N_1113);
xor U1861 (N_1861,N_447,N_624);
and U1862 (N_1862,N_587,N_230);
and U1863 (N_1863,N_1109,N_1195);
or U1864 (N_1864,N_659,N_790);
and U1865 (N_1865,N_322,N_1229);
nor U1866 (N_1866,N_938,N_768);
nand U1867 (N_1867,N_693,N_669);
or U1868 (N_1868,N_142,N_495);
nand U1869 (N_1869,N_497,N_226);
nand U1870 (N_1870,N_467,N_1267);
nor U1871 (N_1871,N_1398,N_1465);
and U1872 (N_1872,N_837,N_1343);
and U1873 (N_1873,N_1471,N_1116);
or U1874 (N_1874,N_555,N_1124);
nand U1875 (N_1875,N_724,N_343);
or U1876 (N_1876,N_192,N_1139);
nand U1877 (N_1877,N_1014,N_1155);
nand U1878 (N_1878,N_289,N_439);
nand U1879 (N_1879,N_1261,N_1430);
nor U1880 (N_1880,N_94,N_180);
and U1881 (N_1881,N_485,N_281);
nand U1882 (N_1882,N_337,N_1081);
and U1883 (N_1883,N_642,N_320);
nor U1884 (N_1884,N_225,N_454);
xor U1885 (N_1885,N_535,N_1281);
and U1886 (N_1886,N_1411,N_1336);
and U1887 (N_1887,N_1390,N_328);
nand U1888 (N_1888,N_1246,N_1441);
and U1889 (N_1889,N_1106,N_481);
nand U1890 (N_1890,N_756,N_706);
nand U1891 (N_1891,N_722,N_1483);
and U1892 (N_1892,N_745,N_335);
xor U1893 (N_1893,N_1387,N_53);
nand U1894 (N_1894,N_834,N_1120);
or U1895 (N_1895,N_813,N_14);
or U1896 (N_1896,N_479,N_1090);
nand U1897 (N_1897,N_1205,N_917);
nor U1898 (N_1898,N_35,N_985);
nor U1899 (N_1899,N_855,N_646);
nor U1900 (N_1900,N_1206,N_93);
nand U1901 (N_1901,N_664,N_382);
nor U1902 (N_1902,N_123,N_137);
and U1903 (N_1903,N_666,N_1438);
xor U1904 (N_1904,N_1247,N_1305);
nor U1905 (N_1905,N_155,N_679);
nand U1906 (N_1906,N_1153,N_743);
nand U1907 (N_1907,N_2,N_176);
or U1908 (N_1908,N_1486,N_1202);
nand U1909 (N_1909,N_317,N_1217);
nor U1910 (N_1910,N_121,N_861);
or U1911 (N_1911,N_206,N_163);
nor U1912 (N_1912,N_1169,N_1097);
and U1913 (N_1913,N_438,N_598);
nor U1914 (N_1914,N_1185,N_735);
nor U1915 (N_1915,N_1252,N_879);
and U1916 (N_1916,N_1027,N_1284);
and U1917 (N_1917,N_904,N_1212);
nor U1918 (N_1918,N_461,N_1404);
and U1919 (N_1919,N_518,N_1346);
nand U1920 (N_1920,N_368,N_933);
nor U1921 (N_1921,N_1302,N_413);
or U1922 (N_1922,N_939,N_86);
nor U1923 (N_1923,N_1364,N_1447);
and U1924 (N_1924,N_114,N_1293);
nor U1925 (N_1925,N_867,N_354);
nand U1926 (N_1926,N_1298,N_219);
or U1927 (N_1927,N_196,N_195);
nand U1928 (N_1928,N_375,N_1086);
or U1929 (N_1929,N_178,N_536);
and U1930 (N_1930,N_817,N_957);
or U1931 (N_1931,N_472,N_1265);
xor U1932 (N_1932,N_967,N_1045);
nor U1933 (N_1933,N_840,N_1231);
nand U1934 (N_1934,N_1384,N_586);
or U1935 (N_1935,N_441,N_1244);
and U1936 (N_1936,N_325,N_538);
or U1937 (N_1937,N_400,N_111);
or U1938 (N_1938,N_1371,N_531);
and U1939 (N_1939,N_1334,N_282);
nor U1940 (N_1940,N_351,N_540);
nor U1941 (N_1941,N_1051,N_1171);
nand U1942 (N_1942,N_385,N_156);
and U1943 (N_1943,N_996,N_1068);
and U1944 (N_1944,N_886,N_1000);
and U1945 (N_1945,N_640,N_170);
or U1946 (N_1946,N_1337,N_394);
nand U1947 (N_1947,N_1088,N_1199);
nand U1948 (N_1948,N_1074,N_303);
nand U1949 (N_1949,N_274,N_372);
xnor U1950 (N_1950,N_21,N_1083);
or U1951 (N_1951,N_102,N_15);
and U1952 (N_1952,N_1007,N_422);
nor U1953 (N_1953,N_697,N_132);
xnor U1954 (N_1954,N_1087,N_1344);
or U1955 (N_1955,N_140,N_1242);
or U1956 (N_1956,N_429,N_1105);
or U1957 (N_1957,N_209,N_498);
and U1958 (N_1958,N_468,N_420);
or U1959 (N_1959,N_781,N_68);
and U1960 (N_1960,N_1396,N_978);
xnor U1961 (N_1961,N_188,N_477);
nor U1962 (N_1962,N_563,N_1470);
xnor U1963 (N_1963,N_66,N_1303);
or U1964 (N_1964,N_278,N_436);
nor U1965 (N_1965,N_409,N_1102);
nor U1966 (N_1966,N_1146,N_973);
nor U1967 (N_1967,N_406,N_491);
or U1968 (N_1968,N_997,N_44);
nor U1969 (N_1969,N_1082,N_313);
and U1970 (N_1970,N_1170,N_13);
xnor U1971 (N_1971,N_1041,N_910);
nand U1972 (N_1972,N_618,N_153);
nand U1973 (N_1973,N_1352,N_381);
nand U1974 (N_1974,N_1254,N_1022);
or U1975 (N_1975,N_1290,N_844);
and U1976 (N_1976,N_546,N_960);
xor U1977 (N_1977,N_884,N_99);
nor U1978 (N_1978,N_17,N_197);
and U1979 (N_1979,N_383,N_609);
nand U1980 (N_1980,N_1313,N_1137);
nor U1981 (N_1981,N_1164,N_815);
nor U1982 (N_1982,N_224,N_391);
and U1983 (N_1983,N_541,N_959);
and U1984 (N_1984,N_761,N_634);
and U1985 (N_1985,N_651,N_913);
nand U1986 (N_1986,N_1314,N_334);
nand U1987 (N_1987,N_1361,N_963);
or U1988 (N_1988,N_858,N_90);
nor U1989 (N_1989,N_528,N_783);
nor U1990 (N_1990,N_300,N_465);
and U1991 (N_1991,N_110,N_902);
and U1992 (N_1992,N_779,N_1010);
and U1993 (N_1993,N_1143,N_1327);
or U1994 (N_1994,N_1099,N_208);
or U1995 (N_1995,N_207,N_769);
nor U1996 (N_1996,N_384,N_1135);
or U1997 (N_1997,N_731,N_1067);
and U1998 (N_1998,N_1215,N_1439);
xnor U1999 (N_1999,N_738,N_1052);
nor U2000 (N_2000,N_554,N_637);
and U2001 (N_2001,N_663,N_1029);
nand U2002 (N_2002,N_809,N_961);
nand U2003 (N_2003,N_597,N_823);
nand U2004 (N_2004,N_811,N_899);
nand U2005 (N_2005,N_583,N_773);
and U2006 (N_2006,N_1363,N_874);
nand U2007 (N_2007,N_739,N_1493);
nor U2008 (N_2008,N_437,N_1151);
nand U2009 (N_2009,N_782,N_1066);
nor U2010 (N_2010,N_1422,N_187);
and U2011 (N_2011,N_488,N_119);
nand U2012 (N_2012,N_1342,N_558);
xor U2013 (N_2013,N_1467,N_1179);
xor U2014 (N_2014,N_1429,N_1056);
nor U2015 (N_2015,N_1131,N_1100);
and U2016 (N_2016,N_1221,N_510);
nand U2017 (N_2017,N_526,N_1241);
nor U2018 (N_2018,N_1026,N_480);
and U2019 (N_2019,N_628,N_1085);
nand U2020 (N_2020,N_1141,N_167);
or U2021 (N_2021,N_87,N_1416);
nor U2022 (N_2022,N_64,N_214);
nand U2023 (N_2023,N_1112,N_1093);
or U2024 (N_2024,N_51,N_459);
or U2025 (N_2025,N_622,N_744);
or U2026 (N_2026,N_1287,N_136);
nor U2027 (N_2027,N_104,N_998);
xor U2028 (N_2028,N_390,N_1357);
nor U2029 (N_2029,N_1362,N_1084);
nand U2030 (N_2030,N_258,N_1080);
or U2031 (N_2031,N_1331,N_1248);
xor U2032 (N_2032,N_1057,N_604);
and U2033 (N_2033,N_942,N_1288);
nor U2034 (N_2034,N_816,N_1176);
and U2035 (N_2035,N_552,N_698);
xnor U2036 (N_2036,N_202,N_4);
xor U2037 (N_2037,N_415,N_1392);
nand U2038 (N_2038,N_1360,N_658);
nor U2039 (N_2039,N_476,N_1355);
nor U2040 (N_2040,N_750,N_1400);
nor U2041 (N_2041,N_891,N_283);
nor U2042 (N_2042,N_1485,N_1379);
and U2043 (N_2043,N_945,N_1260);
and U2044 (N_2044,N_484,N_105);
and U2045 (N_2045,N_131,N_310);
nor U2046 (N_2046,N_117,N_1156);
or U2047 (N_2047,N_831,N_458);
nand U2048 (N_2048,N_1036,N_656);
or U2049 (N_2049,N_160,N_1306);
nor U2050 (N_2050,N_1078,N_792);
and U2051 (N_2051,N_233,N_603);
or U2052 (N_2052,N_1210,N_888);
xnor U2053 (N_2053,N_262,N_446);
nand U2054 (N_2054,N_315,N_97);
or U2055 (N_2055,N_221,N_157);
and U2056 (N_2056,N_841,N_205);
or U2057 (N_2057,N_1012,N_621);
nand U2058 (N_2058,N_108,N_507);
nand U2059 (N_2059,N_427,N_1224);
and U2060 (N_2060,N_760,N_752);
nor U2061 (N_2061,N_41,N_573);
nand U2062 (N_2062,N_503,N_486);
nor U2063 (N_2063,N_1,N_1245);
and U2064 (N_2064,N_846,N_79);
and U2065 (N_2065,N_704,N_509);
or U2066 (N_2066,N_252,N_1456);
nor U2067 (N_2067,N_753,N_284);
nand U2068 (N_2068,N_852,N_1417);
and U2069 (N_2069,N_1098,N_1172);
or U2070 (N_2070,N_444,N_1477);
nand U2071 (N_2071,N_449,N_483);
and U2072 (N_2072,N_983,N_1297);
nor U2073 (N_2073,N_1134,N_952);
nand U2074 (N_2074,N_1276,N_45);
or U2075 (N_2075,N_36,N_259);
or U2076 (N_2076,N_286,N_1111);
and U2077 (N_2077,N_411,N_1228);
and U2078 (N_2078,N_705,N_1167);
and U2079 (N_2079,N_1094,N_1469);
nand U2080 (N_2080,N_584,N_57);
nand U2081 (N_2081,N_742,N_5);
nand U2082 (N_2082,N_1458,N_1058);
or U2083 (N_2083,N_88,N_803);
or U2084 (N_2084,N_445,N_721);
xor U2085 (N_2085,N_620,N_1280);
and U2086 (N_2086,N_971,N_1161);
nand U2087 (N_2087,N_91,N_1043);
nand U2088 (N_2088,N_718,N_1201);
xnor U2089 (N_2089,N_1047,N_1220);
nor U2090 (N_2090,N_363,N_979);
nand U2091 (N_2091,N_923,N_652);
or U2092 (N_2092,N_154,N_962);
or U2093 (N_2093,N_508,N_723);
and U2094 (N_2094,N_227,N_139);
and U2095 (N_2095,N_332,N_850);
xnor U2096 (N_2096,N_1234,N_734);
nor U2097 (N_2097,N_194,N_1223);
or U2098 (N_2098,N_1487,N_231);
nor U2099 (N_2099,N_717,N_548);
and U2100 (N_2100,N_829,N_949);
nor U2101 (N_2101,N_399,N_318);
and U2102 (N_2102,N_860,N_1091);
or U2103 (N_2103,N_1372,N_577);
nor U2104 (N_2104,N_680,N_184);
nand U2105 (N_2105,N_1175,N_838);
nor U2106 (N_2106,N_896,N_62);
and U2107 (N_2107,N_199,N_1233);
nand U2108 (N_2108,N_1250,N_452);
nor U2109 (N_2109,N_593,N_543);
and U2110 (N_2110,N_1182,N_1277);
and U2111 (N_2111,N_865,N_638);
or U2112 (N_2112,N_972,N_314);
nand U2113 (N_2113,N_1114,N_1268);
or U2114 (N_2114,N_694,N_63);
and U2115 (N_2115,N_847,N_512);
or U2116 (N_2116,N_542,N_423);
and U2117 (N_2117,N_635,N_392);
nand U2118 (N_2118,N_1227,N_672);
and U2119 (N_2119,N_610,N_1403);
nor U2120 (N_2120,N_754,N_709);
and U2121 (N_2121,N_175,N_1055);
and U2122 (N_2122,N_1449,N_887);
nand U2123 (N_2123,N_1076,N_285);
xnor U2124 (N_2124,N_134,N_490);
xor U2125 (N_2125,N_1358,N_799);
nor U2126 (N_2126,N_1128,N_499);
nand U2127 (N_2127,N_791,N_398);
nand U2128 (N_2128,N_417,N_222);
xor U2129 (N_2129,N_255,N_122);
and U2130 (N_2130,N_1432,N_419);
or U2131 (N_2131,N_7,N_1177);
and U2132 (N_2132,N_1498,N_827);
nand U2133 (N_2133,N_1490,N_737);
and U2134 (N_2134,N_1257,N_1460);
or U2135 (N_2135,N_741,N_517);
and U2136 (N_2136,N_218,N_1399);
or U2137 (N_2137,N_451,N_948);
and U2138 (N_2138,N_1157,N_936);
or U2139 (N_2139,N_347,N_75);
xnor U2140 (N_2140,N_561,N_359);
nand U2141 (N_2141,N_1095,N_851);
nor U2142 (N_2142,N_1316,N_198);
nor U2143 (N_2143,N_871,N_1044);
or U2144 (N_2144,N_801,N_763);
nor U2145 (N_2145,N_645,N_1148);
nor U2146 (N_2146,N_30,N_43);
or U2147 (N_2147,N_333,N_1283);
nor U2148 (N_2148,N_725,N_297);
nor U2149 (N_2149,N_1325,N_302);
or U2150 (N_2150,N_1286,N_613);
or U2151 (N_2151,N_1282,N_1030);
nor U2152 (N_2152,N_1226,N_982);
nand U2153 (N_2153,N_1178,N_49);
nor U2154 (N_2154,N_32,N_39);
or U2155 (N_2155,N_924,N_487);
and U2156 (N_2156,N_364,N_460);
nor U2157 (N_2157,N_1370,N_944);
xnor U2158 (N_2158,N_701,N_1453);
or U2159 (N_2159,N_853,N_268);
nor U2160 (N_2160,N_185,N_1218);
and U2161 (N_2161,N_665,N_1222);
or U2162 (N_2162,N_627,N_405);
nor U2163 (N_2163,N_42,N_1129);
or U2164 (N_2164,N_3,N_798);
and U2165 (N_2165,N_191,N_1382);
or U2166 (N_2166,N_1216,N_842);
nor U2167 (N_2167,N_649,N_565);
nor U2168 (N_2168,N_95,N_612);
nor U2169 (N_2169,N_469,N_1225);
or U2170 (N_2170,N_189,N_1214);
and U2171 (N_2171,N_560,N_1497);
or U2172 (N_2172,N_273,N_1008);
nor U2173 (N_2173,N_808,N_1473);
and U2174 (N_2174,N_59,N_1365);
and U2175 (N_2175,N_1117,N_934);
nor U2176 (N_2176,N_549,N_1437);
nor U2177 (N_2177,N_515,N_968);
nand U2178 (N_2178,N_898,N_376);
nand U2179 (N_2179,N_885,N_606);
nor U2180 (N_2180,N_279,N_1472);
nand U2181 (N_2181,N_825,N_1270);
nor U2182 (N_2182,N_263,N_1431);
and U2183 (N_2183,N_34,N_138);
nor U2184 (N_2184,N_826,N_1118);
nand U2185 (N_2185,N_987,N_388);
and U2186 (N_2186,N_473,N_1476);
nor U2187 (N_2187,N_1004,N_814);
nand U2188 (N_2188,N_1440,N_599);
or U2189 (N_2189,N_919,N_100);
and U2190 (N_2190,N_271,N_327);
nor U2191 (N_2191,N_76,N_240);
and U2192 (N_2192,N_1323,N_48);
and U2193 (N_2193,N_1039,N_661);
nand U2194 (N_2194,N_572,N_787);
and U2195 (N_2195,N_1463,N_1271);
nor U2196 (N_2196,N_1054,N_1279);
or U2197 (N_2197,N_371,N_590);
and U2198 (N_2198,N_181,N_37);
xnor U2199 (N_2199,N_1162,N_378);
nand U2200 (N_2200,N_1262,N_1479);
or U2201 (N_2201,N_404,N_687);
nor U2202 (N_2202,N_895,N_632);
or U2203 (N_2203,N_537,N_421);
nand U2204 (N_2204,N_615,N_1038);
or U2205 (N_2205,N_519,N_210);
nor U2206 (N_2206,N_1335,N_1354);
or U2207 (N_2207,N_820,N_193);
xnor U2208 (N_2208,N_1168,N_493);
and U2209 (N_2209,N_1299,N_379);
or U2210 (N_2210,N_930,N_453);
nand U2211 (N_2211,N_367,N_1003);
nor U2212 (N_2212,N_241,N_1492);
nor U2213 (N_2213,N_1147,N_246);
or U2214 (N_2214,N_908,N_1136);
nor U2215 (N_2215,N_849,N_591);
nor U2216 (N_2216,N_38,N_203);
or U2217 (N_2217,N_516,N_1115);
or U2218 (N_2218,N_576,N_1213);
nor U2219 (N_2219,N_1209,N_291);
xor U2220 (N_2220,N_670,N_1154);
nand U2221 (N_2221,N_301,N_1285);
nand U2222 (N_2222,N_1317,N_242);
nand U2223 (N_2223,N_173,N_1021);
xor U2224 (N_2224,N_1368,N_854);
or U2225 (N_2225,N_130,N_1243);
or U2226 (N_2226,N_200,N_921);
and U2227 (N_2227,N_186,N_580);
nand U2228 (N_2228,N_424,N_1253);
and U2229 (N_2229,N_812,N_1196);
nor U2230 (N_2230,N_870,N_323);
nand U2231 (N_2231,N_299,N_69);
and U2232 (N_2232,N_1301,N_266);
xnor U2233 (N_2233,N_1294,N_386);
nand U2234 (N_2234,N_1320,N_1251);
or U2235 (N_2235,N_455,N_55);
and U2236 (N_2236,N_1072,N_126);
nand U2237 (N_2237,N_1125,N_1423);
and U2238 (N_2238,N_1173,N_234);
nand U2239 (N_2239,N_1451,N_443);
and U2240 (N_2240,N_568,N_118);
and U2241 (N_2241,N_1442,N_128);
nor U2242 (N_2242,N_641,N_986);
nor U2243 (N_2243,N_457,N_1077);
xor U2244 (N_2244,N_927,N_1339);
nand U2245 (N_2245,N_287,N_65);
or U2246 (N_2246,N_1121,N_1070);
or U2247 (N_2247,N_941,N_1435);
nor U2248 (N_2248,N_342,N_305);
nor U2249 (N_2249,N_928,N_976);
nor U2250 (N_2250,N_609,N_1223);
or U2251 (N_2251,N_1006,N_98);
and U2252 (N_2252,N_814,N_349);
nor U2253 (N_2253,N_285,N_666);
and U2254 (N_2254,N_278,N_1114);
nor U2255 (N_2255,N_1057,N_351);
xnor U2256 (N_2256,N_973,N_1036);
or U2257 (N_2257,N_630,N_1182);
and U2258 (N_2258,N_572,N_1013);
and U2259 (N_2259,N_1045,N_1375);
and U2260 (N_2260,N_8,N_29);
and U2261 (N_2261,N_249,N_687);
and U2262 (N_2262,N_1027,N_1207);
xor U2263 (N_2263,N_542,N_260);
or U2264 (N_2264,N_679,N_81);
or U2265 (N_2265,N_46,N_372);
nand U2266 (N_2266,N_543,N_425);
xnor U2267 (N_2267,N_1442,N_386);
or U2268 (N_2268,N_1113,N_1067);
and U2269 (N_2269,N_784,N_1451);
nand U2270 (N_2270,N_651,N_1163);
xor U2271 (N_2271,N_317,N_1314);
and U2272 (N_2272,N_184,N_832);
or U2273 (N_2273,N_1252,N_675);
nand U2274 (N_2274,N_1189,N_872);
nor U2275 (N_2275,N_373,N_638);
xor U2276 (N_2276,N_5,N_856);
and U2277 (N_2277,N_1135,N_94);
nor U2278 (N_2278,N_528,N_859);
xor U2279 (N_2279,N_561,N_332);
and U2280 (N_2280,N_1053,N_1320);
or U2281 (N_2281,N_92,N_1371);
xnor U2282 (N_2282,N_139,N_1230);
nand U2283 (N_2283,N_896,N_1401);
and U2284 (N_2284,N_1113,N_29);
nand U2285 (N_2285,N_807,N_336);
and U2286 (N_2286,N_1366,N_1334);
nand U2287 (N_2287,N_631,N_432);
or U2288 (N_2288,N_1489,N_416);
nor U2289 (N_2289,N_1193,N_838);
or U2290 (N_2290,N_687,N_1211);
and U2291 (N_2291,N_959,N_614);
nand U2292 (N_2292,N_928,N_464);
and U2293 (N_2293,N_942,N_1299);
xor U2294 (N_2294,N_637,N_1408);
nand U2295 (N_2295,N_137,N_909);
xnor U2296 (N_2296,N_270,N_975);
nor U2297 (N_2297,N_117,N_579);
or U2298 (N_2298,N_796,N_104);
or U2299 (N_2299,N_142,N_849);
or U2300 (N_2300,N_2,N_921);
xor U2301 (N_2301,N_334,N_396);
or U2302 (N_2302,N_1481,N_1384);
and U2303 (N_2303,N_1359,N_208);
nor U2304 (N_2304,N_90,N_1066);
or U2305 (N_2305,N_363,N_1422);
or U2306 (N_2306,N_648,N_152);
nor U2307 (N_2307,N_694,N_1356);
and U2308 (N_2308,N_15,N_697);
nand U2309 (N_2309,N_1091,N_1314);
nand U2310 (N_2310,N_1322,N_452);
and U2311 (N_2311,N_1069,N_1268);
nand U2312 (N_2312,N_1265,N_1036);
or U2313 (N_2313,N_250,N_184);
and U2314 (N_2314,N_1057,N_346);
nand U2315 (N_2315,N_553,N_787);
or U2316 (N_2316,N_352,N_229);
nor U2317 (N_2317,N_158,N_1382);
or U2318 (N_2318,N_493,N_1303);
and U2319 (N_2319,N_261,N_989);
nor U2320 (N_2320,N_278,N_1009);
nand U2321 (N_2321,N_1475,N_144);
or U2322 (N_2322,N_545,N_1246);
and U2323 (N_2323,N_859,N_1466);
nand U2324 (N_2324,N_1027,N_1000);
xnor U2325 (N_2325,N_701,N_377);
and U2326 (N_2326,N_1101,N_1084);
nor U2327 (N_2327,N_20,N_756);
and U2328 (N_2328,N_651,N_841);
and U2329 (N_2329,N_1000,N_979);
or U2330 (N_2330,N_627,N_1120);
nand U2331 (N_2331,N_970,N_1392);
nand U2332 (N_2332,N_1122,N_949);
and U2333 (N_2333,N_477,N_620);
nor U2334 (N_2334,N_1424,N_390);
nor U2335 (N_2335,N_1115,N_503);
and U2336 (N_2336,N_156,N_1060);
nor U2337 (N_2337,N_1278,N_1376);
and U2338 (N_2338,N_189,N_228);
or U2339 (N_2339,N_910,N_1492);
and U2340 (N_2340,N_1203,N_1128);
xnor U2341 (N_2341,N_405,N_860);
and U2342 (N_2342,N_398,N_1327);
or U2343 (N_2343,N_1312,N_1142);
nand U2344 (N_2344,N_1433,N_1232);
or U2345 (N_2345,N_626,N_1453);
nor U2346 (N_2346,N_872,N_401);
and U2347 (N_2347,N_1350,N_613);
nand U2348 (N_2348,N_49,N_1419);
nor U2349 (N_2349,N_1497,N_163);
nand U2350 (N_2350,N_236,N_1064);
nor U2351 (N_2351,N_119,N_1445);
or U2352 (N_2352,N_915,N_1024);
or U2353 (N_2353,N_1076,N_405);
and U2354 (N_2354,N_120,N_18);
nand U2355 (N_2355,N_970,N_681);
and U2356 (N_2356,N_725,N_239);
xor U2357 (N_2357,N_999,N_948);
and U2358 (N_2358,N_627,N_1396);
nor U2359 (N_2359,N_919,N_807);
or U2360 (N_2360,N_455,N_1315);
xnor U2361 (N_2361,N_1077,N_389);
nand U2362 (N_2362,N_111,N_806);
or U2363 (N_2363,N_1155,N_644);
or U2364 (N_2364,N_1382,N_942);
nand U2365 (N_2365,N_674,N_717);
nor U2366 (N_2366,N_1052,N_1398);
and U2367 (N_2367,N_202,N_598);
nor U2368 (N_2368,N_3,N_1098);
nand U2369 (N_2369,N_1163,N_1035);
nor U2370 (N_2370,N_782,N_1432);
and U2371 (N_2371,N_156,N_1349);
xnor U2372 (N_2372,N_587,N_1273);
nor U2373 (N_2373,N_1326,N_682);
and U2374 (N_2374,N_758,N_1323);
and U2375 (N_2375,N_1117,N_284);
xor U2376 (N_2376,N_180,N_1434);
and U2377 (N_2377,N_835,N_752);
nor U2378 (N_2378,N_94,N_869);
nand U2379 (N_2379,N_913,N_675);
xor U2380 (N_2380,N_530,N_1435);
or U2381 (N_2381,N_1356,N_551);
nor U2382 (N_2382,N_774,N_406);
nor U2383 (N_2383,N_1350,N_1421);
nand U2384 (N_2384,N_1188,N_1183);
nand U2385 (N_2385,N_626,N_428);
and U2386 (N_2386,N_277,N_147);
nand U2387 (N_2387,N_325,N_805);
or U2388 (N_2388,N_928,N_1366);
nand U2389 (N_2389,N_89,N_374);
or U2390 (N_2390,N_38,N_399);
xnor U2391 (N_2391,N_396,N_335);
nand U2392 (N_2392,N_149,N_57);
or U2393 (N_2393,N_677,N_1084);
and U2394 (N_2394,N_1289,N_1170);
xor U2395 (N_2395,N_1242,N_617);
nor U2396 (N_2396,N_620,N_596);
nand U2397 (N_2397,N_835,N_1045);
nand U2398 (N_2398,N_1363,N_1321);
nand U2399 (N_2399,N_860,N_1102);
xnor U2400 (N_2400,N_628,N_179);
nor U2401 (N_2401,N_896,N_1036);
and U2402 (N_2402,N_1309,N_695);
or U2403 (N_2403,N_951,N_1311);
and U2404 (N_2404,N_1118,N_894);
xnor U2405 (N_2405,N_593,N_1003);
or U2406 (N_2406,N_35,N_297);
xnor U2407 (N_2407,N_211,N_252);
or U2408 (N_2408,N_616,N_1370);
nand U2409 (N_2409,N_1430,N_447);
and U2410 (N_2410,N_5,N_990);
nor U2411 (N_2411,N_366,N_115);
or U2412 (N_2412,N_1421,N_622);
nor U2413 (N_2413,N_527,N_285);
or U2414 (N_2414,N_603,N_1373);
nor U2415 (N_2415,N_353,N_400);
xor U2416 (N_2416,N_758,N_115);
nor U2417 (N_2417,N_448,N_868);
nand U2418 (N_2418,N_48,N_706);
nor U2419 (N_2419,N_1465,N_1313);
and U2420 (N_2420,N_924,N_702);
and U2421 (N_2421,N_1389,N_184);
xor U2422 (N_2422,N_404,N_1476);
nand U2423 (N_2423,N_1141,N_1424);
and U2424 (N_2424,N_994,N_1387);
or U2425 (N_2425,N_1203,N_1323);
nand U2426 (N_2426,N_993,N_67);
nand U2427 (N_2427,N_581,N_746);
nor U2428 (N_2428,N_131,N_17);
nand U2429 (N_2429,N_750,N_815);
nand U2430 (N_2430,N_1481,N_1294);
nor U2431 (N_2431,N_292,N_1186);
xor U2432 (N_2432,N_1025,N_1287);
and U2433 (N_2433,N_774,N_255);
or U2434 (N_2434,N_476,N_728);
nand U2435 (N_2435,N_28,N_486);
or U2436 (N_2436,N_848,N_35);
or U2437 (N_2437,N_538,N_503);
and U2438 (N_2438,N_1321,N_233);
nand U2439 (N_2439,N_540,N_1037);
nor U2440 (N_2440,N_1387,N_700);
nor U2441 (N_2441,N_1239,N_1437);
and U2442 (N_2442,N_909,N_1272);
or U2443 (N_2443,N_502,N_112);
nand U2444 (N_2444,N_488,N_691);
and U2445 (N_2445,N_697,N_582);
xor U2446 (N_2446,N_785,N_530);
or U2447 (N_2447,N_120,N_229);
or U2448 (N_2448,N_585,N_85);
and U2449 (N_2449,N_883,N_599);
or U2450 (N_2450,N_276,N_1215);
nand U2451 (N_2451,N_1408,N_874);
or U2452 (N_2452,N_892,N_179);
nor U2453 (N_2453,N_49,N_468);
or U2454 (N_2454,N_1015,N_119);
nor U2455 (N_2455,N_1032,N_277);
and U2456 (N_2456,N_40,N_497);
nor U2457 (N_2457,N_1353,N_1398);
nor U2458 (N_2458,N_1461,N_1265);
nand U2459 (N_2459,N_724,N_998);
or U2460 (N_2460,N_712,N_252);
or U2461 (N_2461,N_849,N_96);
and U2462 (N_2462,N_297,N_179);
nor U2463 (N_2463,N_221,N_240);
or U2464 (N_2464,N_497,N_980);
or U2465 (N_2465,N_1261,N_409);
xnor U2466 (N_2466,N_864,N_102);
xnor U2467 (N_2467,N_586,N_0);
nor U2468 (N_2468,N_1180,N_1492);
and U2469 (N_2469,N_1018,N_1235);
and U2470 (N_2470,N_452,N_502);
nor U2471 (N_2471,N_1311,N_828);
xnor U2472 (N_2472,N_1014,N_1411);
nor U2473 (N_2473,N_1224,N_146);
nor U2474 (N_2474,N_357,N_1342);
or U2475 (N_2475,N_511,N_1225);
nand U2476 (N_2476,N_556,N_198);
or U2477 (N_2477,N_1409,N_317);
nor U2478 (N_2478,N_418,N_258);
nor U2479 (N_2479,N_20,N_1101);
and U2480 (N_2480,N_1400,N_545);
nand U2481 (N_2481,N_1117,N_1207);
xor U2482 (N_2482,N_1001,N_981);
xnor U2483 (N_2483,N_124,N_1074);
nor U2484 (N_2484,N_514,N_1381);
nand U2485 (N_2485,N_849,N_668);
xor U2486 (N_2486,N_1075,N_143);
nand U2487 (N_2487,N_1137,N_812);
xnor U2488 (N_2488,N_679,N_1216);
nand U2489 (N_2489,N_1392,N_1325);
or U2490 (N_2490,N_785,N_1005);
and U2491 (N_2491,N_502,N_1220);
and U2492 (N_2492,N_1332,N_973);
nand U2493 (N_2493,N_1099,N_1169);
nand U2494 (N_2494,N_951,N_300);
nor U2495 (N_2495,N_1102,N_937);
or U2496 (N_2496,N_1175,N_521);
and U2497 (N_2497,N_677,N_533);
nor U2498 (N_2498,N_929,N_857);
or U2499 (N_2499,N_502,N_1495);
and U2500 (N_2500,N_3,N_601);
nand U2501 (N_2501,N_109,N_131);
nor U2502 (N_2502,N_1253,N_1217);
and U2503 (N_2503,N_387,N_813);
nand U2504 (N_2504,N_654,N_1299);
or U2505 (N_2505,N_165,N_700);
nor U2506 (N_2506,N_129,N_1118);
xnor U2507 (N_2507,N_1299,N_1431);
xnor U2508 (N_2508,N_1072,N_2);
or U2509 (N_2509,N_983,N_1023);
and U2510 (N_2510,N_627,N_909);
nand U2511 (N_2511,N_441,N_222);
and U2512 (N_2512,N_981,N_126);
nand U2513 (N_2513,N_264,N_979);
nand U2514 (N_2514,N_9,N_1461);
or U2515 (N_2515,N_1226,N_1329);
or U2516 (N_2516,N_886,N_926);
and U2517 (N_2517,N_148,N_1121);
nand U2518 (N_2518,N_437,N_1166);
and U2519 (N_2519,N_1386,N_376);
or U2520 (N_2520,N_1137,N_1198);
or U2521 (N_2521,N_1147,N_1061);
and U2522 (N_2522,N_1480,N_1022);
nand U2523 (N_2523,N_1079,N_1445);
xnor U2524 (N_2524,N_862,N_1357);
and U2525 (N_2525,N_1365,N_1296);
and U2526 (N_2526,N_22,N_229);
nor U2527 (N_2527,N_1172,N_1475);
or U2528 (N_2528,N_407,N_235);
and U2529 (N_2529,N_1062,N_322);
or U2530 (N_2530,N_494,N_504);
nor U2531 (N_2531,N_63,N_1452);
xnor U2532 (N_2532,N_777,N_989);
and U2533 (N_2533,N_141,N_821);
nor U2534 (N_2534,N_570,N_1337);
or U2535 (N_2535,N_287,N_527);
or U2536 (N_2536,N_910,N_1137);
nand U2537 (N_2537,N_1072,N_231);
or U2538 (N_2538,N_1026,N_176);
or U2539 (N_2539,N_748,N_1394);
or U2540 (N_2540,N_602,N_1021);
nor U2541 (N_2541,N_395,N_110);
nor U2542 (N_2542,N_1319,N_841);
or U2543 (N_2543,N_220,N_1258);
and U2544 (N_2544,N_857,N_58);
nor U2545 (N_2545,N_128,N_835);
and U2546 (N_2546,N_537,N_392);
and U2547 (N_2547,N_146,N_283);
and U2548 (N_2548,N_574,N_860);
and U2549 (N_2549,N_153,N_1293);
or U2550 (N_2550,N_634,N_559);
xor U2551 (N_2551,N_1127,N_1481);
and U2552 (N_2552,N_745,N_612);
and U2553 (N_2553,N_1116,N_1268);
and U2554 (N_2554,N_931,N_1243);
and U2555 (N_2555,N_753,N_758);
nor U2556 (N_2556,N_746,N_681);
nor U2557 (N_2557,N_1272,N_630);
nor U2558 (N_2558,N_1222,N_519);
and U2559 (N_2559,N_24,N_552);
and U2560 (N_2560,N_70,N_942);
or U2561 (N_2561,N_907,N_1250);
nor U2562 (N_2562,N_458,N_532);
nand U2563 (N_2563,N_404,N_633);
or U2564 (N_2564,N_259,N_107);
xor U2565 (N_2565,N_1211,N_1344);
nor U2566 (N_2566,N_41,N_1004);
xnor U2567 (N_2567,N_1241,N_446);
and U2568 (N_2568,N_1136,N_225);
and U2569 (N_2569,N_769,N_858);
or U2570 (N_2570,N_1337,N_276);
nor U2571 (N_2571,N_397,N_831);
nor U2572 (N_2572,N_1054,N_782);
nand U2573 (N_2573,N_1088,N_493);
nor U2574 (N_2574,N_499,N_680);
nand U2575 (N_2575,N_384,N_126);
nor U2576 (N_2576,N_1034,N_262);
nand U2577 (N_2577,N_731,N_404);
and U2578 (N_2578,N_693,N_394);
and U2579 (N_2579,N_121,N_1215);
and U2580 (N_2580,N_1276,N_1066);
and U2581 (N_2581,N_1044,N_599);
nand U2582 (N_2582,N_574,N_1219);
or U2583 (N_2583,N_500,N_1023);
and U2584 (N_2584,N_23,N_965);
and U2585 (N_2585,N_335,N_1441);
or U2586 (N_2586,N_1338,N_1310);
nor U2587 (N_2587,N_84,N_1398);
or U2588 (N_2588,N_353,N_766);
or U2589 (N_2589,N_757,N_1230);
and U2590 (N_2590,N_1422,N_891);
nand U2591 (N_2591,N_1072,N_450);
nor U2592 (N_2592,N_174,N_171);
or U2593 (N_2593,N_1452,N_1480);
and U2594 (N_2594,N_1040,N_1395);
and U2595 (N_2595,N_985,N_415);
and U2596 (N_2596,N_335,N_123);
nand U2597 (N_2597,N_257,N_1018);
and U2598 (N_2598,N_1244,N_324);
nor U2599 (N_2599,N_908,N_101);
and U2600 (N_2600,N_1335,N_393);
or U2601 (N_2601,N_599,N_1068);
or U2602 (N_2602,N_1322,N_1363);
or U2603 (N_2603,N_726,N_724);
and U2604 (N_2604,N_207,N_891);
nand U2605 (N_2605,N_229,N_1020);
nand U2606 (N_2606,N_1188,N_25);
and U2607 (N_2607,N_1466,N_461);
nor U2608 (N_2608,N_1209,N_1486);
nand U2609 (N_2609,N_995,N_394);
nand U2610 (N_2610,N_457,N_33);
or U2611 (N_2611,N_33,N_1154);
or U2612 (N_2612,N_721,N_787);
and U2613 (N_2613,N_270,N_1434);
nand U2614 (N_2614,N_182,N_1170);
or U2615 (N_2615,N_1298,N_70);
and U2616 (N_2616,N_286,N_904);
nor U2617 (N_2617,N_951,N_559);
or U2618 (N_2618,N_654,N_509);
nand U2619 (N_2619,N_563,N_335);
nand U2620 (N_2620,N_1105,N_1495);
nand U2621 (N_2621,N_1192,N_1475);
and U2622 (N_2622,N_986,N_205);
and U2623 (N_2623,N_756,N_748);
nand U2624 (N_2624,N_712,N_215);
nor U2625 (N_2625,N_517,N_202);
nor U2626 (N_2626,N_1046,N_1020);
and U2627 (N_2627,N_867,N_620);
nand U2628 (N_2628,N_1464,N_476);
nor U2629 (N_2629,N_195,N_350);
and U2630 (N_2630,N_729,N_1145);
nor U2631 (N_2631,N_668,N_1167);
nand U2632 (N_2632,N_145,N_404);
or U2633 (N_2633,N_1179,N_468);
nor U2634 (N_2634,N_1467,N_818);
nand U2635 (N_2635,N_965,N_1333);
nor U2636 (N_2636,N_219,N_44);
and U2637 (N_2637,N_92,N_81);
or U2638 (N_2638,N_563,N_248);
and U2639 (N_2639,N_1234,N_53);
and U2640 (N_2640,N_42,N_97);
nor U2641 (N_2641,N_466,N_247);
and U2642 (N_2642,N_274,N_840);
or U2643 (N_2643,N_1170,N_1067);
and U2644 (N_2644,N_801,N_202);
nor U2645 (N_2645,N_697,N_104);
or U2646 (N_2646,N_1282,N_1370);
and U2647 (N_2647,N_983,N_934);
xnor U2648 (N_2648,N_1013,N_148);
nor U2649 (N_2649,N_1311,N_319);
xnor U2650 (N_2650,N_506,N_1324);
nand U2651 (N_2651,N_980,N_1297);
nor U2652 (N_2652,N_330,N_437);
nand U2653 (N_2653,N_1192,N_222);
or U2654 (N_2654,N_205,N_1325);
nand U2655 (N_2655,N_243,N_1034);
or U2656 (N_2656,N_1165,N_1140);
or U2657 (N_2657,N_299,N_786);
nor U2658 (N_2658,N_143,N_1278);
nand U2659 (N_2659,N_845,N_983);
or U2660 (N_2660,N_853,N_1153);
nor U2661 (N_2661,N_1424,N_388);
nor U2662 (N_2662,N_785,N_269);
nand U2663 (N_2663,N_763,N_412);
nor U2664 (N_2664,N_338,N_716);
nor U2665 (N_2665,N_1457,N_966);
nand U2666 (N_2666,N_317,N_1482);
nand U2667 (N_2667,N_1080,N_984);
and U2668 (N_2668,N_1322,N_1048);
or U2669 (N_2669,N_610,N_1170);
and U2670 (N_2670,N_1300,N_376);
nor U2671 (N_2671,N_774,N_1211);
nor U2672 (N_2672,N_761,N_1052);
xor U2673 (N_2673,N_521,N_1422);
and U2674 (N_2674,N_1170,N_151);
nand U2675 (N_2675,N_907,N_224);
nor U2676 (N_2676,N_1019,N_1335);
nand U2677 (N_2677,N_637,N_1478);
nor U2678 (N_2678,N_1282,N_248);
and U2679 (N_2679,N_829,N_995);
or U2680 (N_2680,N_268,N_1227);
xnor U2681 (N_2681,N_1402,N_1309);
or U2682 (N_2682,N_1385,N_949);
xnor U2683 (N_2683,N_98,N_27);
nor U2684 (N_2684,N_721,N_562);
nor U2685 (N_2685,N_74,N_978);
and U2686 (N_2686,N_614,N_65);
xnor U2687 (N_2687,N_1492,N_1233);
xor U2688 (N_2688,N_1263,N_79);
xor U2689 (N_2689,N_1086,N_975);
nor U2690 (N_2690,N_227,N_569);
and U2691 (N_2691,N_1182,N_533);
or U2692 (N_2692,N_1250,N_1453);
nand U2693 (N_2693,N_446,N_14);
or U2694 (N_2694,N_466,N_849);
nor U2695 (N_2695,N_361,N_300);
and U2696 (N_2696,N_1226,N_741);
xnor U2697 (N_2697,N_1258,N_787);
xor U2698 (N_2698,N_1059,N_835);
nand U2699 (N_2699,N_787,N_561);
or U2700 (N_2700,N_767,N_561);
or U2701 (N_2701,N_138,N_637);
and U2702 (N_2702,N_130,N_597);
or U2703 (N_2703,N_374,N_477);
nor U2704 (N_2704,N_1358,N_660);
nand U2705 (N_2705,N_1396,N_1153);
or U2706 (N_2706,N_1384,N_31);
nor U2707 (N_2707,N_644,N_41);
and U2708 (N_2708,N_1015,N_464);
nor U2709 (N_2709,N_927,N_1423);
and U2710 (N_2710,N_545,N_257);
nor U2711 (N_2711,N_387,N_1033);
and U2712 (N_2712,N_1410,N_141);
nand U2713 (N_2713,N_1090,N_1232);
or U2714 (N_2714,N_1079,N_206);
or U2715 (N_2715,N_786,N_969);
or U2716 (N_2716,N_360,N_285);
nand U2717 (N_2717,N_260,N_242);
nor U2718 (N_2718,N_756,N_961);
nand U2719 (N_2719,N_846,N_1383);
or U2720 (N_2720,N_759,N_23);
nor U2721 (N_2721,N_865,N_860);
or U2722 (N_2722,N_293,N_1310);
nor U2723 (N_2723,N_925,N_1138);
nand U2724 (N_2724,N_911,N_548);
nand U2725 (N_2725,N_421,N_936);
nand U2726 (N_2726,N_1458,N_1187);
and U2727 (N_2727,N_318,N_1440);
or U2728 (N_2728,N_335,N_800);
nand U2729 (N_2729,N_1246,N_1276);
nor U2730 (N_2730,N_1143,N_97);
nand U2731 (N_2731,N_740,N_1151);
or U2732 (N_2732,N_587,N_78);
nor U2733 (N_2733,N_728,N_1384);
or U2734 (N_2734,N_1400,N_752);
nor U2735 (N_2735,N_309,N_1285);
and U2736 (N_2736,N_484,N_1493);
xor U2737 (N_2737,N_1179,N_381);
nor U2738 (N_2738,N_400,N_562);
nor U2739 (N_2739,N_1342,N_811);
nor U2740 (N_2740,N_1473,N_1062);
nor U2741 (N_2741,N_1057,N_669);
and U2742 (N_2742,N_1032,N_862);
nor U2743 (N_2743,N_414,N_627);
xnor U2744 (N_2744,N_968,N_820);
nor U2745 (N_2745,N_183,N_478);
nor U2746 (N_2746,N_801,N_318);
xnor U2747 (N_2747,N_721,N_764);
nor U2748 (N_2748,N_477,N_1450);
xor U2749 (N_2749,N_385,N_403);
nand U2750 (N_2750,N_16,N_412);
and U2751 (N_2751,N_713,N_712);
nor U2752 (N_2752,N_1278,N_617);
or U2753 (N_2753,N_437,N_325);
and U2754 (N_2754,N_132,N_162);
nor U2755 (N_2755,N_1480,N_1267);
or U2756 (N_2756,N_535,N_559);
and U2757 (N_2757,N_1288,N_744);
and U2758 (N_2758,N_397,N_1087);
nand U2759 (N_2759,N_318,N_930);
and U2760 (N_2760,N_1288,N_2);
xor U2761 (N_2761,N_1472,N_905);
nor U2762 (N_2762,N_376,N_328);
nor U2763 (N_2763,N_643,N_561);
xnor U2764 (N_2764,N_1233,N_432);
xnor U2765 (N_2765,N_837,N_170);
or U2766 (N_2766,N_529,N_1175);
or U2767 (N_2767,N_815,N_1130);
nor U2768 (N_2768,N_390,N_1239);
and U2769 (N_2769,N_1414,N_999);
nor U2770 (N_2770,N_1236,N_1180);
nor U2771 (N_2771,N_789,N_379);
nand U2772 (N_2772,N_1341,N_1033);
nor U2773 (N_2773,N_941,N_655);
nand U2774 (N_2774,N_418,N_656);
nor U2775 (N_2775,N_438,N_315);
nand U2776 (N_2776,N_928,N_247);
nor U2777 (N_2777,N_8,N_735);
or U2778 (N_2778,N_180,N_361);
and U2779 (N_2779,N_1398,N_1343);
nand U2780 (N_2780,N_678,N_638);
nand U2781 (N_2781,N_560,N_1096);
and U2782 (N_2782,N_784,N_209);
and U2783 (N_2783,N_1119,N_1353);
and U2784 (N_2784,N_1130,N_1326);
and U2785 (N_2785,N_1189,N_226);
nand U2786 (N_2786,N_404,N_864);
and U2787 (N_2787,N_899,N_672);
nor U2788 (N_2788,N_553,N_668);
and U2789 (N_2789,N_645,N_304);
nor U2790 (N_2790,N_611,N_220);
or U2791 (N_2791,N_623,N_530);
nand U2792 (N_2792,N_338,N_1164);
nand U2793 (N_2793,N_1076,N_1465);
nor U2794 (N_2794,N_194,N_394);
nand U2795 (N_2795,N_1179,N_910);
nand U2796 (N_2796,N_722,N_884);
and U2797 (N_2797,N_370,N_892);
and U2798 (N_2798,N_1049,N_112);
nand U2799 (N_2799,N_607,N_157);
xnor U2800 (N_2800,N_573,N_103);
or U2801 (N_2801,N_1250,N_648);
nand U2802 (N_2802,N_36,N_1227);
nor U2803 (N_2803,N_1341,N_751);
nand U2804 (N_2804,N_1381,N_801);
nor U2805 (N_2805,N_1064,N_1476);
xor U2806 (N_2806,N_1195,N_1358);
nand U2807 (N_2807,N_1134,N_807);
or U2808 (N_2808,N_124,N_561);
nor U2809 (N_2809,N_23,N_658);
and U2810 (N_2810,N_527,N_1100);
nor U2811 (N_2811,N_1180,N_1049);
xnor U2812 (N_2812,N_536,N_800);
nor U2813 (N_2813,N_64,N_1397);
or U2814 (N_2814,N_24,N_1204);
nand U2815 (N_2815,N_540,N_147);
and U2816 (N_2816,N_342,N_614);
xnor U2817 (N_2817,N_1289,N_1226);
xor U2818 (N_2818,N_1428,N_791);
or U2819 (N_2819,N_1192,N_915);
or U2820 (N_2820,N_1118,N_76);
and U2821 (N_2821,N_1056,N_1072);
or U2822 (N_2822,N_532,N_1357);
and U2823 (N_2823,N_1406,N_843);
or U2824 (N_2824,N_1418,N_1242);
or U2825 (N_2825,N_711,N_1207);
xnor U2826 (N_2826,N_1300,N_770);
or U2827 (N_2827,N_1365,N_64);
nor U2828 (N_2828,N_428,N_275);
nor U2829 (N_2829,N_1009,N_796);
and U2830 (N_2830,N_102,N_552);
and U2831 (N_2831,N_1227,N_1042);
xnor U2832 (N_2832,N_326,N_461);
nor U2833 (N_2833,N_1044,N_209);
or U2834 (N_2834,N_1325,N_557);
nor U2835 (N_2835,N_454,N_1386);
nand U2836 (N_2836,N_1347,N_475);
nor U2837 (N_2837,N_511,N_1121);
xor U2838 (N_2838,N_1015,N_384);
nor U2839 (N_2839,N_775,N_671);
nand U2840 (N_2840,N_1242,N_927);
xnor U2841 (N_2841,N_1371,N_945);
nor U2842 (N_2842,N_240,N_440);
nor U2843 (N_2843,N_946,N_147);
xor U2844 (N_2844,N_627,N_524);
or U2845 (N_2845,N_11,N_1360);
nand U2846 (N_2846,N_1184,N_339);
nor U2847 (N_2847,N_795,N_158);
xor U2848 (N_2848,N_859,N_1237);
nand U2849 (N_2849,N_125,N_510);
xor U2850 (N_2850,N_844,N_1479);
xnor U2851 (N_2851,N_530,N_195);
or U2852 (N_2852,N_865,N_589);
nand U2853 (N_2853,N_848,N_309);
nor U2854 (N_2854,N_518,N_1396);
or U2855 (N_2855,N_1245,N_826);
nand U2856 (N_2856,N_736,N_54);
xnor U2857 (N_2857,N_726,N_260);
or U2858 (N_2858,N_424,N_1163);
nand U2859 (N_2859,N_636,N_503);
or U2860 (N_2860,N_272,N_1101);
and U2861 (N_2861,N_350,N_516);
or U2862 (N_2862,N_851,N_625);
nor U2863 (N_2863,N_153,N_776);
nand U2864 (N_2864,N_1431,N_1460);
nor U2865 (N_2865,N_231,N_931);
and U2866 (N_2866,N_826,N_161);
and U2867 (N_2867,N_1361,N_1110);
and U2868 (N_2868,N_333,N_320);
and U2869 (N_2869,N_1086,N_1157);
nand U2870 (N_2870,N_719,N_582);
nand U2871 (N_2871,N_1247,N_932);
or U2872 (N_2872,N_1371,N_1389);
nand U2873 (N_2873,N_523,N_812);
nand U2874 (N_2874,N_752,N_939);
nor U2875 (N_2875,N_483,N_1005);
nor U2876 (N_2876,N_19,N_229);
or U2877 (N_2877,N_198,N_293);
and U2878 (N_2878,N_1263,N_357);
nor U2879 (N_2879,N_443,N_199);
nand U2880 (N_2880,N_715,N_417);
nor U2881 (N_2881,N_556,N_587);
nand U2882 (N_2882,N_999,N_291);
and U2883 (N_2883,N_796,N_823);
and U2884 (N_2884,N_741,N_1066);
or U2885 (N_2885,N_917,N_733);
or U2886 (N_2886,N_761,N_267);
nor U2887 (N_2887,N_486,N_212);
or U2888 (N_2888,N_1131,N_924);
nand U2889 (N_2889,N_160,N_1058);
or U2890 (N_2890,N_1423,N_1232);
nor U2891 (N_2891,N_866,N_1482);
or U2892 (N_2892,N_1139,N_333);
and U2893 (N_2893,N_688,N_328);
nor U2894 (N_2894,N_1049,N_535);
nand U2895 (N_2895,N_1319,N_633);
nor U2896 (N_2896,N_1449,N_1272);
or U2897 (N_2897,N_1077,N_909);
xnor U2898 (N_2898,N_1162,N_738);
nor U2899 (N_2899,N_905,N_723);
nand U2900 (N_2900,N_711,N_860);
nand U2901 (N_2901,N_1120,N_826);
and U2902 (N_2902,N_92,N_964);
or U2903 (N_2903,N_722,N_1406);
or U2904 (N_2904,N_1229,N_1308);
nand U2905 (N_2905,N_1356,N_259);
nor U2906 (N_2906,N_1026,N_1449);
xor U2907 (N_2907,N_250,N_931);
xnor U2908 (N_2908,N_486,N_1143);
nand U2909 (N_2909,N_1078,N_681);
or U2910 (N_2910,N_1393,N_1333);
nor U2911 (N_2911,N_741,N_525);
nand U2912 (N_2912,N_437,N_1284);
nand U2913 (N_2913,N_1452,N_409);
nand U2914 (N_2914,N_679,N_704);
nor U2915 (N_2915,N_1225,N_1403);
nand U2916 (N_2916,N_705,N_1351);
or U2917 (N_2917,N_700,N_652);
nor U2918 (N_2918,N_616,N_415);
or U2919 (N_2919,N_859,N_1030);
and U2920 (N_2920,N_1275,N_842);
nor U2921 (N_2921,N_71,N_741);
nand U2922 (N_2922,N_1081,N_264);
and U2923 (N_2923,N_160,N_1360);
or U2924 (N_2924,N_840,N_1263);
or U2925 (N_2925,N_728,N_100);
nor U2926 (N_2926,N_884,N_780);
or U2927 (N_2927,N_268,N_1017);
or U2928 (N_2928,N_78,N_911);
or U2929 (N_2929,N_752,N_1051);
or U2930 (N_2930,N_1160,N_450);
or U2931 (N_2931,N_541,N_1406);
and U2932 (N_2932,N_391,N_669);
and U2933 (N_2933,N_1477,N_1118);
nand U2934 (N_2934,N_680,N_425);
nand U2935 (N_2935,N_1179,N_1168);
nand U2936 (N_2936,N_1473,N_97);
nand U2937 (N_2937,N_193,N_904);
or U2938 (N_2938,N_618,N_459);
nand U2939 (N_2939,N_790,N_36);
or U2940 (N_2940,N_1156,N_178);
xor U2941 (N_2941,N_902,N_638);
and U2942 (N_2942,N_1274,N_978);
xor U2943 (N_2943,N_635,N_865);
and U2944 (N_2944,N_196,N_301);
nand U2945 (N_2945,N_1007,N_451);
or U2946 (N_2946,N_98,N_870);
nand U2947 (N_2947,N_334,N_408);
xnor U2948 (N_2948,N_927,N_74);
xor U2949 (N_2949,N_1383,N_708);
nand U2950 (N_2950,N_463,N_1368);
and U2951 (N_2951,N_871,N_1275);
or U2952 (N_2952,N_99,N_655);
and U2953 (N_2953,N_1436,N_395);
nand U2954 (N_2954,N_224,N_638);
xor U2955 (N_2955,N_1145,N_279);
nand U2956 (N_2956,N_1167,N_937);
nand U2957 (N_2957,N_715,N_824);
nand U2958 (N_2958,N_246,N_1229);
nand U2959 (N_2959,N_1343,N_864);
nor U2960 (N_2960,N_799,N_1429);
nand U2961 (N_2961,N_18,N_1488);
nor U2962 (N_2962,N_954,N_1021);
nor U2963 (N_2963,N_487,N_1271);
and U2964 (N_2964,N_469,N_1085);
or U2965 (N_2965,N_586,N_494);
and U2966 (N_2966,N_941,N_1468);
nand U2967 (N_2967,N_765,N_820);
and U2968 (N_2968,N_142,N_548);
nor U2969 (N_2969,N_705,N_875);
or U2970 (N_2970,N_611,N_1260);
and U2971 (N_2971,N_1331,N_1296);
or U2972 (N_2972,N_375,N_83);
and U2973 (N_2973,N_343,N_828);
nor U2974 (N_2974,N_669,N_18);
or U2975 (N_2975,N_914,N_56);
and U2976 (N_2976,N_1262,N_190);
xnor U2977 (N_2977,N_1243,N_273);
nor U2978 (N_2978,N_838,N_1023);
xor U2979 (N_2979,N_920,N_352);
nand U2980 (N_2980,N_856,N_1367);
xor U2981 (N_2981,N_232,N_393);
or U2982 (N_2982,N_1373,N_766);
nand U2983 (N_2983,N_791,N_844);
nor U2984 (N_2984,N_1422,N_82);
xnor U2985 (N_2985,N_697,N_1255);
or U2986 (N_2986,N_1250,N_1298);
nand U2987 (N_2987,N_73,N_1200);
and U2988 (N_2988,N_1250,N_1129);
nor U2989 (N_2989,N_781,N_1066);
and U2990 (N_2990,N_978,N_1195);
nor U2991 (N_2991,N_708,N_1340);
nand U2992 (N_2992,N_703,N_20);
nand U2993 (N_2993,N_633,N_1380);
or U2994 (N_2994,N_34,N_331);
nor U2995 (N_2995,N_881,N_1388);
and U2996 (N_2996,N_1404,N_1050);
and U2997 (N_2997,N_300,N_1111);
nand U2998 (N_2998,N_1329,N_683);
xor U2999 (N_2999,N_833,N_1199);
or U3000 (N_3000,N_1659,N_2222);
xor U3001 (N_3001,N_2450,N_2940);
nor U3002 (N_3002,N_2769,N_1946);
nand U3003 (N_3003,N_2452,N_1976);
or U3004 (N_3004,N_2514,N_1645);
nand U3005 (N_3005,N_2584,N_2245);
and U3006 (N_3006,N_1650,N_1728);
nor U3007 (N_3007,N_2627,N_2290);
nand U3008 (N_3008,N_1817,N_1609);
or U3009 (N_3009,N_1885,N_2443);
nor U3010 (N_3010,N_2480,N_2040);
xnor U3011 (N_3011,N_2505,N_2191);
nand U3012 (N_3012,N_2740,N_2465);
and U3013 (N_3013,N_2432,N_2475);
nand U3014 (N_3014,N_2116,N_1702);
nand U3015 (N_3015,N_2960,N_2555);
and U3016 (N_3016,N_1588,N_1726);
or U3017 (N_3017,N_2814,N_2479);
or U3018 (N_3018,N_2427,N_1804);
or U3019 (N_3019,N_2533,N_2916);
nand U3020 (N_3020,N_2446,N_2905);
and U3021 (N_3021,N_1617,N_2260);
nor U3022 (N_3022,N_2036,N_1908);
nor U3023 (N_3023,N_2108,N_2072);
and U3024 (N_3024,N_1986,N_2504);
or U3025 (N_3025,N_1746,N_1805);
and U3026 (N_3026,N_2351,N_1674);
nand U3027 (N_3027,N_2105,N_2610);
and U3028 (N_3028,N_2244,N_2490);
nor U3029 (N_3029,N_1892,N_1695);
nand U3030 (N_3030,N_1930,N_2546);
or U3031 (N_3031,N_2712,N_2647);
or U3032 (N_3032,N_2941,N_1968);
and U3033 (N_3033,N_1665,N_1918);
and U3034 (N_3034,N_2425,N_2250);
or U3035 (N_3035,N_2795,N_2966);
nor U3036 (N_3036,N_2655,N_1826);
nor U3037 (N_3037,N_2150,N_2551);
nand U3038 (N_3038,N_2032,N_2021);
nand U3039 (N_3039,N_1898,N_1636);
or U3040 (N_3040,N_2558,N_1772);
or U3041 (N_3041,N_1869,N_2217);
nor U3042 (N_3042,N_2713,N_2355);
nor U3043 (N_3043,N_1720,N_2430);
and U3044 (N_3044,N_1597,N_2273);
and U3045 (N_3045,N_2897,N_2020);
or U3046 (N_3046,N_2189,N_1566);
nand U3047 (N_3047,N_2090,N_1630);
and U3048 (N_3048,N_2124,N_2414);
nand U3049 (N_3049,N_2140,N_2748);
or U3050 (N_3050,N_1923,N_2587);
or U3051 (N_3051,N_1935,N_1974);
nor U3052 (N_3052,N_2641,N_1761);
nor U3053 (N_3053,N_1777,N_1823);
and U3054 (N_3054,N_2408,N_2739);
xor U3055 (N_3055,N_2199,N_2606);
xor U3056 (N_3056,N_2709,N_2371);
and U3057 (N_3057,N_2138,N_2939);
or U3058 (N_3058,N_1560,N_1961);
xor U3059 (N_3059,N_2579,N_2074);
nand U3060 (N_3060,N_2007,N_2234);
nor U3061 (N_3061,N_2668,N_2165);
xnor U3062 (N_3062,N_2809,N_2899);
nand U3063 (N_3063,N_2833,N_1768);
and U3064 (N_3064,N_1713,N_2237);
xnor U3065 (N_3065,N_2348,N_2474);
nand U3066 (N_3066,N_1599,N_1792);
and U3067 (N_3067,N_2025,N_2640);
xor U3068 (N_3068,N_2803,N_2413);
or U3069 (N_3069,N_1737,N_2466);
and U3070 (N_3070,N_1529,N_2343);
and U3071 (N_3071,N_2179,N_2110);
xor U3072 (N_3072,N_2580,N_1672);
and U3073 (N_3073,N_2826,N_2318);
nor U3074 (N_3074,N_2213,N_1533);
nand U3075 (N_3075,N_2461,N_2958);
nor U3076 (N_3076,N_2676,N_2562);
nor U3077 (N_3077,N_1510,N_2716);
or U3078 (N_3078,N_1679,N_2780);
nor U3079 (N_3079,N_1558,N_2860);
nor U3080 (N_3080,N_2174,N_1723);
and U3081 (N_3081,N_1606,N_2874);
or U3082 (N_3082,N_2079,N_2394);
nand U3083 (N_3083,N_2919,N_2750);
nor U3084 (N_3084,N_1931,N_2730);
and U3085 (N_3085,N_2064,N_2308);
and U3086 (N_3086,N_2686,N_2291);
nand U3087 (N_3087,N_2554,N_2201);
nor U3088 (N_3088,N_1856,N_2100);
nand U3089 (N_3089,N_2903,N_2783);
or U3090 (N_3090,N_2850,N_2274);
xor U3091 (N_3091,N_2014,N_2926);
and U3092 (N_3092,N_1648,N_2724);
or U3093 (N_3093,N_2873,N_2995);
and U3094 (N_3094,N_1996,N_2653);
nor U3095 (N_3095,N_1812,N_2503);
and U3096 (N_3096,N_1763,N_2332);
xor U3097 (N_3097,N_2018,N_2705);
xnor U3098 (N_3098,N_2876,N_2513);
or U3099 (N_3099,N_2464,N_2870);
nand U3100 (N_3100,N_2359,N_2511);
nor U3101 (N_3101,N_1857,N_2993);
and U3102 (N_3102,N_1766,N_1530);
nand U3103 (N_3103,N_2335,N_1540);
xnor U3104 (N_3104,N_1620,N_2433);
nand U3105 (N_3105,N_1837,N_1552);
nand U3106 (N_3106,N_2798,N_2607);
nor U3107 (N_3107,N_2815,N_2741);
and U3108 (N_3108,N_2577,N_1653);
nor U3109 (N_3109,N_2098,N_1975);
or U3110 (N_3110,N_1685,N_1715);
nor U3111 (N_3111,N_2376,N_2284);
or U3112 (N_3112,N_2133,N_2823);
and U3113 (N_3113,N_1536,N_2434);
nand U3114 (N_3114,N_1534,N_2703);
nor U3115 (N_3115,N_2978,N_2645);
nand U3116 (N_3116,N_1652,N_1760);
or U3117 (N_3117,N_1784,N_1798);
nand U3118 (N_3118,N_1639,N_2779);
or U3119 (N_3119,N_2221,N_2139);
and U3120 (N_3120,N_2114,N_1714);
and U3121 (N_3121,N_2127,N_2917);
xor U3122 (N_3122,N_1683,N_2053);
nor U3123 (N_3123,N_2914,N_2502);
or U3124 (N_3124,N_2373,N_2981);
nor U3125 (N_3125,N_1753,N_1862);
nor U3126 (N_3126,N_2186,N_1513);
or U3127 (N_3127,N_2271,N_2339);
or U3128 (N_3128,N_2008,N_2846);
or U3129 (N_3129,N_1643,N_2661);
nor U3130 (N_3130,N_1988,N_2286);
nor U3131 (N_3131,N_2885,N_2230);
nand U3132 (N_3132,N_2301,N_2596);
nor U3133 (N_3133,N_2386,N_2294);
or U3134 (N_3134,N_1806,N_2871);
nor U3135 (N_3135,N_1596,N_2091);
or U3136 (N_3136,N_1840,N_2964);
nor U3137 (N_3137,N_1854,N_1941);
and U3138 (N_3138,N_2248,N_2422);
or U3139 (N_3139,N_2762,N_2662);
nand U3140 (N_3140,N_2675,N_2188);
and U3141 (N_3141,N_2342,N_2935);
and U3142 (N_3142,N_2509,N_2697);
and U3143 (N_3143,N_2590,N_2855);
or U3144 (N_3144,N_2992,N_2416);
nand U3145 (N_3145,N_2901,N_2298);
nor U3146 (N_3146,N_2977,N_1649);
nand U3147 (N_3147,N_2269,N_2907);
and U3148 (N_3148,N_1591,N_2945);
nor U3149 (N_3149,N_2381,N_2969);
xor U3150 (N_3150,N_2177,N_2089);
nor U3151 (N_3151,N_2297,N_2540);
nand U3152 (N_3152,N_2784,N_2224);
or U3153 (N_3153,N_1911,N_2331);
nor U3154 (N_3154,N_2552,N_2878);
and U3155 (N_3155,N_2481,N_2994);
and U3156 (N_3156,N_2656,N_1570);
and U3157 (N_3157,N_2583,N_2066);
nand U3158 (N_3158,N_2071,N_2470);
and U3159 (N_3159,N_1651,N_2324);
nor U3160 (N_3160,N_2483,N_2956);
nand U3161 (N_3161,N_2785,N_1656);
and U3162 (N_3162,N_2998,N_1776);
xor U3163 (N_3163,N_2435,N_1545);
or U3164 (N_3164,N_1791,N_2962);
nand U3165 (N_3165,N_2868,N_2345);
nand U3166 (N_3166,N_1895,N_1962);
and U3167 (N_3167,N_1842,N_2544);
xnor U3168 (N_3168,N_1644,N_2410);
nand U3169 (N_3169,N_2319,N_2063);
or U3170 (N_3170,N_1500,N_2635);
nand U3171 (N_3171,N_2356,N_2469);
and U3172 (N_3172,N_2953,N_2736);
or U3173 (N_3173,N_2042,N_2375);
and U3174 (N_3174,N_1757,N_1936);
nand U3175 (N_3175,N_2353,N_2488);
or U3176 (N_3176,N_2883,N_2163);
nor U3177 (N_3177,N_2272,N_2758);
xor U3178 (N_3178,N_2158,N_2035);
and U3179 (N_3179,N_2869,N_2918);
and U3180 (N_3180,N_2829,N_2836);
and U3181 (N_3181,N_2218,N_2424);
and U3182 (N_3182,N_1724,N_2787);
nor U3183 (N_3183,N_2537,N_2252);
nand U3184 (N_3184,N_1920,N_2895);
xnor U3185 (N_3185,N_2316,N_2153);
or U3186 (N_3186,N_2262,N_2472);
and U3187 (N_3187,N_2702,N_1511);
and U3188 (N_3188,N_2605,N_2487);
xnor U3189 (N_3189,N_1698,N_2314);
nor U3190 (N_3190,N_2069,N_1820);
nor U3191 (N_3191,N_1957,N_2927);
or U3192 (N_3192,N_2361,N_2698);
or U3193 (N_3193,N_2391,N_2699);
or U3194 (N_3194,N_2211,N_1861);
or U3195 (N_3195,N_2582,N_2445);
nor U3196 (N_3196,N_2543,N_2389);
or U3197 (N_3197,N_1525,N_2832);
and U3198 (N_3198,N_1860,N_2854);
or U3199 (N_3199,N_2838,N_2852);
or U3200 (N_3200,N_2094,N_1825);
or U3201 (N_3201,N_2766,N_2081);
and U3202 (N_3202,N_2911,N_2866);
xnor U3203 (N_3203,N_2499,N_2872);
or U3204 (N_3204,N_2170,N_2970);
xor U3205 (N_3205,N_2048,N_2725);
xor U3206 (N_3206,N_2454,N_1578);
xnor U3207 (N_3207,N_2528,N_1999);
nand U3208 (N_3208,N_2808,N_1811);
and U3209 (N_3209,N_2210,N_2786);
nand U3210 (N_3210,N_2144,N_1501);
and U3211 (N_3211,N_2397,N_1618);
nand U3212 (N_3212,N_2834,N_2660);
and U3213 (N_3213,N_1562,N_2957);
nor U3214 (N_3214,N_1905,N_2457);
nand U3215 (N_3215,N_2323,N_2651);
or U3216 (N_3216,N_2915,N_2396);
or U3217 (N_3217,N_1994,N_2460);
nand U3218 (N_3218,N_1622,N_1956);
xnor U3219 (N_3219,N_1690,N_2898);
or U3220 (N_3220,N_2566,N_1959);
nand U3221 (N_3221,N_2034,N_1575);
or U3222 (N_3222,N_2887,N_1632);
and U3223 (N_3223,N_2849,N_2175);
xor U3224 (N_3224,N_2400,N_2403);
or U3225 (N_3225,N_1933,N_2688);
and U3226 (N_3226,N_2928,N_1789);
and U3227 (N_3227,N_1607,N_1822);
xor U3228 (N_3228,N_2881,N_2774);
or U3229 (N_3229,N_2125,N_2231);
nand U3230 (N_3230,N_2239,N_1693);
or U3231 (N_3231,N_1866,N_2685);
nor U3232 (N_3232,N_2506,N_1754);
or U3233 (N_3233,N_2428,N_1631);
nor U3234 (N_3234,N_1565,N_2087);
and U3235 (N_3235,N_2238,N_2423);
nand U3236 (N_3236,N_2609,N_2659);
or U3237 (N_3237,N_2393,N_2534);
xor U3238 (N_3238,N_2190,N_1716);
and U3239 (N_3239,N_2631,N_1680);
and U3240 (N_3240,N_1557,N_1952);
nand U3241 (N_3241,N_2520,N_1603);
and U3242 (N_3242,N_2029,N_1686);
nor U3243 (N_3243,N_2519,N_2667);
nor U3244 (N_3244,N_2299,N_1912);
nor U3245 (N_3245,N_2406,N_1802);
nand U3246 (N_3246,N_1872,N_2155);
nor U3247 (N_3247,N_2848,N_2997);
and U3248 (N_3248,N_2051,N_2693);
and U3249 (N_3249,N_2492,N_2819);
nand U3250 (N_3250,N_2184,N_1808);
and U3251 (N_3251,N_2575,N_1998);
or U3252 (N_3252,N_2016,N_1663);
or U3253 (N_3253,N_2135,N_2721);
or U3254 (N_3254,N_1752,N_1855);
or U3255 (N_3255,N_1971,N_1559);
nand U3256 (N_3256,N_2954,N_2121);
nand U3257 (N_3257,N_2756,N_2031);
or U3258 (N_3258,N_1980,N_2259);
nor U3259 (N_3259,N_1844,N_2447);
nor U3260 (N_3260,N_1835,N_1934);
or U3261 (N_3261,N_2056,N_2630);
or U3262 (N_3262,N_1735,N_1717);
and U3263 (N_3263,N_1706,N_2824);
nand U3264 (N_3264,N_1646,N_1572);
xnor U3265 (N_3265,N_2530,N_2073);
and U3266 (N_3266,N_2799,N_2482);
xnor U3267 (N_3267,N_2390,N_2597);
and U3268 (N_3268,N_2906,N_2120);
nor U3269 (N_3269,N_1942,N_2126);
or U3270 (N_3270,N_2563,N_2934);
or U3271 (N_3271,N_2524,N_2628);
nor U3272 (N_3272,N_2172,N_2002);
nand U3273 (N_3273,N_1972,N_1523);
nor U3274 (N_3274,N_2160,N_2344);
or U3275 (N_3275,N_1850,N_2060);
or U3276 (N_3276,N_1608,N_1992);
nor U3277 (N_3277,N_1919,N_1582);
nor U3278 (N_3278,N_2159,N_1673);
nand U3279 (N_3279,N_2304,N_1551);
nor U3280 (N_3280,N_1689,N_2652);
and U3281 (N_3281,N_2000,N_2322);
nor U3282 (N_3282,N_2929,N_1793);
nand U3283 (N_3283,N_1878,N_2367);
nor U3284 (N_3284,N_2275,N_2733);
and U3285 (N_3285,N_2019,N_2617);
nor U3286 (N_3286,N_2984,N_2975);
nand U3287 (N_3287,N_2026,N_2560);
or U3288 (N_3288,N_2419,N_2571);
xnor U3289 (N_3289,N_2349,N_2421);
nand U3290 (N_3290,N_2804,N_2167);
and U3291 (N_3291,N_2117,N_2603);
and U3292 (N_3292,N_2489,N_2104);
nor U3293 (N_3293,N_2485,N_2095);
xor U3294 (N_3294,N_1699,N_2681);
or U3295 (N_3295,N_1676,N_2214);
or U3296 (N_3296,N_2658,N_2203);
and U3297 (N_3297,N_2791,N_2076);
or U3298 (N_3298,N_2715,N_2111);
nor U3299 (N_3299,N_1625,N_2145);
nor U3300 (N_3300,N_1696,N_2796);
xnor U3301 (N_3301,N_1989,N_2169);
xnor U3302 (N_3302,N_2204,N_1859);
or U3303 (N_3303,N_1973,N_2388);
xnor U3304 (N_3304,N_2292,N_2276);
and U3305 (N_3305,N_1991,N_1849);
xor U3306 (N_3306,N_2841,N_2147);
and U3307 (N_3307,N_2208,N_1585);
nor U3308 (N_3308,N_2426,N_2828);
and U3309 (N_3309,N_2384,N_1927);
or U3310 (N_3310,N_1883,N_2009);
nand U3311 (N_3311,N_1832,N_1544);
or U3312 (N_3312,N_2746,N_2650);
nor U3313 (N_3313,N_1747,N_2192);
nand U3314 (N_3314,N_2719,N_1939);
or U3315 (N_3315,N_2417,N_2600);
nand U3316 (N_3316,N_2578,N_1697);
nand U3317 (N_3317,N_1796,N_2205);
and U3318 (N_3318,N_2336,N_1561);
or U3319 (N_3319,N_2822,N_2307);
xor U3320 (N_3320,N_1997,N_2831);
or U3321 (N_3321,N_1677,N_2912);
or U3322 (N_3322,N_2023,N_2581);
nand U3323 (N_3323,N_2409,N_2890);
and U3324 (N_3324,N_2951,N_2781);
or U3325 (N_3325,N_1834,N_2991);
nand U3326 (N_3326,N_2080,N_1725);
nand U3327 (N_3327,N_1894,N_2500);
nor U3328 (N_3328,N_2182,N_2083);
and U3329 (N_3329,N_1924,N_2039);
nand U3330 (N_3330,N_2639,N_1521);
nor U3331 (N_3331,N_2696,N_1810);
nand U3332 (N_3332,N_2593,N_1694);
nand U3333 (N_3333,N_1718,N_2102);
nand U3334 (N_3334,N_1587,N_2654);
nor U3335 (N_3335,N_1600,N_2484);
and U3336 (N_3336,N_2541,N_2949);
xnor U3337 (N_3337,N_2556,N_2103);
nand U3338 (N_3338,N_2879,N_1594);
or U3339 (N_3339,N_2197,N_1541);
nand U3340 (N_3340,N_1517,N_2441);
or U3341 (N_3341,N_2088,N_2368);
or U3342 (N_3342,N_2132,N_2200);
nand U3343 (N_3343,N_1688,N_2157);
xnor U3344 (N_3344,N_2086,N_1626);
nor U3345 (N_3345,N_1705,N_2264);
nand U3346 (N_3346,N_2099,N_2550);
nand U3347 (N_3347,N_2363,N_1762);
nand U3348 (N_3348,N_2295,N_2987);
and U3349 (N_3349,N_1567,N_1783);
nor U3350 (N_3350,N_2052,N_2045);
or U3351 (N_3351,N_2706,N_2429);
nor U3352 (N_3352,N_1647,N_2670);
or U3353 (N_3353,N_2494,N_2106);
or U3354 (N_3354,N_1543,N_2471);
xnor U3355 (N_3355,N_2548,N_2119);
or U3356 (N_3356,N_2775,N_2710);
nor U3357 (N_3357,N_2315,N_1756);
or U3358 (N_3358,N_2613,N_1708);
nand U3359 (N_3359,N_2797,N_2764);
nor U3360 (N_3360,N_1584,N_1681);
nor U3361 (N_3361,N_2880,N_1893);
and U3362 (N_3362,N_2875,N_1765);
nand U3363 (N_3363,N_2532,N_2027);
and U3364 (N_3364,N_2924,N_2357);
or U3365 (N_3365,N_2115,N_2877);
nand U3366 (N_3366,N_2082,N_2517);
or U3367 (N_3367,N_2436,N_2801);
nor U3368 (N_3368,N_1848,N_1940);
and U3369 (N_3369,N_2084,N_1890);
nor U3370 (N_3370,N_2112,N_2411);
nor U3371 (N_3371,N_2404,N_1831);
and U3372 (N_3372,N_2235,N_2041);
nand U3373 (N_3373,N_1569,N_1786);
nand U3374 (N_3374,N_2963,N_2621);
or U3375 (N_3375,N_2744,N_2440);
and U3376 (N_3376,N_1583,N_2162);
nand U3377 (N_3377,N_2379,N_1748);
xnor U3378 (N_3378,N_2642,N_2694);
and U3379 (N_3379,N_2501,N_2727);
or U3380 (N_3380,N_2761,N_2392);
or U3381 (N_3381,N_2930,N_2837);
nand U3382 (N_3382,N_2364,N_1669);
nor U3383 (N_3383,N_2033,N_2989);
or U3384 (N_3384,N_2535,N_2477);
nand U3385 (N_3385,N_1751,N_2777);
nor U3386 (N_3386,N_2198,N_2718);
nor U3387 (N_3387,N_2910,N_2844);
xor U3388 (N_3388,N_1982,N_2401);
or U3389 (N_3389,N_2195,N_1514);
nand U3390 (N_3390,N_2176,N_1614);
nand U3391 (N_3391,N_1891,N_2478);
or U3392 (N_3392,N_2825,N_1897);
nor U3393 (N_3393,N_2438,N_2734);
or U3394 (N_3394,N_1902,N_2003);
nand U3395 (N_3395,N_2937,N_1785);
nor U3396 (N_3396,N_1979,N_2399);
nand U3397 (N_3397,N_2944,N_1925);
nand U3398 (N_3398,N_2202,N_2679);
nand U3399 (N_3399,N_2690,N_2212);
nand U3400 (N_3400,N_1661,N_2772);
or U3401 (N_3401,N_2526,N_1819);
nand U3402 (N_3402,N_1836,N_2648);
or U3403 (N_3403,N_2366,N_1660);
nor U3404 (N_3404,N_2270,N_1788);
nand U3405 (N_3405,N_2782,N_1733);
or U3406 (N_3406,N_2143,N_2148);
xor U3407 (N_3407,N_1910,N_2258);
nor U3408 (N_3408,N_1602,N_1616);
nor U3409 (N_3409,N_2946,N_2700);
xnor U3410 (N_3410,N_1749,N_1764);
or U3411 (N_3411,N_1877,N_2277);
nor U3412 (N_3412,N_1712,N_1538);
and U3413 (N_3413,N_2268,N_2037);
nor U3414 (N_3414,N_1884,N_1507);
nor U3415 (N_3415,N_1880,N_1556);
nand U3416 (N_3416,N_2522,N_1990);
nand U3417 (N_3417,N_2305,N_2840);
xor U3418 (N_3418,N_2792,N_2811);
and U3419 (N_3419,N_1830,N_2168);
and U3420 (N_3420,N_1739,N_2129);
xor U3421 (N_3421,N_2687,N_2805);
nand U3422 (N_3422,N_2136,N_1938);
or U3423 (N_3423,N_1829,N_1943);
or U3424 (N_3424,N_1729,N_2227);
nor U3425 (N_3425,N_2771,N_2624);
and U3426 (N_3426,N_2225,N_1955);
and U3427 (N_3427,N_1553,N_2330);
or U3428 (N_3428,N_2952,N_2933);
or U3429 (N_3429,N_1548,N_2623);
or U3430 (N_3430,N_2902,N_2757);
nand U3431 (N_3431,N_2862,N_2346);
nor U3432 (N_3432,N_1816,N_1667);
and U3433 (N_3433,N_2932,N_1947);
nor U3434 (N_3434,N_1611,N_2982);
nand U3435 (N_3435,N_2085,N_2938);
xnor U3436 (N_3436,N_1546,N_2638);
nor U3437 (N_3437,N_2022,N_2439);
or U3438 (N_3438,N_2614,N_1782);
or U3439 (N_3439,N_2886,N_1858);
or U3440 (N_3440,N_2959,N_2853);
or U3441 (N_3441,N_2059,N_1707);
nand U3442 (N_3442,N_1506,N_1985);
or U3443 (N_3443,N_2161,N_2742);
or U3444 (N_3444,N_2857,N_2038);
nand U3445 (N_3445,N_1503,N_2674);
nor U3446 (N_3446,N_2180,N_2588);
nor U3447 (N_3447,N_2515,N_2673);
nand U3448 (N_3448,N_1531,N_2402);
nor U3449 (N_3449,N_2508,N_1547);
xor U3450 (N_3450,N_1948,N_1532);
and U3451 (N_3451,N_2921,N_2545);
or U3452 (N_3452,N_2374,N_1619);
and U3453 (N_3453,N_1900,N_2251);
nand U3454 (N_3454,N_2620,N_2468);
nor U3455 (N_3455,N_1818,N_2711);
nand U3456 (N_3456,N_2768,N_2178);
and U3457 (N_3457,N_2256,N_1519);
or U3458 (N_3458,N_2507,N_2398);
nand U3459 (N_3459,N_2961,N_2325);
or U3460 (N_3460,N_2559,N_1592);
nor U3461 (N_3461,N_2612,N_2456);
and U3462 (N_3462,N_2415,N_1827);
and U3463 (N_3463,N_1509,N_2329);
or U3464 (N_3464,N_1564,N_2570);
or U3465 (N_3465,N_1767,N_1970);
or U3466 (N_3466,N_1522,N_2810);
xnor U3467 (N_3467,N_2619,N_2050);
nand U3468 (N_3468,N_1727,N_2156);
and U3469 (N_3469,N_2473,N_2372);
and U3470 (N_3470,N_2726,N_2173);
nor U3471 (N_3471,N_2776,N_2249);
and U3472 (N_3472,N_1601,N_2451);
nand U3473 (N_3473,N_2677,N_2280);
nor U3474 (N_3474,N_2884,N_1678);
and U3475 (N_3475,N_1527,N_2096);
and U3476 (N_3476,N_2043,N_1516);
nand U3477 (N_3477,N_2701,N_2128);
nand U3478 (N_3478,N_2317,N_1515);
or U3479 (N_3479,N_2134,N_2861);
nor U3480 (N_3480,N_1951,N_1932);
and U3481 (N_3481,N_1847,N_1550);
nand U3482 (N_3482,N_2955,N_1958);
and U3483 (N_3483,N_1605,N_1571);
and U3484 (N_3484,N_2255,N_2044);
and U3485 (N_3485,N_1658,N_1542);
nand U3486 (N_3486,N_1668,N_2947);
nor U3487 (N_3487,N_2818,N_1978);
nand U3488 (N_3488,N_1535,N_1873);
nand U3489 (N_3489,N_2611,N_2263);
nand U3490 (N_3490,N_2215,N_2093);
nor U3491 (N_3491,N_1711,N_2663);
xor U3492 (N_3492,N_1719,N_1833);
nor U3493 (N_3493,N_2707,N_1769);
and U3494 (N_3494,N_2405,N_1773);
nor U3495 (N_3495,N_1654,N_1917);
or U3496 (N_3496,N_2017,N_2141);
nor U3497 (N_3497,N_1744,N_2738);
nand U3498 (N_3498,N_2665,N_2523);
xnor U3499 (N_3499,N_2171,N_1750);
and U3500 (N_3500,N_1967,N_1520);
nand U3501 (N_3501,N_1615,N_2491);
nor U3502 (N_3502,N_2206,N_1730);
nor U3503 (N_3503,N_1964,N_2793);
nor U3504 (N_3504,N_2109,N_2616);
or U3505 (N_3505,N_2193,N_2751);
nor U3506 (N_3506,N_2518,N_2737);
xnor U3507 (N_3507,N_1969,N_2196);
and U3508 (N_3508,N_2598,N_2802);
nand U3509 (N_3509,N_1528,N_2067);
xnor U3510 (N_3510,N_2999,N_2830);
and U3511 (N_3511,N_1809,N_2678);
nor U3512 (N_3512,N_2242,N_2525);
and U3513 (N_3513,N_2643,N_2625);
nand U3514 (N_3514,N_1721,N_2976);
nand U3515 (N_3515,N_1944,N_1886);
nand U3516 (N_3516,N_2257,N_2858);
or U3517 (N_3517,N_1841,N_1613);
nand U3518 (N_3518,N_1666,N_1921);
nor U3519 (N_3519,N_1635,N_1790);
and U3520 (N_3520,N_1505,N_2789);
and U3521 (N_3521,N_2723,N_2006);
nor U3522 (N_3522,N_2637,N_2773);
and U3523 (N_3523,N_2800,N_2985);
and U3524 (N_3524,N_1839,N_1828);
nor U3525 (N_3525,N_2908,N_2010);
nand U3526 (N_3526,N_1853,N_2664);
nor U3527 (N_3527,N_2790,N_2755);
nor U3528 (N_3528,N_2101,N_2236);
xnor U3529 (N_3529,N_2370,N_2567);
nand U3530 (N_3530,N_1655,N_1682);
or U3531 (N_3531,N_2778,N_1815);
nor U3532 (N_3532,N_2122,N_2293);
xor U3533 (N_3533,N_2130,N_1795);
or U3534 (N_3534,N_2974,N_2636);
nor U3535 (N_3535,N_2943,N_1512);
or U3536 (N_3536,N_1758,N_2431);
xor U3537 (N_3537,N_1709,N_2925);
or U3538 (N_3538,N_2568,N_1875);
or U3539 (N_3539,N_2936,N_2005);
or U3540 (N_3540,N_2306,N_1549);
or U3541 (N_3541,N_1906,N_2986);
or U3542 (N_3542,N_2765,N_2971);
and U3543 (N_3543,N_2564,N_2531);
or U3544 (N_3544,N_2747,N_2241);
nand U3545 (N_3545,N_2683,N_2547);
nor U3546 (N_3546,N_2448,N_2219);
nor U3547 (N_3547,N_2498,N_2714);
nand U3548 (N_3548,N_1759,N_2574);
nor U3549 (N_3549,N_2692,N_1662);
nand U3550 (N_3550,N_2618,N_1638);
or U3551 (N_3551,N_2657,N_1604);
nand U3552 (N_3552,N_1977,N_2666);
and U3553 (N_3553,N_2536,N_1914);
and U3554 (N_3554,N_2722,N_2882);
nand U3555 (N_3555,N_2891,N_2302);
nand U3556 (N_3556,N_2486,N_2061);
or U3557 (N_3557,N_2615,N_2839);
nand U3558 (N_3558,N_1870,N_2216);
xnor U3559 (N_3559,N_2247,N_2309);
nand U3560 (N_3560,N_2763,N_1907);
nand U3561 (N_3561,N_2770,N_2350);
and U3562 (N_3562,N_1899,N_1701);
nor U3563 (N_3563,N_2806,N_2437);
xnor U3564 (N_3564,N_2632,N_2463);
nand U3565 (N_3565,N_2360,N_1966);
nor U3566 (N_3566,N_1634,N_2996);
nor U3567 (N_3567,N_2240,N_2728);
nor U3568 (N_3568,N_1641,N_1742);
nor U3569 (N_3569,N_2923,N_2154);
and U3570 (N_3570,N_2704,N_2253);
and U3571 (N_3571,N_2922,N_1963);
nor U3572 (N_3572,N_2538,N_2669);
and U3573 (N_3573,N_2055,N_1580);
and U3574 (N_3574,N_2592,N_2842);
or U3575 (N_3575,N_1589,N_1945);
nor U3576 (N_3576,N_1755,N_2118);
nand U3577 (N_3577,N_2561,N_1612);
nand U3578 (N_3578,N_2752,N_1774);
nor U3579 (N_3579,N_1771,N_2695);
nor U3580 (N_3580,N_1627,N_2759);
and U3581 (N_3581,N_1779,N_2904);
nor U3582 (N_3582,N_2387,N_2226);
nor U3583 (N_3583,N_1590,N_1518);
or U3584 (N_3584,N_2743,N_2028);
or U3585 (N_3585,N_1732,N_2243);
nor U3586 (N_3586,N_2285,N_1965);
and U3587 (N_3587,N_1738,N_2187);
or U3588 (N_3588,N_2950,N_2282);
and U3589 (N_3589,N_1867,N_2672);
nand U3590 (N_3590,N_1539,N_1887);
or U3591 (N_3591,N_1843,N_2289);
nand U3592 (N_3592,N_2968,N_1915);
and U3593 (N_3593,N_1703,N_1995);
nand U3594 (N_3594,N_2151,N_1568);
or U3595 (N_3595,N_2888,N_2228);
nand U3596 (N_3596,N_1577,N_2321);
and U3597 (N_3597,N_1863,N_2113);
or U3598 (N_3598,N_2731,N_1675);
xnor U3599 (N_3599,N_1671,N_1981);
nand U3600 (N_3600,N_2418,N_1610);
nor U3601 (N_3601,N_1807,N_2229);
or U3602 (N_3602,N_1504,N_1799);
or U3603 (N_3603,N_2572,N_2646);
or U3604 (N_3604,N_2209,N_1797);
or U3605 (N_3605,N_2341,N_2980);
or U3606 (N_3606,N_1537,N_2246);
and U3607 (N_3607,N_1864,N_1993);
and U3608 (N_3608,N_2807,N_2812);
or U3609 (N_3609,N_2283,N_1740);
xnor U3610 (N_3610,N_1573,N_2223);
nor U3611 (N_3611,N_2062,N_2011);
or U3612 (N_3612,N_1741,N_1868);
nand U3613 (N_3613,N_2680,N_1984);
xnor U3614 (N_3614,N_1846,N_1657);
or U3615 (N_3615,N_2453,N_2626);
nor U3616 (N_3616,N_1640,N_1949);
and U3617 (N_3617,N_1736,N_2909);
xor U3618 (N_3618,N_2320,N_1954);
or U3619 (N_3619,N_2462,N_2166);
xnor U3620 (N_3620,N_1814,N_2281);
xnor U3621 (N_3621,N_2267,N_2311);
or U3622 (N_3622,N_1621,N_1770);
nand U3623 (N_3623,N_1624,N_1926);
nor U3624 (N_3624,N_1526,N_2867);
nand U3625 (N_3625,N_1983,N_2012);
xor U3626 (N_3626,N_2745,N_1874);
xnor U3627 (N_3627,N_2058,N_2476);
and U3628 (N_3628,N_1845,N_2900);
and U3629 (N_3629,N_2527,N_1824);
xnor U3630 (N_3630,N_1803,N_2068);
nand U3631 (N_3631,N_1642,N_2983);
nor U3632 (N_3632,N_2057,N_2573);
or U3633 (N_3633,N_2516,N_2369);
nor U3634 (N_3634,N_1865,N_2691);
nor U3635 (N_3635,N_1901,N_2092);
xor U3636 (N_3636,N_2864,N_2965);
nor U3637 (N_3637,N_2729,N_2382);
nand U3638 (N_3638,N_2137,N_2449);
or U3639 (N_3639,N_1781,N_2496);
nor U3640 (N_3640,N_2589,N_2279);
nor U3641 (N_3641,N_1916,N_1896);
xor U3642 (N_3642,N_2380,N_2146);
nor U3643 (N_3643,N_1598,N_1731);
and U3644 (N_3644,N_1554,N_2407);
nor U3645 (N_3645,N_2820,N_2720);
nor U3646 (N_3646,N_2682,N_2123);
nand U3647 (N_3647,N_2467,N_2990);
and U3648 (N_3648,N_2300,N_2920);
or U3649 (N_3649,N_2542,N_2337);
xor U3650 (N_3650,N_2767,N_2732);
nand U3651 (N_3651,N_2539,N_2893);
nand U3652 (N_3652,N_2254,N_2065);
xnor U3653 (N_3653,N_1687,N_2181);
and U3654 (N_3654,N_2334,N_1881);
and U3655 (N_3655,N_2591,N_2859);
nand U3656 (N_3656,N_1871,N_1745);
or U3657 (N_3657,N_1574,N_1888);
xnor U3658 (N_3658,N_2358,N_2835);
and U3659 (N_3659,N_1922,N_1628);
nand U3660 (N_3660,N_1778,N_1909);
xnor U3661 (N_3661,N_2972,N_2328);
and U3662 (N_3662,N_1794,N_1852);
nand U3663 (N_3663,N_2967,N_1960);
and U3664 (N_3664,N_2054,N_1879);
nor U3665 (N_3665,N_2553,N_1904);
or U3666 (N_3666,N_2931,N_1928);
xnor U3667 (N_3667,N_2164,N_2015);
and U3668 (N_3668,N_2220,N_1889);
nand U3669 (N_3669,N_2333,N_2816);
and U3670 (N_3670,N_2827,N_2077);
nand U3671 (N_3671,N_1692,N_2586);
nand U3672 (N_3672,N_1524,N_2097);
nand U3673 (N_3673,N_2510,N_2495);
or U3674 (N_3674,N_1700,N_2313);
and U3675 (N_3675,N_2601,N_2892);
nor U3676 (N_3676,N_1710,N_1882);
or U3677 (N_3677,N_2420,N_1743);
or U3678 (N_3678,N_1821,N_2004);
nand U3679 (N_3679,N_2338,N_2629);
nand U3680 (N_3680,N_2856,N_2569);
nor U3681 (N_3681,N_2794,N_2760);
nand U3682 (N_3682,N_1502,N_2385);
nand U3683 (N_3683,N_2754,N_2753);
or U3684 (N_3684,N_2988,N_2265);
and U3685 (N_3685,N_2865,N_2684);
nor U3686 (N_3686,N_2847,N_2497);
nand U3687 (N_3687,N_2383,N_1950);
and U3688 (N_3688,N_2851,N_2232);
and U3689 (N_3689,N_1903,N_2046);
or U3690 (N_3690,N_2412,N_2529);
nor U3691 (N_3691,N_2565,N_2717);
xor U3692 (N_3692,N_2207,N_2512);
or U3693 (N_3693,N_2455,N_2788);
nor U3694 (N_3694,N_2493,N_2149);
nand U3695 (N_3695,N_2142,N_2889);
and U3696 (N_3696,N_2896,N_1987);
nand U3697 (N_3697,N_2622,N_2813);
or U3698 (N_3698,N_2644,N_2576);
nand U3699 (N_3699,N_2131,N_2078);
or U3700 (N_3700,N_2649,N_2030);
and U3701 (N_3701,N_2347,N_1684);
nor U3702 (N_3702,N_2585,N_2288);
nand U3703 (N_3703,N_1623,N_2310);
or U3704 (N_3704,N_2049,N_2261);
nor U3705 (N_3705,N_2863,N_2973);
nor U3706 (N_3706,N_2001,N_2152);
nand U3707 (N_3707,N_2107,N_2671);
nor U3708 (N_3708,N_1937,N_2521);
nor U3709 (N_3709,N_2185,N_2444);
nand U3710 (N_3710,N_1913,N_1563);
nand U3711 (N_3711,N_1664,N_1800);
and U3712 (N_3712,N_1929,N_2979);
or U3713 (N_3713,N_2594,N_2312);
or U3714 (N_3714,N_2362,N_1508);
nand U3715 (N_3715,N_2604,N_1595);
nor U3716 (N_3716,N_2395,N_1734);
xor U3717 (N_3717,N_2377,N_1581);
nand U3718 (N_3718,N_1670,N_2194);
or U3719 (N_3719,N_2843,N_2599);
or U3720 (N_3720,N_2296,N_1576);
nand U3721 (N_3721,N_2365,N_2689);
nor U3722 (N_3722,N_1953,N_2602);
nor U3723 (N_3723,N_2352,N_2354);
nand U3724 (N_3724,N_2303,N_2845);
and U3725 (N_3725,N_1704,N_1555);
nand U3726 (N_3726,N_2749,N_1801);
nand U3727 (N_3727,N_1629,N_2024);
or U3728 (N_3728,N_2634,N_2287);
nand U3729 (N_3729,N_2075,N_2183);
nand U3730 (N_3730,N_2047,N_2327);
nor U3731 (N_3731,N_2549,N_2894);
nand U3732 (N_3732,N_1579,N_2442);
and U3733 (N_3733,N_2070,N_1722);
or U3734 (N_3734,N_2326,N_2013);
or U3735 (N_3735,N_1780,N_1586);
or U3736 (N_3736,N_2913,N_2948);
nand U3737 (N_3737,N_2942,N_2821);
and U3738 (N_3738,N_2278,N_2458);
or U3739 (N_3739,N_2708,N_2459);
and U3740 (N_3740,N_1876,N_2233);
or U3741 (N_3741,N_1787,N_1813);
xor U3742 (N_3742,N_2378,N_1838);
or U3743 (N_3743,N_2633,N_1593);
nand U3744 (N_3744,N_2557,N_1851);
and U3745 (N_3745,N_1691,N_2595);
or U3746 (N_3746,N_2340,N_2608);
xor U3747 (N_3747,N_1775,N_2817);
and U3748 (N_3748,N_2735,N_2266);
nor U3749 (N_3749,N_1633,N_1637);
nor U3750 (N_3750,N_2036,N_1811);
nand U3751 (N_3751,N_2185,N_2964);
nor U3752 (N_3752,N_1709,N_2453);
nor U3753 (N_3753,N_2171,N_2833);
nand U3754 (N_3754,N_1614,N_2864);
or U3755 (N_3755,N_1963,N_2182);
nand U3756 (N_3756,N_2194,N_2364);
or U3757 (N_3757,N_2894,N_1774);
or U3758 (N_3758,N_2640,N_1673);
nand U3759 (N_3759,N_1811,N_1919);
nand U3760 (N_3760,N_2138,N_1588);
and U3761 (N_3761,N_1762,N_2809);
nor U3762 (N_3762,N_2796,N_2409);
and U3763 (N_3763,N_1623,N_2664);
nand U3764 (N_3764,N_2002,N_2226);
or U3765 (N_3765,N_1601,N_2293);
nor U3766 (N_3766,N_2232,N_1985);
nand U3767 (N_3767,N_2630,N_2113);
nor U3768 (N_3768,N_2640,N_2205);
xor U3769 (N_3769,N_2588,N_1745);
nand U3770 (N_3770,N_1882,N_2247);
xnor U3771 (N_3771,N_1979,N_2575);
and U3772 (N_3772,N_1892,N_2814);
nand U3773 (N_3773,N_2329,N_2153);
nor U3774 (N_3774,N_2763,N_1895);
nand U3775 (N_3775,N_1608,N_2595);
xnor U3776 (N_3776,N_1616,N_2049);
xnor U3777 (N_3777,N_2932,N_1957);
nand U3778 (N_3778,N_2543,N_2404);
nor U3779 (N_3779,N_2916,N_2915);
nor U3780 (N_3780,N_1989,N_2927);
nor U3781 (N_3781,N_2090,N_1597);
or U3782 (N_3782,N_2534,N_1922);
nor U3783 (N_3783,N_2312,N_2398);
nand U3784 (N_3784,N_2883,N_2651);
nor U3785 (N_3785,N_1666,N_2471);
or U3786 (N_3786,N_1765,N_1651);
xor U3787 (N_3787,N_2193,N_2619);
or U3788 (N_3788,N_2329,N_2643);
nor U3789 (N_3789,N_2579,N_2998);
and U3790 (N_3790,N_2899,N_2035);
or U3791 (N_3791,N_2358,N_2677);
or U3792 (N_3792,N_2687,N_1956);
nand U3793 (N_3793,N_1687,N_2781);
nand U3794 (N_3794,N_1848,N_1810);
and U3795 (N_3795,N_2320,N_2786);
nor U3796 (N_3796,N_2923,N_2574);
nand U3797 (N_3797,N_2261,N_1693);
nor U3798 (N_3798,N_2566,N_2738);
or U3799 (N_3799,N_2731,N_1835);
or U3800 (N_3800,N_2109,N_2977);
nor U3801 (N_3801,N_2970,N_1933);
nand U3802 (N_3802,N_2154,N_2441);
or U3803 (N_3803,N_2301,N_1773);
nand U3804 (N_3804,N_1752,N_2003);
nand U3805 (N_3805,N_2215,N_1813);
or U3806 (N_3806,N_2122,N_1515);
nor U3807 (N_3807,N_2813,N_2047);
or U3808 (N_3808,N_2467,N_2248);
nor U3809 (N_3809,N_2939,N_1627);
or U3810 (N_3810,N_2229,N_1855);
nor U3811 (N_3811,N_2054,N_1749);
or U3812 (N_3812,N_2102,N_2737);
nand U3813 (N_3813,N_2772,N_2813);
and U3814 (N_3814,N_1790,N_2791);
nor U3815 (N_3815,N_2657,N_1766);
xnor U3816 (N_3816,N_2929,N_2780);
nand U3817 (N_3817,N_2352,N_2178);
nor U3818 (N_3818,N_2484,N_2092);
nor U3819 (N_3819,N_2195,N_2275);
and U3820 (N_3820,N_1876,N_2630);
nor U3821 (N_3821,N_2092,N_2375);
and U3822 (N_3822,N_2478,N_2802);
nand U3823 (N_3823,N_1511,N_2062);
and U3824 (N_3824,N_1811,N_2193);
and U3825 (N_3825,N_1520,N_2467);
nor U3826 (N_3826,N_1631,N_2132);
and U3827 (N_3827,N_1914,N_2939);
and U3828 (N_3828,N_2414,N_2547);
xnor U3829 (N_3829,N_2522,N_2193);
or U3830 (N_3830,N_2089,N_1659);
xor U3831 (N_3831,N_2536,N_2932);
nand U3832 (N_3832,N_1639,N_2415);
nor U3833 (N_3833,N_2612,N_2775);
and U3834 (N_3834,N_1943,N_2775);
xnor U3835 (N_3835,N_2610,N_2904);
nand U3836 (N_3836,N_2813,N_2348);
nor U3837 (N_3837,N_1888,N_2882);
nor U3838 (N_3838,N_1815,N_2979);
xor U3839 (N_3839,N_2708,N_1834);
nor U3840 (N_3840,N_1977,N_1566);
and U3841 (N_3841,N_2105,N_2269);
xor U3842 (N_3842,N_1835,N_2482);
or U3843 (N_3843,N_2819,N_2417);
and U3844 (N_3844,N_2258,N_1960);
or U3845 (N_3845,N_2635,N_2639);
nand U3846 (N_3846,N_2503,N_2771);
or U3847 (N_3847,N_2451,N_1834);
or U3848 (N_3848,N_2076,N_1647);
xor U3849 (N_3849,N_1889,N_2463);
and U3850 (N_3850,N_2888,N_2916);
xor U3851 (N_3851,N_2283,N_2020);
nor U3852 (N_3852,N_2742,N_1809);
nand U3853 (N_3853,N_1976,N_2140);
nor U3854 (N_3854,N_1606,N_2029);
nand U3855 (N_3855,N_1864,N_1576);
or U3856 (N_3856,N_2264,N_2981);
nor U3857 (N_3857,N_1867,N_2199);
nand U3858 (N_3858,N_1907,N_1853);
nor U3859 (N_3859,N_1796,N_1945);
nor U3860 (N_3860,N_1783,N_1582);
xnor U3861 (N_3861,N_1544,N_1552);
or U3862 (N_3862,N_2466,N_1730);
and U3863 (N_3863,N_1648,N_1731);
and U3864 (N_3864,N_2981,N_2171);
xnor U3865 (N_3865,N_1653,N_2772);
nand U3866 (N_3866,N_2774,N_1659);
nor U3867 (N_3867,N_1896,N_2427);
nor U3868 (N_3868,N_2163,N_2037);
nor U3869 (N_3869,N_2945,N_2472);
or U3870 (N_3870,N_2619,N_2631);
and U3871 (N_3871,N_2493,N_1907);
xnor U3872 (N_3872,N_1687,N_2442);
nor U3873 (N_3873,N_2793,N_2101);
nor U3874 (N_3874,N_2507,N_2779);
and U3875 (N_3875,N_2962,N_1566);
and U3876 (N_3876,N_2234,N_1840);
nor U3877 (N_3877,N_2800,N_1656);
or U3878 (N_3878,N_2093,N_2581);
nor U3879 (N_3879,N_2079,N_2933);
and U3880 (N_3880,N_2795,N_1882);
nor U3881 (N_3881,N_1788,N_2722);
nand U3882 (N_3882,N_2824,N_2432);
or U3883 (N_3883,N_2537,N_2406);
and U3884 (N_3884,N_2945,N_1562);
nand U3885 (N_3885,N_2013,N_1714);
xor U3886 (N_3886,N_1880,N_1524);
nand U3887 (N_3887,N_1581,N_2862);
nand U3888 (N_3888,N_2346,N_2009);
or U3889 (N_3889,N_2524,N_2583);
nand U3890 (N_3890,N_2451,N_1520);
or U3891 (N_3891,N_2942,N_2134);
or U3892 (N_3892,N_2330,N_2691);
nand U3893 (N_3893,N_1854,N_1593);
nor U3894 (N_3894,N_2882,N_1863);
and U3895 (N_3895,N_2238,N_1711);
nor U3896 (N_3896,N_1735,N_2643);
or U3897 (N_3897,N_1529,N_2409);
xnor U3898 (N_3898,N_1842,N_2255);
nand U3899 (N_3899,N_1513,N_1530);
or U3900 (N_3900,N_1868,N_2219);
nand U3901 (N_3901,N_2722,N_1541);
or U3902 (N_3902,N_2344,N_2079);
nand U3903 (N_3903,N_1851,N_2727);
nor U3904 (N_3904,N_1579,N_2443);
or U3905 (N_3905,N_2154,N_2664);
or U3906 (N_3906,N_2193,N_2560);
nor U3907 (N_3907,N_2763,N_2056);
nor U3908 (N_3908,N_1642,N_2824);
and U3909 (N_3909,N_2285,N_2891);
or U3910 (N_3910,N_2878,N_2714);
or U3911 (N_3911,N_2981,N_1835);
nor U3912 (N_3912,N_2360,N_1870);
nand U3913 (N_3913,N_2633,N_2189);
and U3914 (N_3914,N_2763,N_1927);
or U3915 (N_3915,N_1743,N_1595);
or U3916 (N_3916,N_1797,N_2201);
nor U3917 (N_3917,N_1564,N_2668);
nand U3918 (N_3918,N_1678,N_2967);
nor U3919 (N_3919,N_2906,N_1856);
and U3920 (N_3920,N_2465,N_2729);
nor U3921 (N_3921,N_1560,N_2542);
or U3922 (N_3922,N_2046,N_2569);
and U3923 (N_3923,N_1915,N_1614);
xnor U3924 (N_3924,N_2313,N_1921);
xnor U3925 (N_3925,N_1702,N_2469);
nand U3926 (N_3926,N_2913,N_2686);
and U3927 (N_3927,N_1964,N_2809);
and U3928 (N_3928,N_2299,N_1651);
and U3929 (N_3929,N_2412,N_2727);
or U3930 (N_3930,N_2869,N_2742);
and U3931 (N_3931,N_2845,N_2158);
nand U3932 (N_3932,N_2645,N_1537);
nand U3933 (N_3933,N_2706,N_2328);
nor U3934 (N_3934,N_1857,N_1599);
nand U3935 (N_3935,N_2511,N_2874);
or U3936 (N_3936,N_2073,N_2669);
nor U3937 (N_3937,N_2913,N_2481);
or U3938 (N_3938,N_2447,N_2644);
and U3939 (N_3939,N_1539,N_2171);
or U3940 (N_3940,N_2385,N_2839);
nand U3941 (N_3941,N_2527,N_2329);
nor U3942 (N_3942,N_1735,N_2363);
nor U3943 (N_3943,N_1852,N_2389);
and U3944 (N_3944,N_2764,N_1768);
or U3945 (N_3945,N_1614,N_1996);
and U3946 (N_3946,N_1986,N_2517);
and U3947 (N_3947,N_1620,N_1721);
or U3948 (N_3948,N_2113,N_2027);
nor U3949 (N_3949,N_1834,N_1642);
nand U3950 (N_3950,N_2606,N_1987);
nor U3951 (N_3951,N_2809,N_1750);
or U3952 (N_3952,N_1545,N_2652);
and U3953 (N_3953,N_2423,N_2180);
nor U3954 (N_3954,N_1989,N_2588);
xor U3955 (N_3955,N_2610,N_1526);
nor U3956 (N_3956,N_1946,N_1543);
nand U3957 (N_3957,N_2200,N_2914);
nand U3958 (N_3958,N_2565,N_2443);
or U3959 (N_3959,N_2426,N_2862);
nor U3960 (N_3960,N_1645,N_1803);
and U3961 (N_3961,N_2192,N_1993);
nor U3962 (N_3962,N_2934,N_2423);
or U3963 (N_3963,N_2665,N_2831);
nor U3964 (N_3964,N_1581,N_2882);
xor U3965 (N_3965,N_2606,N_2286);
nand U3966 (N_3966,N_2719,N_2239);
xor U3967 (N_3967,N_2506,N_2062);
nor U3968 (N_3968,N_2836,N_2786);
and U3969 (N_3969,N_1887,N_2808);
nand U3970 (N_3970,N_2473,N_1678);
nand U3971 (N_3971,N_2341,N_1960);
and U3972 (N_3972,N_1958,N_1923);
nor U3973 (N_3973,N_1921,N_2126);
nor U3974 (N_3974,N_1717,N_2114);
and U3975 (N_3975,N_2434,N_2825);
xnor U3976 (N_3976,N_2984,N_2202);
nand U3977 (N_3977,N_1930,N_2548);
and U3978 (N_3978,N_1753,N_2808);
and U3979 (N_3979,N_1971,N_1987);
nand U3980 (N_3980,N_1894,N_2446);
xor U3981 (N_3981,N_2403,N_1547);
or U3982 (N_3982,N_2828,N_1803);
or U3983 (N_3983,N_2738,N_2589);
nand U3984 (N_3984,N_2091,N_2320);
or U3985 (N_3985,N_2163,N_1848);
or U3986 (N_3986,N_2462,N_2178);
and U3987 (N_3987,N_2060,N_2119);
and U3988 (N_3988,N_1528,N_1907);
nand U3989 (N_3989,N_2029,N_1551);
nor U3990 (N_3990,N_2983,N_2092);
or U3991 (N_3991,N_2709,N_1811);
or U3992 (N_3992,N_2941,N_2580);
xor U3993 (N_3993,N_1846,N_1574);
or U3994 (N_3994,N_2417,N_2403);
and U3995 (N_3995,N_1584,N_1769);
nand U3996 (N_3996,N_2584,N_2929);
nand U3997 (N_3997,N_1809,N_2861);
nand U3998 (N_3998,N_1806,N_1716);
or U3999 (N_3999,N_2041,N_2319);
nor U4000 (N_4000,N_1981,N_1811);
and U4001 (N_4001,N_1593,N_2977);
nor U4002 (N_4002,N_2668,N_1502);
xor U4003 (N_4003,N_2930,N_1936);
or U4004 (N_4004,N_2441,N_2421);
or U4005 (N_4005,N_2360,N_1912);
or U4006 (N_4006,N_2165,N_2340);
nand U4007 (N_4007,N_2820,N_1693);
or U4008 (N_4008,N_1814,N_2586);
and U4009 (N_4009,N_2198,N_1528);
xnor U4010 (N_4010,N_2946,N_1756);
xor U4011 (N_4011,N_2374,N_2558);
or U4012 (N_4012,N_2639,N_2696);
nor U4013 (N_4013,N_2039,N_2108);
nor U4014 (N_4014,N_2071,N_2660);
nor U4015 (N_4015,N_2653,N_1654);
nand U4016 (N_4016,N_1598,N_2216);
nand U4017 (N_4017,N_2937,N_1916);
xnor U4018 (N_4018,N_2910,N_2675);
and U4019 (N_4019,N_1803,N_1823);
or U4020 (N_4020,N_2244,N_2325);
or U4021 (N_4021,N_1660,N_1656);
or U4022 (N_4022,N_2329,N_1558);
nor U4023 (N_4023,N_2482,N_2749);
and U4024 (N_4024,N_1853,N_2843);
nand U4025 (N_4025,N_2686,N_2165);
or U4026 (N_4026,N_2606,N_1704);
nor U4027 (N_4027,N_2615,N_1882);
xor U4028 (N_4028,N_2905,N_2347);
or U4029 (N_4029,N_2147,N_2086);
nand U4030 (N_4030,N_2658,N_2680);
nor U4031 (N_4031,N_1534,N_2568);
nor U4032 (N_4032,N_2641,N_2329);
or U4033 (N_4033,N_2747,N_1727);
nor U4034 (N_4034,N_2710,N_1519);
xor U4035 (N_4035,N_2697,N_1925);
xnor U4036 (N_4036,N_1944,N_2564);
or U4037 (N_4037,N_1584,N_2544);
and U4038 (N_4038,N_2975,N_2242);
and U4039 (N_4039,N_2531,N_2316);
nor U4040 (N_4040,N_2220,N_1973);
nand U4041 (N_4041,N_2659,N_1798);
nand U4042 (N_4042,N_2278,N_2168);
and U4043 (N_4043,N_2511,N_2876);
and U4044 (N_4044,N_2011,N_2340);
or U4045 (N_4045,N_1528,N_1604);
and U4046 (N_4046,N_2969,N_1658);
nand U4047 (N_4047,N_2306,N_2801);
nor U4048 (N_4048,N_2691,N_2866);
or U4049 (N_4049,N_2105,N_1832);
nand U4050 (N_4050,N_2551,N_2775);
or U4051 (N_4051,N_1525,N_2306);
and U4052 (N_4052,N_1517,N_2797);
nand U4053 (N_4053,N_2314,N_2936);
and U4054 (N_4054,N_1998,N_1760);
and U4055 (N_4055,N_2730,N_2279);
nor U4056 (N_4056,N_1631,N_2949);
and U4057 (N_4057,N_2095,N_2426);
nand U4058 (N_4058,N_2436,N_2279);
nand U4059 (N_4059,N_1514,N_2741);
or U4060 (N_4060,N_2373,N_2656);
nor U4061 (N_4061,N_2924,N_2286);
nand U4062 (N_4062,N_2036,N_1538);
nor U4063 (N_4063,N_2080,N_2147);
xor U4064 (N_4064,N_2916,N_2674);
nor U4065 (N_4065,N_2271,N_2095);
and U4066 (N_4066,N_1619,N_2098);
nand U4067 (N_4067,N_2515,N_2602);
xor U4068 (N_4068,N_2880,N_1736);
xor U4069 (N_4069,N_2927,N_1950);
and U4070 (N_4070,N_2388,N_2902);
nand U4071 (N_4071,N_1927,N_1568);
nor U4072 (N_4072,N_2769,N_2742);
and U4073 (N_4073,N_2047,N_1547);
and U4074 (N_4074,N_2707,N_2546);
or U4075 (N_4075,N_1940,N_1727);
and U4076 (N_4076,N_2882,N_2771);
or U4077 (N_4077,N_1859,N_2384);
and U4078 (N_4078,N_1904,N_1644);
or U4079 (N_4079,N_2965,N_1572);
nor U4080 (N_4080,N_2106,N_2323);
and U4081 (N_4081,N_2838,N_2823);
or U4082 (N_4082,N_1840,N_2036);
nor U4083 (N_4083,N_2984,N_2927);
nor U4084 (N_4084,N_2434,N_2381);
and U4085 (N_4085,N_2163,N_1811);
nor U4086 (N_4086,N_2054,N_1774);
nand U4087 (N_4087,N_2415,N_1803);
nand U4088 (N_4088,N_2695,N_2113);
or U4089 (N_4089,N_1581,N_1946);
and U4090 (N_4090,N_2778,N_2075);
and U4091 (N_4091,N_2408,N_2791);
or U4092 (N_4092,N_2985,N_2433);
and U4093 (N_4093,N_1812,N_1711);
nor U4094 (N_4094,N_2344,N_2129);
nand U4095 (N_4095,N_2108,N_1584);
nand U4096 (N_4096,N_2365,N_2961);
and U4097 (N_4097,N_1529,N_1810);
and U4098 (N_4098,N_2155,N_2542);
or U4099 (N_4099,N_1519,N_1605);
and U4100 (N_4100,N_2626,N_2894);
or U4101 (N_4101,N_2750,N_2976);
nor U4102 (N_4102,N_2413,N_1891);
nor U4103 (N_4103,N_2727,N_2812);
nor U4104 (N_4104,N_2895,N_2588);
nand U4105 (N_4105,N_2918,N_1950);
or U4106 (N_4106,N_1569,N_2362);
nand U4107 (N_4107,N_2844,N_1871);
or U4108 (N_4108,N_2229,N_2340);
nor U4109 (N_4109,N_2301,N_1557);
and U4110 (N_4110,N_1760,N_2925);
nand U4111 (N_4111,N_2662,N_1917);
nand U4112 (N_4112,N_1803,N_1890);
and U4113 (N_4113,N_2724,N_2091);
and U4114 (N_4114,N_2090,N_1533);
or U4115 (N_4115,N_1740,N_2959);
nand U4116 (N_4116,N_2848,N_1701);
nor U4117 (N_4117,N_1923,N_2543);
nor U4118 (N_4118,N_2943,N_1507);
and U4119 (N_4119,N_1692,N_1911);
nand U4120 (N_4120,N_1840,N_2926);
nand U4121 (N_4121,N_2400,N_1918);
nor U4122 (N_4122,N_1972,N_2204);
or U4123 (N_4123,N_2354,N_2122);
or U4124 (N_4124,N_2806,N_1840);
and U4125 (N_4125,N_2189,N_1571);
or U4126 (N_4126,N_2824,N_2383);
nor U4127 (N_4127,N_2971,N_1875);
and U4128 (N_4128,N_2300,N_1955);
and U4129 (N_4129,N_2093,N_2323);
nand U4130 (N_4130,N_1906,N_1958);
xor U4131 (N_4131,N_2358,N_1999);
and U4132 (N_4132,N_2095,N_1792);
nor U4133 (N_4133,N_2376,N_2666);
or U4134 (N_4134,N_2457,N_1893);
nor U4135 (N_4135,N_1502,N_1696);
nand U4136 (N_4136,N_2684,N_2713);
xnor U4137 (N_4137,N_1793,N_2323);
and U4138 (N_4138,N_2876,N_2178);
nor U4139 (N_4139,N_2615,N_2655);
nand U4140 (N_4140,N_1841,N_2032);
nor U4141 (N_4141,N_2115,N_2673);
or U4142 (N_4142,N_2129,N_2834);
and U4143 (N_4143,N_2516,N_2771);
and U4144 (N_4144,N_2293,N_2483);
nand U4145 (N_4145,N_2792,N_1681);
or U4146 (N_4146,N_1531,N_2765);
nand U4147 (N_4147,N_2530,N_2206);
nand U4148 (N_4148,N_2504,N_2997);
nor U4149 (N_4149,N_2756,N_2392);
nor U4150 (N_4150,N_1611,N_2446);
nand U4151 (N_4151,N_1857,N_1852);
and U4152 (N_4152,N_2509,N_1899);
xor U4153 (N_4153,N_2149,N_1707);
nand U4154 (N_4154,N_2646,N_2782);
nand U4155 (N_4155,N_1680,N_2188);
and U4156 (N_4156,N_2169,N_2077);
nand U4157 (N_4157,N_2593,N_2735);
nand U4158 (N_4158,N_2248,N_1550);
nand U4159 (N_4159,N_1851,N_2269);
and U4160 (N_4160,N_2722,N_2837);
nor U4161 (N_4161,N_2212,N_2261);
or U4162 (N_4162,N_2431,N_2765);
or U4163 (N_4163,N_2873,N_1694);
and U4164 (N_4164,N_2987,N_1609);
xor U4165 (N_4165,N_2678,N_2533);
and U4166 (N_4166,N_2861,N_1834);
or U4167 (N_4167,N_2007,N_1597);
and U4168 (N_4168,N_2276,N_1928);
nand U4169 (N_4169,N_2343,N_2757);
xnor U4170 (N_4170,N_1513,N_1618);
nor U4171 (N_4171,N_2450,N_2560);
and U4172 (N_4172,N_1885,N_1721);
nor U4173 (N_4173,N_2230,N_2643);
xnor U4174 (N_4174,N_2072,N_1580);
or U4175 (N_4175,N_1680,N_2295);
and U4176 (N_4176,N_1866,N_1836);
xnor U4177 (N_4177,N_2000,N_2930);
or U4178 (N_4178,N_2331,N_2278);
nand U4179 (N_4179,N_2912,N_2586);
nor U4180 (N_4180,N_2080,N_2685);
nor U4181 (N_4181,N_2494,N_2429);
nand U4182 (N_4182,N_1521,N_2227);
or U4183 (N_4183,N_2682,N_2861);
and U4184 (N_4184,N_2085,N_2828);
nor U4185 (N_4185,N_1704,N_2659);
nand U4186 (N_4186,N_2463,N_2871);
nand U4187 (N_4187,N_2988,N_2444);
or U4188 (N_4188,N_2809,N_1881);
nand U4189 (N_4189,N_2231,N_1500);
or U4190 (N_4190,N_1739,N_1756);
or U4191 (N_4191,N_2128,N_2722);
nor U4192 (N_4192,N_2477,N_2302);
and U4193 (N_4193,N_2685,N_2696);
or U4194 (N_4194,N_2903,N_2358);
nand U4195 (N_4195,N_2160,N_1632);
xor U4196 (N_4196,N_2750,N_1882);
nand U4197 (N_4197,N_1770,N_2561);
nand U4198 (N_4198,N_1732,N_2697);
nand U4199 (N_4199,N_2435,N_2962);
or U4200 (N_4200,N_2542,N_2772);
nor U4201 (N_4201,N_2294,N_1705);
nand U4202 (N_4202,N_2205,N_1999);
nor U4203 (N_4203,N_1792,N_2524);
nor U4204 (N_4204,N_2383,N_2044);
or U4205 (N_4205,N_2339,N_1959);
nor U4206 (N_4206,N_2577,N_1753);
nand U4207 (N_4207,N_2182,N_2916);
nand U4208 (N_4208,N_2467,N_1984);
xnor U4209 (N_4209,N_1560,N_1518);
or U4210 (N_4210,N_2877,N_2055);
and U4211 (N_4211,N_2305,N_2204);
and U4212 (N_4212,N_2119,N_1594);
and U4213 (N_4213,N_2461,N_1690);
nand U4214 (N_4214,N_1669,N_1550);
nor U4215 (N_4215,N_2582,N_2172);
and U4216 (N_4216,N_2976,N_2712);
nand U4217 (N_4217,N_1967,N_2274);
or U4218 (N_4218,N_1572,N_2628);
or U4219 (N_4219,N_2989,N_1871);
nand U4220 (N_4220,N_2995,N_2430);
nand U4221 (N_4221,N_2066,N_1943);
nor U4222 (N_4222,N_2781,N_2522);
nor U4223 (N_4223,N_2198,N_2822);
nand U4224 (N_4224,N_2658,N_1600);
and U4225 (N_4225,N_1659,N_2928);
or U4226 (N_4226,N_2300,N_2900);
or U4227 (N_4227,N_2375,N_2063);
or U4228 (N_4228,N_2061,N_2616);
nand U4229 (N_4229,N_2734,N_1714);
and U4230 (N_4230,N_2930,N_2873);
or U4231 (N_4231,N_2455,N_2692);
nand U4232 (N_4232,N_1991,N_2682);
and U4233 (N_4233,N_1914,N_1901);
and U4234 (N_4234,N_1985,N_2630);
or U4235 (N_4235,N_1731,N_1501);
xor U4236 (N_4236,N_2115,N_2575);
nand U4237 (N_4237,N_2871,N_2650);
nor U4238 (N_4238,N_2728,N_1757);
xor U4239 (N_4239,N_1557,N_2002);
nor U4240 (N_4240,N_2444,N_1796);
or U4241 (N_4241,N_1602,N_2949);
nor U4242 (N_4242,N_1551,N_2071);
nand U4243 (N_4243,N_2730,N_2746);
nor U4244 (N_4244,N_2558,N_2827);
or U4245 (N_4245,N_2230,N_2581);
or U4246 (N_4246,N_1824,N_1750);
and U4247 (N_4247,N_2763,N_2141);
and U4248 (N_4248,N_2369,N_2444);
nor U4249 (N_4249,N_1778,N_2780);
and U4250 (N_4250,N_2813,N_2887);
nor U4251 (N_4251,N_2876,N_2303);
nor U4252 (N_4252,N_2672,N_2626);
nand U4253 (N_4253,N_2363,N_2013);
xor U4254 (N_4254,N_1851,N_2214);
nand U4255 (N_4255,N_2192,N_2937);
and U4256 (N_4256,N_2311,N_1752);
and U4257 (N_4257,N_1958,N_2981);
and U4258 (N_4258,N_2464,N_2585);
or U4259 (N_4259,N_2702,N_1940);
nand U4260 (N_4260,N_1653,N_2157);
nand U4261 (N_4261,N_2387,N_1686);
nor U4262 (N_4262,N_2229,N_2197);
nor U4263 (N_4263,N_2549,N_2011);
nor U4264 (N_4264,N_2844,N_1775);
or U4265 (N_4265,N_2382,N_2750);
or U4266 (N_4266,N_2971,N_1537);
nand U4267 (N_4267,N_1919,N_2043);
and U4268 (N_4268,N_2534,N_2700);
or U4269 (N_4269,N_2836,N_1586);
or U4270 (N_4270,N_1821,N_2864);
or U4271 (N_4271,N_2120,N_1641);
nand U4272 (N_4272,N_1838,N_1536);
and U4273 (N_4273,N_2524,N_1546);
and U4274 (N_4274,N_2746,N_2415);
or U4275 (N_4275,N_2695,N_2204);
and U4276 (N_4276,N_2502,N_2470);
or U4277 (N_4277,N_2762,N_1676);
xnor U4278 (N_4278,N_2583,N_2496);
and U4279 (N_4279,N_1543,N_2993);
xnor U4280 (N_4280,N_2759,N_2165);
and U4281 (N_4281,N_2627,N_1704);
and U4282 (N_4282,N_2508,N_2334);
nand U4283 (N_4283,N_2749,N_2788);
and U4284 (N_4284,N_1897,N_2680);
nand U4285 (N_4285,N_1521,N_2377);
nor U4286 (N_4286,N_1943,N_2251);
nand U4287 (N_4287,N_2500,N_2656);
xnor U4288 (N_4288,N_2856,N_1917);
and U4289 (N_4289,N_1748,N_2444);
nand U4290 (N_4290,N_2018,N_2834);
nor U4291 (N_4291,N_2186,N_2688);
and U4292 (N_4292,N_2694,N_2486);
nor U4293 (N_4293,N_1940,N_2605);
and U4294 (N_4294,N_2975,N_2260);
nand U4295 (N_4295,N_2706,N_1982);
nor U4296 (N_4296,N_2981,N_1584);
or U4297 (N_4297,N_2205,N_1934);
or U4298 (N_4298,N_1737,N_2081);
nor U4299 (N_4299,N_2905,N_2685);
nand U4300 (N_4300,N_1763,N_1814);
and U4301 (N_4301,N_1716,N_1822);
nor U4302 (N_4302,N_2235,N_2609);
and U4303 (N_4303,N_1823,N_1686);
nand U4304 (N_4304,N_1790,N_1767);
and U4305 (N_4305,N_1987,N_2236);
nand U4306 (N_4306,N_1810,N_2474);
xor U4307 (N_4307,N_2471,N_2325);
or U4308 (N_4308,N_1591,N_1798);
nor U4309 (N_4309,N_2790,N_1951);
or U4310 (N_4310,N_2300,N_1566);
or U4311 (N_4311,N_1997,N_1629);
nand U4312 (N_4312,N_2492,N_1584);
and U4313 (N_4313,N_2942,N_1561);
nor U4314 (N_4314,N_2652,N_2399);
and U4315 (N_4315,N_1605,N_1771);
or U4316 (N_4316,N_2026,N_1642);
or U4317 (N_4317,N_1767,N_1659);
or U4318 (N_4318,N_1707,N_2749);
nor U4319 (N_4319,N_2343,N_1746);
xnor U4320 (N_4320,N_1654,N_2038);
and U4321 (N_4321,N_2380,N_2302);
and U4322 (N_4322,N_2874,N_2814);
nor U4323 (N_4323,N_2280,N_2061);
and U4324 (N_4324,N_2800,N_1945);
and U4325 (N_4325,N_1560,N_1755);
nor U4326 (N_4326,N_2560,N_2134);
xor U4327 (N_4327,N_1835,N_2367);
nand U4328 (N_4328,N_2107,N_1901);
and U4329 (N_4329,N_2780,N_2594);
and U4330 (N_4330,N_2052,N_1757);
nand U4331 (N_4331,N_2319,N_2481);
xor U4332 (N_4332,N_2573,N_1857);
nor U4333 (N_4333,N_1954,N_1828);
nand U4334 (N_4334,N_2765,N_2756);
or U4335 (N_4335,N_2785,N_1861);
and U4336 (N_4336,N_2532,N_1841);
nor U4337 (N_4337,N_1636,N_1997);
or U4338 (N_4338,N_1583,N_2377);
xnor U4339 (N_4339,N_1635,N_2912);
nand U4340 (N_4340,N_1961,N_1511);
and U4341 (N_4341,N_2776,N_1918);
nand U4342 (N_4342,N_1621,N_2057);
or U4343 (N_4343,N_1553,N_1613);
nor U4344 (N_4344,N_2068,N_2157);
and U4345 (N_4345,N_2596,N_2720);
nor U4346 (N_4346,N_2248,N_2692);
xnor U4347 (N_4347,N_1685,N_1878);
and U4348 (N_4348,N_2138,N_2305);
nand U4349 (N_4349,N_1544,N_1700);
and U4350 (N_4350,N_2487,N_1776);
nor U4351 (N_4351,N_1872,N_2829);
nand U4352 (N_4352,N_1942,N_2083);
or U4353 (N_4353,N_2797,N_2636);
or U4354 (N_4354,N_2575,N_1943);
or U4355 (N_4355,N_1560,N_1785);
nand U4356 (N_4356,N_2108,N_2624);
nor U4357 (N_4357,N_1825,N_2979);
nand U4358 (N_4358,N_1914,N_2989);
nand U4359 (N_4359,N_1585,N_1987);
and U4360 (N_4360,N_1911,N_2503);
or U4361 (N_4361,N_2485,N_1917);
and U4362 (N_4362,N_2482,N_2034);
and U4363 (N_4363,N_2553,N_2524);
nor U4364 (N_4364,N_2840,N_2899);
or U4365 (N_4365,N_2188,N_1983);
nor U4366 (N_4366,N_2355,N_2950);
and U4367 (N_4367,N_1600,N_2825);
or U4368 (N_4368,N_2506,N_1720);
nand U4369 (N_4369,N_1586,N_1822);
nand U4370 (N_4370,N_2801,N_1770);
or U4371 (N_4371,N_2721,N_2702);
or U4372 (N_4372,N_1503,N_2386);
or U4373 (N_4373,N_1718,N_2274);
or U4374 (N_4374,N_2790,N_1619);
or U4375 (N_4375,N_1877,N_1873);
nor U4376 (N_4376,N_1534,N_2362);
nand U4377 (N_4377,N_2563,N_2612);
or U4378 (N_4378,N_2522,N_1682);
nand U4379 (N_4379,N_2931,N_2708);
and U4380 (N_4380,N_1535,N_1926);
nand U4381 (N_4381,N_2340,N_2086);
and U4382 (N_4382,N_1789,N_1849);
nand U4383 (N_4383,N_2869,N_1793);
or U4384 (N_4384,N_2027,N_2862);
nor U4385 (N_4385,N_2724,N_2356);
nand U4386 (N_4386,N_1871,N_2984);
nor U4387 (N_4387,N_2658,N_2971);
nand U4388 (N_4388,N_2073,N_2984);
nand U4389 (N_4389,N_1970,N_1563);
nor U4390 (N_4390,N_1804,N_1953);
or U4391 (N_4391,N_2718,N_2639);
and U4392 (N_4392,N_2778,N_1863);
nand U4393 (N_4393,N_2537,N_2973);
nand U4394 (N_4394,N_1538,N_2541);
xnor U4395 (N_4395,N_2625,N_1898);
and U4396 (N_4396,N_2756,N_1649);
or U4397 (N_4397,N_2063,N_1527);
nand U4398 (N_4398,N_2684,N_2992);
or U4399 (N_4399,N_1790,N_1828);
or U4400 (N_4400,N_2743,N_2562);
nand U4401 (N_4401,N_2990,N_2878);
nand U4402 (N_4402,N_1990,N_2626);
or U4403 (N_4403,N_2646,N_2708);
xnor U4404 (N_4404,N_2611,N_1908);
or U4405 (N_4405,N_2923,N_2880);
nor U4406 (N_4406,N_2035,N_2332);
nand U4407 (N_4407,N_2758,N_1670);
nand U4408 (N_4408,N_1841,N_2533);
and U4409 (N_4409,N_2325,N_2433);
nand U4410 (N_4410,N_1503,N_2894);
nand U4411 (N_4411,N_1801,N_2156);
nand U4412 (N_4412,N_1725,N_2320);
nand U4413 (N_4413,N_2952,N_2052);
nand U4414 (N_4414,N_1731,N_1717);
nand U4415 (N_4415,N_2271,N_1686);
or U4416 (N_4416,N_1524,N_2145);
nand U4417 (N_4417,N_2767,N_1946);
nand U4418 (N_4418,N_1583,N_1812);
and U4419 (N_4419,N_2214,N_2629);
or U4420 (N_4420,N_2595,N_2228);
or U4421 (N_4421,N_2050,N_2095);
or U4422 (N_4422,N_2873,N_2541);
and U4423 (N_4423,N_1516,N_1910);
nand U4424 (N_4424,N_2724,N_2372);
xnor U4425 (N_4425,N_2827,N_2212);
or U4426 (N_4426,N_1807,N_2957);
or U4427 (N_4427,N_2773,N_2834);
nand U4428 (N_4428,N_2316,N_2375);
nand U4429 (N_4429,N_2100,N_1718);
or U4430 (N_4430,N_1934,N_2141);
nand U4431 (N_4431,N_1984,N_2706);
xor U4432 (N_4432,N_1617,N_2892);
xor U4433 (N_4433,N_1677,N_1773);
nor U4434 (N_4434,N_2302,N_2815);
nand U4435 (N_4435,N_1994,N_2066);
or U4436 (N_4436,N_1542,N_2205);
nand U4437 (N_4437,N_2624,N_2002);
or U4438 (N_4438,N_2175,N_1940);
and U4439 (N_4439,N_2480,N_2957);
and U4440 (N_4440,N_1619,N_2118);
xor U4441 (N_4441,N_2097,N_1631);
and U4442 (N_4442,N_2699,N_2987);
nor U4443 (N_4443,N_1519,N_2978);
nand U4444 (N_4444,N_2073,N_2031);
nor U4445 (N_4445,N_1780,N_2302);
nand U4446 (N_4446,N_2936,N_2242);
nand U4447 (N_4447,N_2944,N_2654);
nor U4448 (N_4448,N_2333,N_2630);
or U4449 (N_4449,N_2702,N_2092);
xnor U4450 (N_4450,N_2807,N_1535);
xnor U4451 (N_4451,N_2452,N_2335);
or U4452 (N_4452,N_2728,N_1502);
and U4453 (N_4453,N_1773,N_2225);
xnor U4454 (N_4454,N_2509,N_2895);
and U4455 (N_4455,N_1557,N_2415);
and U4456 (N_4456,N_2347,N_2101);
or U4457 (N_4457,N_2960,N_2232);
nor U4458 (N_4458,N_2012,N_1656);
nor U4459 (N_4459,N_2983,N_2484);
nor U4460 (N_4460,N_2545,N_1886);
nor U4461 (N_4461,N_2403,N_1720);
nand U4462 (N_4462,N_2850,N_2361);
or U4463 (N_4463,N_2406,N_1844);
nand U4464 (N_4464,N_2139,N_2348);
xor U4465 (N_4465,N_2374,N_1828);
and U4466 (N_4466,N_2897,N_1572);
nand U4467 (N_4467,N_1514,N_2426);
nand U4468 (N_4468,N_2296,N_2088);
nor U4469 (N_4469,N_2980,N_2068);
and U4470 (N_4470,N_2492,N_2139);
and U4471 (N_4471,N_2459,N_2993);
or U4472 (N_4472,N_1623,N_1772);
nand U4473 (N_4473,N_1587,N_1870);
nor U4474 (N_4474,N_2591,N_2933);
and U4475 (N_4475,N_2088,N_2820);
and U4476 (N_4476,N_1998,N_2319);
nand U4477 (N_4477,N_2506,N_2378);
or U4478 (N_4478,N_1909,N_2764);
xor U4479 (N_4479,N_2148,N_1916);
nor U4480 (N_4480,N_1958,N_2996);
nand U4481 (N_4481,N_2655,N_1534);
nor U4482 (N_4482,N_2815,N_2554);
and U4483 (N_4483,N_1769,N_1967);
or U4484 (N_4484,N_2500,N_2780);
nor U4485 (N_4485,N_1979,N_2649);
or U4486 (N_4486,N_2313,N_2455);
nor U4487 (N_4487,N_2381,N_2378);
nand U4488 (N_4488,N_2174,N_2069);
nor U4489 (N_4489,N_2053,N_2217);
xor U4490 (N_4490,N_2019,N_1863);
nor U4491 (N_4491,N_1950,N_2525);
or U4492 (N_4492,N_1990,N_1882);
and U4493 (N_4493,N_2804,N_2545);
and U4494 (N_4494,N_2101,N_2744);
or U4495 (N_4495,N_2096,N_2606);
xnor U4496 (N_4496,N_1726,N_2289);
nor U4497 (N_4497,N_2563,N_1690);
or U4498 (N_4498,N_1976,N_1833);
or U4499 (N_4499,N_2016,N_1933);
or U4500 (N_4500,N_3779,N_4219);
nand U4501 (N_4501,N_3241,N_3460);
or U4502 (N_4502,N_3987,N_4408);
and U4503 (N_4503,N_3323,N_4329);
xor U4504 (N_4504,N_3286,N_3840);
and U4505 (N_4505,N_3956,N_3978);
nor U4506 (N_4506,N_3683,N_3681);
nor U4507 (N_4507,N_4280,N_3447);
xnor U4508 (N_4508,N_3642,N_4295);
nand U4509 (N_4509,N_4416,N_3743);
and U4510 (N_4510,N_4396,N_3467);
or U4511 (N_4511,N_3153,N_4303);
nand U4512 (N_4512,N_3227,N_4201);
nand U4513 (N_4513,N_4334,N_3019);
nor U4514 (N_4514,N_3870,N_3098);
nor U4515 (N_4515,N_3458,N_3672);
and U4516 (N_4516,N_3992,N_4022);
or U4517 (N_4517,N_3977,N_4174);
and U4518 (N_4518,N_4037,N_3424);
nand U4519 (N_4519,N_3583,N_4133);
xnor U4520 (N_4520,N_4134,N_3169);
xor U4521 (N_4521,N_4002,N_3664);
nand U4522 (N_4522,N_3637,N_4340);
or U4523 (N_4523,N_3552,N_3224);
or U4524 (N_4524,N_4228,N_3395);
and U4525 (N_4525,N_3167,N_3414);
nor U4526 (N_4526,N_4252,N_3079);
nor U4527 (N_4527,N_4194,N_3633);
nor U4528 (N_4528,N_4302,N_4316);
nor U4529 (N_4529,N_3644,N_4063);
and U4530 (N_4530,N_3916,N_4333);
or U4531 (N_4531,N_4138,N_4311);
or U4532 (N_4532,N_3708,N_3666);
xnor U4533 (N_4533,N_3898,N_3364);
and U4534 (N_4534,N_3184,N_3839);
and U4535 (N_4535,N_3686,N_3551);
xor U4536 (N_4536,N_3385,N_3125);
xor U4537 (N_4537,N_3721,N_4075);
nor U4538 (N_4538,N_3906,N_3472);
and U4539 (N_4539,N_3556,N_3021);
or U4540 (N_4540,N_4341,N_3288);
and U4541 (N_4541,N_4042,N_4442);
and U4542 (N_4542,N_3762,N_4413);
nor U4543 (N_4543,N_3040,N_3730);
and U4544 (N_4544,N_3541,N_4218);
nor U4545 (N_4545,N_4166,N_4149);
or U4546 (N_4546,N_3381,N_4446);
nand U4547 (N_4547,N_3090,N_3028);
nand U4548 (N_4548,N_3111,N_4198);
or U4549 (N_4549,N_4139,N_4088);
nand U4550 (N_4550,N_4006,N_3256);
and U4551 (N_4551,N_3067,N_3187);
nand U4552 (N_4552,N_3397,N_3896);
nor U4553 (N_4553,N_3305,N_4077);
nand U4554 (N_4554,N_4026,N_3759);
and U4555 (N_4555,N_3426,N_4065);
and U4556 (N_4556,N_3110,N_3947);
and U4557 (N_4557,N_4232,N_3737);
nor U4558 (N_4558,N_3131,N_4010);
nand U4559 (N_4559,N_3190,N_3081);
nand U4560 (N_4560,N_3588,N_4122);
nand U4561 (N_4561,N_3272,N_3676);
nor U4562 (N_4562,N_3830,N_3496);
or U4563 (N_4563,N_3781,N_3359);
nand U4564 (N_4564,N_4444,N_4168);
and U4565 (N_4565,N_4216,N_3826);
or U4566 (N_4566,N_4058,N_3157);
or U4567 (N_4567,N_4241,N_4235);
and U4568 (N_4568,N_4143,N_3173);
and U4569 (N_4569,N_4220,N_3736);
xnor U4570 (N_4570,N_4369,N_3941);
xor U4571 (N_4571,N_3452,N_4274);
or U4572 (N_4572,N_3542,N_4182);
xnor U4573 (N_4573,N_4244,N_4494);
nor U4574 (N_4574,N_4205,N_4181);
and U4575 (N_4575,N_3907,N_4357);
nor U4576 (N_4576,N_3832,N_3069);
and U4577 (N_4577,N_4074,N_3035);
and U4578 (N_4578,N_3309,N_3599);
xor U4579 (N_4579,N_3484,N_3236);
nand U4580 (N_4580,N_3611,N_3905);
nand U4581 (N_4581,N_3124,N_3852);
nor U4582 (N_4582,N_3334,N_4150);
nand U4583 (N_4583,N_4217,N_4269);
or U4584 (N_4584,N_4435,N_3917);
or U4585 (N_4585,N_4136,N_3194);
xnor U4586 (N_4586,N_4422,N_3927);
and U4587 (N_4587,N_3833,N_4488);
nor U4588 (N_4588,N_3457,N_3842);
nor U4589 (N_4589,N_3471,N_4251);
nand U4590 (N_4590,N_4083,N_3527);
nand U4591 (N_4591,N_3219,N_3738);
and U4592 (N_4592,N_3147,N_3324);
nor U4593 (N_4593,N_4439,N_3586);
nor U4594 (N_4594,N_4076,N_3796);
and U4595 (N_4595,N_4484,N_3445);
nor U4596 (N_4596,N_4306,N_3281);
nor U4597 (N_4597,N_3198,N_3469);
nor U4598 (N_4598,N_4170,N_4210);
nor U4599 (N_4599,N_4095,N_3546);
and U4600 (N_4600,N_3902,N_4257);
xor U4601 (N_4601,N_4445,N_4278);
xnor U4602 (N_4602,N_3192,N_4381);
xor U4603 (N_4603,N_3861,N_3411);
and U4604 (N_4604,N_3302,N_3365);
nand U4605 (N_4605,N_3101,N_3126);
or U4606 (N_4606,N_3981,N_3547);
and U4607 (N_4607,N_3922,N_4009);
nor U4608 (N_4608,N_3073,N_4367);
or U4609 (N_4609,N_3604,N_3133);
and U4610 (N_4610,N_3972,N_3529);
nand U4611 (N_4611,N_3712,N_3605);
and U4612 (N_4612,N_3888,N_3382);
xor U4613 (N_4613,N_3439,N_3944);
nand U4614 (N_4614,N_3825,N_4068);
nor U4615 (N_4615,N_3294,N_3119);
nor U4616 (N_4616,N_3435,N_4346);
and U4617 (N_4617,N_3361,N_3874);
nand U4618 (N_4618,N_3549,N_3699);
nand U4619 (N_4619,N_3910,N_3348);
nand U4620 (N_4620,N_4188,N_3572);
and U4621 (N_4621,N_3533,N_3744);
nor U4622 (N_4622,N_4116,N_4014);
xnor U4623 (N_4623,N_3495,N_4052);
nor U4624 (N_4624,N_3798,N_3873);
nand U4625 (N_4625,N_3061,N_3008);
xnor U4626 (N_4626,N_3024,N_4415);
or U4627 (N_4627,N_3389,N_3540);
and U4628 (N_4628,N_3363,N_4067);
and U4629 (N_4629,N_4144,N_3568);
or U4630 (N_4630,N_3836,N_3523);
nor U4631 (N_4631,N_4394,N_4270);
and U4632 (N_4632,N_3399,N_3973);
xor U4633 (N_4633,N_4079,N_4043);
nor U4634 (N_4634,N_3319,N_3171);
xnor U4635 (N_4635,N_3632,N_3850);
nand U4636 (N_4636,N_3006,N_3161);
nor U4637 (N_4637,N_3786,N_4094);
nor U4638 (N_4638,N_4467,N_3204);
or U4639 (N_4639,N_3165,N_3827);
nand U4640 (N_4640,N_4392,N_3601);
and U4641 (N_4641,N_4407,N_3369);
xnor U4642 (N_4642,N_3525,N_3170);
nor U4643 (N_4643,N_3876,N_3217);
nor U4644 (N_4644,N_4045,N_4493);
nand U4645 (N_4645,N_3403,N_4487);
xor U4646 (N_4646,N_4363,N_3859);
or U4647 (N_4647,N_3433,N_3974);
xnor U4648 (N_4648,N_4403,N_4382);
or U4649 (N_4649,N_3934,N_3889);
nor U4650 (N_4650,N_4418,N_3473);
nor U4651 (N_4651,N_3921,N_3453);
or U4652 (N_4652,N_3657,N_3490);
or U4653 (N_4653,N_3392,N_3329);
or U4654 (N_4654,N_3248,N_3384);
or U4655 (N_4655,N_3690,N_4160);
or U4656 (N_4656,N_3314,N_3176);
nand U4657 (N_4657,N_3985,N_4425);
nor U4658 (N_4658,N_4368,N_4365);
nand U4659 (N_4659,N_3937,N_3474);
nand U4660 (N_4660,N_3865,N_3007);
or U4661 (N_4661,N_4126,N_3650);
xnor U4662 (N_4662,N_3229,N_3624);
nand U4663 (N_4663,N_3596,N_3506);
and U4664 (N_4664,N_4383,N_4154);
nor U4665 (N_4665,N_4214,N_3347);
or U4666 (N_4666,N_3320,N_3018);
nand U4667 (N_4667,N_3951,N_4438);
or U4668 (N_4668,N_4236,N_4495);
or U4669 (N_4669,N_3087,N_3408);
or U4670 (N_4670,N_4261,N_3052);
xor U4671 (N_4671,N_3429,N_3327);
and U4672 (N_4672,N_4080,N_3544);
nand U4673 (N_4673,N_4350,N_3567);
and U4674 (N_4674,N_3141,N_3520);
or U4675 (N_4675,N_4127,N_3377);
nand U4676 (N_4676,N_4344,N_3005);
nand U4677 (N_4677,N_3846,N_4040);
or U4678 (N_4678,N_3036,N_3579);
and U4679 (N_4679,N_4061,N_3986);
or U4680 (N_4680,N_3501,N_3116);
and U4681 (N_4681,N_3012,N_4410);
and U4682 (N_4682,N_3724,N_3380);
or U4683 (N_4683,N_3335,N_3741);
nand U4684 (N_4684,N_3488,N_4414);
xor U4685 (N_4685,N_3763,N_3162);
nor U4686 (N_4686,N_4498,N_3585);
and U4687 (N_4687,N_3441,N_3869);
and U4688 (N_4688,N_4480,N_4356);
and U4689 (N_4689,N_3145,N_4400);
nand U4690 (N_4690,N_4243,N_3750);
nor U4691 (N_4691,N_4451,N_3393);
and U4692 (N_4692,N_4049,N_4229);
nor U4693 (N_4693,N_4455,N_3310);
and U4694 (N_4694,N_3056,N_3748);
and U4695 (N_4695,N_3107,N_4212);
nand U4696 (N_4696,N_4427,N_4059);
or U4697 (N_4697,N_4288,N_3104);
or U4698 (N_4698,N_3963,N_4245);
or U4699 (N_4699,N_3267,N_4390);
or U4700 (N_4700,N_4070,N_4342);
nand U4701 (N_4701,N_3451,N_3275);
and U4702 (N_4702,N_3802,N_4432);
nor U4703 (N_4703,N_4175,N_3867);
and U4704 (N_4704,N_4277,N_4405);
nor U4705 (N_4705,N_3514,N_3276);
xor U4706 (N_4706,N_3476,N_3534);
nand U4707 (N_4707,N_3793,N_4215);
xnor U4708 (N_4708,N_3623,N_3720);
and U4709 (N_4709,N_4440,N_3371);
or U4710 (N_4710,N_4283,N_3622);
nor U4711 (N_4711,N_3918,N_4273);
or U4712 (N_4712,N_3091,N_3909);
or U4713 (N_4713,N_3423,N_3791);
or U4714 (N_4714,N_3487,N_3290);
or U4715 (N_4715,N_3716,N_3971);
and U4716 (N_4716,N_3123,N_3819);
or U4717 (N_4717,N_4072,N_3853);
and U4718 (N_4718,N_4366,N_4130);
or U4719 (N_4719,N_3270,N_3448);
xnor U4720 (N_4720,N_4259,N_4299);
nor U4721 (N_4721,N_3203,N_3769);
nor U4722 (N_4722,N_4486,N_3422);
nor U4723 (N_4723,N_4370,N_3128);
or U4724 (N_4724,N_3696,N_4128);
nand U4725 (N_4725,N_3331,N_3625);
and U4726 (N_4726,N_4179,N_3428);
or U4727 (N_4727,N_4066,N_3231);
nand U4728 (N_4728,N_3402,N_3265);
and U4729 (N_4729,N_3687,N_4264);
nand U4730 (N_4730,N_4073,N_4330);
nand U4731 (N_4731,N_4465,N_3560);
xor U4732 (N_4732,N_4475,N_4349);
nor U4733 (N_4733,N_4424,N_3945);
nor U4734 (N_4734,N_4098,N_3230);
xor U4735 (N_4735,N_3463,N_3046);
nand U4736 (N_4736,N_3077,N_3245);
and U4737 (N_4737,N_4419,N_4352);
nand U4738 (N_4738,N_3880,N_3096);
nand U4739 (N_4739,N_3595,N_4148);
and U4740 (N_4740,N_3026,N_3148);
and U4741 (N_4741,N_3692,N_3868);
nand U4742 (N_4742,N_4391,N_3780);
or U4743 (N_4743,N_3099,N_4000);
or U4744 (N_4744,N_4158,N_3935);
or U4745 (N_4745,N_4092,N_3015);
and U4746 (N_4746,N_3160,N_3903);
nand U4747 (N_4747,N_4393,N_3790);
nor U4748 (N_4748,N_3651,N_3718);
or U4749 (N_4749,N_4267,N_4119);
nand U4750 (N_4750,N_3197,N_3706);
or U4751 (N_4751,N_3114,N_3214);
and U4752 (N_4752,N_4191,N_4053);
and U4753 (N_4753,N_3800,N_4018);
and U4754 (N_4754,N_3232,N_3001);
nor U4755 (N_4755,N_3654,N_4492);
nor U4756 (N_4756,N_3185,N_4448);
and U4757 (N_4757,N_3698,N_4108);
nand U4758 (N_4758,N_3703,N_3419);
and U4759 (N_4759,N_4199,N_4189);
and U4760 (N_4760,N_3901,N_3949);
nor U4761 (N_4761,N_3795,N_3996);
or U4762 (N_4762,N_4019,N_3892);
nand U4763 (N_4763,N_4490,N_4031);
and U4764 (N_4764,N_3845,N_4239);
nor U4765 (N_4765,N_4025,N_3695);
or U4766 (N_4766,N_3349,N_4204);
and U4767 (N_4767,N_3031,N_3979);
and U4768 (N_4768,N_4271,N_3299);
nand U4769 (N_4769,N_3784,N_4300);
nand U4770 (N_4770,N_4282,N_4208);
nand U4771 (N_4771,N_3911,N_3884);
nor U4772 (N_4772,N_3834,N_3273);
or U4773 (N_4773,N_4101,N_4055);
or U4774 (N_4774,N_3117,N_4473);
and U4775 (N_4775,N_3094,N_3237);
nand U4776 (N_4776,N_3924,N_3044);
or U4777 (N_4777,N_3895,N_3225);
and U4778 (N_4778,N_3083,N_3966);
or U4779 (N_4779,N_3038,N_4472);
xor U4780 (N_4780,N_4364,N_3837);
nor U4781 (N_4781,N_3166,N_3020);
nor U4782 (N_4782,N_3564,N_3844);
nor U4783 (N_4783,N_3866,N_3089);
nand U4784 (N_4784,N_3831,N_3930);
nor U4785 (N_4785,N_3952,N_4436);
or U4786 (N_4786,N_4443,N_3756);
nand U4787 (N_4787,N_4355,N_3242);
nand U4788 (N_4788,N_3548,N_3082);
or U4789 (N_4789,N_3565,N_3068);
nand U4790 (N_4790,N_3912,N_3500);
or U4791 (N_4791,N_4331,N_3456);
nor U4792 (N_4792,N_4082,N_4041);
and U4793 (N_4793,N_3617,N_3358);
or U4794 (N_4794,N_4423,N_3396);
nor U4795 (N_4795,N_3355,N_3758);
nand U4796 (N_4796,N_3112,N_3969);
and U4797 (N_4797,N_3958,N_3444);
xnor U4798 (N_4798,N_3285,N_4089);
nor U4799 (N_4799,N_3156,N_3801);
and U4800 (N_4800,N_4429,N_3612);
nor U4801 (N_4801,N_3155,N_3394);
nor U4802 (N_4802,N_3813,N_3120);
xor U4803 (N_4803,N_4290,N_4406);
or U4804 (N_4804,N_4338,N_4348);
nor U4805 (N_4805,N_4113,N_4304);
nand U4806 (N_4806,N_3693,N_3961);
or U4807 (N_4807,N_3461,N_3339);
or U4808 (N_4808,N_4325,N_3266);
and U4809 (N_4809,N_3691,N_3530);
nor U4810 (N_4810,N_3726,N_3032);
nand U4811 (N_4811,N_3561,N_3881);
nor U4812 (N_4812,N_3278,N_3477);
nor U4813 (N_4813,N_3600,N_3747);
nand U4814 (N_4814,N_4001,N_3598);
nor U4815 (N_4815,N_3218,N_3356);
or U4816 (N_4816,N_3602,N_3746);
and U4817 (N_4817,N_4461,N_4362);
nand U4818 (N_4818,N_3516,N_3072);
xor U4819 (N_4819,N_4376,N_3988);
nand U4820 (N_4820,N_4032,N_3936);
nor U4821 (N_4821,N_3057,N_3550);
nor U4822 (N_4822,N_4140,N_4012);
and U4823 (N_4823,N_4151,N_4110);
nor U4824 (N_4824,N_3480,N_3191);
or U4825 (N_4825,N_4434,N_3647);
nand U4826 (N_4826,N_4230,N_3189);
nand U4827 (N_4827,N_3250,N_3725);
nor U4828 (N_4828,N_3606,N_3158);
and U4829 (N_4829,N_4377,N_4275);
xor U4830 (N_4830,N_3658,N_4293);
nand U4831 (N_4831,N_4183,N_4029);
and U4832 (N_4832,N_3163,N_4156);
nand U4833 (N_4833,N_3140,N_3254);
and U4834 (N_4834,N_4141,N_3055);
nor U4835 (N_4835,N_3920,N_3263);
and U4836 (N_4836,N_4456,N_3238);
and U4837 (N_4837,N_3159,N_4231);
and U4838 (N_4838,N_3584,N_3528);
nor U4839 (N_4839,N_4057,N_3482);
nor U4840 (N_4840,N_4421,N_3931);
or U4841 (N_4841,N_3841,N_3298);
nand U4842 (N_4842,N_3345,N_4114);
or U4843 (N_4843,N_3566,N_3206);
xnor U4844 (N_4844,N_3130,N_4260);
and U4845 (N_4845,N_4353,N_4384);
or U4846 (N_4846,N_4211,N_3915);
nor U4847 (N_4847,N_3492,N_3221);
nor U4848 (N_4848,N_3661,N_4086);
nand U4849 (N_4849,N_4386,N_3209);
and U4850 (N_4850,N_3416,N_3614);
nor U4851 (N_4851,N_3401,N_4142);
or U4852 (N_4852,N_3127,N_3521);
nor U4853 (N_4853,N_4279,N_3200);
or U4854 (N_4854,N_4431,N_4466);
or U4855 (N_4855,N_4004,N_3406);
and U4856 (N_4856,N_3731,N_4102);
nor U4857 (N_4857,N_3732,N_3092);
xor U4858 (N_4858,N_3249,N_4437);
or U4859 (N_4859,N_4310,N_4285);
nor U4860 (N_4860,N_4469,N_4048);
and U4861 (N_4861,N_4308,N_3631);
nor U4862 (N_4862,N_3220,N_4447);
nor U4863 (N_4863,N_4294,N_4450);
or U4864 (N_4864,N_3353,N_3054);
nor U4865 (N_4865,N_3244,N_4103);
or U4866 (N_4866,N_3485,N_3715);
or U4867 (N_4867,N_3053,N_3771);
nor U4868 (N_4868,N_3000,N_3269);
nor U4869 (N_4869,N_3727,N_3372);
and U4870 (N_4870,N_3878,N_4327);
nand U4871 (N_4871,N_4233,N_3591);
and U4872 (N_4872,N_3427,N_3593);
and U4873 (N_4873,N_3885,N_4096);
and U4874 (N_4874,N_3048,N_3667);
nor U4875 (N_4875,N_3459,N_4497);
nor U4876 (N_4876,N_3875,N_4246);
nor U4877 (N_4877,N_3291,N_3438);
nor U4878 (N_4878,N_4054,N_3627);
nor U4879 (N_4879,N_4195,N_3177);
nor U4880 (N_4880,N_3086,N_3014);
and U4881 (N_4881,N_4281,N_4258);
nor U4882 (N_4882,N_3538,N_3789);
xnor U4883 (N_4883,N_3150,N_3103);
and U4884 (N_4884,N_4343,N_3526);
or U4885 (N_4885,N_3649,N_3663);
or U4886 (N_4886,N_3948,N_3284);
and U4887 (N_4887,N_3351,N_3362);
nor U4888 (N_4888,N_3172,N_4153);
and U4889 (N_4889,N_4301,N_3494);
nor U4890 (N_4890,N_3900,N_3659);
xor U4891 (N_4891,N_3803,N_3264);
nand U4892 (N_4892,N_3388,N_3734);
nand U4893 (N_4893,N_3047,N_3709);
nand U4894 (N_4894,N_3199,N_3431);
nand U4895 (N_4895,N_3558,N_3222);
or U4896 (N_4896,N_3455,N_3811);
or U4897 (N_4897,N_3149,N_3675);
nand U4898 (N_4898,N_4132,N_3437);
nand U4899 (N_4899,N_3976,N_3761);
xor U4900 (N_4900,N_3407,N_3955);
nand U4901 (N_4901,N_3146,N_4309);
and U4902 (N_4902,N_3168,N_3645);
and U4903 (N_4903,N_4115,N_3300);
nand U4904 (N_4904,N_3325,N_3060);
xnor U4905 (N_4905,N_3694,N_3188);
and U4906 (N_4906,N_4359,N_3757);
nor U4907 (N_4907,N_3857,N_4206);
or U4908 (N_4908,N_4173,N_4155);
and U4909 (N_4909,N_3838,N_3536);
or U4910 (N_4910,N_4389,N_3717);
and U4911 (N_4911,N_3809,N_3289);
and U4912 (N_4912,N_3739,N_3806);
nand U4913 (N_4913,N_4387,N_3823);
nand U4914 (N_4914,N_3352,N_4047);
nand U4915 (N_4915,N_4091,N_3366);
nand U4916 (N_4916,N_4378,N_3573);
nor U4917 (N_4917,N_3860,N_3704);
nor U4918 (N_4918,N_4135,N_3822);
and U4919 (N_4919,N_3084,N_4499);
nor U4920 (N_4920,N_3665,N_3923);
nand U4921 (N_4921,N_4249,N_3563);
nand U4922 (N_4922,N_4192,N_4137);
nand U4923 (N_4923,N_3233,N_3680);
and U4924 (N_4924,N_3260,N_3387);
and U4925 (N_4925,N_3999,N_3466);
nor U4926 (N_4926,N_3807,N_3701);
nor U4927 (N_4927,N_4412,N_4462);
nand U4928 (N_4928,N_3571,N_3373);
xor U4929 (N_4929,N_3093,N_3328);
or U4930 (N_4930,N_3179,N_4147);
nand U4931 (N_4931,N_3505,N_3629);
nor U4932 (N_4932,N_3797,N_3064);
xnor U4933 (N_4933,N_3735,N_4162);
nor U4934 (N_4934,N_3071,N_3280);
xor U4935 (N_4935,N_3783,N_3995);
or U4936 (N_4936,N_3531,N_3940);
or U4937 (N_4937,N_3821,N_4064);
nand U4938 (N_4938,N_3926,N_3702);
nand U4939 (N_4939,N_3478,N_3315);
or U4940 (N_4940,N_4207,N_3368);
and U4941 (N_4941,N_4307,N_3182);
and U4942 (N_4942,N_4380,N_4324);
nor U4943 (N_4943,N_3522,N_4008);
nand U4944 (N_4944,N_3722,N_4268);
nor U4945 (N_4945,N_3297,N_3929);
nand U4946 (N_4946,N_3656,N_4417);
nor U4947 (N_4947,N_3980,N_4404);
or U4948 (N_4948,N_4225,N_4409);
nor U4949 (N_4949,N_4453,N_3287);
nand U4950 (N_4950,N_4374,N_3848);
and U4951 (N_4951,N_4109,N_3023);
or U4952 (N_4952,N_3178,N_3535);
nand U4953 (N_4953,N_3251,N_3764);
nor U4954 (N_4954,N_3894,N_3043);
or U4955 (N_4955,N_3343,N_3113);
and U4956 (N_4956,N_3223,N_3829);
and U4957 (N_4957,N_3740,N_3507);
nand U4958 (N_4958,N_3378,N_4056);
nor U4959 (N_4959,N_3076,N_3618);
and U4960 (N_4960,N_4118,N_4167);
or U4961 (N_4961,N_4123,N_3211);
or U4962 (N_4962,N_3333,N_4003);
or U4963 (N_4963,N_3555,N_3933);
xor U4964 (N_4964,N_3639,N_4388);
and U4965 (N_4965,N_4203,N_3041);
and U4966 (N_4966,N_4452,N_3193);
nor U4967 (N_4967,N_3835,N_3446);
nor U4968 (N_4968,N_3879,N_3375);
and U4969 (N_4969,N_3134,N_3643);
nor U4970 (N_4970,N_3578,N_4265);
or U4971 (N_4971,N_3982,N_3843);
nand U4972 (N_4972,N_4491,N_3964);
nor U4973 (N_4973,N_4069,N_4196);
and U4974 (N_4974,N_3886,N_3410);
nand U4975 (N_4975,N_3313,N_3713);
nand U4976 (N_4976,N_3050,N_3409);
nor U4977 (N_4977,N_3619,N_3205);
and U4978 (N_4978,N_3246,N_3174);
nor U4979 (N_4979,N_3653,N_4030);
nand U4980 (N_4980,N_4016,N_3095);
nand U4981 (N_4981,N_4379,N_4193);
nand U4982 (N_4982,N_3818,N_4411);
or U4983 (N_4983,N_3805,N_3186);
nand U4984 (N_4984,N_3752,N_3760);
nand U4985 (N_4985,N_3420,N_4081);
nor U4986 (N_4986,N_4313,N_4420);
nand U4987 (N_4987,N_3684,N_4399);
and U4988 (N_4988,N_4090,N_3671);
or U4989 (N_4989,N_3854,N_3518);
nand U4990 (N_4990,N_3367,N_4477);
or U4991 (N_4991,N_4426,N_3201);
nand U4992 (N_4992,N_3776,N_4152);
nand U4993 (N_4993,N_3181,N_3151);
nand U4994 (N_4994,N_4371,N_3468);
or U4995 (N_4995,N_3577,N_4197);
nand U4996 (N_4996,N_3804,N_4397);
nor U4997 (N_4997,N_3858,N_3129);
nand U4998 (N_4998,N_4255,N_3662);
nand U4999 (N_4999,N_4328,N_3212);
xor U5000 (N_5000,N_3493,N_4186);
and U5001 (N_5001,N_4161,N_4020);
or U5002 (N_5002,N_3062,N_3183);
and U5003 (N_5003,N_3322,N_3983);
and U5004 (N_5004,N_3855,N_4460);
xnor U5005 (N_5005,N_3465,N_3863);
nor U5006 (N_5006,N_3210,N_3580);
or U5007 (N_5007,N_3379,N_3570);
nand U5008 (N_5008,N_3346,N_3425);
nand U5009 (N_5009,N_4213,N_3962);
nor U5010 (N_5010,N_3959,N_3820);
or U5011 (N_5011,N_3648,N_3404);
xnor U5012 (N_5012,N_3688,N_3646);
nor U5013 (N_5013,N_3051,N_3135);
xnor U5014 (N_5014,N_3862,N_4483);
nor U5015 (N_5015,N_4100,N_3939);
xor U5016 (N_5016,N_3754,N_3772);
or U5017 (N_5017,N_3960,N_3308);
nor U5018 (N_5018,N_3215,N_3677);
xnor U5019 (N_5019,N_3295,N_4479);
and U5020 (N_5020,N_3226,N_4062);
nor U5021 (N_5021,N_3851,N_3318);
nand U5022 (N_5022,N_3228,N_4470);
and U5023 (N_5023,N_4385,N_3828);
and U5024 (N_5024,N_3635,N_3768);
and U5025 (N_5025,N_3705,N_3258);
nor U5026 (N_5026,N_4458,N_3432);
and U5027 (N_5027,N_3942,N_3011);
nor U5028 (N_5028,N_3626,N_3849);
nor U5029 (N_5029,N_4117,N_3418);
or U5030 (N_5030,N_3136,N_3815);
and U5031 (N_5031,N_4360,N_4209);
or U5032 (N_5032,N_4454,N_4250);
and U5033 (N_5033,N_4221,N_3872);
nor U5034 (N_5034,N_3042,N_4335);
nand U5035 (N_5035,N_4165,N_4084);
nor U5036 (N_5036,N_3271,N_3543);
nand U5037 (N_5037,N_4430,N_3301);
or U5038 (N_5038,N_4222,N_3033);
and U5039 (N_5039,N_4428,N_3239);
nand U5040 (N_5040,N_4289,N_3943);
and U5041 (N_5041,N_3016,N_3512);
and U5042 (N_5042,N_4305,N_3787);
nand U5043 (N_5043,N_4449,N_4373);
nor U5044 (N_5044,N_3357,N_3890);
nor U5045 (N_5045,N_3312,N_3252);
nor U5046 (N_5046,N_3714,N_3669);
or U5047 (N_5047,N_3470,N_3668);
and U5048 (N_5048,N_4286,N_3109);
or U5049 (N_5049,N_4071,N_3679);
or U5050 (N_5050,N_3799,N_3587);
nor U5051 (N_5051,N_3321,N_3581);
nor U5052 (N_5052,N_3519,N_3010);
nand U5053 (N_5053,N_4256,N_3088);
xnor U5054 (N_5054,N_4272,N_3443);
nand U5055 (N_5055,N_3508,N_4478);
nand U5056 (N_5056,N_4481,N_3652);
nand U5057 (N_5057,N_3785,N_4121);
nand U5058 (N_5058,N_3682,N_4332);
nor U5059 (N_5059,N_4011,N_3817);
and U5060 (N_5060,N_4489,N_4184);
nor U5061 (N_5061,N_3773,N_3967);
xor U5062 (N_5062,N_4051,N_3576);
nand U5063 (N_5063,N_3597,N_3070);
xnor U5064 (N_5064,N_3279,N_3932);
and U5065 (N_5065,N_3138,N_3034);
nand U5066 (N_5066,N_4253,N_3337);
xor U5067 (N_5067,N_3481,N_4202);
and U5068 (N_5068,N_3749,N_3017);
xor U5069 (N_5069,N_3569,N_3144);
and U5070 (N_5070,N_3350,N_4145);
nor U5071 (N_5071,N_4463,N_3066);
or U5072 (N_5072,N_3592,N_4007);
nand U5073 (N_5073,N_4180,N_4292);
and U5074 (N_5074,N_4457,N_3513);
nand U5075 (N_5075,N_3794,N_3537);
or U5076 (N_5076,N_3950,N_3511);
and U5077 (N_5077,N_3882,N_3274);
and U5078 (N_5078,N_3953,N_4078);
nor U5079 (N_5079,N_3607,N_3243);
nand U5080 (N_5080,N_4185,N_4023);
and U5081 (N_5081,N_3022,N_3774);
nor U5082 (N_5082,N_3697,N_3938);
nand U5083 (N_5083,N_4087,N_3253);
xnor U5084 (N_5084,N_3058,N_4319);
nor U5085 (N_5085,N_3891,N_4314);
nand U5086 (N_5086,N_3390,N_3984);
nor U5087 (N_5087,N_3234,N_4224);
nand U5088 (N_5088,N_3304,N_4169);
and U5089 (N_5089,N_4226,N_4125);
nand U5090 (N_5090,N_3195,N_4336);
or U5091 (N_5091,N_3499,N_3998);
xor U5092 (N_5092,N_3700,N_3386);
and U5093 (N_5093,N_4120,N_3913);
nand U5094 (N_5094,N_3317,N_3118);
or U5095 (N_5095,N_4223,N_3989);
nand U5096 (N_5096,N_3589,N_4298);
nand U5097 (N_5097,N_4320,N_3609);
and U5098 (N_5098,N_3914,N_3332);
xor U5099 (N_5099,N_4441,N_3994);
xor U5100 (N_5100,N_4358,N_4402);
and U5101 (N_5101,N_3608,N_3678);
or U5102 (N_5102,N_3616,N_3925);
nand U5103 (N_5103,N_3282,N_3808);
xor U5104 (N_5104,N_3792,N_4046);
or U5105 (N_5105,N_4178,N_4044);
nor U5106 (N_5106,N_3075,N_4005);
nand U5107 (N_5107,N_4482,N_4021);
nand U5108 (N_5108,N_3483,N_3504);
and U5109 (N_5109,N_3122,N_4395);
nor U5110 (N_5110,N_4159,N_3143);
or U5111 (N_5111,N_4190,N_3968);
nor U5112 (N_5112,N_3603,N_3449);
and U5113 (N_5113,N_3590,N_3400);
nor U5114 (N_5114,N_4291,N_3027);
and U5115 (N_5115,N_3670,N_3856);
nor U5116 (N_5116,N_3594,N_4106);
xor U5117 (N_5117,N_4099,N_4459);
nor U5118 (N_5118,N_4361,N_3311);
and U5119 (N_5119,N_3137,N_3660);
nand U5120 (N_5120,N_3037,N_4326);
nor U5121 (N_5121,N_4085,N_4024);
and U5122 (N_5122,N_4227,N_3341);
nor U5123 (N_5123,N_4287,N_3376);
xnor U5124 (N_5124,N_4237,N_4093);
nor U5125 (N_5125,N_3412,N_3919);
or U5126 (N_5126,N_3342,N_4107);
and U5127 (N_5127,N_3788,N_3154);
and U5128 (N_5128,N_3202,N_3338);
xor U5129 (N_5129,N_3991,N_3059);
nor U5130 (N_5130,N_3509,N_3562);
nor U5131 (N_5131,N_3306,N_3553);
nand U5132 (N_5132,N_4033,N_4104);
nor U5133 (N_5133,N_3899,N_3975);
and U5134 (N_5134,N_3078,N_3503);
nand U5135 (N_5135,N_3132,N_3711);
nor U5136 (N_5136,N_3778,N_3610);
nand U5137 (N_5137,N_4187,N_4315);
nor U5138 (N_5138,N_3782,N_3770);
or U5139 (N_5139,N_4254,N_3970);
or U5140 (N_5140,N_4323,N_3296);
nand U5141 (N_5141,N_3063,N_4284);
nor U5142 (N_5142,N_3142,N_3641);
and U5143 (N_5143,N_3723,N_3454);
nor U5144 (N_5144,N_3640,N_4297);
or U5145 (N_5145,N_3085,N_3340);
and U5146 (N_5146,N_3954,N_4238);
xor U5147 (N_5147,N_4296,N_3775);
and U5148 (N_5148,N_3100,N_3489);
or U5149 (N_5149,N_3957,N_4345);
and U5150 (N_5150,N_3436,N_3755);
and U5151 (N_5151,N_3559,N_4375);
nor U5152 (N_5152,N_3307,N_4263);
xnor U5153 (N_5153,N_3004,N_4177);
or U5154 (N_5154,N_3498,N_4013);
and U5155 (N_5155,N_3440,N_4015);
or U5156 (N_5156,N_3636,N_3097);
xnor U5157 (N_5157,N_3261,N_3719);
and U5158 (N_5158,N_3908,N_3383);
nor U5159 (N_5159,N_3421,N_3620);
nand U5160 (N_5160,N_3316,N_4322);
nor U5161 (N_5161,N_3216,N_3777);
xnor U5162 (N_5162,N_3326,N_4050);
nand U5163 (N_5163,N_3344,N_3030);
nand U5164 (N_5164,N_3398,N_4468);
nor U5165 (N_5165,N_4247,N_3767);
and U5166 (N_5166,N_3152,N_4398);
xor U5167 (N_5167,N_4034,N_4347);
or U5168 (N_5168,N_3883,N_4017);
or U5169 (N_5169,N_3336,N_3479);
nor U5170 (N_5170,N_4351,N_3106);
nor U5171 (N_5171,N_3121,N_4112);
and U5172 (N_5172,N_3283,N_3430);
nand U5173 (N_5173,N_3074,N_3532);
nand U5174 (N_5174,N_3517,N_4172);
nor U5175 (N_5175,N_3893,N_3707);
nand U5176 (N_5176,N_3904,N_4372);
or U5177 (N_5177,N_3655,N_4401);
or U5178 (N_5178,N_4234,N_3877);
and U5179 (N_5179,N_3557,N_3766);
or U5180 (N_5180,N_4200,N_3928);
or U5181 (N_5181,N_3293,N_3751);
and U5182 (N_5182,N_3450,N_3442);
xnor U5183 (N_5183,N_3235,N_3268);
and U5184 (N_5184,N_3080,N_3729);
nand U5185 (N_5185,N_3824,N_4485);
nor U5186 (N_5186,N_3049,N_3303);
and U5187 (N_5187,N_3621,N_3745);
xor U5188 (N_5188,N_4317,N_3065);
nor U5189 (N_5189,N_3582,N_3816);
or U5190 (N_5190,N_3009,N_4240);
or U5191 (N_5191,N_3180,N_4496);
nand U5192 (N_5192,N_3993,N_3330);
and U5193 (N_5193,N_3897,N_3257);
nor U5194 (N_5194,N_3689,N_4464);
nor U5195 (N_5195,N_3887,N_4060);
or U5196 (N_5196,N_3374,N_3196);
nor U5197 (N_5197,N_3262,N_3391);
and U5198 (N_5198,N_4028,N_3417);
xor U5199 (N_5199,N_3965,N_4476);
or U5200 (N_5200,N_3997,N_3628);
nor U5201 (N_5201,N_3370,N_3360);
nor U5202 (N_5202,N_3545,N_4105);
and U5203 (N_5203,N_3292,N_3108);
or U5204 (N_5204,N_3515,N_4312);
nor U5205 (N_5205,N_4248,N_3864);
or U5206 (N_5206,N_4433,N_4036);
or U5207 (N_5207,N_3102,N_4131);
nand U5208 (N_5208,N_4163,N_3491);
or U5209 (N_5209,N_3255,N_3025);
and U5210 (N_5210,N_3615,N_4321);
nor U5211 (N_5211,N_4242,N_4276);
and U5212 (N_5212,N_3039,N_3554);
and U5213 (N_5213,N_3208,N_3524);
nand U5214 (N_5214,N_3539,N_3003);
nand U5215 (N_5215,N_3105,N_4171);
nand U5216 (N_5216,N_3240,N_3674);
xor U5217 (N_5217,N_4176,N_3002);
or U5218 (N_5218,N_3673,N_3115);
nor U5219 (N_5219,N_3462,N_3510);
nor U5220 (N_5220,N_3405,N_3634);
and U5221 (N_5221,N_3575,N_3413);
or U5222 (N_5222,N_3638,N_3354);
or U5223 (N_5223,N_3812,N_4039);
nor U5224 (N_5224,N_3742,N_3810);
nor U5225 (N_5225,N_3728,N_4337);
and U5226 (N_5226,N_4027,N_3464);
nand U5227 (N_5227,N_3415,N_3990);
or U5228 (N_5228,N_3613,N_3207);
nor U5229 (N_5229,N_4471,N_3175);
and U5230 (N_5230,N_3434,N_4111);
nor U5231 (N_5231,N_3753,N_4157);
nor U5232 (N_5232,N_3259,N_3765);
nand U5233 (N_5233,N_3847,N_4262);
or U5234 (N_5234,N_3710,N_4474);
nor U5235 (N_5235,N_3814,N_4318);
nand U5236 (N_5236,N_4124,N_4164);
nor U5237 (N_5237,N_3029,N_4097);
nor U5238 (N_5238,N_3247,N_3164);
nor U5239 (N_5239,N_4354,N_3574);
nand U5240 (N_5240,N_3502,N_3497);
or U5241 (N_5241,N_3475,N_3013);
nor U5242 (N_5242,N_3871,N_3946);
nand U5243 (N_5243,N_4266,N_4035);
and U5244 (N_5244,N_4038,N_3045);
or U5245 (N_5245,N_3733,N_3486);
nand U5246 (N_5246,N_3630,N_3213);
nor U5247 (N_5247,N_3685,N_3277);
and U5248 (N_5248,N_4339,N_4146);
nand U5249 (N_5249,N_3139,N_4129);
and U5250 (N_5250,N_4286,N_3803);
and U5251 (N_5251,N_3338,N_3931);
nand U5252 (N_5252,N_3522,N_3544);
nor U5253 (N_5253,N_3412,N_4097);
or U5254 (N_5254,N_4096,N_3505);
and U5255 (N_5255,N_3815,N_4190);
and U5256 (N_5256,N_3980,N_4217);
or U5257 (N_5257,N_3417,N_3256);
nor U5258 (N_5258,N_3371,N_3506);
or U5259 (N_5259,N_3226,N_3012);
nor U5260 (N_5260,N_3895,N_4069);
and U5261 (N_5261,N_4228,N_4119);
nand U5262 (N_5262,N_4330,N_3558);
nand U5263 (N_5263,N_3406,N_3212);
or U5264 (N_5264,N_3057,N_4469);
or U5265 (N_5265,N_3241,N_3866);
nor U5266 (N_5266,N_3014,N_3597);
nor U5267 (N_5267,N_4442,N_3191);
and U5268 (N_5268,N_3815,N_4491);
or U5269 (N_5269,N_3752,N_3808);
nor U5270 (N_5270,N_3482,N_4276);
and U5271 (N_5271,N_4060,N_3046);
and U5272 (N_5272,N_4022,N_4060);
and U5273 (N_5273,N_3635,N_3132);
and U5274 (N_5274,N_3320,N_3568);
or U5275 (N_5275,N_3269,N_4177);
or U5276 (N_5276,N_4130,N_4313);
nand U5277 (N_5277,N_4427,N_3839);
and U5278 (N_5278,N_4231,N_3302);
or U5279 (N_5279,N_4034,N_3699);
xnor U5280 (N_5280,N_3617,N_4339);
or U5281 (N_5281,N_3022,N_4146);
nor U5282 (N_5282,N_4470,N_3925);
and U5283 (N_5283,N_3682,N_3121);
and U5284 (N_5284,N_3136,N_4343);
or U5285 (N_5285,N_3356,N_3406);
xnor U5286 (N_5286,N_3501,N_3282);
xnor U5287 (N_5287,N_4100,N_4253);
nand U5288 (N_5288,N_4072,N_4178);
and U5289 (N_5289,N_4127,N_4223);
nor U5290 (N_5290,N_4358,N_3257);
and U5291 (N_5291,N_3363,N_3721);
nor U5292 (N_5292,N_3931,N_3357);
nand U5293 (N_5293,N_3699,N_4112);
and U5294 (N_5294,N_3917,N_3193);
and U5295 (N_5295,N_4408,N_3488);
nor U5296 (N_5296,N_4024,N_3368);
xnor U5297 (N_5297,N_3291,N_3718);
nand U5298 (N_5298,N_3951,N_3591);
and U5299 (N_5299,N_3318,N_4315);
or U5300 (N_5300,N_3046,N_3798);
nor U5301 (N_5301,N_4080,N_4388);
and U5302 (N_5302,N_3723,N_3203);
nor U5303 (N_5303,N_4308,N_4484);
and U5304 (N_5304,N_4300,N_3513);
and U5305 (N_5305,N_3554,N_3585);
nor U5306 (N_5306,N_4383,N_3978);
or U5307 (N_5307,N_3729,N_3212);
nor U5308 (N_5308,N_3993,N_3713);
or U5309 (N_5309,N_3237,N_3454);
nand U5310 (N_5310,N_3515,N_3364);
and U5311 (N_5311,N_3221,N_3550);
nor U5312 (N_5312,N_4432,N_3188);
nor U5313 (N_5313,N_4214,N_3690);
and U5314 (N_5314,N_4317,N_3970);
nand U5315 (N_5315,N_3221,N_3036);
xor U5316 (N_5316,N_3217,N_3938);
and U5317 (N_5317,N_3974,N_4070);
nor U5318 (N_5318,N_3538,N_4226);
and U5319 (N_5319,N_3820,N_3204);
or U5320 (N_5320,N_3054,N_3986);
or U5321 (N_5321,N_3122,N_3970);
and U5322 (N_5322,N_3738,N_3941);
and U5323 (N_5323,N_4327,N_3588);
and U5324 (N_5324,N_3194,N_3154);
nand U5325 (N_5325,N_4348,N_3286);
and U5326 (N_5326,N_3008,N_4080);
nand U5327 (N_5327,N_4477,N_3140);
and U5328 (N_5328,N_3923,N_3597);
nand U5329 (N_5329,N_4455,N_3916);
nand U5330 (N_5330,N_3084,N_3069);
and U5331 (N_5331,N_3225,N_4399);
nand U5332 (N_5332,N_4340,N_3598);
and U5333 (N_5333,N_3636,N_3643);
nor U5334 (N_5334,N_4026,N_3267);
and U5335 (N_5335,N_3803,N_4473);
nor U5336 (N_5336,N_4269,N_4475);
nor U5337 (N_5337,N_3666,N_4397);
xor U5338 (N_5338,N_3604,N_3548);
nor U5339 (N_5339,N_3784,N_3003);
nor U5340 (N_5340,N_3101,N_3285);
nand U5341 (N_5341,N_4318,N_3087);
nand U5342 (N_5342,N_3816,N_3131);
or U5343 (N_5343,N_4086,N_4061);
or U5344 (N_5344,N_4126,N_3020);
xnor U5345 (N_5345,N_4128,N_4168);
or U5346 (N_5346,N_4363,N_3815);
or U5347 (N_5347,N_4204,N_4491);
nor U5348 (N_5348,N_3515,N_4427);
and U5349 (N_5349,N_4044,N_4497);
and U5350 (N_5350,N_3912,N_3907);
nand U5351 (N_5351,N_3841,N_3753);
and U5352 (N_5352,N_4172,N_4338);
nand U5353 (N_5353,N_4443,N_4076);
nor U5354 (N_5354,N_4213,N_4366);
or U5355 (N_5355,N_3182,N_3227);
xnor U5356 (N_5356,N_4014,N_4231);
nand U5357 (N_5357,N_4041,N_3048);
xor U5358 (N_5358,N_4415,N_3689);
or U5359 (N_5359,N_4348,N_4313);
nand U5360 (N_5360,N_3396,N_3224);
nor U5361 (N_5361,N_4005,N_3571);
nand U5362 (N_5362,N_3246,N_3680);
and U5363 (N_5363,N_4291,N_3481);
or U5364 (N_5364,N_3672,N_4379);
nand U5365 (N_5365,N_4042,N_3773);
nor U5366 (N_5366,N_3364,N_4105);
or U5367 (N_5367,N_4317,N_3854);
and U5368 (N_5368,N_4013,N_3794);
nor U5369 (N_5369,N_4102,N_4416);
nand U5370 (N_5370,N_3727,N_4053);
and U5371 (N_5371,N_3220,N_3033);
nor U5372 (N_5372,N_3423,N_3788);
and U5373 (N_5373,N_3759,N_3065);
xor U5374 (N_5374,N_3601,N_3405);
or U5375 (N_5375,N_3254,N_3366);
or U5376 (N_5376,N_4334,N_4044);
nand U5377 (N_5377,N_3510,N_4192);
or U5378 (N_5378,N_3773,N_4013);
or U5379 (N_5379,N_3140,N_3897);
xor U5380 (N_5380,N_4139,N_3615);
nor U5381 (N_5381,N_3320,N_3602);
nor U5382 (N_5382,N_3816,N_4282);
nor U5383 (N_5383,N_3997,N_4063);
nand U5384 (N_5384,N_4298,N_3678);
nand U5385 (N_5385,N_3510,N_3891);
and U5386 (N_5386,N_4295,N_3498);
nor U5387 (N_5387,N_3443,N_3537);
or U5388 (N_5388,N_4226,N_4289);
or U5389 (N_5389,N_3943,N_4101);
or U5390 (N_5390,N_3475,N_3346);
and U5391 (N_5391,N_4056,N_3584);
or U5392 (N_5392,N_4238,N_3169);
nor U5393 (N_5393,N_4284,N_3059);
nand U5394 (N_5394,N_3569,N_4016);
nand U5395 (N_5395,N_3051,N_3298);
nor U5396 (N_5396,N_3747,N_4052);
or U5397 (N_5397,N_3113,N_3645);
xor U5398 (N_5398,N_4311,N_3452);
nand U5399 (N_5399,N_3478,N_3148);
and U5400 (N_5400,N_3978,N_4135);
nor U5401 (N_5401,N_4478,N_3610);
nor U5402 (N_5402,N_3542,N_3461);
and U5403 (N_5403,N_4026,N_3333);
nand U5404 (N_5404,N_3008,N_3779);
or U5405 (N_5405,N_3806,N_3727);
xor U5406 (N_5406,N_3107,N_3777);
nand U5407 (N_5407,N_4322,N_3089);
xnor U5408 (N_5408,N_3024,N_4499);
and U5409 (N_5409,N_4339,N_3095);
or U5410 (N_5410,N_4110,N_4440);
nor U5411 (N_5411,N_4228,N_3726);
and U5412 (N_5412,N_3369,N_4360);
nor U5413 (N_5413,N_4338,N_4006);
or U5414 (N_5414,N_3954,N_3204);
nor U5415 (N_5415,N_3317,N_4222);
or U5416 (N_5416,N_3580,N_3937);
nand U5417 (N_5417,N_4220,N_3728);
nor U5418 (N_5418,N_4024,N_4463);
nand U5419 (N_5419,N_3115,N_3060);
xnor U5420 (N_5420,N_3205,N_4127);
xnor U5421 (N_5421,N_3463,N_4105);
nor U5422 (N_5422,N_3062,N_4079);
or U5423 (N_5423,N_3318,N_3553);
nor U5424 (N_5424,N_3610,N_4499);
nand U5425 (N_5425,N_3284,N_4207);
or U5426 (N_5426,N_4348,N_3673);
nand U5427 (N_5427,N_4274,N_4286);
and U5428 (N_5428,N_3895,N_3169);
and U5429 (N_5429,N_4309,N_3170);
and U5430 (N_5430,N_3391,N_3194);
or U5431 (N_5431,N_4396,N_4021);
or U5432 (N_5432,N_4201,N_3200);
and U5433 (N_5433,N_3454,N_3467);
and U5434 (N_5434,N_4054,N_4024);
nor U5435 (N_5435,N_3091,N_3372);
or U5436 (N_5436,N_3787,N_3273);
nand U5437 (N_5437,N_4055,N_3972);
nand U5438 (N_5438,N_4126,N_4419);
nor U5439 (N_5439,N_4322,N_4229);
or U5440 (N_5440,N_3766,N_4362);
nand U5441 (N_5441,N_4384,N_3707);
nand U5442 (N_5442,N_3207,N_4345);
xor U5443 (N_5443,N_3103,N_3285);
nand U5444 (N_5444,N_3773,N_3374);
or U5445 (N_5445,N_4123,N_4415);
nor U5446 (N_5446,N_3486,N_3081);
or U5447 (N_5447,N_3789,N_4006);
nor U5448 (N_5448,N_4441,N_3232);
or U5449 (N_5449,N_3961,N_4006);
and U5450 (N_5450,N_4172,N_3673);
and U5451 (N_5451,N_3037,N_3861);
nor U5452 (N_5452,N_3197,N_3297);
or U5453 (N_5453,N_3514,N_3679);
nor U5454 (N_5454,N_3615,N_4293);
and U5455 (N_5455,N_3954,N_4458);
nand U5456 (N_5456,N_3055,N_3930);
nand U5457 (N_5457,N_3809,N_3208);
nor U5458 (N_5458,N_3701,N_3198);
nand U5459 (N_5459,N_3792,N_4314);
or U5460 (N_5460,N_4246,N_3895);
or U5461 (N_5461,N_3012,N_4216);
nand U5462 (N_5462,N_3229,N_4495);
and U5463 (N_5463,N_4360,N_4191);
nand U5464 (N_5464,N_3894,N_3948);
nand U5465 (N_5465,N_3325,N_3594);
or U5466 (N_5466,N_4073,N_4212);
nor U5467 (N_5467,N_4004,N_3983);
nand U5468 (N_5468,N_3620,N_4092);
and U5469 (N_5469,N_3643,N_3333);
and U5470 (N_5470,N_3459,N_3684);
nand U5471 (N_5471,N_3626,N_3430);
xnor U5472 (N_5472,N_3375,N_4307);
nand U5473 (N_5473,N_3182,N_4375);
or U5474 (N_5474,N_4223,N_3448);
nor U5475 (N_5475,N_3701,N_3928);
nand U5476 (N_5476,N_3431,N_4465);
and U5477 (N_5477,N_3586,N_3347);
nor U5478 (N_5478,N_3869,N_4465);
nor U5479 (N_5479,N_3573,N_3717);
and U5480 (N_5480,N_3086,N_3008);
or U5481 (N_5481,N_3754,N_3782);
and U5482 (N_5482,N_4257,N_3172);
and U5483 (N_5483,N_4138,N_3794);
and U5484 (N_5484,N_3873,N_3191);
nor U5485 (N_5485,N_3670,N_3878);
and U5486 (N_5486,N_3485,N_3523);
or U5487 (N_5487,N_3698,N_4175);
nor U5488 (N_5488,N_4027,N_3419);
nand U5489 (N_5489,N_4346,N_3689);
nand U5490 (N_5490,N_3969,N_3028);
xor U5491 (N_5491,N_3018,N_4466);
and U5492 (N_5492,N_3688,N_3604);
xor U5493 (N_5493,N_3566,N_3392);
xnor U5494 (N_5494,N_4077,N_3927);
nor U5495 (N_5495,N_4070,N_4414);
nor U5496 (N_5496,N_3160,N_4077);
or U5497 (N_5497,N_3665,N_4230);
and U5498 (N_5498,N_3797,N_3979);
nand U5499 (N_5499,N_3499,N_3373);
or U5500 (N_5500,N_3981,N_3312);
nand U5501 (N_5501,N_4122,N_3751);
xnor U5502 (N_5502,N_3308,N_4114);
or U5503 (N_5503,N_3635,N_3852);
nor U5504 (N_5504,N_3085,N_3320);
or U5505 (N_5505,N_4198,N_4285);
and U5506 (N_5506,N_4311,N_4381);
nor U5507 (N_5507,N_3253,N_3505);
or U5508 (N_5508,N_3096,N_4185);
or U5509 (N_5509,N_3229,N_3998);
and U5510 (N_5510,N_4093,N_4190);
nand U5511 (N_5511,N_3174,N_3440);
nor U5512 (N_5512,N_3883,N_3461);
nor U5513 (N_5513,N_3522,N_3230);
nand U5514 (N_5514,N_3530,N_4384);
and U5515 (N_5515,N_3897,N_3990);
nand U5516 (N_5516,N_3121,N_3889);
xor U5517 (N_5517,N_3322,N_3954);
and U5518 (N_5518,N_3801,N_3248);
or U5519 (N_5519,N_3602,N_3711);
and U5520 (N_5520,N_4067,N_4469);
nor U5521 (N_5521,N_4331,N_3868);
and U5522 (N_5522,N_3534,N_4178);
xor U5523 (N_5523,N_3318,N_3719);
and U5524 (N_5524,N_4103,N_3642);
and U5525 (N_5525,N_3315,N_3934);
and U5526 (N_5526,N_4252,N_3053);
nand U5527 (N_5527,N_3491,N_3410);
and U5528 (N_5528,N_3926,N_3839);
nand U5529 (N_5529,N_3613,N_4260);
or U5530 (N_5530,N_3111,N_3261);
nand U5531 (N_5531,N_3993,N_3359);
nand U5532 (N_5532,N_3875,N_3039);
or U5533 (N_5533,N_3294,N_3696);
or U5534 (N_5534,N_4396,N_4406);
nor U5535 (N_5535,N_3843,N_3511);
nor U5536 (N_5536,N_4273,N_3901);
nor U5537 (N_5537,N_3844,N_4445);
or U5538 (N_5538,N_3207,N_3907);
or U5539 (N_5539,N_4261,N_4341);
nand U5540 (N_5540,N_3610,N_3847);
and U5541 (N_5541,N_4390,N_3673);
xor U5542 (N_5542,N_3316,N_3759);
nor U5543 (N_5543,N_3813,N_3103);
or U5544 (N_5544,N_4334,N_3583);
xor U5545 (N_5545,N_4024,N_3877);
or U5546 (N_5546,N_3392,N_3168);
nor U5547 (N_5547,N_4382,N_4204);
nor U5548 (N_5548,N_4450,N_3964);
or U5549 (N_5549,N_3178,N_3588);
nand U5550 (N_5550,N_4472,N_3774);
and U5551 (N_5551,N_3810,N_3620);
nor U5552 (N_5552,N_4192,N_4214);
and U5553 (N_5553,N_3719,N_3414);
nor U5554 (N_5554,N_4033,N_3020);
nor U5555 (N_5555,N_4199,N_3588);
or U5556 (N_5556,N_4404,N_3750);
and U5557 (N_5557,N_3951,N_3277);
and U5558 (N_5558,N_4319,N_4304);
nand U5559 (N_5559,N_4176,N_4272);
nand U5560 (N_5560,N_3220,N_3656);
nand U5561 (N_5561,N_3150,N_4232);
or U5562 (N_5562,N_3453,N_3577);
nor U5563 (N_5563,N_3465,N_3092);
nand U5564 (N_5564,N_4137,N_3383);
nor U5565 (N_5565,N_3904,N_3900);
and U5566 (N_5566,N_3466,N_3897);
and U5567 (N_5567,N_3270,N_3143);
nand U5568 (N_5568,N_4349,N_4489);
and U5569 (N_5569,N_4062,N_4182);
or U5570 (N_5570,N_3595,N_4038);
nor U5571 (N_5571,N_4078,N_3952);
xor U5572 (N_5572,N_4047,N_3678);
nand U5573 (N_5573,N_3495,N_4158);
and U5574 (N_5574,N_3352,N_3753);
nand U5575 (N_5575,N_4274,N_3489);
nor U5576 (N_5576,N_4192,N_3614);
nor U5577 (N_5577,N_4430,N_3662);
nor U5578 (N_5578,N_3670,N_3890);
and U5579 (N_5579,N_4019,N_4309);
or U5580 (N_5580,N_4181,N_4045);
or U5581 (N_5581,N_3145,N_4368);
or U5582 (N_5582,N_3398,N_4246);
and U5583 (N_5583,N_3306,N_3095);
nor U5584 (N_5584,N_3695,N_3759);
nand U5585 (N_5585,N_3343,N_3960);
nor U5586 (N_5586,N_3380,N_3695);
or U5587 (N_5587,N_3154,N_3310);
xor U5588 (N_5588,N_4034,N_4193);
or U5589 (N_5589,N_3231,N_3476);
nand U5590 (N_5590,N_3255,N_4217);
nand U5591 (N_5591,N_3074,N_3268);
nor U5592 (N_5592,N_3719,N_4056);
nor U5593 (N_5593,N_4104,N_4361);
xor U5594 (N_5594,N_3783,N_3977);
nor U5595 (N_5595,N_4490,N_3364);
nor U5596 (N_5596,N_3894,N_4046);
and U5597 (N_5597,N_3717,N_4094);
nand U5598 (N_5598,N_3275,N_4179);
nand U5599 (N_5599,N_3963,N_4019);
nand U5600 (N_5600,N_3180,N_3050);
and U5601 (N_5601,N_4091,N_4211);
nand U5602 (N_5602,N_4289,N_3309);
xnor U5603 (N_5603,N_4433,N_3131);
or U5604 (N_5604,N_3120,N_3174);
or U5605 (N_5605,N_4293,N_4439);
or U5606 (N_5606,N_4072,N_3216);
and U5607 (N_5607,N_4036,N_3918);
and U5608 (N_5608,N_4085,N_4455);
or U5609 (N_5609,N_3762,N_4399);
nand U5610 (N_5610,N_3442,N_3227);
xnor U5611 (N_5611,N_3695,N_3151);
or U5612 (N_5612,N_3785,N_3880);
nand U5613 (N_5613,N_3532,N_3320);
or U5614 (N_5614,N_3812,N_3325);
xnor U5615 (N_5615,N_3279,N_3053);
and U5616 (N_5616,N_4435,N_3339);
nand U5617 (N_5617,N_3125,N_3216);
nor U5618 (N_5618,N_4243,N_4152);
nor U5619 (N_5619,N_4058,N_3132);
and U5620 (N_5620,N_3844,N_4276);
xnor U5621 (N_5621,N_3382,N_3017);
and U5622 (N_5622,N_3639,N_3170);
or U5623 (N_5623,N_3106,N_3502);
nor U5624 (N_5624,N_3497,N_3492);
nor U5625 (N_5625,N_3238,N_3861);
and U5626 (N_5626,N_3381,N_3356);
or U5627 (N_5627,N_3508,N_3254);
nand U5628 (N_5628,N_3412,N_4350);
or U5629 (N_5629,N_3304,N_3120);
nand U5630 (N_5630,N_3769,N_4073);
and U5631 (N_5631,N_3885,N_4072);
nand U5632 (N_5632,N_3547,N_3170);
nor U5633 (N_5633,N_3506,N_3523);
nor U5634 (N_5634,N_3961,N_3987);
and U5635 (N_5635,N_4424,N_4311);
or U5636 (N_5636,N_3807,N_3005);
or U5637 (N_5637,N_3072,N_4283);
nand U5638 (N_5638,N_3103,N_4263);
or U5639 (N_5639,N_4221,N_3589);
nand U5640 (N_5640,N_4088,N_3852);
nor U5641 (N_5641,N_3705,N_3061);
nor U5642 (N_5642,N_4038,N_4332);
nor U5643 (N_5643,N_3382,N_4099);
nor U5644 (N_5644,N_3718,N_3288);
or U5645 (N_5645,N_3181,N_3422);
and U5646 (N_5646,N_3549,N_3843);
nand U5647 (N_5647,N_3049,N_3826);
nand U5648 (N_5648,N_3767,N_3484);
nand U5649 (N_5649,N_3127,N_4257);
nor U5650 (N_5650,N_3625,N_4336);
or U5651 (N_5651,N_3723,N_3705);
or U5652 (N_5652,N_4403,N_3891);
or U5653 (N_5653,N_4237,N_4230);
or U5654 (N_5654,N_3037,N_4253);
nor U5655 (N_5655,N_4407,N_3800);
nand U5656 (N_5656,N_4368,N_3638);
nand U5657 (N_5657,N_3118,N_3271);
nor U5658 (N_5658,N_4302,N_3300);
nor U5659 (N_5659,N_3004,N_3863);
and U5660 (N_5660,N_3463,N_4299);
or U5661 (N_5661,N_3093,N_3830);
or U5662 (N_5662,N_4192,N_3224);
and U5663 (N_5663,N_4466,N_3096);
and U5664 (N_5664,N_3236,N_3199);
and U5665 (N_5665,N_3971,N_3822);
nor U5666 (N_5666,N_4336,N_4343);
or U5667 (N_5667,N_3062,N_4408);
or U5668 (N_5668,N_3983,N_3318);
or U5669 (N_5669,N_3139,N_3340);
or U5670 (N_5670,N_3029,N_4213);
nor U5671 (N_5671,N_3469,N_3680);
or U5672 (N_5672,N_4230,N_4027);
nor U5673 (N_5673,N_4012,N_3714);
nor U5674 (N_5674,N_4038,N_4026);
or U5675 (N_5675,N_3320,N_3216);
and U5676 (N_5676,N_4245,N_3962);
nand U5677 (N_5677,N_3605,N_3555);
nand U5678 (N_5678,N_4058,N_3824);
or U5679 (N_5679,N_3934,N_3437);
nand U5680 (N_5680,N_3397,N_3214);
nor U5681 (N_5681,N_4313,N_3535);
or U5682 (N_5682,N_4116,N_3051);
nor U5683 (N_5683,N_4396,N_4336);
xnor U5684 (N_5684,N_3101,N_4371);
nand U5685 (N_5685,N_3935,N_4343);
or U5686 (N_5686,N_4222,N_4258);
nor U5687 (N_5687,N_3835,N_3983);
nand U5688 (N_5688,N_4057,N_3042);
nand U5689 (N_5689,N_3436,N_3704);
xnor U5690 (N_5690,N_3660,N_3360);
or U5691 (N_5691,N_3351,N_3503);
or U5692 (N_5692,N_3560,N_4421);
nand U5693 (N_5693,N_4155,N_4137);
nor U5694 (N_5694,N_4353,N_3808);
nor U5695 (N_5695,N_3347,N_4197);
nand U5696 (N_5696,N_4395,N_4455);
nand U5697 (N_5697,N_4122,N_3079);
and U5698 (N_5698,N_4070,N_3408);
or U5699 (N_5699,N_3058,N_4348);
and U5700 (N_5700,N_4114,N_4129);
xnor U5701 (N_5701,N_3798,N_3041);
and U5702 (N_5702,N_3274,N_4378);
nor U5703 (N_5703,N_3767,N_3495);
nand U5704 (N_5704,N_3130,N_3795);
nand U5705 (N_5705,N_3602,N_3213);
nand U5706 (N_5706,N_3109,N_3136);
or U5707 (N_5707,N_3720,N_3627);
nand U5708 (N_5708,N_4109,N_3915);
xor U5709 (N_5709,N_3903,N_3574);
nand U5710 (N_5710,N_4029,N_4280);
nand U5711 (N_5711,N_4232,N_3354);
and U5712 (N_5712,N_3755,N_3444);
or U5713 (N_5713,N_4102,N_4232);
nor U5714 (N_5714,N_3569,N_3900);
or U5715 (N_5715,N_3407,N_4165);
or U5716 (N_5716,N_3948,N_3624);
nor U5717 (N_5717,N_3321,N_3850);
nor U5718 (N_5718,N_4307,N_3641);
xor U5719 (N_5719,N_3955,N_3626);
nor U5720 (N_5720,N_4244,N_3389);
and U5721 (N_5721,N_3438,N_3514);
nand U5722 (N_5722,N_3612,N_3971);
nand U5723 (N_5723,N_3273,N_3338);
and U5724 (N_5724,N_3603,N_4114);
nand U5725 (N_5725,N_4339,N_3894);
nand U5726 (N_5726,N_3465,N_4236);
xnor U5727 (N_5727,N_3911,N_4069);
and U5728 (N_5728,N_3166,N_4134);
nand U5729 (N_5729,N_4271,N_3290);
xor U5730 (N_5730,N_4155,N_3643);
nor U5731 (N_5731,N_3305,N_3429);
nor U5732 (N_5732,N_3796,N_3785);
nor U5733 (N_5733,N_4252,N_3113);
or U5734 (N_5734,N_3321,N_3277);
and U5735 (N_5735,N_3288,N_3314);
and U5736 (N_5736,N_4038,N_3061);
nor U5737 (N_5737,N_4030,N_3812);
nor U5738 (N_5738,N_3225,N_3853);
or U5739 (N_5739,N_3950,N_3651);
nor U5740 (N_5740,N_3873,N_3645);
nor U5741 (N_5741,N_4248,N_3449);
xnor U5742 (N_5742,N_4090,N_3686);
nor U5743 (N_5743,N_3974,N_3693);
nor U5744 (N_5744,N_3962,N_4133);
nand U5745 (N_5745,N_3846,N_3902);
and U5746 (N_5746,N_4438,N_3545);
and U5747 (N_5747,N_4381,N_4459);
and U5748 (N_5748,N_4441,N_3902);
or U5749 (N_5749,N_4163,N_4036);
or U5750 (N_5750,N_3305,N_4493);
nand U5751 (N_5751,N_4152,N_3757);
xor U5752 (N_5752,N_3975,N_3950);
xor U5753 (N_5753,N_3675,N_3940);
and U5754 (N_5754,N_4303,N_4357);
and U5755 (N_5755,N_3139,N_4360);
and U5756 (N_5756,N_4012,N_3010);
nor U5757 (N_5757,N_4018,N_3921);
nor U5758 (N_5758,N_3891,N_3150);
nand U5759 (N_5759,N_3841,N_3230);
or U5760 (N_5760,N_4038,N_4062);
or U5761 (N_5761,N_3204,N_3231);
nand U5762 (N_5762,N_3433,N_3256);
and U5763 (N_5763,N_3108,N_3671);
nor U5764 (N_5764,N_3215,N_3020);
nand U5765 (N_5765,N_4332,N_3934);
and U5766 (N_5766,N_3031,N_3622);
nor U5767 (N_5767,N_3988,N_3742);
xor U5768 (N_5768,N_3711,N_3835);
nor U5769 (N_5769,N_3896,N_3177);
nor U5770 (N_5770,N_4014,N_3329);
and U5771 (N_5771,N_3800,N_3786);
and U5772 (N_5772,N_3826,N_4323);
nor U5773 (N_5773,N_4169,N_4157);
nor U5774 (N_5774,N_3938,N_3761);
or U5775 (N_5775,N_3080,N_4297);
nand U5776 (N_5776,N_3610,N_3162);
nor U5777 (N_5777,N_4019,N_3257);
nor U5778 (N_5778,N_4140,N_3880);
nand U5779 (N_5779,N_3226,N_3289);
nand U5780 (N_5780,N_4026,N_4363);
nand U5781 (N_5781,N_4165,N_4255);
nand U5782 (N_5782,N_3449,N_4050);
nand U5783 (N_5783,N_3264,N_4278);
or U5784 (N_5784,N_3766,N_3135);
or U5785 (N_5785,N_3393,N_4422);
nand U5786 (N_5786,N_3255,N_3961);
or U5787 (N_5787,N_3726,N_4346);
nand U5788 (N_5788,N_3491,N_3594);
and U5789 (N_5789,N_3315,N_4328);
or U5790 (N_5790,N_3073,N_4487);
nor U5791 (N_5791,N_4321,N_4133);
nor U5792 (N_5792,N_4321,N_4384);
nor U5793 (N_5793,N_4374,N_3174);
and U5794 (N_5794,N_3367,N_3929);
xnor U5795 (N_5795,N_4250,N_3082);
nor U5796 (N_5796,N_3159,N_3198);
or U5797 (N_5797,N_3594,N_3869);
nand U5798 (N_5798,N_3328,N_3016);
nor U5799 (N_5799,N_3589,N_3424);
and U5800 (N_5800,N_4366,N_3812);
or U5801 (N_5801,N_3186,N_3371);
and U5802 (N_5802,N_3540,N_3193);
xnor U5803 (N_5803,N_3957,N_3034);
nand U5804 (N_5804,N_3721,N_3624);
or U5805 (N_5805,N_3188,N_3894);
or U5806 (N_5806,N_3935,N_3065);
nand U5807 (N_5807,N_3190,N_3075);
and U5808 (N_5808,N_3432,N_4177);
or U5809 (N_5809,N_3792,N_4435);
nor U5810 (N_5810,N_3243,N_4208);
and U5811 (N_5811,N_4061,N_3946);
or U5812 (N_5812,N_3168,N_4027);
nor U5813 (N_5813,N_3350,N_3234);
and U5814 (N_5814,N_4351,N_4249);
nor U5815 (N_5815,N_3499,N_4218);
nor U5816 (N_5816,N_3823,N_4344);
and U5817 (N_5817,N_3347,N_4456);
nor U5818 (N_5818,N_4234,N_3079);
nor U5819 (N_5819,N_3435,N_3028);
nor U5820 (N_5820,N_4457,N_4173);
xnor U5821 (N_5821,N_3608,N_3375);
and U5822 (N_5822,N_3502,N_3147);
nand U5823 (N_5823,N_4455,N_3792);
or U5824 (N_5824,N_3458,N_3922);
or U5825 (N_5825,N_3918,N_4372);
or U5826 (N_5826,N_3304,N_4186);
nor U5827 (N_5827,N_3525,N_3658);
or U5828 (N_5828,N_3069,N_3271);
or U5829 (N_5829,N_3016,N_3867);
nand U5830 (N_5830,N_3648,N_3673);
and U5831 (N_5831,N_3116,N_3557);
xnor U5832 (N_5832,N_3205,N_3827);
nor U5833 (N_5833,N_3955,N_3435);
or U5834 (N_5834,N_3330,N_3567);
nor U5835 (N_5835,N_4281,N_4245);
or U5836 (N_5836,N_3405,N_4074);
nor U5837 (N_5837,N_3502,N_3423);
and U5838 (N_5838,N_3324,N_3801);
and U5839 (N_5839,N_3850,N_3878);
and U5840 (N_5840,N_4259,N_4295);
xor U5841 (N_5841,N_4354,N_4125);
and U5842 (N_5842,N_3286,N_3818);
or U5843 (N_5843,N_3420,N_3398);
nor U5844 (N_5844,N_3704,N_3950);
nor U5845 (N_5845,N_4031,N_4140);
nand U5846 (N_5846,N_3651,N_3434);
and U5847 (N_5847,N_3435,N_3293);
nor U5848 (N_5848,N_4445,N_3392);
nand U5849 (N_5849,N_3778,N_3152);
and U5850 (N_5850,N_3632,N_3732);
or U5851 (N_5851,N_3945,N_3502);
nand U5852 (N_5852,N_3432,N_3769);
nand U5853 (N_5853,N_4370,N_4336);
or U5854 (N_5854,N_4137,N_3535);
or U5855 (N_5855,N_4338,N_4005);
xnor U5856 (N_5856,N_3976,N_3275);
nor U5857 (N_5857,N_4390,N_4125);
or U5858 (N_5858,N_3097,N_3918);
and U5859 (N_5859,N_3106,N_3012);
nor U5860 (N_5860,N_4254,N_3812);
or U5861 (N_5861,N_3192,N_3534);
or U5862 (N_5862,N_3220,N_3224);
xnor U5863 (N_5863,N_3827,N_3360);
and U5864 (N_5864,N_3508,N_3229);
or U5865 (N_5865,N_3226,N_3785);
or U5866 (N_5866,N_4233,N_4290);
nand U5867 (N_5867,N_3936,N_3504);
or U5868 (N_5868,N_3225,N_3735);
and U5869 (N_5869,N_3085,N_3682);
nor U5870 (N_5870,N_4271,N_4023);
nand U5871 (N_5871,N_3415,N_3365);
and U5872 (N_5872,N_3057,N_3159);
xor U5873 (N_5873,N_3943,N_3514);
and U5874 (N_5874,N_3854,N_3989);
or U5875 (N_5875,N_3644,N_3538);
and U5876 (N_5876,N_3662,N_3821);
and U5877 (N_5877,N_3529,N_3725);
and U5878 (N_5878,N_4056,N_3780);
or U5879 (N_5879,N_3764,N_3936);
or U5880 (N_5880,N_3491,N_3111);
nor U5881 (N_5881,N_3484,N_4405);
and U5882 (N_5882,N_3848,N_3839);
nor U5883 (N_5883,N_3278,N_4459);
or U5884 (N_5884,N_4197,N_3978);
xor U5885 (N_5885,N_3361,N_3908);
and U5886 (N_5886,N_3856,N_3181);
nand U5887 (N_5887,N_4450,N_3728);
nand U5888 (N_5888,N_3240,N_3089);
nor U5889 (N_5889,N_3057,N_3145);
nand U5890 (N_5890,N_3160,N_3535);
and U5891 (N_5891,N_4029,N_4332);
or U5892 (N_5892,N_4407,N_3420);
nand U5893 (N_5893,N_3972,N_3394);
nand U5894 (N_5894,N_3622,N_4034);
nand U5895 (N_5895,N_4064,N_3235);
nor U5896 (N_5896,N_3327,N_4101);
nor U5897 (N_5897,N_4250,N_4332);
or U5898 (N_5898,N_4161,N_3446);
nor U5899 (N_5899,N_4224,N_4457);
nor U5900 (N_5900,N_4283,N_4125);
nand U5901 (N_5901,N_3198,N_3703);
xnor U5902 (N_5902,N_4443,N_3459);
or U5903 (N_5903,N_3922,N_3042);
xnor U5904 (N_5904,N_3970,N_3542);
xnor U5905 (N_5905,N_3889,N_3304);
and U5906 (N_5906,N_4071,N_4342);
nor U5907 (N_5907,N_4438,N_4359);
or U5908 (N_5908,N_3245,N_4068);
nor U5909 (N_5909,N_3375,N_4086);
or U5910 (N_5910,N_3577,N_3154);
or U5911 (N_5911,N_4373,N_4484);
and U5912 (N_5912,N_4353,N_3434);
xor U5913 (N_5913,N_3914,N_3039);
nor U5914 (N_5914,N_3897,N_3945);
and U5915 (N_5915,N_3936,N_3663);
and U5916 (N_5916,N_3846,N_3993);
nor U5917 (N_5917,N_4308,N_3807);
or U5918 (N_5918,N_4032,N_3352);
nor U5919 (N_5919,N_3104,N_3935);
or U5920 (N_5920,N_4278,N_3893);
nor U5921 (N_5921,N_4418,N_4434);
xor U5922 (N_5922,N_3728,N_3964);
nand U5923 (N_5923,N_3859,N_3897);
nor U5924 (N_5924,N_3734,N_3808);
and U5925 (N_5925,N_4254,N_4215);
nor U5926 (N_5926,N_4303,N_4266);
nand U5927 (N_5927,N_3645,N_3283);
nor U5928 (N_5928,N_3196,N_4348);
nand U5929 (N_5929,N_3480,N_3288);
nand U5930 (N_5930,N_4111,N_3674);
or U5931 (N_5931,N_3309,N_4245);
nand U5932 (N_5932,N_3537,N_3279);
nand U5933 (N_5933,N_3111,N_4099);
nand U5934 (N_5934,N_3914,N_4066);
nor U5935 (N_5935,N_3147,N_4435);
or U5936 (N_5936,N_4093,N_4412);
or U5937 (N_5937,N_4380,N_3799);
and U5938 (N_5938,N_4037,N_4137);
and U5939 (N_5939,N_4049,N_4314);
or U5940 (N_5940,N_3050,N_3068);
nor U5941 (N_5941,N_3141,N_3460);
and U5942 (N_5942,N_3606,N_3285);
or U5943 (N_5943,N_3770,N_3386);
or U5944 (N_5944,N_3219,N_3472);
or U5945 (N_5945,N_3678,N_3035);
nand U5946 (N_5946,N_4289,N_4397);
nand U5947 (N_5947,N_3550,N_3200);
and U5948 (N_5948,N_3448,N_3858);
nor U5949 (N_5949,N_3384,N_4019);
nor U5950 (N_5950,N_3398,N_4329);
nor U5951 (N_5951,N_3710,N_3314);
nor U5952 (N_5952,N_3780,N_4302);
nand U5953 (N_5953,N_3653,N_4301);
nor U5954 (N_5954,N_3603,N_4457);
nand U5955 (N_5955,N_3453,N_4418);
nor U5956 (N_5956,N_3514,N_3875);
nor U5957 (N_5957,N_4285,N_3627);
or U5958 (N_5958,N_4442,N_3021);
or U5959 (N_5959,N_3191,N_3576);
nor U5960 (N_5960,N_4469,N_3072);
and U5961 (N_5961,N_4134,N_3602);
xor U5962 (N_5962,N_3759,N_3271);
nand U5963 (N_5963,N_3786,N_3134);
nand U5964 (N_5964,N_3982,N_4141);
nor U5965 (N_5965,N_3428,N_3440);
and U5966 (N_5966,N_3711,N_3284);
nor U5967 (N_5967,N_4151,N_3774);
xor U5968 (N_5968,N_4072,N_3258);
nand U5969 (N_5969,N_3532,N_4114);
and U5970 (N_5970,N_3417,N_4217);
or U5971 (N_5971,N_3685,N_4127);
nand U5972 (N_5972,N_3688,N_3111);
and U5973 (N_5973,N_4093,N_4298);
nand U5974 (N_5974,N_3359,N_3875);
xor U5975 (N_5975,N_4166,N_3798);
or U5976 (N_5976,N_3755,N_3369);
and U5977 (N_5977,N_4172,N_4175);
nand U5978 (N_5978,N_3139,N_3299);
xor U5979 (N_5979,N_3273,N_3414);
or U5980 (N_5980,N_3571,N_4425);
nor U5981 (N_5981,N_3441,N_4255);
and U5982 (N_5982,N_4308,N_3799);
or U5983 (N_5983,N_3801,N_4052);
and U5984 (N_5984,N_4066,N_3789);
nand U5985 (N_5985,N_3437,N_3831);
nand U5986 (N_5986,N_4315,N_3000);
nand U5987 (N_5987,N_3944,N_4462);
or U5988 (N_5988,N_3853,N_3957);
and U5989 (N_5989,N_4279,N_4330);
nand U5990 (N_5990,N_3448,N_4289);
and U5991 (N_5991,N_4046,N_3779);
or U5992 (N_5992,N_3735,N_3906);
nand U5993 (N_5993,N_3988,N_3306);
and U5994 (N_5994,N_3055,N_3745);
or U5995 (N_5995,N_3652,N_3421);
nand U5996 (N_5996,N_4230,N_4431);
nand U5997 (N_5997,N_4190,N_3963);
nand U5998 (N_5998,N_3691,N_3292);
nor U5999 (N_5999,N_4253,N_3010);
nand U6000 (N_6000,N_5991,N_5453);
or U6001 (N_6001,N_5314,N_5512);
or U6002 (N_6002,N_5874,N_5196);
xor U6003 (N_6003,N_4542,N_5933);
or U6004 (N_6004,N_5842,N_5264);
nand U6005 (N_6005,N_5496,N_5797);
and U6006 (N_6006,N_5862,N_5714);
and U6007 (N_6007,N_4764,N_5455);
nor U6008 (N_6008,N_5403,N_5103);
nor U6009 (N_6009,N_5989,N_4709);
and U6010 (N_6010,N_5972,N_5609);
nor U6011 (N_6011,N_5800,N_5720);
nand U6012 (N_6012,N_5883,N_5508);
nand U6013 (N_6013,N_5821,N_4794);
nor U6014 (N_6014,N_5974,N_4776);
nand U6015 (N_6015,N_5456,N_4703);
nand U6016 (N_6016,N_4511,N_5876);
and U6017 (N_6017,N_5979,N_4697);
or U6018 (N_6018,N_5430,N_5451);
or U6019 (N_6019,N_5546,N_5768);
and U6020 (N_6020,N_5412,N_4926);
and U6021 (N_6021,N_5008,N_5581);
nand U6022 (N_6022,N_4646,N_5481);
nor U6023 (N_6023,N_5914,N_4716);
or U6024 (N_6024,N_5203,N_5676);
nor U6025 (N_6025,N_5149,N_5510);
xor U6026 (N_6026,N_5856,N_5330);
nand U6027 (N_6027,N_4550,N_5003);
nor U6028 (N_6028,N_5640,N_5025);
and U6029 (N_6029,N_5966,N_4955);
nor U6030 (N_6030,N_4717,N_5529);
nor U6031 (N_6031,N_5279,N_4607);
nand U6032 (N_6032,N_4623,N_5897);
and U6033 (N_6033,N_5464,N_5034);
and U6034 (N_6034,N_4500,N_5225);
nor U6035 (N_6035,N_5488,N_5076);
nor U6036 (N_6036,N_5892,N_4959);
or U6037 (N_6037,N_5328,N_5185);
nand U6038 (N_6038,N_4835,N_5202);
or U6039 (N_6039,N_5891,N_4973);
nor U6040 (N_6040,N_5498,N_5490);
and U6041 (N_6041,N_4958,N_4611);
nor U6042 (N_6042,N_5472,N_4521);
and U6043 (N_6043,N_5391,N_4605);
nand U6044 (N_6044,N_5716,N_4830);
nor U6045 (N_6045,N_5290,N_5251);
and U6046 (N_6046,N_5492,N_5411);
nand U6047 (N_6047,N_5593,N_5358);
or U6048 (N_6048,N_5127,N_5918);
nand U6049 (N_6049,N_4633,N_4555);
nand U6050 (N_6050,N_4674,N_4564);
and U6051 (N_6051,N_4723,N_4897);
and U6052 (N_6052,N_5701,N_5383);
nand U6053 (N_6053,N_4933,N_5980);
nor U6054 (N_6054,N_5155,N_5572);
nor U6055 (N_6055,N_5617,N_5793);
and U6056 (N_6056,N_5938,N_4597);
and U6057 (N_6057,N_5882,N_4778);
nor U6058 (N_6058,N_4600,N_4894);
and U6059 (N_6059,N_4781,N_4843);
nor U6060 (N_6060,N_5514,N_4968);
and U6061 (N_6061,N_4601,N_4745);
and U6062 (N_6062,N_5486,N_5469);
and U6063 (N_6063,N_4667,N_4957);
and U6064 (N_6064,N_4532,N_5881);
nand U6065 (N_6065,N_5880,N_4841);
nor U6066 (N_6066,N_5532,N_5098);
and U6067 (N_6067,N_5106,N_5295);
nand U6068 (N_6068,N_5243,N_5211);
nand U6069 (N_6069,N_4617,N_5347);
and U6070 (N_6070,N_4788,N_5585);
nand U6071 (N_6071,N_5135,N_5960);
and U6072 (N_6072,N_5148,N_4922);
or U6073 (N_6073,N_5958,N_5592);
nor U6074 (N_6074,N_5485,N_5725);
and U6075 (N_6075,N_4707,N_4828);
or U6076 (N_6076,N_4834,N_4874);
nor U6077 (N_6077,N_5166,N_4867);
or U6078 (N_6078,N_5582,N_4662);
nand U6079 (N_6079,N_5482,N_4851);
or U6080 (N_6080,N_4577,N_4816);
nand U6081 (N_6081,N_5493,N_4995);
nor U6082 (N_6082,N_5107,N_4685);
nor U6083 (N_6083,N_5915,N_4935);
xor U6084 (N_6084,N_4702,N_5740);
or U6085 (N_6085,N_5712,N_5332);
nand U6086 (N_6086,N_5888,N_5682);
nor U6087 (N_6087,N_5679,N_5401);
or U6088 (N_6088,N_5010,N_4932);
nand U6089 (N_6089,N_5598,N_5305);
or U6090 (N_6090,N_4963,N_5303);
and U6091 (N_6091,N_5755,N_5470);
and U6092 (N_6092,N_4584,N_5925);
xor U6093 (N_6093,N_5045,N_5084);
nand U6094 (N_6094,N_5365,N_5758);
nand U6095 (N_6095,N_5535,N_4883);
xor U6096 (N_6096,N_5519,N_5757);
and U6097 (N_6097,N_5928,N_5537);
nand U6098 (N_6098,N_5431,N_4814);
nor U6099 (N_6099,N_4525,N_5605);
nor U6100 (N_6100,N_5936,N_5904);
nor U6101 (N_6101,N_4836,N_4575);
nor U6102 (N_6102,N_5688,N_5088);
or U6103 (N_6103,N_4630,N_4668);
nand U6104 (N_6104,N_5929,N_4684);
or U6105 (N_6105,N_4665,N_5600);
nand U6106 (N_6106,N_5452,N_4798);
or U6107 (N_6107,N_4724,N_4733);
or U6108 (N_6108,N_5300,N_4947);
nand U6109 (N_6109,N_4711,N_4658);
or U6110 (N_6110,N_4567,N_5380);
or U6111 (N_6111,N_5967,N_5908);
nor U6112 (N_6112,N_5566,N_5041);
and U6113 (N_6113,N_4654,N_5689);
xor U6114 (N_6114,N_5497,N_4990);
and U6115 (N_6115,N_4868,N_5082);
nand U6116 (N_6116,N_4616,N_5371);
or U6117 (N_6117,N_5746,N_5425);
nand U6118 (N_6118,N_4850,N_5143);
and U6119 (N_6119,N_5723,N_5810);
nand U6120 (N_6120,N_5263,N_5559);
nor U6121 (N_6121,N_5217,N_4965);
nand U6122 (N_6122,N_5174,N_4948);
and U6123 (N_6123,N_5931,N_5717);
or U6124 (N_6124,N_4857,N_4978);
nand U6125 (N_6125,N_5941,N_5257);
nor U6126 (N_6126,N_5176,N_5028);
nand U6127 (N_6127,N_5130,N_5551);
or U6128 (N_6128,N_5139,N_5816);
or U6129 (N_6129,N_5618,N_4692);
xnor U6130 (N_6130,N_4679,N_4604);
nand U6131 (N_6131,N_5584,N_4648);
and U6132 (N_6132,N_5164,N_5602);
nand U6133 (N_6133,N_5752,N_4576);
or U6134 (N_6134,N_5942,N_5169);
nor U6135 (N_6135,N_4505,N_5457);
nand U6136 (N_6136,N_5554,N_5361);
or U6137 (N_6137,N_5927,N_4678);
nand U6138 (N_6138,N_4865,N_4939);
and U6139 (N_6139,N_4722,N_5553);
nor U6140 (N_6140,N_4910,N_5696);
or U6141 (N_6141,N_4520,N_5691);
and U6142 (N_6142,N_5400,N_5359);
nand U6143 (N_6143,N_5090,N_5138);
nor U6144 (N_6144,N_4853,N_4903);
nand U6145 (N_6145,N_5051,N_5092);
or U6146 (N_6146,N_5930,N_5655);
and U6147 (N_6147,N_5626,N_5327);
xnor U6148 (N_6148,N_5760,N_5170);
xnor U6149 (N_6149,N_5099,N_4921);
and U6150 (N_6150,N_5561,N_5248);
or U6151 (N_6151,N_5624,N_5053);
nor U6152 (N_6152,N_5483,N_4615);
or U6153 (N_6153,N_5236,N_5031);
or U6154 (N_6154,N_4636,N_5309);
and U6155 (N_6155,N_5595,N_5132);
nor U6156 (N_6156,N_5009,N_5635);
and U6157 (N_6157,N_5230,N_4608);
nor U6158 (N_6158,N_4971,N_5188);
xnor U6159 (N_6159,N_5748,N_4975);
and U6160 (N_6160,N_5987,N_4758);
nor U6161 (N_6161,N_4821,N_5830);
or U6162 (N_6162,N_4770,N_5619);
and U6163 (N_6163,N_5476,N_4522);
nand U6164 (N_6164,N_5794,N_4765);
nor U6165 (N_6165,N_5580,N_5413);
and U6166 (N_6166,N_5069,N_4704);
or U6167 (N_6167,N_5840,N_4647);
nand U6168 (N_6168,N_5956,N_5161);
nor U6169 (N_6169,N_5732,N_5377);
nand U6170 (N_6170,N_5479,N_5474);
and U6171 (N_6171,N_5146,N_4751);
nand U6172 (N_6172,N_4671,N_4889);
or U6173 (N_6173,N_5190,N_4817);
or U6174 (N_6174,N_5843,N_5072);
nor U6175 (N_6175,N_5766,N_4811);
nor U6176 (N_6176,N_5920,N_4873);
nor U6177 (N_6177,N_5407,N_5478);
nor U6178 (N_6178,N_5799,N_5017);
xor U6179 (N_6179,N_5875,N_5737);
nor U6180 (N_6180,N_4730,N_4902);
and U6181 (N_6181,N_5722,N_5978);
or U6182 (N_6182,N_4527,N_4824);
nor U6183 (N_6183,N_5890,N_4536);
nand U6184 (N_6184,N_5256,N_5742);
and U6185 (N_6185,N_5707,N_5286);
nor U6186 (N_6186,N_5750,N_5007);
or U6187 (N_6187,N_5375,N_4944);
nand U6188 (N_6188,N_5633,N_4560);
nor U6189 (N_6189,N_4643,N_4918);
or U6190 (N_6190,N_5321,N_5306);
and U6191 (N_6191,N_5692,N_5563);
or U6192 (N_6192,N_5808,N_5822);
nand U6193 (N_6193,N_5167,N_5871);
nor U6194 (N_6194,N_5477,N_5513);
nand U6195 (N_6195,N_5657,N_5531);
nor U6196 (N_6196,N_4710,N_4559);
nor U6197 (N_6197,N_4988,N_5664);
or U6198 (N_6198,N_5005,N_5675);
nor U6199 (N_6199,N_5181,N_5302);
and U6200 (N_6200,N_5289,N_5694);
nand U6201 (N_6201,N_5448,N_5674);
and U6202 (N_6202,N_5858,N_4856);
nor U6203 (N_6203,N_5705,N_4657);
or U6204 (N_6204,N_4913,N_4732);
or U6205 (N_6205,N_4610,N_5160);
nor U6206 (N_6206,N_4507,N_5686);
nand U6207 (N_6207,N_4984,N_5050);
xnor U6208 (N_6208,N_5061,N_5992);
and U6209 (N_6209,N_5839,N_5643);
or U6210 (N_6210,N_5133,N_4695);
nor U6211 (N_6211,N_4529,N_5636);
nor U6212 (N_6212,N_5437,N_4742);
xor U6213 (N_6213,N_4693,N_5011);
nor U6214 (N_6214,N_5278,N_5199);
nand U6215 (N_6215,N_5975,N_5173);
or U6216 (N_6216,N_4720,N_5648);
or U6217 (N_6217,N_4991,N_5820);
nand U6218 (N_6218,N_5893,N_5128);
and U6219 (N_6219,N_4681,N_5708);
or U6220 (N_6220,N_4721,N_4712);
or U6221 (N_6221,N_4736,N_5790);
nor U6222 (N_6222,N_5733,N_4534);
and U6223 (N_6223,N_4892,N_5193);
and U6224 (N_6224,N_5518,N_5706);
nor U6225 (N_6225,N_5153,N_5734);
xor U6226 (N_6226,N_5670,N_5634);
nand U6227 (N_6227,N_5432,N_5015);
nor U6228 (N_6228,N_5102,N_5877);
nand U6229 (N_6229,N_5204,N_5183);
nor U6230 (N_6230,N_5039,N_5104);
and U6231 (N_6231,N_4649,N_5591);
nor U6232 (N_6232,N_5272,N_5885);
xnor U6233 (N_6233,N_5861,N_5271);
nor U6234 (N_6234,N_5285,N_5063);
nand U6235 (N_6235,N_5525,N_4760);
and U6236 (N_6236,N_5949,N_5604);
and U6237 (N_6237,N_5228,N_4980);
and U6238 (N_6238,N_5982,N_5651);
and U6239 (N_6239,N_4785,N_4791);
nand U6240 (N_6240,N_5724,N_5048);
nor U6241 (N_6241,N_5868,N_5662);
or U6242 (N_6242,N_5433,N_5629);
nor U6243 (N_6243,N_5703,N_4666);
nor U6244 (N_6244,N_5612,N_5276);
and U6245 (N_6245,N_4516,N_4951);
or U6246 (N_6246,N_4734,N_5976);
and U6247 (N_6247,N_5122,N_4741);
xor U6248 (N_6248,N_4718,N_5487);
or U6249 (N_6249,N_5774,N_5838);
nand U6250 (N_6250,N_4727,N_5252);
or U6251 (N_6251,N_5036,N_5847);
nand U6252 (N_6252,N_5350,N_4923);
nor U6253 (N_6253,N_5653,N_4673);
and U6254 (N_6254,N_5564,N_5834);
nand U6255 (N_6255,N_5998,N_5690);
nand U6256 (N_6256,N_4927,N_5959);
xnor U6257 (N_6257,N_4763,N_4936);
nand U6258 (N_6258,N_5113,N_5419);
and U6259 (N_6259,N_5325,N_4793);
or U6260 (N_6260,N_5610,N_5237);
nor U6261 (N_6261,N_5282,N_5587);
or U6262 (N_6262,N_5940,N_4840);
or U6263 (N_6263,N_4848,N_4938);
nor U6264 (N_6264,N_5484,N_5806);
or U6265 (N_6265,N_5515,N_5192);
and U6266 (N_6266,N_5846,N_5783);
nor U6267 (N_6267,N_5089,N_5521);
or U6268 (N_6268,N_4744,N_5895);
nand U6269 (N_6269,N_5913,N_4967);
nor U6270 (N_6270,N_4638,N_4640);
and U6271 (N_6271,N_4925,N_5024);
nand U6272 (N_6272,N_5280,N_5659);
nor U6273 (N_6273,N_5268,N_4854);
xor U6274 (N_6274,N_5394,N_5091);
nand U6275 (N_6275,N_5136,N_5150);
xnor U6276 (N_6276,N_5338,N_5438);
nor U6277 (N_6277,N_5503,N_5771);
nor U6278 (N_6278,N_5466,N_4872);
and U6279 (N_6279,N_4799,N_5825);
nand U6280 (N_6280,N_5500,N_5417);
nand U6281 (N_6281,N_5086,N_4627);
nand U6282 (N_6282,N_5555,N_4642);
or U6283 (N_6283,N_4737,N_5850);
nand U6284 (N_6284,N_5596,N_5579);
nor U6285 (N_6285,N_5832,N_5534);
or U6286 (N_6286,N_5898,N_5265);
nor U6287 (N_6287,N_5067,N_5423);
xnor U6288 (N_6288,N_5544,N_5094);
xor U6289 (N_6289,N_5260,N_5741);
nand U6290 (N_6290,N_5349,N_5985);
nand U6291 (N_6291,N_5126,N_4795);
or U6292 (N_6292,N_4598,N_5056);
nand U6293 (N_6293,N_5058,N_4682);
xor U6294 (N_6294,N_5462,N_5022);
nor U6295 (N_6295,N_4829,N_5189);
and U6296 (N_6296,N_5526,N_5761);
xnor U6297 (N_6297,N_5951,N_4761);
nor U6298 (N_6298,N_4573,N_5953);
or U6299 (N_6299,N_5680,N_5334);
nor U6300 (N_6300,N_4904,N_5569);
or U6301 (N_6301,N_5616,N_5198);
or U6302 (N_6302,N_4878,N_4808);
nor U6303 (N_6303,N_5630,N_4628);
nand U6304 (N_6304,N_5855,N_5753);
nand U6305 (N_6305,N_4837,N_5502);
nor U6306 (N_6306,N_5772,N_4592);
nor U6307 (N_6307,N_5152,N_5886);
nor U6308 (N_6308,N_5678,N_5499);
and U6309 (N_6309,N_4637,N_5731);
nor U6310 (N_6310,N_5578,N_5522);
xor U6311 (N_6311,N_4864,N_4772);
or U6312 (N_6312,N_4691,N_5288);
nor U6313 (N_6313,N_4541,N_5379);
and U6314 (N_6314,N_5550,N_5887);
nor U6315 (N_6315,N_5854,N_4786);
and U6316 (N_6316,N_5267,N_5818);
xnor U6317 (N_6317,N_4538,N_5191);
xnor U6318 (N_6318,N_4566,N_5646);
nor U6319 (N_6319,N_4509,N_5787);
or U6320 (N_6320,N_5351,N_5157);
and U6321 (N_6321,N_4981,N_5932);
or U6322 (N_6322,N_5934,N_5418);
or U6323 (N_6323,N_5789,N_5239);
and U6324 (N_6324,N_5187,N_5410);
and U6325 (N_6325,N_4940,N_4782);
or U6326 (N_6326,N_4999,N_4546);
xnor U6327 (N_6327,N_4802,N_5661);
and U6328 (N_6328,N_5156,N_5607);
and U6329 (N_6329,N_5516,N_4634);
nor U6330 (N_6330,N_4590,N_5627);
nor U6331 (N_6331,N_5356,N_4937);
and U6332 (N_6332,N_5815,N_5027);
nand U6333 (N_6333,N_5971,N_5826);
or U6334 (N_6334,N_5226,N_4934);
nor U6335 (N_6335,N_5620,N_5125);
nand U6336 (N_6336,N_5172,N_5819);
nor U6337 (N_6337,N_4888,N_5804);
and U6338 (N_6338,N_5200,N_4930);
nor U6339 (N_6339,N_5909,N_5223);
nor U6340 (N_6340,N_4982,N_5345);
xnor U6341 (N_6341,N_5320,N_4747);
nand U6342 (N_6342,N_4757,N_4832);
nand U6343 (N_6343,N_4537,N_5450);
xnor U6344 (N_6344,N_5853,N_4557);
or U6345 (N_6345,N_5786,N_5404);
nand U6346 (N_6346,N_4543,N_5700);
xor U6347 (N_6347,N_4900,N_4645);
or U6348 (N_6348,N_5283,N_5037);
or U6349 (N_6349,N_5044,N_5744);
nand U6350 (N_6350,N_4533,N_4725);
or U6351 (N_6351,N_4920,N_4881);
nand U6352 (N_6352,N_5023,N_4544);
and U6353 (N_6353,N_5475,N_5154);
nor U6354 (N_6354,N_5736,N_5219);
or U6355 (N_6355,N_4952,N_5129);
nand U6356 (N_6356,N_5970,N_5611);
nor U6357 (N_6357,N_5355,N_5020);
nor U6358 (N_6358,N_5939,N_5363);
nand U6359 (N_6359,N_5628,N_5182);
and U6360 (N_6360,N_5296,N_5745);
or U6361 (N_6361,N_5030,N_5241);
nand U6362 (N_6362,N_4582,N_5709);
nor U6363 (N_6363,N_5637,N_4804);
nand U6364 (N_6364,N_5052,N_5147);
and U6365 (N_6365,N_5727,N_5726);
nor U6366 (N_6366,N_5310,N_4513);
and U6367 (N_6367,N_5428,N_4596);
or U6368 (N_6368,N_5112,N_5335);
or U6369 (N_6369,N_5762,N_5242);
nor U6370 (N_6370,N_5207,N_5507);
and U6371 (N_6371,N_4964,N_5851);
nor U6372 (N_6372,N_5767,N_4983);
xnor U6373 (N_6373,N_4746,N_5719);
xor U6374 (N_6374,N_4552,N_5536);
nand U6375 (N_6375,N_4539,N_5070);
and U6376 (N_6376,N_5054,N_4606);
or U6377 (N_6377,N_4972,N_5669);
and U6378 (N_6378,N_5171,N_5543);
and U6379 (N_6379,N_5001,N_5270);
nand U6380 (N_6380,N_5458,N_4801);
or U6381 (N_6381,N_4992,N_5728);
or U6382 (N_6382,N_5258,N_5828);
nor U6383 (N_6383,N_5159,N_5867);
xor U6384 (N_6384,N_5197,N_4528);
nor U6385 (N_6385,N_5965,N_5119);
nor U6386 (N_6386,N_5623,N_5575);
or U6387 (N_6387,N_4631,N_5685);
and U6388 (N_6388,N_5527,N_5683);
nand U6389 (N_6389,N_5552,N_4869);
xor U6390 (N_6390,N_4663,N_5573);
nor U6391 (N_6391,N_4563,N_5990);
or U6392 (N_6392,N_5903,N_5331);
nor U6393 (N_6393,N_4916,N_4943);
or U6394 (N_6394,N_5057,N_4842);
nor U6395 (N_6395,N_5528,N_5866);
and U6396 (N_6396,N_5699,N_5947);
and U6397 (N_6397,N_4813,N_5195);
nor U6398 (N_6398,N_5955,N_5567);
nand U6399 (N_6399,N_5151,N_5381);
or U6400 (N_6400,N_5046,N_4797);
or U6401 (N_6401,N_5344,N_5795);
nand U6402 (N_6402,N_5354,N_5163);
or U6403 (N_6403,N_5333,N_5221);
and U6404 (N_6404,N_5074,N_4735);
and U6405 (N_6405,N_4531,N_4558);
or U6406 (N_6406,N_4928,N_5548);
nand U6407 (N_6407,N_5583,N_5827);
nor U6408 (N_6408,N_4508,N_5281);
and U6409 (N_6409,N_5775,N_5963);
nand U6410 (N_6410,N_4635,N_4510);
or U6411 (N_6411,N_5565,N_5779);
or U6412 (N_6412,N_5390,N_4807);
and U6413 (N_6413,N_5663,N_5341);
or U6414 (N_6414,N_4659,N_5711);
nor U6415 (N_6415,N_5879,N_5625);
and U6416 (N_6416,N_5446,N_5601);
and U6417 (N_6417,N_5704,N_4749);
nor U6418 (N_6418,N_5441,N_5118);
nor U6419 (N_6419,N_5545,N_4986);
nor U6420 (N_6420,N_5549,N_4979);
nor U6421 (N_6421,N_4549,N_5899);
nand U6422 (N_6422,N_4554,N_5117);
or U6423 (N_6423,N_4858,N_4783);
and U6424 (N_6424,N_5615,N_5336);
xor U6425 (N_6425,N_5777,N_5317);
or U6426 (N_6426,N_5710,N_4766);
and U6427 (N_6427,N_5184,N_5426);
and U6428 (N_6428,N_4846,N_4650);
nor U6429 (N_6429,N_5468,N_5429);
nand U6430 (N_6430,N_5560,N_5644);
or U6431 (N_6431,N_5638,N_5801);
nor U6432 (N_6432,N_4890,N_4547);
nor U6433 (N_6433,N_4880,N_5049);
and U6434 (N_6434,N_5393,N_4886);
and U6435 (N_6435,N_4803,N_4595);
and U6436 (N_6436,N_5220,N_5062);
or U6437 (N_6437,N_5218,N_5864);
nor U6438 (N_6438,N_5353,N_5729);
and U6439 (N_6439,N_5250,N_5209);
or U6440 (N_6440,N_5443,N_5673);
xor U6441 (N_6441,N_5238,N_5162);
nor U6442 (N_6442,N_5253,N_4523);
nand U6443 (N_6443,N_5323,N_5409);
nand U6444 (N_6444,N_5594,N_5340);
and U6445 (N_6445,N_5080,N_5542);
or U6446 (N_6446,N_5145,N_5981);
and U6447 (N_6447,N_5570,N_5603);
nand U6448 (N_6448,N_5274,N_5889);
xor U6449 (N_6449,N_4676,N_4587);
nand U6450 (N_6450,N_4540,N_5420);
nor U6451 (N_6451,N_4911,N_4954);
or U6452 (N_6452,N_4530,N_4977);
nand U6453 (N_6453,N_4572,N_5459);
nor U6454 (N_6454,N_5695,N_5684);
and U6455 (N_6455,N_5697,N_5465);
or U6456 (N_6456,N_5568,N_5988);
nor U6457 (N_6457,N_5713,N_4729);
xor U6458 (N_6458,N_5614,N_5780);
and U6459 (N_6459,N_5399,N_5964);
and U6460 (N_6460,N_5240,N_4652);
or U6461 (N_6461,N_5042,N_5158);
xor U6462 (N_6462,N_5342,N_5389);
nor U6463 (N_6463,N_5852,N_5759);
nand U6464 (N_6464,N_5460,N_4579);
nor U6465 (N_6465,N_5756,N_5259);
nand U6466 (N_6466,N_4743,N_4519);
or U6467 (N_6467,N_5116,N_5357);
and U6468 (N_6468,N_4621,N_4775);
nand U6469 (N_6469,N_4784,N_5523);
or U6470 (N_6470,N_4626,N_5739);
or U6471 (N_6471,N_5060,N_4792);
nor U6472 (N_6472,N_4614,N_4998);
nand U6473 (N_6473,N_5805,N_4893);
nor U6474 (N_6474,N_5366,N_5026);
xor U6475 (N_6475,N_5702,N_5785);
nand U6476 (N_6476,N_5231,N_5922);
or U6477 (N_6477,N_5299,N_4655);
nor U6478 (N_6478,N_4960,N_4518);
and U6479 (N_6479,N_5943,N_5859);
nand U6480 (N_6480,N_4683,N_5422);
nand U6481 (N_6481,N_5919,N_5807);
nand U6482 (N_6482,N_5654,N_5995);
and U6483 (N_6483,N_5445,N_4501);
nand U6484 (N_6484,N_5002,N_5304);
and U6485 (N_6485,N_5994,N_5083);
or U6486 (N_6486,N_5235,N_4641);
nor U6487 (N_6487,N_4812,N_5473);
or U6488 (N_6488,N_5520,N_4844);
nand U6489 (N_6489,N_4594,N_5574);
nand U6490 (N_6490,N_4545,N_4517);
nor U6491 (N_6491,N_4987,N_5408);
nand U6492 (N_6492,N_5370,N_5539);
nand U6493 (N_6493,N_4871,N_5923);
and U6494 (N_6494,N_5926,N_4580);
nand U6495 (N_6495,N_5910,N_4612);
and U6496 (N_6496,N_5079,N_4970);
and U6497 (N_6497,N_5016,N_5384);
nand U6498 (N_6498,N_5912,N_4561);
nor U6499 (N_6499,N_5811,N_5809);
nand U6500 (N_6500,N_5447,N_5033);
and U6501 (N_6501,N_4669,N_5547);
nor U6502 (N_6502,N_5364,N_4512);
nand U6503 (N_6503,N_5900,N_5687);
and U6504 (N_6504,N_5261,N_4653);
or U6505 (N_6505,N_5878,N_4591);
nand U6506 (N_6506,N_4706,N_5266);
nand U6507 (N_6507,N_5095,N_5019);
nor U6508 (N_6508,N_5763,N_4941);
nand U6509 (N_6509,N_5298,N_4570);
and U6510 (N_6510,N_4670,N_5905);
xnor U6511 (N_6511,N_5368,N_5764);
nand U6512 (N_6512,N_5667,N_5140);
or U6513 (N_6513,N_5329,N_4514);
or U6514 (N_6514,N_5018,N_4578);
nor U6515 (N_6515,N_5463,N_5081);
nor U6516 (N_6516,N_4588,N_5071);
nand U6517 (N_6517,N_5059,N_4779);
and U6518 (N_6518,N_5836,N_5319);
and U6519 (N_6519,N_5421,N_4924);
nand U6520 (N_6520,N_5123,N_5954);
or U6521 (N_6521,N_5109,N_4661);
nand U6522 (N_6522,N_5124,N_5316);
or U6523 (N_6523,N_4680,N_5093);
nor U6524 (N_6524,N_4855,N_4796);
nor U6525 (N_6525,N_5747,N_5901);
or U6526 (N_6526,N_4603,N_5222);
nor U6527 (N_6527,N_4849,N_5427);
and U6528 (N_6528,N_4585,N_5829);
and U6529 (N_6529,N_5206,N_5844);
xnor U6530 (N_6530,N_4672,N_4901);
or U6531 (N_6531,N_4805,N_5315);
and U6532 (N_6532,N_4863,N_4847);
nor U6533 (N_6533,N_4879,N_4884);
or U6534 (N_6534,N_4862,N_5986);
or U6535 (N_6535,N_4945,N_5823);
xnor U6536 (N_6536,N_5273,N_5754);
or U6537 (N_6537,N_5778,N_5194);
nand U6538 (N_6538,N_5773,N_5935);
nand U6539 (N_6539,N_5577,N_4950);
nor U6540 (N_6540,N_5414,N_4571);
nand U6541 (N_6541,N_4825,N_5835);
nor U6542 (N_6542,N_5374,N_5533);
or U6543 (N_6543,N_5012,N_5751);
nor U6544 (N_6544,N_5229,N_5115);
and U6545 (N_6545,N_5632,N_4726);
or U6546 (N_6546,N_4620,N_5945);
or U6547 (N_6547,N_5352,N_5906);
or U6548 (N_6548,N_5255,N_5969);
xor U6549 (N_6549,N_5291,N_5948);
and U6550 (N_6550,N_5517,N_4997);
or U6551 (N_6551,N_5491,N_4750);
and U6552 (N_6552,N_4899,N_5562);
or U6553 (N_6553,N_4506,N_4905);
nor U6554 (N_6554,N_5111,N_5035);
and U6555 (N_6555,N_5666,N_4574);
or U6556 (N_6556,N_5137,N_5066);
nand U6557 (N_6557,N_5524,N_5467);
nand U6558 (N_6558,N_5902,N_4502);
nand U6559 (N_6559,N_5444,N_4713);
nand U6560 (N_6560,N_4974,N_5781);
nand U6561 (N_6561,N_5262,N_5275);
or U6562 (N_6562,N_5402,N_4976);
or U6563 (N_6563,N_4827,N_5378);
nor U6564 (N_6564,N_5180,N_5884);
nand U6565 (N_6565,N_4861,N_5681);
or U6566 (N_6566,N_4688,N_5658);
nor U6567 (N_6567,N_4762,N_5131);
and U6568 (N_6568,N_5973,N_5308);
or U6569 (N_6569,N_5110,N_5907);
or U6570 (N_6570,N_4565,N_4946);
or U6571 (N_6571,N_4870,N_5896);
and U6572 (N_6572,N_4551,N_5813);
xnor U6573 (N_6573,N_4553,N_5436);
or U6574 (N_6574,N_5064,N_5134);
or U6575 (N_6575,N_5397,N_5645);
nand U6576 (N_6576,N_5435,N_5269);
nor U6577 (N_6577,N_4524,N_4852);
nor U6578 (N_6578,N_4752,N_4819);
xor U6579 (N_6579,N_4929,N_5065);
nand U6580 (N_6580,N_5511,N_4714);
nand U6581 (N_6581,N_5178,N_5246);
nand U6582 (N_6582,N_5944,N_5738);
and U6583 (N_6583,N_5043,N_4877);
nand U6584 (N_6584,N_5997,N_4823);
nor U6585 (N_6585,N_5208,N_4664);
nand U6586 (N_6586,N_4891,N_5590);
or U6587 (N_6587,N_5597,N_4767);
nand U6588 (N_6588,N_5557,N_4906);
nand U6589 (N_6589,N_4860,N_4756);
and U6590 (N_6590,N_4622,N_5294);
nand U6591 (N_6591,N_4694,N_5824);
nor U6592 (N_6592,N_5040,N_5769);
nand U6593 (N_6593,N_5946,N_5586);
or U6594 (N_6594,N_5073,N_5872);
and U6595 (N_6595,N_5077,N_4810);
nor U6596 (N_6596,N_4609,N_5216);
nand U6597 (N_6597,N_5372,N_4822);
xnor U6598 (N_6598,N_5993,N_4568);
and U6599 (N_6599,N_5911,N_4993);
nand U6600 (N_6600,N_4583,N_5100);
and U6601 (N_6601,N_4768,N_5916);
nand U6602 (N_6602,N_4740,N_4701);
nand U6603 (N_6603,N_4787,N_4777);
nand U6604 (N_6604,N_4866,N_4618);
nand U6605 (N_6605,N_5952,N_5849);
or U6606 (N_6606,N_5589,N_4696);
and U6607 (N_6607,N_5504,N_5087);
or U6608 (N_6608,N_5957,N_4629);
nor U6609 (N_6609,N_5075,N_4826);
and U6610 (N_6610,N_5141,N_5245);
nor U6611 (N_6611,N_5405,N_5622);
nor U6612 (N_6612,N_5765,N_4908);
or U6613 (N_6613,N_5501,N_5540);
nand U6614 (N_6614,N_5006,N_4586);
and U6615 (N_6615,N_4833,N_5313);
xor U6616 (N_6616,N_5114,N_4912);
xnor U6617 (N_6617,N_4731,N_5870);
nor U6618 (N_6618,N_5984,N_5977);
xor U6619 (N_6619,N_5494,N_5406);
and U6620 (N_6620,N_5398,N_4660);
nor U6621 (N_6621,N_4914,N_5677);
nor U6622 (N_6622,N_4593,N_5671);
nand U6623 (N_6623,N_4896,N_5311);
xnor U6624 (N_6624,N_5788,N_4898);
nor U6625 (N_6625,N_5047,N_5287);
nand U6626 (N_6626,N_4526,N_5385);
and U6627 (N_6627,N_5665,N_5078);
nor U6628 (N_6628,N_5085,N_4942);
nand U6629 (N_6629,N_5186,N_5014);
and U6630 (N_6630,N_4675,N_4515);
or U6631 (N_6631,N_5224,N_5348);
or U6632 (N_6632,N_4953,N_5312);
nand U6633 (N_6633,N_5558,N_5029);
and U6634 (N_6634,N_5606,N_5917);
xnor U6635 (N_6635,N_4773,N_5434);
xor U6636 (N_6636,N_5210,N_5776);
nand U6637 (N_6637,N_4589,N_5021);
nand U6638 (N_6638,N_5440,N_4624);
nor U6639 (N_6639,N_5297,N_4705);
nand U6640 (N_6640,N_5845,N_4800);
or U6641 (N_6641,N_5326,N_5831);
nor U6642 (N_6642,N_5770,N_5869);
xnor U6643 (N_6643,N_5004,N_5292);
xnor U6644 (N_6644,N_4774,N_5538);
nand U6645 (N_6645,N_5343,N_5232);
or U6646 (N_6646,N_5505,N_4686);
nor U6647 (N_6647,N_5865,N_5791);
xnor U6648 (N_6648,N_5608,N_4989);
nand U6649 (N_6649,N_5227,N_5307);
xor U6650 (N_6650,N_5803,N_4548);
nand U6651 (N_6651,N_5439,N_5937);
nand U6652 (N_6652,N_4882,N_5096);
nand U6653 (N_6653,N_5812,N_5376);
xnor U6654 (N_6654,N_4728,N_4845);
nand U6655 (N_6655,N_4949,N_5735);
and U6656 (N_6656,N_5120,N_5599);
nor U6657 (N_6657,N_4917,N_5894);
nand U6658 (N_6658,N_5848,N_5798);
or U6659 (N_6659,N_5387,N_4699);
nor U6660 (N_6660,N_5863,N_5647);
and U6661 (N_6661,N_5175,N_5013);
nor U6662 (N_6662,N_4820,N_5841);
nor U6663 (N_6663,N_4969,N_4931);
and U6664 (N_6664,N_5244,N_5718);
nand U6665 (N_6665,N_5424,N_4994);
nand U6666 (N_6666,N_5924,N_5715);
nand U6667 (N_6667,N_4907,N_5214);
xor U6668 (N_6668,N_5382,N_4831);
nand U6669 (N_6669,N_5293,N_5471);
or U6670 (N_6670,N_5212,N_5416);
and U6671 (N_6671,N_5983,N_5032);
and U6672 (N_6672,N_4748,N_5301);
nand U6673 (N_6673,N_5495,N_4644);
or U6674 (N_6674,N_5461,N_4677);
nand U6675 (N_6675,N_4895,N_4619);
xor U6676 (N_6676,N_5068,N_5621);
xor U6677 (N_6677,N_5000,N_5950);
xnor U6678 (N_6678,N_4504,N_4719);
or U6679 (N_6679,N_4738,N_4687);
nor U6680 (N_6680,N_5177,N_5873);
nor U6681 (N_6681,N_5055,N_4639);
nor U6682 (N_6682,N_5360,N_5668);
nor U6683 (N_6683,N_4966,N_5247);
nand U6684 (N_6684,N_4789,N_5962);
xnor U6685 (N_6685,N_5833,N_4632);
and U6686 (N_6686,N_4599,N_5784);
nand U6687 (N_6687,N_5318,N_5506);
xor U6688 (N_6688,N_4556,N_4715);
or U6689 (N_6689,N_4780,N_5641);
or U6690 (N_6690,N_4700,N_5346);
nor U6691 (N_6691,N_5165,N_5489);
nor U6692 (N_6692,N_5392,N_4859);
nand U6693 (N_6693,N_4753,N_5693);
and U6694 (N_6694,N_5038,N_4885);
and U6695 (N_6695,N_5205,N_5660);
and U6696 (N_6696,N_5254,N_4656);
and U6697 (N_6697,N_5215,N_5571);
or U6698 (N_6698,N_5362,N_5556);
nor U6699 (N_6699,N_4790,N_5108);
nor U6700 (N_6700,N_5802,N_5588);
and U6701 (N_6701,N_5277,N_5249);
or U6702 (N_6702,N_4806,N_4562);
nor U6703 (N_6703,N_5576,N_4915);
and U6704 (N_6704,N_4581,N_4689);
xor U6705 (N_6705,N_5698,N_5968);
nor U6706 (N_6706,N_5442,N_5837);
nand U6707 (N_6707,N_4919,N_5796);
or U6708 (N_6708,N_5179,N_5792);
or U6709 (N_6709,N_5814,N_5168);
xnor U6710 (N_6710,N_5650,N_5649);
or U6711 (N_6711,N_4818,N_4739);
nor U6712 (N_6712,N_5337,N_5782);
or U6713 (N_6713,N_4602,N_5743);
and U6714 (N_6714,N_5921,N_5101);
or U6715 (N_6715,N_4535,N_5652);
nor U6716 (N_6716,N_5388,N_5730);
nand U6717 (N_6717,N_5656,N_4961);
nand U6718 (N_6718,N_4690,N_4876);
and U6719 (N_6719,N_5386,N_5857);
or U6720 (N_6720,N_4962,N_5631);
nor U6721 (N_6721,N_5144,N_5322);
or U6722 (N_6722,N_5234,N_5449);
nor U6723 (N_6723,N_4956,N_5639);
xor U6724 (N_6724,N_5415,N_5817);
nor U6725 (N_6725,N_5373,N_4909);
nor U6726 (N_6726,N_5996,N_5860);
nor U6727 (N_6727,N_5284,N_5541);
nor U6728 (N_6728,N_5749,N_4613);
and U6729 (N_6729,N_5233,N_5509);
and U6730 (N_6730,N_5369,N_5339);
or U6731 (N_6731,N_4771,N_5367);
nor U6732 (N_6732,N_4996,N_5480);
nor U6733 (N_6733,N_5105,N_5213);
and U6734 (N_6734,N_4769,N_5142);
nor U6735 (N_6735,N_5613,N_4815);
nand U6736 (N_6736,N_4887,N_4809);
and U6737 (N_6737,N_5201,N_5121);
and U6738 (N_6738,N_4754,N_5672);
nand U6739 (N_6739,N_4698,N_5530);
or U6740 (N_6740,N_4503,N_4985);
and U6741 (N_6741,N_4875,N_5396);
xor U6742 (N_6742,N_4838,N_5324);
and U6743 (N_6743,N_4625,N_5097);
xnor U6744 (N_6744,N_5454,N_4759);
nor U6745 (N_6745,N_5961,N_5395);
and U6746 (N_6746,N_4651,N_4839);
and U6747 (N_6747,N_4755,N_5999);
nand U6748 (N_6748,N_5642,N_5721);
nor U6749 (N_6749,N_4708,N_4569);
or U6750 (N_6750,N_4555,N_5930);
xnor U6751 (N_6751,N_5661,N_5642);
nand U6752 (N_6752,N_5740,N_5745);
and U6753 (N_6753,N_5728,N_4889);
nand U6754 (N_6754,N_5011,N_5672);
nand U6755 (N_6755,N_5634,N_4971);
nand U6756 (N_6756,N_5554,N_4514);
xor U6757 (N_6757,N_5668,N_5818);
nor U6758 (N_6758,N_4630,N_5223);
nand U6759 (N_6759,N_5138,N_5685);
or U6760 (N_6760,N_5853,N_5950);
nor U6761 (N_6761,N_4739,N_5328);
nor U6762 (N_6762,N_5876,N_5430);
or U6763 (N_6763,N_4856,N_5293);
and U6764 (N_6764,N_5829,N_4881);
and U6765 (N_6765,N_5679,N_4709);
and U6766 (N_6766,N_4640,N_5005);
and U6767 (N_6767,N_4531,N_5264);
and U6768 (N_6768,N_4523,N_5275);
nand U6769 (N_6769,N_5350,N_5272);
and U6770 (N_6770,N_5452,N_5530);
xor U6771 (N_6771,N_5972,N_5152);
or U6772 (N_6772,N_5644,N_5672);
nand U6773 (N_6773,N_4694,N_5634);
and U6774 (N_6774,N_5734,N_5816);
xnor U6775 (N_6775,N_5767,N_5505);
nor U6776 (N_6776,N_4532,N_4557);
or U6777 (N_6777,N_5022,N_5972);
nor U6778 (N_6778,N_5298,N_5699);
nor U6779 (N_6779,N_4527,N_5468);
nand U6780 (N_6780,N_5479,N_5575);
nor U6781 (N_6781,N_5598,N_4943);
nand U6782 (N_6782,N_4825,N_5958);
nor U6783 (N_6783,N_5531,N_4650);
nor U6784 (N_6784,N_5586,N_5449);
nor U6785 (N_6785,N_5857,N_5902);
nor U6786 (N_6786,N_5983,N_5456);
nand U6787 (N_6787,N_5764,N_4701);
and U6788 (N_6788,N_5382,N_5910);
and U6789 (N_6789,N_4575,N_4609);
nand U6790 (N_6790,N_5512,N_5666);
or U6791 (N_6791,N_5174,N_4704);
or U6792 (N_6792,N_5232,N_5642);
nand U6793 (N_6793,N_5178,N_5271);
nor U6794 (N_6794,N_5490,N_5380);
nand U6795 (N_6795,N_5140,N_5289);
or U6796 (N_6796,N_4523,N_5805);
nor U6797 (N_6797,N_4811,N_5093);
nand U6798 (N_6798,N_5920,N_5810);
nand U6799 (N_6799,N_5878,N_5422);
nor U6800 (N_6800,N_5796,N_5337);
xor U6801 (N_6801,N_4758,N_5887);
and U6802 (N_6802,N_5129,N_4512);
nor U6803 (N_6803,N_5842,N_5494);
nand U6804 (N_6804,N_5735,N_5415);
nand U6805 (N_6805,N_4726,N_5176);
and U6806 (N_6806,N_5470,N_5413);
xor U6807 (N_6807,N_5799,N_4814);
nand U6808 (N_6808,N_4648,N_5555);
xnor U6809 (N_6809,N_5374,N_5065);
nor U6810 (N_6810,N_5505,N_5330);
and U6811 (N_6811,N_4625,N_5109);
nor U6812 (N_6812,N_5030,N_5364);
nor U6813 (N_6813,N_4553,N_5449);
nor U6814 (N_6814,N_5224,N_5701);
and U6815 (N_6815,N_5352,N_5582);
and U6816 (N_6816,N_4620,N_5781);
xnor U6817 (N_6817,N_4931,N_5007);
and U6818 (N_6818,N_4973,N_5398);
and U6819 (N_6819,N_4615,N_5589);
or U6820 (N_6820,N_4994,N_4859);
and U6821 (N_6821,N_5860,N_5567);
or U6822 (N_6822,N_4579,N_5185);
or U6823 (N_6823,N_5050,N_5039);
and U6824 (N_6824,N_5633,N_5692);
nand U6825 (N_6825,N_5801,N_5004);
nor U6826 (N_6826,N_4704,N_4689);
nor U6827 (N_6827,N_4947,N_4844);
xor U6828 (N_6828,N_5403,N_4612);
or U6829 (N_6829,N_5150,N_5138);
nand U6830 (N_6830,N_5313,N_4883);
nand U6831 (N_6831,N_5113,N_5405);
and U6832 (N_6832,N_4921,N_4570);
nor U6833 (N_6833,N_5195,N_5115);
or U6834 (N_6834,N_4526,N_4537);
nor U6835 (N_6835,N_5829,N_5315);
nor U6836 (N_6836,N_5225,N_5036);
nand U6837 (N_6837,N_5365,N_5459);
nand U6838 (N_6838,N_5577,N_5821);
nand U6839 (N_6839,N_5082,N_4876);
and U6840 (N_6840,N_5665,N_5728);
nand U6841 (N_6841,N_5477,N_5050);
nand U6842 (N_6842,N_5375,N_4957);
or U6843 (N_6843,N_5530,N_5756);
or U6844 (N_6844,N_5192,N_4947);
and U6845 (N_6845,N_5511,N_5262);
or U6846 (N_6846,N_5761,N_5599);
or U6847 (N_6847,N_5988,N_5453);
nand U6848 (N_6848,N_4597,N_5175);
xnor U6849 (N_6849,N_4713,N_5803);
and U6850 (N_6850,N_5604,N_5628);
and U6851 (N_6851,N_5793,N_5194);
and U6852 (N_6852,N_5118,N_5771);
or U6853 (N_6853,N_5793,N_5756);
and U6854 (N_6854,N_4585,N_5258);
nand U6855 (N_6855,N_5572,N_5530);
xnor U6856 (N_6856,N_5884,N_4707);
or U6857 (N_6857,N_5484,N_4955);
nor U6858 (N_6858,N_5574,N_5084);
and U6859 (N_6859,N_5500,N_5073);
nor U6860 (N_6860,N_5121,N_5955);
and U6861 (N_6861,N_4803,N_5897);
and U6862 (N_6862,N_5560,N_5410);
xor U6863 (N_6863,N_5506,N_5134);
nor U6864 (N_6864,N_5911,N_5896);
or U6865 (N_6865,N_4547,N_5009);
nor U6866 (N_6866,N_5689,N_5162);
xnor U6867 (N_6867,N_4990,N_5390);
nand U6868 (N_6868,N_4791,N_4831);
and U6869 (N_6869,N_5242,N_4736);
and U6870 (N_6870,N_4823,N_5400);
or U6871 (N_6871,N_5681,N_5556);
xor U6872 (N_6872,N_5081,N_5114);
and U6873 (N_6873,N_5897,N_5204);
nand U6874 (N_6874,N_4592,N_4685);
xnor U6875 (N_6875,N_4950,N_4768);
nor U6876 (N_6876,N_5087,N_5103);
nand U6877 (N_6877,N_5659,N_5640);
or U6878 (N_6878,N_5958,N_5556);
or U6879 (N_6879,N_4865,N_5277);
and U6880 (N_6880,N_5508,N_5444);
nand U6881 (N_6881,N_5216,N_4571);
nor U6882 (N_6882,N_5143,N_5653);
or U6883 (N_6883,N_4969,N_5804);
or U6884 (N_6884,N_5939,N_4828);
nor U6885 (N_6885,N_5879,N_4959);
and U6886 (N_6886,N_5826,N_4992);
and U6887 (N_6887,N_5956,N_5504);
and U6888 (N_6888,N_4544,N_5938);
or U6889 (N_6889,N_5634,N_4659);
or U6890 (N_6890,N_4719,N_4886);
and U6891 (N_6891,N_5666,N_4681);
or U6892 (N_6892,N_5308,N_5835);
nor U6893 (N_6893,N_5145,N_4518);
nand U6894 (N_6894,N_5149,N_5208);
nor U6895 (N_6895,N_5607,N_5966);
nor U6896 (N_6896,N_5887,N_5042);
nor U6897 (N_6897,N_4650,N_5980);
or U6898 (N_6898,N_4870,N_5461);
or U6899 (N_6899,N_4672,N_5053);
nor U6900 (N_6900,N_5566,N_5157);
xnor U6901 (N_6901,N_5930,N_4722);
nor U6902 (N_6902,N_4828,N_5122);
nor U6903 (N_6903,N_4955,N_4681);
nor U6904 (N_6904,N_4876,N_5579);
and U6905 (N_6905,N_5914,N_5922);
or U6906 (N_6906,N_4694,N_4927);
and U6907 (N_6907,N_5794,N_4522);
nand U6908 (N_6908,N_5084,N_5800);
or U6909 (N_6909,N_4918,N_4553);
and U6910 (N_6910,N_5687,N_5773);
nand U6911 (N_6911,N_4563,N_5352);
nor U6912 (N_6912,N_5150,N_4924);
nand U6913 (N_6913,N_4923,N_5436);
nand U6914 (N_6914,N_5853,N_5793);
and U6915 (N_6915,N_5600,N_4677);
nor U6916 (N_6916,N_4630,N_5347);
nand U6917 (N_6917,N_4638,N_5552);
nor U6918 (N_6918,N_5917,N_5411);
nand U6919 (N_6919,N_5152,N_5368);
xor U6920 (N_6920,N_5259,N_5312);
and U6921 (N_6921,N_5056,N_4976);
and U6922 (N_6922,N_5497,N_5440);
or U6923 (N_6923,N_4947,N_4746);
nor U6924 (N_6924,N_5098,N_5026);
and U6925 (N_6925,N_5322,N_5030);
or U6926 (N_6926,N_5378,N_5628);
and U6927 (N_6927,N_5200,N_4641);
nor U6928 (N_6928,N_5548,N_5706);
nor U6929 (N_6929,N_4772,N_5095);
and U6930 (N_6930,N_5990,N_5379);
or U6931 (N_6931,N_5084,N_5691);
and U6932 (N_6932,N_4828,N_4895);
and U6933 (N_6933,N_5947,N_5036);
nand U6934 (N_6934,N_5436,N_5847);
or U6935 (N_6935,N_5294,N_5158);
nand U6936 (N_6936,N_5107,N_5301);
or U6937 (N_6937,N_5762,N_5897);
nor U6938 (N_6938,N_5184,N_5361);
nor U6939 (N_6939,N_5416,N_5052);
xor U6940 (N_6940,N_5026,N_5544);
nor U6941 (N_6941,N_4815,N_4550);
nand U6942 (N_6942,N_5964,N_5114);
or U6943 (N_6943,N_5030,N_5904);
nor U6944 (N_6944,N_5997,N_5345);
and U6945 (N_6945,N_5747,N_5912);
and U6946 (N_6946,N_5425,N_4988);
or U6947 (N_6947,N_5836,N_4685);
and U6948 (N_6948,N_5972,N_5675);
xnor U6949 (N_6949,N_5726,N_5788);
nand U6950 (N_6950,N_5141,N_4625);
or U6951 (N_6951,N_5830,N_5483);
and U6952 (N_6952,N_4823,N_5597);
nor U6953 (N_6953,N_5439,N_5998);
nand U6954 (N_6954,N_4830,N_5898);
or U6955 (N_6955,N_5502,N_4577);
or U6956 (N_6956,N_4924,N_4994);
or U6957 (N_6957,N_4712,N_5282);
xor U6958 (N_6958,N_4947,N_5827);
nand U6959 (N_6959,N_4516,N_5815);
or U6960 (N_6960,N_5612,N_5977);
nand U6961 (N_6961,N_4942,N_5542);
and U6962 (N_6962,N_5511,N_4822);
nand U6963 (N_6963,N_5348,N_4947);
or U6964 (N_6964,N_5157,N_4616);
or U6965 (N_6965,N_5737,N_5220);
nor U6966 (N_6966,N_4675,N_4762);
and U6967 (N_6967,N_5516,N_4500);
nor U6968 (N_6968,N_4656,N_5099);
nand U6969 (N_6969,N_5438,N_4749);
or U6970 (N_6970,N_5208,N_4610);
or U6971 (N_6971,N_5632,N_5163);
nand U6972 (N_6972,N_5511,N_4895);
nor U6973 (N_6973,N_5225,N_5481);
and U6974 (N_6974,N_4746,N_5070);
and U6975 (N_6975,N_4669,N_5085);
or U6976 (N_6976,N_5431,N_5112);
nor U6977 (N_6977,N_5292,N_5097);
and U6978 (N_6978,N_4849,N_5137);
nor U6979 (N_6979,N_5015,N_5494);
or U6980 (N_6980,N_5917,N_4994);
nor U6981 (N_6981,N_5783,N_4975);
or U6982 (N_6982,N_5816,N_5780);
nand U6983 (N_6983,N_5245,N_4704);
or U6984 (N_6984,N_4775,N_5824);
nand U6985 (N_6985,N_5197,N_5873);
nor U6986 (N_6986,N_5747,N_5955);
xor U6987 (N_6987,N_4939,N_5549);
xnor U6988 (N_6988,N_4937,N_5180);
and U6989 (N_6989,N_5780,N_5793);
nand U6990 (N_6990,N_5546,N_5488);
or U6991 (N_6991,N_5436,N_5933);
nor U6992 (N_6992,N_4837,N_5233);
nand U6993 (N_6993,N_5749,N_4706);
nand U6994 (N_6994,N_4558,N_4569);
nor U6995 (N_6995,N_5062,N_5988);
nor U6996 (N_6996,N_4813,N_4987);
or U6997 (N_6997,N_4548,N_5673);
or U6998 (N_6998,N_5038,N_4569);
and U6999 (N_6999,N_5301,N_5344);
nand U7000 (N_7000,N_5725,N_5643);
nand U7001 (N_7001,N_5785,N_5648);
and U7002 (N_7002,N_5347,N_4563);
or U7003 (N_7003,N_4915,N_4559);
or U7004 (N_7004,N_4732,N_4612);
and U7005 (N_7005,N_4953,N_4549);
xor U7006 (N_7006,N_4921,N_5117);
or U7007 (N_7007,N_5268,N_5926);
nor U7008 (N_7008,N_5401,N_5240);
and U7009 (N_7009,N_4668,N_5596);
nor U7010 (N_7010,N_4765,N_5102);
nand U7011 (N_7011,N_4746,N_5555);
xnor U7012 (N_7012,N_4516,N_5376);
xnor U7013 (N_7013,N_5332,N_5611);
or U7014 (N_7014,N_5924,N_4877);
nand U7015 (N_7015,N_5646,N_4977);
and U7016 (N_7016,N_5334,N_5640);
or U7017 (N_7017,N_5207,N_5263);
nor U7018 (N_7018,N_5242,N_5979);
or U7019 (N_7019,N_5816,N_4744);
nor U7020 (N_7020,N_5571,N_5433);
nand U7021 (N_7021,N_5129,N_4769);
or U7022 (N_7022,N_5857,N_4805);
nor U7023 (N_7023,N_5810,N_4733);
nand U7024 (N_7024,N_4514,N_5719);
nor U7025 (N_7025,N_5032,N_5702);
nor U7026 (N_7026,N_4712,N_5181);
nor U7027 (N_7027,N_5187,N_4768);
nand U7028 (N_7028,N_5608,N_4954);
nor U7029 (N_7029,N_5143,N_5952);
nor U7030 (N_7030,N_5133,N_4652);
nor U7031 (N_7031,N_5788,N_4505);
or U7032 (N_7032,N_4992,N_5459);
nand U7033 (N_7033,N_5164,N_4964);
and U7034 (N_7034,N_5580,N_5567);
xnor U7035 (N_7035,N_5179,N_5419);
and U7036 (N_7036,N_5113,N_4893);
and U7037 (N_7037,N_4858,N_4914);
and U7038 (N_7038,N_5189,N_5494);
nand U7039 (N_7039,N_5068,N_4857);
nor U7040 (N_7040,N_4951,N_4673);
xor U7041 (N_7041,N_5950,N_5240);
xnor U7042 (N_7042,N_4638,N_5713);
or U7043 (N_7043,N_5254,N_4602);
and U7044 (N_7044,N_4593,N_4859);
nor U7045 (N_7045,N_5333,N_5673);
nor U7046 (N_7046,N_5933,N_5654);
and U7047 (N_7047,N_5537,N_4826);
nand U7048 (N_7048,N_5443,N_4536);
nand U7049 (N_7049,N_4717,N_5055);
and U7050 (N_7050,N_5946,N_5115);
or U7051 (N_7051,N_5220,N_5024);
nor U7052 (N_7052,N_5752,N_5079);
nor U7053 (N_7053,N_5836,N_4891);
nor U7054 (N_7054,N_4738,N_4554);
or U7055 (N_7055,N_4614,N_4553);
or U7056 (N_7056,N_5673,N_4788);
nand U7057 (N_7057,N_5843,N_4953);
nor U7058 (N_7058,N_5977,N_5242);
or U7059 (N_7059,N_5077,N_5996);
or U7060 (N_7060,N_5538,N_4708);
nor U7061 (N_7061,N_5558,N_4785);
nand U7062 (N_7062,N_5625,N_5034);
nor U7063 (N_7063,N_5215,N_5818);
and U7064 (N_7064,N_5998,N_5710);
and U7065 (N_7065,N_4702,N_5179);
nor U7066 (N_7066,N_5057,N_4632);
nand U7067 (N_7067,N_5318,N_5205);
or U7068 (N_7068,N_5890,N_4945);
and U7069 (N_7069,N_5927,N_4961);
nand U7070 (N_7070,N_5497,N_4938);
xnor U7071 (N_7071,N_5695,N_4544);
or U7072 (N_7072,N_5669,N_4988);
nor U7073 (N_7073,N_5874,N_5056);
nor U7074 (N_7074,N_4909,N_5931);
and U7075 (N_7075,N_5814,N_5134);
and U7076 (N_7076,N_5555,N_5259);
xnor U7077 (N_7077,N_4855,N_4631);
xor U7078 (N_7078,N_4728,N_4904);
nor U7079 (N_7079,N_4686,N_5797);
or U7080 (N_7080,N_4640,N_5661);
and U7081 (N_7081,N_4540,N_4989);
or U7082 (N_7082,N_5087,N_5722);
and U7083 (N_7083,N_5815,N_5684);
nand U7084 (N_7084,N_5775,N_5324);
nand U7085 (N_7085,N_5420,N_4896);
and U7086 (N_7086,N_4821,N_5194);
nand U7087 (N_7087,N_5389,N_5651);
nor U7088 (N_7088,N_4828,N_4864);
nor U7089 (N_7089,N_4881,N_5236);
nand U7090 (N_7090,N_4699,N_5601);
nand U7091 (N_7091,N_5751,N_5054);
or U7092 (N_7092,N_5073,N_5503);
or U7093 (N_7093,N_4698,N_5374);
nand U7094 (N_7094,N_5796,N_5903);
nand U7095 (N_7095,N_5852,N_5038);
and U7096 (N_7096,N_4933,N_5698);
nand U7097 (N_7097,N_4519,N_4640);
nor U7098 (N_7098,N_5015,N_5074);
nand U7099 (N_7099,N_5070,N_5833);
and U7100 (N_7100,N_4966,N_5723);
xnor U7101 (N_7101,N_5829,N_5338);
nor U7102 (N_7102,N_4572,N_4994);
nor U7103 (N_7103,N_4514,N_5733);
or U7104 (N_7104,N_4774,N_5061);
and U7105 (N_7105,N_4532,N_5192);
or U7106 (N_7106,N_4576,N_4943);
nand U7107 (N_7107,N_5150,N_5727);
or U7108 (N_7108,N_4715,N_5559);
nor U7109 (N_7109,N_5799,N_4987);
nor U7110 (N_7110,N_4739,N_5721);
nor U7111 (N_7111,N_5447,N_5448);
nor U7112 (N_7112,N_4837,N_5187);
nand U7113 (N_7113,N_5809,N_4590);
nand U7114 (N_7114,N_4889,N_4852);
nor U7115 (N_7115,N_5996,N_5019);
nand U7116 (N_7116,N_4584,N_4713);
nand U7117 (N_7117,N_4675,N_4524);
xnor U7118 (N_7118,N_5498,N_5741);
and U7119 (N_7119,N_5794,N_4822);
xnor U7120 (N_7120,N_4829,N_5907);
nand U7121 (N_7121,N_5922,N_4771);
or U7122 (N_7122,N_5619,N_5588);
nor U7123 (N_7123,N_5874,N_4607);
or U7124 (N_7124,N_5777,N_5719);
or U7125 (N_7125,N_4641,N_5548);
and U7126 (N_7126,N_5947,N_5640);
and U7127 (N_7127,N_5107,N_5197);
nand U7128 (N_7128,N_5158,N_5699);
nor U7129 (N_7129,N_5215,N_4810);
or U7130 (N_7130,N_5557,N_4849);
or U7131 (N_7131,N_5365,N_4839);
xor U7132 (N_7132,N_4766,N_4586);
or U7133 (N_7133,N_5076,N_5574);
and U7134 (N_7134,N_5387,N_5805);
nand U7135 (N_7135,N_5441,N_4560);
or U7136 (N_7136,N_5369,N_5289);
nand U7137 (N_7137,N_5878,N_4720);
nand U7138 (N_7138,N_5378,N_5874);
or U7139 (N_7139,N_5945,N_5885);
nand U7140 (N_7140,N_4504,N_5500);
and U7141 (N_7141,N_5682,N_4765);
or U7142 (N_7142,N_5379,N_4620);
and U7143 (N_7143,N_4783,N_4595);
xor U7144 (N_7144,N_5508,N_5588);
or U7145 (N_7145,N_4984,N_5914);
nand U7146 (N_7146,N_5048,N_4896);
nor U7147 (N_7147,N_5986,N_4796);
and U7148 (N_7148,N_4703,N_4620);
xor U7149 (N_7149,N_4521,N_5948);
nor U7150 (N_7150,N_5233,N_5761);
xnor U7151 (N_7151,N_4896,N_5655);
xor U7152 (N_7152,N_5878,N_5075);
and U7153 (N_7153,N_5380,N_4814);
nand U7154 (N_7154,N_4819,N_5864);
nand U7155 (N_7155,N_5858,N_4910);
or U7156 (N_7156,N_5372,N_5488);
nor U7157 (N_7157,N_5355,N_4942);
nor U7158 (N_7158,N_5643,N_5776);
or U7159 (N_7159,N_5684,N_4799);
or U7160 (N_7160,N_5979,N_4547);
nand U7161 (N_7161,N_5974,N_5206);
or U7162 (N_7162,N_4777,N_5358);
nor U7163 (N_7163,N_5758,N_5607);
nor U7164 (N_7164,N_5739,N_4823);
nor U7165 (N_7165,N_4906,N_4845);
or U7166 (N_7166,N_4954,N_5017);
and U7167 (N_7167,N_4656,N_5725);
and U7168 (N_7168,N_4937,N_5798);
or U7169 (N_7169,N_4687,N_4827);
and U7170 (N_7170,N_5874,N_4842);
xnor U7171 (N_7171,N_5371,N_5289);
nor U7172 (N_7172,N_5343,N_5366);
and U7173 (N_7173,N_5420,N_4955);
and U7174 (N_7174,N_5508,N_4911);
nand U7175 (N_7175,N_4774,N_5323);
or U7176 (N_7176,N_4993,N_4908);
nand U7177 (N_7177,N_4588,N_5987);
nor U7178 (N_7178,N_5562,N_5174);
and U7179 (N_7179,N_5956,N_5115);
nor U7180 (N_7180,N_4566,N_5529);
and U7181 (N_7181,N_4649,N_5526);
nand U7182 (N_7182,N_4642,N_5311);
or U7183 (N_7183,N_5837,N_5240);
and U7184 (N_7184,N_5554,N_4825);
nand U7185 (N_7185,N_5271,N_5889);
nand U7186 (N_7186,N_4654,N_5283);
nor U7187 (N_7187,N_5942,N_5894);
and U7188 (N_7188,N_5002,N_4611);
or U7189 (N_7189,N_4760,N_4989);
nor U7190 (N_7190,N_4564,N_5770);
xnor U7191 (N_7191,N_4502,N_5365);
nor U7192 (N_7192,N_4917,N_4729);
or U7193 (N_7193,N_4673,N_5753);
xor U7194 (N_7194,N_5718,N_5286);
xor U7195 (N_7195,N_5149,N_5532);
nand U7196 (N_7196,N_5044,N_4682);
and U7197 (N_7197,N_5908,N_4637);
xor U7198 (N_7198,N_5393,N_5379);
nor U7199 (N_7199,N_5555,N_4656);
or U7200 (N_7200,N_5921,N_5528);
xor U7201 (N_7201,N_5065,N_5705);
nor U7202 (N_7202,N_5219,N_5677);
and U7203 (N_7203,N_4951,N_5339);
nand U7204 (N_7204,N_5212,N_5583);
and U7205 (N_7205,N_4567,N_5325);
or U7206 (N_7206,N_5590,N_5470);
nand U7207 (N_7207,N_4951,N_5776);
and U7208 (N_7208,N_4813,N_5394);
or U7209 (N_7209,N_4524,N_5949);
nand U7210 (N_7210,N_5118,N_4916);
nor U7211 (N_7211,N_4819,N_4603);
and U7212 (N_7212,N_4845,N_5213);
and U7213 (N_7213,N_4600,N_5729);
or U7214 (N_7214,N_4602,N_5278);
or U7215 (N_7215,N_5558,N_5148);
nand U7216 (N_7216,N_5204,N_4972);
and U7217 (N_7217,N_5368,N_5241);
or U7218 (N_7218,N_5479,N_4883);
xnor U7219 (N_7219,N_4619,N_4875);
and U7220 (N_7220,N_5980,N_5680);
and U7221 (N_7221,N_5852,N_5877);
or U7222 (N_7222,N_5985,N_5203);
and U7223 (N_7223,N_5958,N_5231);
and U7224 (N_7224,N_5279,N_5449);
and U7225 (N_7225,N_5256,N_5004);
or U7226 (N_7226,N_4686,N_4905);
nand U7227 (N_7227,N_5548,N_4710);
nor U7228 (N_7228,N_5683,N_5374);
and U7229 (N_7229,N_5784,N_5456);
nand U7230 (N_7230,N_5582,N_5184);
and U7231 (N_7231,N_5979,N_5666);
or U7232 (N_7232,N_4890,N_5638);
nor U7233 (N_7233,N_4549,N_4506);
nand U7234 (N_7234,N_5112,N_5244);
xnor U7235 (N_7235,N_5533,N_5822);
or U7236 (N_7236,N_5473,N_5041);
nor U7237 (N_7237,N_5411,N_5714);
xnor U7238 (N_7238,N_5537,N_4875);
and U7239 (N_7239,N_4870,N_5657);
nand U7240 (N_7240,N_5558,N_5498);
nand U7241 (N_7241,N_5124,N_5763);
nand U7242 (N_7242,N_4577,N_5533);
nor U7243 (N_7243,N_5277,N_5651);
nand U7244 (N_7244,N_4821,N_5642);
nand U7245 (N_7245,N_4664,N_5498);
and U7246 (N_7246,N_5490,N_5529);
and U7247 (N_7247,N_5212,N_4799);
or U7248 (N_7248,N_4895,N_4820);
or U7249 (N_7249,N_4709,N_4828);
nand U7250 (N_7250,N_5686,N_5895);
xor U7251 (N_7251,N_5025,N_4980);
or U7252 (N_7252,N_5919,N_4742);
or U7253 (N_7253,N_4509,N_4877);
xnor U7254 (N_7254,N_5668,N_5380);
and U7255 (N_7255,N_4593,N_5373);
and U7256 (N_7256,N_4695,N_5151);
or U7257 (N_7257,N_4719,N_4685);
or U7258 (N_7258,N_5837,N_4915);
nand U7259 (N_7259,N_5763,N_5277);
nand U7260 (N_7260,N_5174,N_5556);
nand U7261 (N_7261,N_5578,N_5072);
nand U7262 (N_7262,N_4640,N_5263);
nand U7263 (N_7263,N_4976,N_4737);
and U7264 (N_7264,N_5723,N_5399);
nand U7265 (N_7265,N_4886,N_4726);
or U7266 (N_7266,N_5837,N_5933);
nor U7267 (N_7267,N_5588,N_4567);
or U7268 (N_7268,N_5865,N_5514);
nand U7269 (N_7269,N_5563,N_5110);
nor U7270 (N_7270,N_5221,N_4613);
or U7271 (N_7271,N_5380,N_4601);
nor U7272 (N_7272,N_5055,N_5744);
and U7273 (N_7273,N_4533,N_5032);
nand U7274 (N_7274,N_5882,N_4541);
and U7275 (N_7275,N_5209,N_4533);
nor U7276 (N_7276,N_5072,N_4516);
nor U7277 (N_7277,N_4596,N_5669);
nand U7278 (N_7278,N_4713,N_5535);
and U7279 (N_7279,N_4872,N_5170);
and U7280 (N_7280,N_4656,N_4578);
or U7281 (N_7281,N_5540,N_5651);
or U7282 (N_7282,N_4516,N_4800);
xnor U7283 (N_7283,N_5844,N_4914);
nor U7284 (N_7284,N_4697,N_5325);
nand U7285 (N_7285,N_4557,N_5834);
nand U7286 (N_7286,N_5624,N_5283);
and U7287 (N_7287,N_5008,N_4819);
and U7288 (N_7288,N_5975,N_5709);
nor U7289 (N_7289,N_5177,N_5100);
or U7290 (N_7290,N_5274,N_4818);
nand U7291 (N_7291,N_5089,N_5965);
and U7292 (N_7292,N_4539,N_4735);
nand U7293 (N_7293,N_5808,N_5852);
nand U7294 (N_7294,N_5436,N_4534);
nor U7295 (N_7295,N_5110,N_4793);
and U7296 (N_7296,N_4551,N_5485);
xnor U7297 (N_7297,N_4808,N_5346);
nand U7298 (N_7298,N_5656,N_5887);
xnor U7299 (N_7299,N_4997,N_5801);
and U7300 (N_7300,N_5933,N_5011);
and U7301 (N_7301,N_5410,N_5962);
nor U7302 (N_7302,N_5458,N_5289);
or U7303 (N_7303,N_5002,N_5506);
or U7304 (N_7304,N_5617,N_4800);
or U7305 (N_7305,N_5938,N_4734);
or U7306 (N_7306,N_4851,N_4597);
or U7307 (N_7307,N_4753,N_5180);
xor U7308 (N_7308,N_4944,N_5106);
xor U7309 (N_7309,N_5534,N_4711);
or U7310 (N_7310,N_5557,N_4874);
nand U7311 (N_7311,N_4564,N_5527);
and U7312 (N_7312,N_5851,N_5913);
or U7313 (N_7313,N_5043,N_5273);
or U7314 (N_7314,N_5867,N_5410);
xor U7315 (N_7315,N_5793,N_5100);
nand U7316 (N_7316,N_5515,N_4731);
or U7317 (N_7317,N_5973,N_5758);
nor U7318 (N_7318,N_5350,N_5767);
nand U7319 (N_7319,N_5256,N_4768);
or U7320 (N_7320,N_4976,N_5157);
nor U7321 (N_7321,N_5828,N_5605);
or U7322 (N_7322,N_5450,N_4752);
nand U7323 (N_7323,N_5062,N_5151);
nor U7324 (N_7324,N_5523,N_5004);
nand U7325 (N_7325,N_5011,N_5041);
nor U7326 (N_7326,N_5538,N_4769);
nor U7327 (N_7327,N_4781,N_5694);
or U7328 (N_7328,N_5739,N_4716);
nor U7329 (N_7329,N_5925,N_5700);
or U7330 (N_7330,N_5663,N_5367);
nand U7331 (N_7331,N_5425,N_5330);
and U7332 (N_7332,N_5314,N_4528);
xnor U7333 (N_7333,N_4878,N_4636);
and U7334 (N_7334,N_5269,N_5748);
nor U7335 (N_7335,N_4586,N_4948);
or U7336 (N_7336,N_4504,N_5347);
xnor U7337 (N_7337,N_5856,N_5255);
xnor U7338 (N_7338,N_4946,N_5973);
nand U7339 (N_7339,N_5209,N_5571);
and U7340 (N_7340,N_5367,N_4565);
nand U7341 (N_7341,N_5432,N_5841);
or U7342 (N_7342,N_5463,N_5094);
or U7343 (N_7343,N_5148,N_5231);
xnor U7344 (N_7344,N_5025,N_5752);
and U7345 (N_7345,N_5916,N_5727);
nor U7346 (N_7346,N_5066,N_4890);
nor U7347 (N_7347,N_5941,N_5699);
or U7348 (N_7348,N_4847,N_5445);
xor U7349 (N_7349,N_4588,N_5323);
nand U7350 (N_7350,N_4512,N_4893);
and U7351 (N_7351,N_4958,N_5009);
nor U7352 (N_7352,N_5730,N_5935);
xor U7353 (N_7353,N_4654,N_5418);
xor U7354 (N_7354,N_5532,N_4685);
or U7355 (N_7355,N_4843,N_5589);
and U7356 (N_7356,N_5134,N_5114);
or U7357 (N_7357,N_5713,N_4824);
nor U7358 (N_7358,N_4786,N_4573);
nand U7359 (N_7359,N_4758,N_5391);
nor U7360 (N_7360,N_5827,N_5613);
and U7361 (N_7361,N_5085,N_4832);
nand U7362 (N_7362,N_5494,N_4888);
xnor U7363 (N_7363,N_4525,N_5882);
nor U7364 (N_7364,N_5875,N_5600);
nand U7365 (N_7365,N_5253,N_4786);
nand U7366 (N_7366,N_5331,N_5615);
and U7367 (N_7367,N_4955,N_5521);
and U7368 (N_7368,N_5750,N_5372);
and U7369 (N_7369,N_4835,N_5935);
nand U7370 (N_7370,N_5451,N_5758);
or U7371 (N_7371,N_4871,N_5368);
nor U7372 (N_7372,N_5370,N_5610);
nand U7373 (N_7373,N_4697,N_5055);
nand U7374 (N_7374,N_5731,N_5127);
nand U7375 (N_7375,N_5692,N_5836);
or U7376 (N_7376,N_5209,N_4812);
or U7377 (N_7377,N_5708,N_4518);
nand U7378 (N_7378,N_5681,N_5756);
nor U7379 (N_7379,N_5252,N_5664);
and U7380 (N_7380,N_5054,N_5882);
xnor U7381 (N_7381,N_4949,N_5361);
xor U7382 (N_7382,N_5254,N_5458);
nor U7383 (N_7383,N_5513,N_4557);
nand U7384 (N_7384,N_5524,N_5383);
nor U7385 (N_7385,N_5015,N_5991);
xnor U7386 (N_7386,N_5710,N_5989);
or U7387 (N_7387,N_4950,N_4574);
nand U7388 (N_7388,N_4700,N_4849);
nand U7389 (N_7389,N_4538,N_4829);
or U7390 (N_7390,N_5118,N_5583);
nor U7391 (N_7391,N_4724,N_4795);
and U7392 (N_7392,N_5822,N_5315);
xor U7393 (N_7393,N_5563,N_5007);
xnor U7394 (N_7394,N_5961,N_5197);
nand U7395 (N_7395,N_4694,N_4827);
nand U7396 (N_7396,N_5421,N_4896);
or U7397 (N_7397,N_5967,N_4995);
nor U7398 (N_7398,N_4838,N_5445);
nor U7399 (N_7399,N_4759,N_5374);
or U7400 (N_7400,N_5090,N_4945);
nand U7401 (N_7401,N_4589,N_5124);
and U7402 (N_7402,N_5483,N_5135);
nor U7403 (N_7403,N_5713,N_4806);
or U7404 (N_7404,N_5956,N_4858);
or U7405 (N_7405,N_5829,N_5741);
nor U7406 (N_7406,N_4798,N_5346);
and U7407 (N_7407,N_5049,N_5525);
or U7408 (N_7408,N_5870,N_5993);
and U7409 (N_7409,N_5324,N_5335);
xnor U7410 (N_7410,N_4766,N_5580);
nor U7411 (N_7411,N_4646,N_5725);
nor U7412 (N_7412,N_4991,N_5491);
nand U7413 (N_7413,N_5468,N_5519);
xnor U7414 (N_7414,N_4929,N_4960);
nand U7415 (N_7415,N_4712,N_5015);
xor U7416 (N_7416,N_5419,N_5314);
or U7417 (N_7417,N_5369,N_5190);
and U7418 (N_7418,N_5296,N_5972);
nand U7419 (N_7419,N_5703,N_4616);
and U7420 (N_7420,N_5528,N_5736);
or U7421 (N_7421,N_4997,N_4730);
or U7422 (N_7422,N_5389,N_5533);
nor U7423 (N_7423,N_5558,N_4619);
nor U7424 (N_7424,N_5567,N_4750);
nand U7425 (N_7425,N_4845,N_4884);
and U7426 (N_7426,N_5845,N_5878);
xor U7427 (N_7427,N_5991,N_5636);
nand U7428 (N_7428,N_4570,N_4575);
and U7429 (N_7429,N_5578,N_5007);
xor U7430 (N_7430,N_5666,N_4608);
xor U7431 (N_7431,N_5652,N_4776);
and U7432 (N_7432,N_4824,N_4572);
or U7433 (N_7433,N_4554,N_5700);
nand U7434 (N_7434,N_5932,N_5062);
and U7435 (N_7435,N_5268,N_4726);
nand U7436 (N_7436,N_5141,N_5056);
or U7437 (N_7437,N_5019,N_4996);
or U7438 (N_7438,N_5120,N_5354);
or U7439 (N_7439,N_5328,N_4613);
and U7440 (N_7440,N_5040,N_5963);
nand U7441 (N_7441,N_5597,N_5897);
and U7442 (N_7442,N_5245,N_4985);
nand U7443 (N_7443,N_4628,N_5657);
nand U7444 (N_7444,N_5550,N_4511);
and U7445 (N_7445,N_4952,N_4707);
nand U7446 (N_7446,N_5805,N_5147);
nor U7447 (N_7447,N_4969,N_5015);
and U7448 (N_7448,N_5493,N_5434);
and U7449 (N_7449,N_5659,N_4879);
nand U7450 (N_7450,N_5820,N_5977);
nand U7451 (N_7451,N_5392,N_4855);
and U7452 (N_7452,N_5881,N_5379);
and U7453 (N_7453,N_5777,N_5786);
or U7454 (N_7454,N_5549,N_4954);
or U7455 (N_7455,N_5161,N_5852);
xor U7456 (N_7456,N_4932,N_5476);
nor U7457 (N_7457,N_4545,N_5100);
and U7458 (N_7458,N_5317,N_5383);
and U7459 (N_7459,N_5699,N_5128);
nand U7460 (N_7460,N_4683,N_5908);
and U7461 (N_7461,N_5762,N_5133);
xor U7462 (N_7462,N_5930,N_4892);
xor U7463 (N_7463,N_5695,N_5373);
and U7464 (N_7464,N_4531,N_4554);
nor U7465 (N_7465,N_5810,N_5149);
nor U7466 (N_7466,N_4868,N_5442);
xor U7467 (N_7467,N_5305,N_5422);
and U7468 (N_7468,N_4831,N_4882);
or U7469 (N_7469,N_5719,N_5770);
and U7470 (N_7470,N_5937,N_5900);
nand U7471 (N_7471,N_4591,N_4761);
nand U7472 (N_7472,N_4587,N_4632);
nand U7473 (N_7473,N_4640,N_5230);
nand U7474 (N_7474,N_4649,N_5288);
nand U7475 (N_7475,N_5332,N_4614);
or U7476 (N_7476,N_5056,N_5350);
or U7477 (N_7477,N_5318,N_5911);
and U7478 (N_7478,N_5454,N_4851);
nand U7479 (N_7479,N_4816,N_5480);
nand U7480 (N_7480,N_4872,N_4659);
nor U7481 (N_7481,N_5401,N_4858);
nor U7482 (N_7482,N_5627,N_4621);
and U7483 (N_7483,N_5827,N_5132);
nand U7484 (N_7484,N_4513,N_4913);
nor U7485 (N_7485,N_5898,N_5621);
nand U7486 (N_7486,N_5623,N_5748);
nor U7487 (N_7487,N_5758,N_5959);
nand U7488 (N_7488,N_5758,N_5449);
xnor U7489 (N_7489,N_4522,N_5885);
nand U7490 (N_7490,N_5921,N_5251);
and U7491 (N_7491,N_4702,N_5252);
xor U7492 (N_7492,N_5683,N_4625);
nor U7493 (N_7493,N_5438,N_5910);
and U7494 (N_7494,N_4601,N_5109);
xnor U7495 (N_7495,N_5533,N_5278);
nand U7496 (N_7496,N_5520,N_5539);
nor U7497 (N_7497,N_4783,N_5047);
or U7498 (N_7498,N_5609,N_4998);
and U7499 (N_7499,N_4622,N_4963);
or U7500 (N_7500,N_6808,N_7241);
nand U7501 (N_7501,N_7111,N_7369);
nor U7502 (N_7502,N_7313,N_6827);
xor U7503 (N_7503,N_6675,N_6847);
or U7504 (N_7504,N_6903,N_6050);
or U7505 (N_7505,N_6452,N_6739);
nand U7506 (N_7506,N_6367,N_7475);
nand U7507 (N_7507,N_6942,N_6843);
and U7508 (N_7508,N_6248,N_7028);
xnor U7509 (N_7509,N_7181,N_6465);
or U7510 (N_7510,N_7389,N_6812);
nand U7511 (N_7511,N_7092,N_7271);
or U7512 (N_7512,N_7007,N_6447);
nand U7513 (N_7513,N_6134,N_7406);
and U7514 (N_7514,N_6947,N_6585);
nor U7515 (N_7515,N_6940,N_7094);
xnor U7516 (N_7516,N_7299,N_7414);
nor U7517 (N_7517,N_7168,N_6271);
nor U7518 (N_7518,N_6058,N_7477);
and U7519 (N_7519,N_6820,N_6784);
and U7520 (N_7520,N_6118,N_6000);
or U7521 (N_7521,N_6354,N_6706);
nor U7522 (N_7522,N_6399,N_7073);
nor U7523 (N_7523,N_6573,N_6148);
xnor U7524 (N_7524,N_6082,N_6147);
or U7525 (N_7525,N_7067,N_6306);
or U7526 (N_7526,N_7180,N_7485);
nand U7527 (N_7527,N_6873,N_7176);
nor U7528 (N_7528,N_6772,N_6714);
nor U7529 (N_7529,N_6830,N_7309);
or U7530 (N_7530,N_7050,N_6881);
and U7531 (N_7531,N_6021,N_7266);
nand U7532 (N_7532,N_6020,N_6995);
xnor U7533 (N_7533,N_6123,N_6298);
nor U7534 (N_7534,N_6076,N_6190);
or U7535 (N_7535,N_7471,N_6448);
or U7536 (N_7536,N_7053,N_7203);
nand U7537 (N_7537,N_7156,N_6192);
or U7538 (N_7538,N_7441,N_7044);
nand U7539 (N_7539,N_6136,N_7012);
nand U7540 (N_7540,N_6799,N_6958);
or U7541 (N_7541,N_7341,N_6682);
and U7542 (N_7542,N_7136,N_7319);
nor U7543 (N_7543,N_6727,N_6900);
or U7544 (N_7544,N_6960,N_6048);
or U7545 (N_7545,N_6894,N_7242);
xnor U7546 (N_7546,N_7106,N_7404);
nand U7547 (N_7547,N_6583,N_6909);
or U7548 (N_7548,N_6009,N_6911);
or U7549 (N_7549,N_6528,N_6420);
or U7550 (N_7550,N_6987,N_6033);
or U7551 (N_7551,N_7324,N_6029);
xnor U7552 (N_7552,N_7353,N_7129);
and U7553 (N_7553,N_7010,N_6926);
nand U7554 (N_7554,N_6760,N_6007);
and U7555 (N_7555,N_6416,N_6219);
and U7556 (N_7556,N_6150,N_6487);
or U7557 (N_7557,N_6652,N_7030);
or U7558 (N_7558,N_6647,N_7009);
or U7559 (N_7559,N_7470,N_7461);
nand U7560 (N_7560,N_6746,N_7458);
or U7561 (N_7561,N_7302,N_6563);
nand U7562 (N_7562,N_7356,N_7188);
and U7563 (N_7563,N_6197,N_7000);
or U7564 (N_7564,N_6419,N_6196);
nor U7565 (N_7565,N_6172,N_6656);
and U7566 (N_7566,N_7339,N_6941);
and U7567 (N_7567,N_6587,N_6855);
nand U7568 (N_7568,N_6501,N_6993);
and U7569 (N_7569,N_6923,N_6616);
nor U7570 (N_7570,N_6520,N_7005);
and U7571 (N_7571,N_6054,N_6317);
xor U7572 (N_7572,N_6034,N_6715);
or U7573 (N_7573,N_7175,N_6445);
and U7574 (N_7574,N_6291,N_6829);
or U7575 (N_7575,N_7371,N_7059);
xnor U7576 (N_7576,N_6260,N_7365);
or U7577 (N_7577,N_7442,N_6632);
and U7578 (N_7578,N_6906,N_6622);
or U7579 (N_7579,N_6166,N_6879);
nand U7580 (N_7580,N_7400,N_7103);
nor U7581 (N_7581,N_7446,N_6188);
nand U7582 (N_7582,N_7427,N_6691);
nand U7583 (N_7583,N_7114,N_6561);
nand U7584 (N_7584,N_6098,N_7417);
and U7585 (N_7585,N_7056,N_6513);
nand U7586 (N_7586,N_6815,N_6075);
xor U7587 (N_7587,N_6731,N_6154);
nand U7588 (N_7588,N_6878,N_7373);
and U7589 (N_7589,N_6686,N_7047);
nand U7590 (N_7590,N_6174,N_7318);
or U7591 (N_7591,N_6981,N_7454);
nor U7592 (N_7592,N_7394,N_6552);
nand U7593 (N_7593,N_6112,N_6488);
nor U7594 (N_7594,N_6766,N_6756);
nand U7595 (N_7595,N_7230,N_7143);
nand U7596 (N_7596,N_7322,N_6945);
or U7597 (N_7597,N_7054,N_7431);
nor U7598 (N_7598,N_6948,N_6822);
or U7599 (N_7599,N_6544,N_6730);
nand U7600 (N_7600,N_6685,N_6200);
nor U7601 (N_7601,N_6162,N_7061);
nand U7602 (N_7602,N_7002,N_7126);
nand U7603 (N_7603,N_6968,N_6755);
or U7604 (N_7604,N_7447,N_6998);
nand U7605 (N_7605,N_6574,N_6964);
and U7606 (N_7606,N_7307,N_6687);
nor U7607 (N_7607,N_6074,N_6592);
or U7608 (N_7608,N_6439,N_6762);
nor U7609 (N_7609,N_6671,N_6626);
and U7610 (N_7610,N_7069,N_6594);
or U7611 (N_7611,N_6156,N_6710);
and U7612 (N_7612,N_7121,N_7088);
nand U7613 (N_7613,N_7193,N_6599);
xor U7614 (N_7614,N_7274,N_6584);
nor U7615 (N_7615,N_7240,N_6179);
and U7616 (N_7616,N_7004,N_6153);
and U7617 (N_7617,N_6523,N_6289);
and U7618 (N_7618,N_6704,N_6937);
and U7619 (N_7619,N_6231,N_6272);
or U7620 (N_7620,N_7185,N_7418);
and U7621 (N_7621,N_7253,N_7478);
nor U7622 (N_7622,N_7452,N_7157);
nor U7623 (N_7623,N_6598,N_6888);
nand U7624 (N_7624,N_6770,N_6208);
or U7625 (N_7625,N_6159,N_7158);
or U7626 (N_7626,N_6230,N_7084);
nor U7627 (N_7627,N_6660,N_6758);
nand U7628 (N_7628,N_6538,N_7236);
or U7629 (N_7629,N_6553,N_7104);
nand U7630 (N_7630,N_6546,N_7306);
nand U7631 (N_7631,N_6170,N_6176);
xor U7632 (N_7632,N_6117,N_6434);
and U7633 (N_7633,N_7419,N_7037);
and U7634 (N_7634,N_6576,N_6939);
xnor U7635 (N_7635,N_6044,N_7448);
and U7636 (N_7636,N_6525,N_7423);
nand U7637 (N_7637,N_6071,N_6446);
or U7638 (N_7638,N_6883,N_7166);
nand U7639 (N_7639,N_6910,N_7277);
or U7640 (N_7640,N_6678,N_7382);
or U7641 (N_7641,N_6423,N_6454);
nor U7642 (N_7642,N_6751,N_6902);
or U7643 (N_7643,N_7496,N_6030);
or U7644 (N_7644,N_7314,N_6719);
and U7645 (N_7645,N_6823,N_6807);
nand U7646 (N_7646,N_6703,N_6612);
and U7647 (N_7647,N_7378,N_6386);
or U7648 (N_7648,N_6411,N_7479);
and U7649 (N_7649,N_6657,N_7125);
nand U7650 (N_7650,N_6177,N_7410);
xnor U7651 (N_7651,N_6066,N_6346);
nand U7652 (N_7652,N_6341,N_6249);
or U7653 (N_7653,N_7215,N_7021);
nor U7654 (N_7654,N_7492,N_7364);
xor U7655 (N_7655,N_7097,N_6936);
or U7656 (N_7656,N_6314,N_6173);
nand U7657 (N_7657,N_7337,N_7467);
xnor U7658 (N_7658,N_6433,N_6845);
nor U7659 (N_7659,N_7110,N_6957);
and U7660 (N_7660,N_7335,N_7233);
or U7661 (N_7661,N_6068,N_6108);
or U7662 (N_7662,N_6677,N_6056);
or U7663 (N_7663,N_6429,N_6253);
nand U7664 (N_7664,N_6398,N_6466);
and U7665 (N_7665,N_6654,N_6359);
and U7666 (N_7666,N_6426,N_7334);
or U7667 (N_7667,N_7395,N_6524);
and U7668 (N_7668,N_7172,N_6099);
nand U7669 (N_7669,N_7312,N_7279);
and U7670 (N_7670,N_6861,N_7015);
and U7671 (N_7671,N_6522,N_7433);
nor U7672 (N_7672,N_6832,N_6593);
and U7673 (N_7673,N_7023,N_7331);
and U7674 (N_7674,N_6921,N_7098);
and U7675 (N_7675,N_6158,N_7301);
and U7676 (N_7676,N_6498,N_7354);
or U7677 (N_7677,N_6182,N_6540);
nor U7678 (N_7678,N_6672,N_6613);
nand U7679 (N_7679,N_6178,N_6326);
or U7680 (N_7680,N_6803,N_6602);
xor U7681 (N_7681,N_6167,N_7255);
and U7682 (N_7682,N_6623,N_6745);
and U7683 (N_7683,N_7208,N_6673);
xnor U7684 (N_7684,N_7330,N_7495);
nor U7685 (N_7685,N_6798,N_7090);
xnor U7686 (N_7686,N_7042,N_7179);
or U7687 (N_7687,N_6103,N_7049);
nand U7688 (N_7688,N_6813,N_6251);
and U7689 (N_7689,N_7304,N_6637);
nor U7690 (N_7690,N_6336,N_6383);
and U7691 (N_7691,N_7064,N_7290);
xor U7692 (N_7692,N_6826,N_6155);
nand U7693 (N_7693,N_6031,N_7192);
and U7694 (N_7694,N_6045,N_6581);
nor U7695 (N_7695,N_6129,N_7041);
and U7696 (N_7696,N_7439,N_7018);
or U7697 (N_7697,N_6478,N_6436);
nor U7698 (N_7698,N_6629,N_6535);
and U7699 (N_7699,N_6287,N_6662);
or U7700 (N_7700,N_6787,N_7093);
or U7701 (N_7701,N_6116,N_6290);
xor U7702 (N_7702,N_7276,N_6062);
and U7703 (N_7703,N_6709,N_7288);
nand U7704 (N_7704,N_6925,N_6791);
and U7705 (N_7705,N_7183,N_7197);
nand U7706 (N_7706,N_6224,N_6839);
nand U7707 (N_7707,N_6049,N_6037);
or U7708 (N_7708,N_7194,N_6181);
nor U7709 (N_7709,N_7155,N_7117);
or U7710 (N_7710,N_6027,N_6320);
or U7711 (N_7711,N_7095,N_6226);
and U7712 (N_7712,N_6459,N_6198);
and U7713 (N_7713,N_7174,N_6644);
nor U7714 (N_7714,N_7296,N_6476);
nor U7715 (N_7715,N_6761,N_6774);
or U7716 (N_7716,N_7162,N_7430);
or U7717 (N_7717,N_7191,N_7469);
and U7718 (N_7718,N_6018,N_7115);
or U7719 (N_7719,N_6352,N_7038);
and U7720 (N_7720,N_6024,N_6254);
or U7721 (N_7721,N_6299,N_7150);
or U7722 (N_7722,N_6413,N_6779);
and U7723 (N_7723,N_6504,N_6880);
or U7724 (N_7724,N_6972,N_6281);
and U7725 (N_7725,N_6577,N_6959);
or U7726 (N_7726,N_6139,N_6407);
or U7727 (N_7727,N_6956,N_6014);
and U7728 (N_7728,N_6418,N_6953);
nor U7729 (N_7729,N_7380,N_6624);
xnor U7730 (N_7730,N_6405,N_7344);
xnor U7731 (N_7731,N_6194,N_6935);
or U7732 (N_7732,N_6651,N_7317);
nand U7733 (N_7733,N_7426,N_6328);
or U7734 (N_7734,N_6676,N_6350);
xor U7735 (N_7735,N_6640,N_6424);
and U7736 (N_7736,N_6195,N_6381);
and U7737 (N_7737,N_7286,N_6060);
and U7738 (N_7738,N_6296,N_7247);
and U7739 (N_7739,N_7078,N_7081);
nand U7740 (N_7740,N_7167,N_7292);
nor U7741 (N_7741,N_6580,N_6143);
and U7742 (N_7742,N_7029,N_6639);
and U7743 (N_7743,N_6617,N_7220);
or U7744 (N_7744,N_7403,N_7333);
and U7745 (N_7745,N_6858,N_6451);
or U7746 (N_7746,N_7281,N_6674);
nand U7747 (N_7747,N_6893,N_6087);
nand U7748 (N_7748,N_6868,N_6363);
nand U7749 (N_7749,N_6047,N_6063);
nand U7750 (N_7750,N_7248,N_6518);
and U7751 (N_7751,N_6978,N_6396);
and U7752 (N_7752,N_6737,N_7351);
and U7753 (N_7753,N_7204,N_6088);
or U7754 (N_7754,N_6521,N_7466);
or U7755 (N_7755,N_7130,N_7421);
xnor U7756 (N_7756,N_7184,N_6729);
xor U7757 (N_7757,N_7284,N_6467);
and U7758 (N_7758,N_6023,N_6963);
nand U7759 (N_7759,N_6241,N_6876);
nor U7760 (N_7760,N_7374,N_7034);
xor U7761 (N_7761,N_6505,N_6951);
xnor U7762 (N_7762,N_7264,N_6851);
xnor U7763 (N_7763,N_6242,N_6468);
or U7764 (N_7764,N_6754,N_6450);
and U7765 (N_7765,N_6889,N_6526);
nor U7766 (N_7766,N_7295,N_7391);
or U7767 (N_7767,N_6223,N_6109);
nand U7768 (N_7768,N_7428,N_6225);
nand U7769 (N_7769,N_6286,N_7138);
nor U7770 (N_7770,N_7213,N_6252);
and U7771 (N_7771,N_7108,N_6015);
and U7772 (N_7772,N_6236,N_6274);
xor U7773 (N_7773,N_6740,N_7152);
nand U7774 (N_7774,N_7127,N_6205);
or U7775 (N_7775,N_6543,N_6991);
and U7776 (N_7776,N_7209,N_6872);
nand U7777 (N_7777,N_6119,N_6469);
or U7778 (N_7778,N_7057,N_6933);
nor U7779 (N_7779,N_6856,N_7082);
nand U7780 (N_7780,N_6705,N_7463);
nand U7781 (N_7781,N_6759,N_6841);
and U7782 (N_7782,N_6069,N_7457);
xor U7783 (N_7783,N_6428,N_6595);
xor U7784 (N_7784,N_6897,N_7462);
or U7785 (N_7785,N_7298,N_7385);
or U7786 (N_7786,N_6137,N_6749);
or U7787 (N_7787,N_6510,N_6268);
nor U7788 (N_7788,N_6800,N_6794);
and U7789 (N_7789,N_7397,N_6548);
nand U7790 (N_7790,N_6221,N_6276);
nand U7791 (N_7791,N_6569,N_7133);
nor U7792 (N_7792,N_6128,N_7486);
nor U7793 (N_7793,N_6920,N_6517);
xnor U7794 (N_7794,N_6261,N_6421);
nor U7795 (N_7795,N_6683,N_6578);
or U7796 (N_7796,N_7392,N_6722);
or U7797 (N_7797,N_7438,N_7372);
and U7798 (N_7798,N_7216,N_7122);
or U7799 (N_7799,N_7480,N_6091);
or U7800 (N_7800,N_6366,N_7214);
nand U7801 (N_7801,N_6619,N_6508);
nor U7802 (N_7802,N_6701,N_6022);
xor U7803 (N_7803,N_6110,N_6896);
or U7804 (N_7804,N_6011,N_7390);
nand U7805 (N_7805,N_6734,N_6319);
nand U7806 (N_7806,N_6885,N_6202);
nand U7807 (N_7807,N_6372,N_6688);
or U7808 (N_7808,N_7338,N_6771);
nand U7809 (N_7809,N_6782,N_6204);
nand U7810 (N_7810,N_6887,N_6892);
or U7811 (N_7811,N_6057,N_6643);
xor U7812 (N_7812,N_6401,N_6360);
and U7813 (N_7813,N_6470,N_7013);
and U7814 (N_7814,N_6625,N_7109);
and U7815 (N_7815,N_6975,N_7280);
nand U7816 (N_7816,N_6788,N_6562);
and U7817 (N_7817,N_6008,N_7405);
or U7818 (N_7818,N_6690,N_6485);
and U7819 (N_7819,N_6615,N_7261);
nor U7820 (N_7820,N_6406,N_7226);
and U7821 (N_7821,N_6663,N_6560);
xor U7822 (N_7822,N_6131,N_6275);
or U7823 (N_7823,N_6438,N_6618);
or U7824 (N_7824,N_6149,N_6785);
and U7825 (N_7825,N_6353,N_7416);
or U7826 (N_7826,N_7198,N_6984);
and U7827 (N_7827,N_6209,N_6541);
or U7828 (N_7828,N_6748,N_6515);
and U7829 (N_7829,N_7259,N_6309);
or U7830 (N_7830,N_6871,N_6781);
and U7831 (N_7831,N_6141,N_6596);
or U7832 (N_7832,N_7003,N_6665);
nor U7833 (N_7833,N_6816,N_7011);
xor U7834 (N_7834,N_6097,N_7346);
nor U7835 (N_7835,N_6977,N_6012);
xor U7836 (N_7836,N_6111,N_6554);
nand U7837 (N_7837,N_6973,N_6831);
nand U7838 (N_7838,N_6404,N_6232);
or U7839 (N_7839,N_7362,N_6486);
or U7840 (N_7840,N_6165,N_6990);
xor U7841 (N_7841,N_6104,N_6567);
nand U7842 (N_7842,N_6575,N_7258);
xor U7843 (N_7843,N_7490,N_7178);
nor U7844 (N_7844,N_6453,N_6240);
and U7845 (N_7845,N_6073,N_6928);
and U7846 (N_7846,N_6443,N_6989);
and U7847 (N_7847,N_6850,N_6101);
nor U7848 (N_7848,N_6979,N_6093);
nor U7849 (N_7849,N_6283,N_6122);
nand U7850 (N_7850,N_7221,N_6742);
nand U7851 (N_7851,N_6475,N_7497);
or U7852 (N_7852,N_6915,N_7119);
nand U7853 (N_7853,N_6713,N_7205);
or U7854 (N_7854,N_6113,N_6806);
nand U7855 (N_7855,N_7349,N_6245);
nor U7856 (N_7856,N_7422,N_6650);
or U7857 (N_7857,N_6493,N_7498);
nand U7858 (N_7858,N_7336,N_7164);
nand U7859 (N_7859,N_6400,N_7275);
and U7860 (N_7860,N_6456,N_7291);
nand U7861 (N_7861,N_6222,N_6345);
nor U7862 (N_7862,N_6218,N_6065);
or U7863 (N_7863,N_6321,N_7083);
nor U7864 (N_7864,N_6130,N_6938);
nand U7865 (N_7865,N_6497,N_6262);
xnor U7866 (N_7866,N_7432,N_6708);
and U7867 (N_7867,N_6792,N_6600);
nand U7868 (N_7868,N_6532,N_7161);
nand U7869 (N_7869,N_6944,N_6330);
or U7870 (N_7870,N_6661,N_6768);
and U7871 (N_7871,N_6233,N_6107);
or U7872 (N_7872,N_6536,N_6934);
nand U7873 (N_7873,N_7376,N_6971);
nor U7874 (N_7874,N_6607,N_7315);
and U7875 (N_7875,N_6636,N_6085);
xor U7876 (N_7876,N_6904,N_6482);
or U7877 (N_7877,N_7375,N_6606);
or U7878 (N_7878,N_7272,N_6999);
nand U7879 (N_7879,N_6899,N_6988);
or U7880 (N_7880,N_6234,N_6358);
nand U7881 (N_7881,N_6125,N_6735);
or U7882 (N_7882,N_7357,N_6763);
nand U7883 (N_7883,N_6946,N_7408);
nor U7884 (N_7884,N_6982,N_6862);
nor U7885 (N_7885,N_6343,N_6059);
and U7886 (N_7886,N_6821,N_7483);
and U7887 (N_7887,N_6696,N_6891);
or U7888 (N_7888,N_6002,N_7355);
and U7889 (N_7889,N_6649,N_7060);
nor U7890 (N_7890,N_7252,N_6474);
or U7891 (N_7891,N_7032,N_6444);
or U7892 (N_7892,N_6414,N_6187);
or U7893 (N_7893,N_6601,N_6670);
nor U7894 (N_7894,N_6724,N_6203);
nor U7895 (N_7895,N_6417,N_6611);
nand U7896 (N_7896,N_7434,N_6288);
and U7897 (N_7897,N_6503,N_7345);
nor U7898 (N_7898,N_6371,N_6431);
and U7899 (N_7899,N_6913,N_6375);
and U7900 (N_7900,N_6974,N_6409);
or U7901 (N_7901,N_7407,N_7238);
or U7902 (N_7902,N_7347,N_6259);
and U7903 (N_7903,N_7019,N_6531);
nor U7904 (N_7904,N_7107,N_6916);
nor U7905 (N_7905,N_6064,N_7300);
nor U7906 (N_7906,N_7250,N_6095);
and U7907 (N_7907,N_6094,N_7024);
and U7908 (N_7908,N_6983,N_7366);
nand U7909 (N_7909,N_6461,N_6492);
xor U7910 (N_7910,N_6322,N_7112);
or U7911 (N_7911,N_6385,N_6356);
and U7912 (N_7912,N_7245,N_6929);
nor U7913 (N_7913,N_6627,N_7293);
nor U7914 (N_7914,N_6080,N_6707);
and U7915 (N_7915,N_6216,N_6457);
or U7916 (N_7916,N_7035,N_7232);
or U7917 (N_7917,N_7223,N_6537);
nand U7918 (N_7918,N_6645,N_6115);
xor U7919 (N_7919,N_7268,N_7260);
and U7920 (N_7920,N_6040,N_6684);
and U7921 (N_7921,N_6695,N_6310);
nand U7922 (N_7922,N_7171,N_7487);
and U7923 (N_7923,N_6519,N_7144);
xor U7924 (N_7924,N_6114,N_6171);
or U7925 (N_7925,N_7285,N_6667);
or U7926 (N_7926,N_7388,N_7101);
or U7927 (N_7927,N_7451,N_6490);
or U7928 (N_7928,N_6316,N_6185);
nand U7929 (N_7929,N_6952,N_7071);
nand U7930 (N_7930,N_6848,N_6379);
nor U7931 (N_7931,N_7160,N_6392);
and U7932 (N_7932,N_6516,N_6324);
nor U7933 (N_7933,N_6303,N_6403);
and U7934 (N_7934,N_6373,N_6266);
or U7935 (N_7935,N_7066,N_7476);
or U7936 (N_7936,N_6752,N_6874);
nor U7937 (N_7937,N_6042,N_6698);
or U7938 (N_7938,N_7320,N_7459);
nand U7939 (N_7939,N_7048,N_6693);
and U7940 (N_7940,N_6484,N_6702);
xor U7941 (N_7941,N_6086,N_6043);
nor U7942 (N_7942,N_6864,N_6284);
xor U7943 (N_7943,N_7128,N_6603);
or U7944 (N_7944,N_6743,N_6610);
nor U7945 (N_7945,N_6238,N_6680);
nand U7946 (N_7946,N_6364,N_7257);
and U7947 (N_7947,N_7008,N_7140);
nand U7948 (N_7948,N_7100,N_6228);
nand U7949 (N_7949,N_6757,N_6175);
xor U7950 (N_7950,N_6295,N_6529);
or U7951 (N_7951,N_7332,N_6494);
or U7952 (N_7952,N_6070,N_6302);
or U7953 (N_7953,N_6186,N_6912);
nand U7954 (N_7954,N_6697,N_6747);
nand U7955 (N_7955,N_6917,N_6332);
or U7956 (N_7956,N_6801,N_7225);
nor U7957 (N_7957,N_6716,N_6135);
xor U7958 (N_7958,N_7381,N_6315);
nor U7959 (N_7959,N_6163,N_7363);
and U7960 (N_7960,N_6395,N_6837);
or U7961 (N_7961,N_7358,N_6633);
and U7962 (N_7962,N_7249,N_6997);
and U7963 (N_7963,N_6870,N_7246);
xor U7964 (N_7964,N_6437,N_6374);
nand U7965 (N_7965,N_6700,N_6199);
or U7966 (N_7966,N_7440,N_6214);
or U7967 (N_7967,N_7170,N_7411);
xnor U7968 (N_7968,N_6986,N_6384);
nor U7969 (N_7969,N_6124,N_6140);
or U7970 (N_7970,N_7142,N_6846);
and U7971 (N_7971,N_6083,N_6402);
and U7972 (N_7972,N_6293,N_6530);
nand U7973 (N_7973,N_6327,N_6255);
nand U7974 (N_7974,N_6246,N_7413);
or U7975 (N_7975,N_6863,N_6767);
or U7976 (N_7976,N_6072,N_6144);
or U7977 (N_7977,N_7025,N_7494);
and U7978 (N_7978,N_6814,N_7489);
and U7979 (N_7979,N_6985,N_6160);
and U7980 (N_7980,N_7200,N_7022);
nand U7981 (N_7981,N_7244,N_6961);
nand U7982 (N_7982,N_6765,N_7465);
nor U7983 (N_7983,N_7352,N_6010);
or U7984 (N_7984,N_6570,N_6355);
nor U7985 (N_7985,N_7415,N_7474);
xor U7986 (N_7986,N_6970,N_6338);
or U7987 (N_7987,N_7177,N_6263);
nor U7988 (N_7988,N_6631,N_7287);
nand U7989 (N_7989,N_7072,N_6499);
nand U7990 (N_7990,N_7113,N_6164);
nand U7991 (N_7991,N_6718,N_7350);
nor U7992 (N_7992,N_7055,N_7086);
nand U7993 (N_7993,N_6005,N_6733);
or U7994 (N_7994,N_7243,N_7173);
nand U7995 (N_7995,N_6919,N_7062);
nand U7996 (N_7996,N_7137,N_6491);
nand U7997 (N_7997,N_7368,N_6282);
nor U7998 (N_7998,N_7063,N_7045);
nand U7999 (N_7999,N_6854,N_7085);
nor U8000 (N_8000,N_6053,N_6509);
nand U8001 (N_8001,N_6728,N_6559);
and U8002 (N_8002,N_6455,N_6308);
nand U8003 (N_8003,N_6753,N_7096);
nand U8004 (N_8004,N_6250,N_6720);
xnor U8005 (N_8005,N_6828,N_6669);
and U8006 (N_8006,N_6390,N_6067);
nor U8007 (N_8007,N_7269,N_6323);
or U8008 (N_8008,N_6001,N_6084);
or U8009 (N_8009,N_6277,N_6052);
and U8010 (N_8010,N_6329,N_6930);
or U8011 (N_8011,N_6025,N_6480);
or U8012 (N_8012,N_6955,N_7124);
nand U8013 (N_8013,N_7052,N_6557);
or U8014 (N_8014,N_7484,N_6723);
or U8015 (N_8015,N_6582,N_7263);
and U8016 (N_8016,N_6646,N_7154);
or U8017 (N_8017,N_7464,N_6805);
nand U8018 (N_8018,N_6539,N_7196);
nor U8019 (N_8019,N_7120,N_6655);
nand U8020 (N_8020,N_7282,N_6502);
or U8021 (N_8021,N_7224,N_7383);
or U8022 (N_8022,N_6013,N_6996);
xor U8023 (N_8023,N_6852,N_7283);
and U8024 (N_8024,N_6555,N_6511);
and U8025 (N_8025,N_7014,N_6589);
or U8026 (N_8026,N_6796,N_7135);
and U8027 (N_8027,N_6435,N_6427);
nor U8028 (N_8028,N_7343,N_7348);
xnor U8029 (N_8029,N_6220,N_6608);
nand U8030 (N_8030,N_6679,N_6449);
and U8031 (N_8031,N_6918,N_6797);
or U8032 (N_8032,N_6412,N_6668);
and U8033 (N_8033,N_7031,N_6500);
and U8034 (N_8034,N_7270,N_6351);
nand U8035 (N_8035,N_6967,N_6388);
or U8036 (N_8036,N_7169,N_6778);
nor U8037 (N_8037,N_7326,N_6368);
and U8038 (N_8038,N_7328,N_6965);
or U8039 (N_8039,N_6859,N_6408);
or U8040 (N_8040,N_6003,N_6256);
and U8041 (N_8041,N_6496,N_7325);
nor U8042 (N_8042,N_6422,N_6463);
xnor U8043 (N_8043,N_6630,N_6635);
nor U8044 (N_8044,N_6464,N_7099);
or U8045 (N_8045,N_7409,N_6096);
or U8046 (N_8046,N_7231,N_6382);
nor U8047 (N_8047,N_7199,N_6440);
and U8048 (N_8048,N_6634,N_6394);
xor U8049 (N_8049,N_7189,N_6041);
and U8050 (N_8050,N_6994,N_7303);
or U8051 (N_8051,N_6962,N_6736);
or U8052 (N_8052,N_6483,N_6389);
or U8053 (N_8053,N_6458,N_7190);
nor U8054 (N_8054,N_6473,N_6750);
and U8055 (N_8055,N_6699,N_6032);
nor U8056 (N_8056,N_6365,N_7265);
xnor U8057 (N_8057,N_7444,N_6092);
nand U8058 (N_8058,N_7070,N_7212);
nand U8059 (N_8059,N_6370,N_7134);
xor U8060 (N_8060,N_6247,N_7033);
nor U8061 (N_8061,N_6397,N_7132);
nor U8062 (N_8062,N_6802,N_6725);
or U8063 (N_8063,N_6620,N_6331);
or U8064 (N_8064,N_6304,N_6783);
and U8065 (N_8065,N_7080,N_6922);
and U8066 (N_8066,N_6628,N_7206);
nand U8067 (N_8067,N_6307,N_6264);
nand U8068 (N_8068,N_6090,N_6833);
nand U8069 (N_8069,N_7429,N_6362);
nor U8070 (N_8070,N_7493,N_6151);
nand U8071 (N_8071,N_7043,N_7254);
or U8072 (N_8072,N_6775,N_6605);
xor U8073 (N_8073,N_6089,N_6258);
nand U8074 (N_8074,N_6278,N_7436);
or U8075 (N_8075,N_6764,N_6132);
xor U8076 (N_8076,N_6931,N_6217);
nor U8077 (N_8077,N_6035,N_6777);
nand U8078 (N_8078,N_7068,N_6908);
nor U8079 (N_8079,N_6689,N_6865);
or U8080 (N_8080,N_7482,N_7146);
or U8081 (N_8081,N_6168,N_6694);
or U8082 (N_8082,N_6609,N_6744);
nand U8083 (N_8083,N_6120,N_7229);
nand U8084 (N_8084,N_6191,N_7201);
or U8085 (N_8085,N_6169,N_6442);
and U8086 (N_8086,N_6717,N_6506);
nor U8087 (N_8087,N_7402,N_6377);
or U8088 (N_8088,N_7386,N_7256);
nand U8089 (N_8089,N_7420,N_6793);
nand U8090 (N_8090,N_7491,N_6325);
or U8091 (N_8091,N_7151,N_6206);
and U8092 (N_8092,N_6545,N_6857);
xnor U8093 (N_8093,N_7384,N_7001);
nand U8094 (N_8094,N_6376,N_7468);
nor U8095 (N_8095,N_6586,N_6597);
xnor U8096 (N_8096,N_7087,N_6591);
or U8097 (N_8097,N_6549,N_6495);
nand U8098 (N_8098,N_7443,N_7340);
or U8099 (N_8099,N_6590,N_6305);
xor U8100 (N_8100,N_6653,N_6138);
xnor U8101 (N_8101,N_6507,N_6193);
nor U8102 (N_8102,N_6051,N_6969);
xnor U8103 (N_8103,N_7217,N_7163);
nand U8104 (N_8104,N_6239,N_7449);
nand U8105 (N_8105,N_6213,N_7308);
and U8106 (N_8106,N_7305,N_6301);
nand U8107 (N_8107,N_6215,N_6542);
or U8108 (N_8108,N_6227,N_7329);
and U8109 (N_8109,N_7396,N_6026);
and U8110 (N_8110,N_7219,N_7262);
xor U8111 (N_8111,N_6378,N_6838);
and U8112 (N_8112,N_6349,N_6721);
xor U8113 (N_8113,N_7058,N_7316);
nor U8114 (N_8114,N_6534,N_6681);
or U8115 (N_8115,N_6471,N_7359);
nor U8116 (N_8116,N_7401,N_7202);
and U8117 (N_8117,N_6924,N_6621);
or U8118 (N_8118,N_7153,N_6312);
nor U8119 (N_8119,N_6393,N_7020);
nor U8120 (N_8120,N_6901,N_7273);
and U8121 (N_8121,N_7102,N_6339);
nor U8122 (N_8122,N_6267,N_6882);
nand U8123 (N_8123,N_7323,N_6257);
or U8124 (N_8124,N_7499,N_6361);
xor U8125 (N_8125,N_6292,N_6666);
nand U8126 (N_8126,N_7234,N_7222);
nor U8127 (N_8127,N_6790,N_7294);
and U8128 (N_8128,N_6479,N_7218);
nor U8129 (N_8129,N_6280,N_6142);
and U8130 (N_8130,N_6836,N_6126);
or U8131 (N_8131,N_6212,N_6809);
nand U8132 (N_8132,N_7379,N_7187);
nand U8133 (N_8133,N_6441,N_6875);
or U8134 (N_8134,N_6571,N_7039);
or U8135 (N_8135,N_6462,N_6297);
or U8136 (N_8136,N_6568,N_7393);
nand U8137 (N_8137,N_7139,N_6614);
nand U8138 (N_8138,N_6430,N_6004);
and U8139 (N_8139,N_6078,N_6489);
xnor U8140 (N_8140,N_7207,N_6237);
or U8141 (N_8141,N_7488,N_6773);
and U8142 (N_8142,N_6907,N_6391);
nor U8143 (N_8143,N_7377,N_7182);
nand U8144 (N_8144,N_6133,N_6932);
nor U8145 (N_8145,N_6834,N_7267);
nor U8146 (N_8146,N_6337,N_6157);
nor U8147 (N_8147,N_6300,N_7460);
or U8148 (N_8148,N_6334,N_6895);
or U8149 (N_8149,N_6357,N_6006);
nor U8150 (N_8150,N_6077,N_7472);
xnor U8151 (N_8151,N_6547,N_7089);
and U8152 (N_8152,N_6642,N_7435);
nand U8153 (N_8153,N_7437,N_6664);
nor U8154 (N_8154,N_6804,N_7310);
or U8155 (N_8155,N_6340,N_6776);
nor U8156 (N_8156,N_7026,N_6558);
and U8157 (N_8157,N_7145,N_6318);
xnor U8158 (N_8158,N_6565,N_6914);
or U8159 (N_8159,N_6243,N_6824);
or U8160 (N_8160,N_6269,N_7148);
and U8161 (N_8161,N_6732,N_7105);
or U8162 (N_8162,N_7076,N_6949);
nand U8163 (N_8163,N_6481,N_6853);
nor U8164 (N_8164,N_6886,N_6410);
or U8165 (N_8165,N_7425,N_6992);
nor U8166 (N_8166,N_6976,N_7424);
and U8167 (N_8167,N_7450,N_7165);
and U8168 (N_8168,N_7091,N_6180);
or U8169 (N_8169,N_6789,N_7017);
or U8170 (N_8170,N_7445,N_6344);
nand U8171 (N_8171,N_7360,N_6810);
nand U8172 (N_8172,N_6795,N_7116);
or U8173 (N_8173,N_7453,N_7040);
and U8174 (N_8174,N_7079,N_6604);
and U8175 (N_8175,N_6311,N_6100);
and U8176 (N_8176,N_6564,N_7327);
and U8177 (N_8177,N_7370,N_6161);
or U8178 (N_8178,N_6387,N_6380);
nor U8179 (N_8179,N_6235,N_7289);
nor U8180 (N_8180,N_6313,N_7147);
and U8181 (N_8181,N_6127,N_6189);
nor U8182 (N_8182,N_6369,N_6638);
or U8183 (N_8183,N_6285,N_6835);
and U8184 (N_8184,N_6183,N_6333);
and U8185 (N_8185,N_7278,N_6818);
or U8186 (N_8186,N_7251,N_6533);
nor U8187 (N_8187,N_6244,N_7456);
xnor U8188 (N_8188,N_6966,N_6869);
nor U8189 (N_8189,N_6152,N_6184);
nand U8190 (N_8190,N_6572,N_6512);
and U8191 (N_8191,N_6641,N_6036);
or U8192 (N_8192,N_6207,N_6566);
xnor U8193 (N_8193,N_6866,N_6211);
or U8194 (N_8194,N_7227,N_6229);
or U8195 (N_8195,N_6884,N_6106);
nor U8196 (N_8196,N_6648,N_6105);
xor U8197 (N_8197,N_6780,N_6726);
nor U8198 (N_8198,N_7046,N_6954);
and U8199 (N_8199,N_7195,N_6860);
and U8200 (N_8200,N_6588,N_7455);
and U8201 (N_8201,N_6477,N_7027);
or U8202 (N_8202,N_6038,N_6028);
or U8203 (N_8203,N_6898,N_6817);
nor U8204 (N_8204,N_7412,N_6472);
or U8205 (N_8205,N_6867,N_7074);
nor U8206 (N_8206,N_6712,N_7077);
or U8207 (N_8207,N_6079,N_6342);
nor U8208 (N_8208,N_6551,N_6145);
and U8209 (N_8209,N_6017,N_6811);
nor U8210 (N_8210,N_6016,N_6335);
or U8211 (N_8211,N_6950,N_6769);
nand U8212 (N_8212,N_6081,N_6741);
or U8213 (N_8213,N_6294,N_7321);
xor U8214 (N_8214,N_7342,N_7159);
and U8215 (N_8215,N_6527,N_6556);
nor U8216 (N_8216,N_7131,N_7006);
nor U8217 (N_8217,N_7118,N_6347);
xor U8218 (N_8218,N_7211,N_7016);
or U8219 (N_8219,N_6943,N_6039);
and U8220 (N_8220,N_6711,N_7237);
nand U8221 (N_8221,N_7473,N_7075);
and U8222 (N_8222,N_6905,N_6825);
and U8223 (N_8223,N_6658,N_7123);
and U8224 (N_8224,N_6786,N_6877);
and U8225 (N_8225,N_6270,N_6046);
or U8226 (N_8226,N_6102,N_6659);
nand U8227 (N_8227,N_7065,N_6210);
nor U8228 (N_8228,N_6849,N_7149);
nor U8229 (N_8229,N_7235,N_6844);
nand U8230 (N_8230,N_7398,N_6980);
nand U8231 (N_8231,N_6579,N_7186);
nor U8232 (N_8232,N_6201,N_6019);
nand U8233 (N_8233,N_7141,N_6055);
and U8234 (N_8234,N_6425,N_6514);
xor U8235 (N_8235,N_6415,N_7228);
nand U8236 (N_8236,N_6550,N_6840);
and U8237 (N_8237,N_6273,N_7210);
and U8238 (N_8238,N_6146,N_7399);
or U8239 (N_8239,N_7361,N_7239);
or U8240 (N_8240,N_6927,N_6348);
or U8241 (N_8241,N_6265,N_7311);
nand U8242 (N_8242,N_7036,N_7367);
and U8243 (N_8243,N_6842,N_6121);
and U8244 (N_8244,N_7481,N_7297);
xnor U8245 (N_8245,N_6460,N_6692);
or U8246 (N_8246,N_6432,N_6061);
nand U8247 (N_8247,N_6890,N_6738);
nor U8248 (N_8248,N_7387,N_7051);
nor U8249 (N_8249,N_6819,N_6279);
nor U8250 (N_8250,N_7293,N_6791);
and U8251 (N_8251,N_6812,N_6680);
xnor U8252 (N_8252,N_6780,N_7251);
nand U8253 (N_8253,N_6932,N_7474);
nand U8254 (N_8254,N_6098,N_6305);
and U8255 (N_8255,N_7365,N_7237);
or U8256 (N_8256,N_6932,N_6354);
or U8257 (N_8257,N_6168,N_7082);
nand U8258 (N_8258,N_6451,N_6538);
nor U8259 (N_8259,N_7017,N_7311);
xor U8260 (N_8260,N_6674,N_6810);
or U8261 (N_8261,N_6757,N_6913);
nor U8262 (N_8262,N_7021,N_6207);
nor U8263 (N_8263,N_6454,N_7484);
and U8264 (N_8264,N_6203,N_6592);
or U8265 (N_8265,N_6055,N_6626);
nor U8266 (N_8266,N_6269,N_6879);
xnor U8267 (N_8267,N_6962,N_6861);
and U8268 (N_8268,N_6989,N_7356);
nand U8269 (N_8269,N_6065,N_7184);
or U8270 (N_8270,N_6189,N_6549);
and U8271 (N_8271,N_6459,N_7141);
and U8272 (N_8272,N_7029,N_6254);
xnor U8273 (N_8273,N_7121,N_7332);
xor U8274 (N_8274,N_7489,N_7335);
nand U8275 (N_8275,N_7342,N_6995);
nor U8276 (N_8276,N_6058,N_6363);
or U8277 (N_8277,N_6529,N_6576);
nand U8278 (N_8278,N_6223,N_7188);
nor U8279 (N_8279,N_7356,N_6789);
or U8280 (N_8280,N_7069,N_7266);
and U8281 (N_8281,N_6892,N_6931);
nor U8282 (N_8282,N_6023,N_7304);
and U8283 (N_8283,N_6787,N_7295);
and U8284 (N_8284,N_7023,N_7346);
and U8285 (N_8285,N_6711,N_6525);
nand U8286 (N_8286,N_6284,N_7412);
and U8287 (N_8287,N_7326,N_6812);
or U8288 (N_8288,N_7117,N_6386);
and U8289 (N_8289,N_6244,N_6605);
nor U8290 (N_8290,N_7194,N_6567);
nor U8291 (N_8291,N_6366,N_7081);
nand U8292 (N_8292,N_7349,N_7182);
and U8293 (N_8293,N_7058,N_6410);
nor U8294 (N_8294,N_7306,N_6121);
and U8295 (N_8295,N_6220,N_7268);
nand U8296 (N_8296,N_6281,N_7131);
nor U8297 (N_8297,N_6961,N_7013);
or U8298 (N_8298,N_6644,N_6796);
nand U8299 (N_8299,N_6053,N_6780);
nand U8300 (N_8300,N_6423,N_6511);
nor U8301 (N_8301,N_6362,N_6828);
and U8302 (N_8302,N_6711,N_6655);
or U8303 (N_8303,N_7408,N_6322);
nand U8304 (N_8304,N_7321,N_6404);
nand U8305 (N_8305,N_6371,N_7442);
or U8306 (N_8306,N_7335,N_6647);
nor U8307 (N_8307,N_6907,N_6176);
and U8308 (N_8308,N_7304,N_6513);
xor U8309 (N_8309,N_6990,N_6904);
or U8310 (N_8310,N_6456,N_7190);
nor U8311 (N_8311,N_7433,N_7026);
nand U8312 (N_8312,N_7100,N_6597);
or U8313 (N_8313,N_7001,N_6810);
or U8314 (N_8314,N_6440,N_6851);
and U8315 (N_8315,N_6418,N_6127);
nor U8316 (N_8316,N_7211,N_7207);
nand U8317 (N_8317,N_6870,N_6791);
or U8318 (N_8318,N_6039,N_6135);
xor U8319 (N_8319,N_6702,N_7374);
and U8320 (N_8320,N_6970,N_7213);
xnor U8321 (N_8321,N_6608,N_6180);
or U8322 (N_8322,N_6290,N_7147);
and U8323 (N_8323,N_6355,N_7187);
and U8324 (N_8324,N_6804,N_6783);
or U8325 (N_8325,N_6232,N_7337);
or U8326 (N_8326,N_7122,N_6306);
nor U8327 (N_8327,N_7141,N_6355);
and U8328 (N_8328,N_6372,N_7038);
and U8329 (N_8329,N_6432,N_6834);
and U8330 (N_8330,N_6541,N_7421);
and U8331 (N_8331,N_6858,N_6829);
or U8332 (N_8332,N_6833,N_6449);
xnor U8333 (N_8333,N_7314,N_6669);
nor U8334 (N_8334,N_7002,N_6487);
and U8335 (N_8335,N_7481,N_6089);
nand U8336 (N_8336,N_7110,N_6530);
and U8337 (N_8337,N_7038,N_6972);
or U8338 (N_8338,N_6844,N_6520);
nor U8339 (N_8339,N_6560,N_7242);
nor U8340 (N_8340,N_6387,N_6626);
and U8341 (N_8341,N_7284,N_7422);
nor U8342 (N_8342,N_6171,N_6201);
nand U8343 (N_8343,N_6507,N_6757);
nor U8344 (N_8344,N_6943,N_6613);
or U8345 (N_8345,N_6063,N_6809);
nand U8346 (N_8346,N_7186,N_6030);
nor U8347 (N_8347,N_7184,N_6132);
or U8348 (N_8348,N_7038,N_6766);
nand U8349 (N_8349,N_6998,N_7344);
nand U8350 (N_8350,N_6044,N_6505);
nand U8351 (N_8351,N_7256,N_7252);
or U8352 (N_8352,N_6778,N_6221);
nand U8353 (N_8353,N_6973,N_6814);
and U8354 (N_8354,N_6948,N_6151);
nand U8355 (N_8355,N_6517,N_6747);
nor U8356 (N_8356,N_7225,N_7029);
or U8357 (N_8357,N_6945,N_6228);
nor U8358 (N_8358,N_6379,N_6101);
nor U8359 (N_8359,N_7157,N_6907);
xor U8360 (N_8360,N_7475,N_7424);
nor U8361 (N_8361,N_6356,N_7327);
nor U8362 (N_8362,N_7080,N_6212);
and U8363 (N_8363,N_6682,N_7085);
and U8364 (N_8364,N_6872,N_6386);
or U8365 (N_8365,N_7070,N_7483);
nor U8366 (N_8366,N_7422,N_6777);
nor U8367 (N_8367,N_7284,N_7007);
nand U8368 (N_8368,N_7143,N_7040);
nand U8369 (N_8369,N_6982,N_6521);
nand U8370 (N_8370,N_7273,N_6976);
nor U8371 (N_8371,N_6422,N_6304);
nor U8372 (N_8372,N_6172,N_7219);
or U8373 (N_8373,N_7406,N_7104);
or U8374 (N_8374,N_6446,N_6129);
nand U8375 (N_8375,N_6452,N_6442);
nor U8376 (N_8376,N_6490,N_7226);
nor U8377 (N_8377,N_7107,N_6592);
nor U8378 (N_8378,N_7000,N_6240);
and U8379 (N_8379,N_7330,N_6476);
nand U8380 (N_8380,N_6443,N_6976);
and U8381 (N_8381,N_7420,N_6068);
nand U8382 (N_8382,N_7281,N_6264);
nor U8383 (N_8383,N_6032,N_7278);
or U8384 (N_8384,N_7126,N_6644);
nor U8385 (N_8385,N_6943,N_6406);
nor U8386 (N_8386,N_6092,N_6172);
nand U8387 (N_8387,N_6249,N_6335);
or U8388 (N_8388,N_6902,N_6025);
nor U8389 (N_8389,N_7487,N_7414);
or U8390 (N_8390,N_6099,N_6056);
or U8391 (N_8391,N_6028,N_6112);
or U8392 (N_8392,N_6123,N_6647);
and U8393 (N_8393,N_6735,N_6861);
or U8394 (N_8394,N_6704,N_6081);
and U8395 (N_8395,N_6944,N_6137);
nand U8396 (N_8396,N_7209,N_7164);
nor U8397 (N_8397,N_6074,N_7344);
xnor U8398 (N_8398,N_6295,N_6715);
and U8399 (N_8399,N_6960,N_7439);
or U8400 (N_8400,N_6313,N_6154);
nand U8401 (N_8401,N_6405,N_7481);
and U8402 (N_8402,N_6017,N_7352);
or U8403 (N_8403,N_6577,N_6239);
or U8404 (N_8404,N_7288,N_6535);
or U8405 (N_8405,N_7453,N_6257);
xnor U8406 (N_8406,N_6029,N_6064);
nand U8407 (N_8407,N_6909,N_7064);
or U8408 (N_8408,N_6679,N_6490);
nor U8409 (N_8409,N_6844,N_6988);
nor U8410 (N_8410,N_6498,N_6717);
nor U8411 (N_8411,N_7473,N_6646);
nor U8412 (N_8412,N_7139,N_6801);
nand U8413 (N_8413,N_6086,N_7475);
nand U8414 (N_8414,N_6037,N_7011);
or U8415 (N_8415,N_7334,N_6413);
and U8416 (N_8416,N_7360,N_6581);
nand U8417 (N_8417,N_6779,N_6331);
nand U8418 (N_8418,N_6934,N_6595);
nand U8419 (N_8419,N_6656,N_6883);
nand U8420 (N_8420,N_6462,N_6729);
nand U8421 (N_8421,N_6296,N_6302);
nor U8422 (N_8422,N_6929,N_6238);
and U8423 (N_8423,N_6259,N_7227);
nand U8424 (N_8424,N_7150,N_6692);
nor U8425 (N_8425,N_6746,N_7040);
and U8426 (N_8426,N_6628,N_7490);
nand U8427 (N_8427,N_6355,N_6065);
and U8428 (N_8428,N_6844,N_7389);
and U8429 (N_8429,N_7463,N_7255);
nand U8430 (N_8430,N_7240,N_6573);
and U8431 (N_8431,N_6416,N_6720);
nor U8432 (N_8432,N_6765,N_6284);
or U8433 (N_8433,N_6200,N_7226);
nand U8434 (N_8434,N_7456,N_6521);
xor U8435 (N_8435,N_6543,N_7080);
or U8436 (N_8436,N_7360,N_6872);
and U8437 (N_8437,N_7247,N_7308);
and U8438 (N_8438,N_7202,N_6996);
nand U8439 (N_8439,N_6968,N_6217);
and U8440 (N_8440,N_7335,N_6710);
xor U8441 (N_8441,N_6833,N_6519);
or U8442 (N_8442,N_6696,N_7197);
nand U8443 (N_8443,N_7426,N_6470);
and U8444 (N_8444,N_7053,N_7353);
nor U8445 (N_8445,N_7237,N_6127);
or U8446 (N_8446,N_7382,N_6080);
xnor U8447 (N_8447,N_6422,N_6839);
or U8448 (N_8448,N_6886,N_6710);
nor U8449 (N_8449,N_7055,N_6257);
xor U8450 (N_8450,N_7000,N_7208);
nand U8451 (N_8451,N_6545,N_6088);
nor U8452 (N_8452,N_6227,N_6090);
and U8453 (N_8453,N_6644,N_6499);
nand U8454 (N_8454,N_6882,N_6469);
nor U8455 (N_8455,N_6733,N_7484);
nor U8456 (N_8456,N_6424,N_6288);
and U8457 (N_8457,N_6360,N_7069);
nor U8458 (N_8458,N_6069,N_6525);
nand U8459 (N_8459,N_6598,N_6728);
nor U8460 (N_8460,N_7299,N_7013);
xor U8461 (N_8461,N_6680,N_7139);
and U8462 (N_8462,N_6317,N_7003);
nor U8463 (N_8463,N_7037,N_7476);
xor U8464 (N_8464,N_6749,N_6822);
xor U8465 (N_8465,N_6589,N_7253);
nor U8466 (N_8466,N_6132,N_6580);
and U8467 (N_8467,N_6214,N_6933);
xnor U8468 (N_8468,N_6448,N_6280);
nor U8469 (N_8469,N_6707,N_6845);
nor U8470 (N_8470,N_7340,N_6546);
nand U8471 (N_8471,N_7277,N_7028);
nor U8472 (N_8472,N_6407,N_7428);
and U8473 (N_8473,N_6994,N_7015);
nor U8474 (N_8474,N_6661,N_6575);
and U8475 (N_8475,N_6140,N_6338);
or U8476 (N_8476,N_6190,N_6104);
or U8477 (N_8477,N_6443,N_6811);
or U8478 (N_8478,N_7314,N_6224);
nor U8479 (N_8479,N_7156,N_7470);
and U8480 (N_8480,N_6170,N_7357);
or U8481 (N_8481,N_6061,N_7372);
or U8482 (N_8482,N_6182,N_7106);
nor U8483 (N_8483,N_7456,N_7151);
nand U8484 (N_8484,N_6244,N_6145);
nand U8485 (N_8485,N_6466,N_7335);
or U8486 (N_8486,N_6330,N_6796);
nor U8487 (N_8487,N_6253,N_6329);
nor U8488 (N_8488,N_7022,N_7258);
or U8489 (N_8489,N_6132,N_6505);
nor U8490 (N_8490,N_6833,N_6347);
nor U8491 (N_8491,N_6556,N_6351);
xnor U8492 (N_8492,N_7178,N_6327);
nor U8493 (N_8493,N_7477,N_6391);
nor U8494 (N_8494,N_6498,N_7035);
xnor U8495 (N_8495,N_6864,N_6791);
nor U8496 (N_8496,N_6504,N_6097);
and U8497 (N_8497,N_6837,N_6086);
nand U8498 (N_8498,N_7441,N_7382);
and U8499 (N_8499,N_6286,N_7288);
or U8500 (N_8500,N_6291,N_6392);
and U8501 (N_8501,N_6210,N_7161);
nor U8502 (N_8502,N_6130,N_6404);
or U8503 (N_8503,N_6948,N_7339);
or U8504 (N_8504,N_6575,N_7466);
and U8505 (N_8505,N_7467,N_6168);
nor U8506 (N_8506,N_6142,N_7320);
nand U8507 (N_8507,N_6641,N_6751);
and U8508 (N_8508,N_6558,N_6889);
nand U8509 (N_8509,N_6876,N_6243);
nor U8510 (N_8510,N_6347,N_6622);
nor U8511 (N_8511,N_6732,N_6584);
nand U8512 (N_8512,N_6533,N_6669);
nand U8513 (N_8513,N_6799,N_6987);
or U8514 (N_8514,N_6330,N_6140);
or U8515 (N_8515,N_6125,N_7333);
and U8516 (N_8516,N_7117,N_6947);
and U8517 (N_8517,N_7398,N_7157);
and U8518 (N_8518,N_7105,N_7086);
or U8519 (N_8519,N_6568,N_7383);
nand U8520 (N_8520,N_7426,N_7497);
nor U8521 (N_8521,N_7060,N_6299);
nand U8522 (N_8522,N_6432,N_6062);
or U8523 (N_8523,N_7432,N_6422);
nand U8524 (N_8524,N_6985,N_6692);
nand U8525 (N_8525,N_7029,N_6992);
nor U8526 (N_8526,N_7246,N_6935);
nor U8527 (N_8527,N_6029,N_6638);
nand U8528 (N_8528,N_6688,N_7456);
and U8529 (N_8529,N_7467,N_7193);
nand U8530 (N_8530,N_6022,N_7298);
or U8531 (N_8531,N_7431,N_7468);
and U8532 (N_8532,N_6247,N_6765);
or U8533 (N_8533,N_7044,N_6118);
nor U8534 (N_8534,N_6996,N_6524);
and U8535 (N_8535,N_6929,N_6563);
nor U8536 (N_8536,N_6832,N_7230);
or U8537 (N_8537,N_6980,N_6135);
nand U8538 (N_8538,N_6190,N_7342);
nor U8539 (N_8539,N_6853,N_7186);
and U8540 (N_8540,N_7270,N_7134);
and U8541 (N_8541,N_6132,N_7119);
and U8542 (N_8542,N_7081,N_6166);
xnor U8543 (N_8543,N_7280,N_6316);
nor U8544 (N_8544,N_6314,N_6009);
nand U8545 (N_8545,N_7145,N_6185);
nand U8546 (N_8546,N_6696,N_6426);
nor U8547 (N_8547,N_6947,N_6786);
or U8548 (N_8548,N_7472,N_6045);
nand U8549 (N_8549,N_6437,N_6204);
and U8550 (N_8550,N_7373,N_6624);
or U8551 (N_8551,N_6602,N_6001);
or U8552 (N_8552,N_7332,N_6309);
nand U8553 (N_8553,N_6159,N_6552);
nor U8554 (N_8554,N_6111,N_6727);
or U8555 (N_8555,N_6689,N_7424);
or U8556 (N_8556,N_7057,N_6975);
nand U8557 (N_8557,N_7005,N_7399);
xnor U8558 (N_8558,N_7000,N_6615);
and U8559 (N_8559,N_6559,N_6551);
and U8560 (N_8560,N_6532,N_7188);
nand U8561 (N_8561,N_6510,N_6108);
xor U8562 (N_8562,N_7331,N_6459);
nand U8563 (N_8563,N_6488,N_6204);
or U8564 (N_8564,N_6763,N_6755);
and U8565 (N_8565,N_6031,N_7440);
or U8566 (N_8566,N_6882,N_6255);
or U8567 (N_8567,N_6161,N_7181);
or U8568 (N_8568,N_6864,N_6922);
nand U8569 (N_8569,N_6352,N_7394);
or U8570 (N_8570,N_6381,N_6601);
and U8571 (N_8571,N_7262,N_6945);
or U8572 (N_8572,N_6543,N_6483);
and U8573 (N_8573,N_6037,N_6263);
xor U8574 (N_8574,N_6809,N_7069);
or U8575 (N_8575,N_6979,N_7179);
or U8576 (N_8576,N_6519,N_6609);
xnor U8577 (N_8577,N_6124,N_7284);
or U8578 (N_8578,N_6509,N_6778);
and U8579 (N_8579,N_7343,N_6842);
nand U8580 (N_8580,N_6600,N_6944);
nor U8581 (N_8581,N_6146,N_6528);
or U8582 (N_8582,N_6044,N_7209);
nor U8583 (N_8583,N_7435,N_6706);
nand U8584 (N_8584,N_6864,N_6452);
nor U8585 (N_8585,N_6263,N_6570);
and U8586 (N_8586,N_7386,N_6658);
nand U8587 (N_8587,N_6300,N_6138);
nor U8588 (N_8588,N_7440,N_7451);
nand U8589 (N_8589,N_7112,N_6671);
or U8590 (N_8590,N_6969,N_6589);
nand U8591 (N_8591,N_6960,N_7457);
nor U8592 (N_8592,N_6156,N_7044);
nand U8593 (N_8593,N_7174,N_6469);
and U8594 (N_8594,N_6195,N_6252);
nor U8595 (N_8595,N_7251,N_7487);
nand U8596 (N_8596,N_7450,N_6306);
or U8597 (N_8597,N_7023,N_6699);
and U8598 (N_8598,N_6272,N_6247);
or U8599 (N_8599,N_7306,N_7087);
nand U8600 (N_8600,N_6452,N_7162);
and U8601 (N_8601,N_6769,N_6063);
and U8602 (N_8602,N_6814,N_6769);
and U8603 (N_8603,N_7298,N_7062);
nor U8604 (N_8604,N_6302,N_7432);
nand U8605 (N_8605,N_7056,N_6228);
and U8606 (N_8606,N_6839,N_7281);
and U8607 (N_8607,N_6809,N_6659);
nand U8608 (N_8608,N_6325,N_6670);
nand U8609 (N_8609,N_6385,N_7155);
nor U8610 (N_8610,N_6025,N_6939);
and U8611 (N_8611,N_6076,N_6783);
nor U8612 (N_8612,N_6227,N_7149);
and U8613 (N_8613,N_7009,N_6127);
or U8614 (N_8614,N_6269,N_6171);
nand U8615 (N_8615,N_6287,N_7344);
nand U8616 (N_8616,N_7166,N_6971);
or U8617 (N_8617,N_6753,N_7305);
and U8618 (N_8618,N_7198,N_6632);
xnor U8619 (N_8619,N_6551,N_7126);
nor U8620 (N_8620,N_6161,N_6209);
nor U8621 (N_8621,N_6267,N_6801);
and U8622 (N_8622,N_7442,N_7169);
or U8623 (N_8623,N_6960,N_7303);
nand U8624 (N_8624,N_6811,N_7142);
nand U8625 (N_8625,N_6417,N_6690);
and U8626 (N_8626,N_6465,N_6070);
nand U8627 (N_8627,N_6211,N_6101);
xor U8628 (N_8628,N_6618,N_6830);
xor U8629 (N_8629,N_6607,N_6007);
nor U8630 (N_8630,N_6284,N_7330);
and U8631 (N_8631,N_7042,N_6148);
xor U8632 (N_8632,N_6428,N_7351);
or U8633 (N_8633,N_6265,N_7183);
nand U8634 (N_8634,N_7112,N_7200);
and U8635 (N_8635,N_6288,N_6795);
or U8636 (N_8636,N_6029,N_6189);
or U8637 (N_8637,N_7338,N_6900);
and U8638 (N_8638,N_7245,N_6998);
nand U8639 (N_8639,N_6822,N_6661);
or U8640 (N_8640,N_7032,N_6781);
xnor U8641 (N_8641,N_7124,N_7144);
nor U8642 (N_8642,N_7491,N_6219);
and U8643 (N_8643,N_6987,N_7252);
xor U8644 (N_8644,N_6404,N_6525);
or U8645 (N_8645,N_6271,N_7208);
or U8646 (N_8646,N_6730,N_6477);
or U8647 (N_8647,N_6479,N_6493);
or U8648 (N_8648,N_6959,N_6731);
nor U8649 (N_8649,N_6877,N_6466);
xor U8650 (N_8650,N_7083,N_7275);
or U8651 (N_8651,N_6810,N_6138);
nand U8652 (N_8652,N_7352,N_6075);
or U8653 (N_8653,N_6431,N_6118);
and U8654 (N_8654,N_6148,N_6976);
nand U8655 (N_8655,N_6952,N_7319);
nor U8656 (N_8656,N_6710,N_7139);
nor U8657 (N_8657,N_6966,N_6273);
nor U8658 (N_8658,N_7022,N_6314);
and U8659 (N_8659,N_7226,N_6518);
and U8660 (N_8660,N_6043,N_7117);
or U8661 (N_8661,N_7096,N_7444);
or U8662 (N_8662,N_7496,N_6757);
or U8663 (N_8663,N_7179,N_7400);
nand U8664 (N_8664,N_6907,N_7452);
or U8665 (N_8665,N_7412,N_7142);
and U8666 (N_8666,N_7005,N_6068);
and U8667 (N_8667,N_6865,N_6838);
xnor U8668 (N_8668,N_7476,N_6922);
nand U8669 (N_8669,N_6864,N_6084);
nand U8670 (N_8670,N_6585,N_6332);
nor U8671 (N_8671,N_7310,N_6857);
or U8672 (N_8672,N_6087,N_7351);
and U8673 (N_8673,N_6816,N_6494);
xnor U8674 (N_8674,N_7098,N_7285);
nor U8675 (N_8675,N_6083,N_6599);
or U8676 (N_8676,N_7172,N_7128);
or U8677 (N_8677,N_6613,N_7446);
or U8678 (N_8678,N_6998,N_6953);
or U8679 (N_8679,N_6460,N_7491);
nor U8680 (N_8680,N_6250,N_7472);
and U8681 (N_8681,N_7137,N_6330);
nand U8682 (N_8682,N_6092,N_6705);
nand U8683 (N_8683,N_6869,N_6746);
and U8684 (N_8684,N_6570,N_7141);
nand U8685 (N_8685,N_6893,N_7048);
nand U8686 (N_8686,N_7014,N_6874);
and U8687 (N_8687,N_7091,N_6591);
or U8688 (N_8688,N_6482,N_7322);
nand U8689 (N_8689,N_6360,N_6471);
nand U8690 (N_8690,N_7234,N_6617);
or U8691 (N_8691,N_6694,N_6449);
nor U8692 (N_8692,N_6234,N_6643);
xor U8693 (N_8693,N_6434,N_6534);
nand U8694 (N_8694,N_6039,N_7084);
nor U8695 (N_8695,N_7014,N_6110);
nor U8696 (N_8696,N_6665,N_6838);
xor U8697 (N_8697,N_6282,N_7450);
nor U8698 (N_8698,N_7296,N_6275);
nor U8699 (N_8699,N_6363,N_7411);
or U8700 (N_8700,N_6732,N_6564);
or U8701 (N_8701,N_6105,N_6238);
nand U8702 (N_8702,N_6426,N_7350);
nand U8703 (N_8703,N_6031,N_7056);
and U8704 (N_8704,N_6535,N_7299);
xnor U8705 (N_8705,N_6549,N_6469);
or U8706 (N_8706,N_6862,N_6568);
or U8707 (N_8707,N_6993,N_6886);
nor U8708 (N_8708,N_6055,N_6341);
nor U8709 (N_8709,N_6676,N_7225);
nand U8710 (N_8710,N_6646,N_6497);
and U8711 (N_8711,N_6384,N_7258);
and U8712 (N_8712,N_6797,N_7261);
nand U8713 (N_8713,N_6066,N_6009);
and U8714 (N_8714,N_6828,N_6249);
xnor U8715 (N_8715,N_7462,N_6920);
nor U8716 (N_8716,N_6586,N_6433);
nor U8717 (N_8717,N_7243,N_7216);
or U8718 (N_8718,N_6443,N_7019);
nor U8719 (N_8719,N_6428,N_7287);
or U8720 (N_8720,N_6344,N_7414);
xor U8721 (N_8721,N_6490,N_6807);
nor U8722 (N_8722,N_6265,N_6908);
nand U8723 (N_8723,N_6708,N_7499);
xor U8724 (N_8724,N_6068,N_6218);
nor U8725 (N_8725,N_7159,N_7104);
nand U8726 (N_8726,N_6193,N_6217);
or U8727 (N_8727,N_7371,N_6147);
or U8728 (N_8728,N_6939,N_6700);
or U8729 (N_8729,N_7396,N_6873);
nand U8730 (N_8730,N_6426,N_7144);
or U8731 (N_8731,N_7070,N_6803);
and U8732 (N_8732,N_7263,N_6447);
and U8733 (N_8733,N_6177,N_7131);
nor U8734 (N_8734,N_6831,N_7371);
and U8735 (N_8735,N_7487,N_6071);
nor U8736 (N_8736,N_7365,N_6342);
nor U8737 (N_8737,N_6776,N_7290);
nor U8738 (N_8738,N_6600,N_7483);
and U8739 (N_8739,N_6121,N_7456);
or U8740 (N_8740,N_6744,N_7126);
or U8741 (N_8741,N_7248,N_6105);
or U8742 (N_8742,N_6730,N_6258);
nor U8743 (N_8743,N_6275,N_7174);
or U8744 (N_8744,N_6996,N_6573);
or U8745 (N_8745,N_6517,N_7103);
nand U8746 (N_8746,N_7016,N_6721);
nor U8747 (N_8747,N_6519,N_7337);
and U8748 (N_8748,N_6806,N_7389);
or U8749 (N_8749,N_6213,N_6061);
or U8750 (N_8750,N_6083,N_6634);
or U8751 (N_8751,N_6754,N_6670);
xor U8752 (N_8752,N_6148,N_6553);
xor U8753 (N_8753,N_7491,N_6923);
or U8754 (N_8754,N_7342,N_7434);
nand U8755 (N_8755,N_6279,N_7377);
and U8756 (N_8756,N_6964,N_6050);
nand U8757 (N_8757,N_6507,N_6009);
nor U8758 (N_8758,N_6643,N_6644);
nor U8759 (N_8759,N_6919,N_7042);
nand U8760 (N_8760,N_6037,N_6209);
and U8761 (N_8761,N_6051,N_6976);
xnor U8762 (N_8762,N_6209,N_6290);
or U8763 (N_8763,N_6420,N_6573);
nor U8764 (N_8764,N_7087,N_7444);
nand U8765 (N_8765,N_6873,N_7277);
nor U8766 (N_8766,N_7279,N_7489);
nand U8767 (N_8767,N_7151,N_6583);
and U8768 (N_8768,N_6960,N_6853);
and U8769 (N_8769,N_6187,N_6423);
nor U8770 (N_8770,N_6746,N_6301);
and U8771 (N_8771,N_6294,N_6046);
xnor U8772 (N_8772,N_6742,N_7397);
nor U8773 (N_8773,N_6958,N_6671);
nor U8774 (N_8774,N_6249,N_6495);
nand U8775 (N_8775,N_6782,N_7334);
xnor U8776 (N_8776,N_6500,N_7231);
and U8777 (N_8777,N_6285,N_7305);
nor U8778 (N_8778,N_6729,N_7066);
and U8779 (N_8779,N_6477,N_6617);
nor U8780 (N_8780,N_6189,N_7062);
nor U8781 (N_8781,N_6164,N_6702);
and U8782 (N_8782,N_7273,N_6559);
or U8783 (N_8783,N_6638,N_7427);
and U8784 (N_8784,N_6677,N_6495);
nor U8785 (N_8785,N_7057,N_7206);
nand U8786 (N_8786,N_6239,N_6054);
nor U8787 (N_8787,N_6975,N_7073);
nor U8788 (N_8788,N_7454,N_6883);
or U8789 (N_8789,N_6329,N_6618);
nand U8790 (N_8790,N_6976,N_7264);
or U8791 (N_8791,N_6898,N_6859);
nand U8792 (N_8792,N_6367,N_7285);
nand U8793 (N_8793,N_6303,N_6356);
nor U8794 (N_8794,N_7006,N_7327);
or U8795 (N_8795,N_6256,N_6140);
or U8796 (N_8796,N_6588,N_6151);
xnor U8797 (N_8797,N_6652,N_6037);
nor U8798 (N_8798,N_7237,N_7386);
or U8799 (N_8799,N_7007,N_6216);
xnor U8800 (N_8800,N_7128,N_6671);
nand U8801 (N_8801,N_6005,N_6695);
and U8802 (N_8802,N_6550,N_6439);
nand U8803 (N_8803,N_6470,N_6887);
or U8804 (N_8804,N_6443,N_7146);
or U8805 (N_8805,N_6170,N_7098);
xor U8806 (N_8806,N_6346,N_7052);
and U8807 (N_8807,N_7003,N_7429);
nand U8808 (N_8808,N_7201,N_6764);
nor U8809 (N_8809,N_7279,N_6822);
nand U8810 (N_8810,N_7272,N_7216);
and U8811 (N_8811,N_7307,N_7224);
nor U8812 (N_8812,N_7044,N_6393);
or U8813 (N_8813,N_6562,N_7375);
nand U8814 (N_8814,N_6321,N_6706);
and U8815 (N_8815,N_7328,N_6529);
xnor U8816 (N_8816,N_7075,N_7153);
and U8817 (N_8817,N_7060,N_6432);
nor U8818 (N_8818,N_6581,N_6444);
nand U8819 (N_8819,N_6137,N_7278);
nand U8820 (N_8820,N_6942,N_6607);
and U8821 (N_8821,N_6678,N_6189);
nor U8822 (N_8822,N_6307,N_6315);
xor U8823 (N_8823,N_6469,N_6132);
nor U8824 (N_8824,N_6005,N_6775);
nand U8825 (N_8825,N_7272,N_6025);
nand U8826 (N_8826,N_6485,N_6038);
and U8827 (N_8827,N_6761,N_6676);
or U8828 (N_8828,N_6163,N_6288);
nand U8829 (N_8829,N_7217,N_7086);
or U8830 (N_8830,N_7472,N_7112);
or U8831 (N_8831,N_6449,N_6728);
and U8832 (N_8832,N_6461,N_6361);
nand U8833 (N_8833,N_6736,N_6934);
nor U8834 (N_8834,N_6511,N_6926);
nand U8835 (N_8835,N_6788,N_6685);
xnor U8836 (N_8836,N_6930,N_7137);
nand U8837 (N_8837,N_6156,N_6784);
or U8838 (N_8838,N_6766,N_6829);
xor U8839 (N_8839,N_6860,N_6339);
nor U8840 (N_8840,N_7267,N_6777);
nor U8841 (N_8841,N_6043,N_6235);
nor U8842 (N_8842,N_6195,N_7179);
and U8843 (N_8843,N_6558,N_6131);
nor U8844 (N_8844,N_6492,N_6677);
and U8845 (N_8845,N_6002,N_6734);
nand U8846 (N_8846,N_6966,N_7299);
nor U8847 (N_8847,N_6015,N_6294);
nand U8848 (N_8848,N_7028,N_6947);
and U8849 (N_8849,N_7087,N_6938);
or U8850 (N_8850,N_7368,N_6742);
and U8851 (N_8851,N_6615,N_7179);
and U8852 (N_8852,N_7326,N_6548);
nand U8853 (N_8853,N_7468,N_6181);
nand U8854 (N_8854,N_6927,N_6015);
xnor U8855 (N_8855,N_7130,N_6733);
xor U8856 (N_8856,N_6787,N_6574);
or U8857 (N_8857,N_7286,N_6794);
xor U8858 (N_8858,N_6489,N_7179);
nor U8859 (N_8859,N_7055,N_7174);
and U8860 (N_8860,N_6144,N_6400);
nand U8861 (N_8861,N_7261,N_7243);
nor U8862 (N_8862,N_7329,N_6961);
nor U8863 (N_8863,N_6762,N_7002);
and U8864 (N_8864,N_7375,N_7479);
nor U8865 (N_8865,N_6938,N_7450);
or U8866 (N_8866,N_6180,N_6068);
and U8867 (N_8867,N_6288,N_6534);
or U8868 (N_8868,N_7432,N_6387);
or U8869 (N_8869,N_6955,N_6800);
and U8870 (N_8870,N_6936,N_6670);
nand U8871 (N_8871,N_6811,N_6668);
and U8872 (N_8872,N_6323,N_6575);
nand U8873 (N_8873,N_6275,N_7104);
nand U8874 (N_8874,N_7427,N_6081);
nand U8875 (N_8875,N_7112,N_6330);
or U8876 (N_8876,N_7038,N_6161);
and U8877 (N_8877,N_6918,N_6381);
or U8878 (N_8878,N_6046,N_6574);
and U8879 (N_8879,N_6368,N_6541);
nand U8880 (N_8880,N_7169,N_6759);
xnor U8881 (N_8881,N_7089,N_7222);
or U8882 (N_8882,N_6685,N_6454);
or U8883 (N_8883,N_6438,N_6352);
nor U8884 (N_8884,N_6985,N_7408);
nand U8885 (N_8885,N_6255,N_6726);
xnor U8886 (N_8886,N_6031,N_6119);
and U8887 (N_8887,N_6758,N_6150);
xnor U8888 (N_8888,N_6204,N_7475);
or U8889 (N_8889,N_6495,N_6818);
nor U8890 (N_8890,N_6495,N_6486);
or U8891 (N_8891,N_7259,N_6177);
and U8892 (N_8892,N_6552,N_7253);
nand U8893 (N_8893,N_6411,N_6146);
nor U8894 (N_8894,N_7453,N_6597);
or U8895 (N_8895,N_7310,N_7168);
or U8896 (N_8896,N_7261,N_6291);
and U8897 (N_8897,N_7096,N_6665);
or U8898 (N_8898,N_7238,N_7437);
and U8899 (N_8899,N_7342,N_7073);
or U8900 (N_8900,N_6386,N_6037);
or U8901 (N_8901,N_7499,N_6823);
or U8902 (N_8902,N_6827,N_7277);
and U8903 (N_8903,N_6649,N_7012);
xor U8904 (N_8904,N_7321,N_7007);
and U8905 (N_8905,N_7212,N_6083);
or U8906 (N_8906,N_6487,N_6418);
xnor U8907 (N_8907,N_7129,N_6570);
and U8908 (N_8908,N_6726,N_6730);
nor U8909 (N_8909,N_6857,N_6163);
nand U8910 (N_8910,N_6743,N_6276);
and U8911 (N_8911,N_7445,N_7077);
xnor U8912 (N_8912,N_6442,N_7111);
nor U8913 (N_8913,N_6833,N_6465);
nand U8914 (N_8914,N_7039,N_6803);
nand U8915 (N_8915,N_6385,N_6682);
or U8916 (N_8916,N_7417,N_7159);
nand U8917 (N_8917,N_6984,N_6411);
and U8918 (N_8918,N_6999,N_6113);
or U8919 (N_8919,N_6030,N_7046);
nor U8920 (N_8920,N_6401,N_6493);
nor U8921 (N_8921,N_6413,N_6172);
or U8922 (N_8922,N_6208,N_7015);
and U8923 (N_8923,N_7487,N_6737);
or U8924 (N_8924,N_6520,N_6158);
nor U8925 (N_8925,N_6106,N_6621);
or U8926 (N_8926,N_6493,N_7020);
nand U8927 (N_8927,N_7216,N_6661);
xor U8928 (N_8928,N_6695,N_6263);
nor U8929 (N_8929,N_6446,N_7196);
nand U8930 (N_8930,N_7388,N_6836);
nor U8931 (N_8931,N_6437,N_6929);
nand U8932 (N_8932,N_7158,N_6687);
or U8933 (N_8933,N_6163,N_6794);
and U8934 (N_8934,N_6103,N_6673);
or U8935 (N_8935,N_6466,N_6003);
and U8936 (N_8936,N_6424,N_7283);
nor U8937 (N_8937,N_6802,N_6871);
xor U8938 (N_8938,N_6922,N_6144);
nand U8939 (N_8939,N_7370,N_7299);
and U8940 (N_8940,N_7109,N_7189);
or U8941 (N_8941,N_6269,N_6552);
nor U8942 (N_8942,N_6773,N_6275);
nor U8943 (N_8943,N_6174,N_6885);
nor U8944 (N_8944,N_6103,N_6449);
nand U8945 (N_8945,N_6392,N_7458);
or U8946 (N_8946,N_6726,N_6794);
or U8947 (N_8947,N_7264,N_6226);
nand U8948 (N_8948,N_6588,N_7362);
nor U8949 (N_8949,N_7396,N_6149);
or U8950 (N_8950,N_7436,N_7382);
xor U8951 (N_8951,N_6591,N_7191);
and U8952 (N_8952,N_6721,N_6637);
nor U8953 (N_8953,N_6690,N_6452);
or U8954 (N_8954,N_6873,N_6232);
nand U8955 (N_8955,N_6692,N_6690);
nand U8956 (N_8956,N_6783,N_7200);
and U8957 (N_8957,N_6056,N_6367);
or U8958 (N_8958,N_7208,N_6613);
nand U8959 (N_8959,N_6472,N_7155);
and U8960 (N_8960,N_7417,N_6390);
nor U8961 (N_8961,N_7190,N_7015);
and U8962 (N_8962,N_6848,N_6881);
and U8963 (N_8963,N_6283,N_7183);
and U8964 (N_8964,N_7035,N_6064);
and U8965 (N_8965,N_7238,N_6595);
and U8966 (N_8966,N_6429,N_7020);
xor U8967 (N_8967,N_6525,N_7388);
nand U8968 (N_8968,N_6032,N_6536);
nand U8969 (N_8969,N_6538,N_6592);
nand U8970 (N_8970,N_7377,N_6839);
nand U8971 (N_8971,N_6814,N_6670);
xor U8972 (N_8972,N_7301,N_6085);
or U8973 (N_8973,N_6028,N_6133);
and U8974 (N_8974,N_6965,N_7419);
nor U8975 (N_8975,N_6347,N_6025);
and U8976 (N_8976,N_6040,N_6018);
or U8977 (N_8977,N_6516,N_7022);
nor U8978 (N_8978,N_6208,N_6311);
and U8979 (N_8979,N_6485,N_6455);
or U8980 (N_8980,N_6001,N_6439);
and U8981 (N_8981,N_7384,N_6325);
or U8982 (N_8982,N_7180,N_7494);
or U8983 (N_8983,N_6772,N_6364);
and U8984 (N_8984,N_6278,N_6680);
and U8985 (N_8985,N_6211,N_6059);
or U8986 (N_8986,N_6727,N_7290);
xor U8987 (N_8987,N_6522,N_7225);
nand U8988 (N_8988,N_7004,N_6759);
or U8989 (N_8989,N_7099,N_6638);
nor U8990 (N_8990,N_6798,N_7462);
and U8991 (N_8991,N_7094,N_6532);
and U8992 (N_8992,N_7132,N_7239);
nor U8993 (N_8993,N_6162,N_6530);
xnor U8994 (N_8994,N_7495,N_6342);
xor U8995 (N_8995,N_6801,N_7238);
and U8996 (N_8996,N_6863,N_6430);
nor U8997 (N_8997,N_6243,N_7009);
and U8998 (N_8998,N_6244,N_6553);
or U8999 (N_8999,N_6944,N_6529);
nand U9000 (N_9000,N_8847,N_8901);
nor U9001 (N_9001,N_8304,N_8657);
xnor U9002 (N_9002,N_8969,N_8573);
xnor U9003 (N_9003,N_8717,N_8272);
nand U9004 (N_9004,N_8312,N_8943);
or U9005 (N_9005,N_8523,N_7852);
and U9006 (N_9006,N_7970,N_8986);
or U9007 (N_9007,N_8331,N_7542);
nor U9008 (N_9008,N_8037,N_7574);
nand U9009 (N_9009,N_8200,N_8402);
xnor U9010 (N_9010,N_8317,N_8359);
nand U9011 (N_9011,N_8622,N_8192);
and U9012 (N_9012,N_7725,N_8298);
and U9013 (N_9013,N_8881,N_7677);
or U9014 (N_9014,N_8821,N_7810);
or U9015 (N_9015,N_8929,N_7534);
nand U9016 (N_9016,N_7536,N_7906);
nor U9017 (N_9017,N_7535,N_7537);
and U9018 (N_9018,N_7638,N_8062);
nand U9019 (N_9019,N_8020,N_8355);
nand U9020 (N_9020,N_8188,N_8285);
or U9021 (N_9021,N_7885,N_7686);
and U9022 (N_9022,N_8341,N_7629);
nor U9023 (N_9023,N_7606,N_8547);
and U9024 (N_9024,N_7901,N_8320);
xor U9025 (N_9025,N_8809,N_7708);
nand U9026 (N_9026,N_8505,N_8787);
or U9027 (N_9027,N_7648,N_7655);
or U9028 (N_9028,N_8759,N_7914);
xnor U9029 (N_9029,N_7526,N_8146);
nor U9030 (N_9030,N_8437,N_7944);
or U9031 (N_9031,N_7531,N_8159);
and U9032 (N_9032,N_7704,N_8665);
and U9033 (N_9033,N_8870,N_7987);
xor U9034 (N_9034,N_7821,N_8125);
nand U9035 (N_9035,N_8052,N_8281);
or U9036 (N_9036,N_7774,N_8956);
and U9037 (N_9037,N_8963,N_8033);
and U9038 (N_9038,N_8395,N_8598);
nor U9039 (N_9039,N_7501,N_8132);
nand U9040 (N_9040,N_8295,N_8543);
or U9041 (N_9041,N_8512,N_7862);
nor U9042 (N_9042,N_7771,N_8330);
nand U9043 (N_9043,N_8376,N_7886);
or U9044 (N_9044,N_8303,N_7660);
or U9045 (N_9045,N_7718,N_8444);
nand U9046 (N_9046,N_8055,N_8568);
and U9047 (N_9047,N_7520,N_8154);
or U9048 (N_9048,N_8264,N_8038);
or U9049 (N_9049,N_8096,N_7833);
or U9050 (N_9050,N_8633,N_8489);
and U9051 (N_9051,N_8643,N_8750);
nand U9052 (N_9052,N_7637,N_8930);
nand U9053 (N_9053,N_8455,N_8953);
nand U9054 (N_9054,N_8228,N_8701);
nor U9055 (N_9055,N_8250,N_7974);
nand U9056 (N_9056,N_8648,N_8908);
nand U9057 (N_9057,N_8808,N_8994);
and U9058 (N_9058,N_7892,N_8528);
nor U9059 (N_9059,N_8388,N_8110);
and U9060 (N_9060,N_7891,N_8619);
and U9061 (N_9061,N_8190,N_8689);
or U9062 (N_9062,N_8253,N_7767);
and U9063 (N_9063,N_8477,N_8466);
and U9064 (N_9064,N_8269,N_7807);
nor U9065 (N_9065,N_7759,N_8906);
xnor U9066 (N_9066,N_8004,N_7935);
nor U9067 (N_9067,N_8191,N_8117);
nor U9068 (N_9068,N_7750,N_8488);
nor U9069 (N_9069,N_8168,N_7888);
xnor U9070 (N_9070,N_8555,N_8197);
or U9071 (N_9071,N_8060,N_8240);
nor U9072 (N_9072,N_7741,N_8058);
or U9073 (N_9073,N_7973,N_8100);
or U9074 (N_9074,N_8121,N_8671);
nand U9075 (N_9075,N_8591,N_8091);
nand U9076 (N_9076,N_7634,N_8327);
nor U9077 (N_9077,N_8995,N_8283);
or U9078 (N_9078,N_8570,N_7972);
and U9079 (N_9079,N_7978,N_7786);
nor U9080 (N_9080,N_8583,N_7778);
and U9081 (N_9081,N_8845,N_8380);
or U9082 (N_9082,N_8438,N_8003);
nand U9083 (N_9083,N_7919,N_8127);
or U9084 (N_9084,N_8765,N_8844);
nand U9085 (N_9085,N_8079,N_8075);
or U9086 (N_9086,N_7632,N_8469);
and U9087 (N_9087,N_7670,N_8928);
xor U9088 (N_9088,N_7986,N_7793);
and U9089 (N_9089,N_8763,N_7685);
nand U9090 (N_9090,N_8500,N_8603);
xnor U9091 (N_9091,N_7755,N_7934);
or U9092 (N_9092,N_8369,N_8288);
xnor U9093 (N_9093,N_7905,N_8138);
xor U9094 (N_9094,N_8397,N_7931);
or U9095 (N_9095,N_8920,N_8804);
xnor U9096 (N_9096,N_8467,N_7925);
and U9097 (N_9097,N_8178,N_8034);
and U9098 (N_9098,N_7761,N_7819);
and U9099 (N_9099,N_8051,N_8365);
or U9100 (N_9100,N_8954,N_7969);
or U9101 (N_9101,N_7651,N_8483);
nand U9102 (N_9102,N_8268,N_8875);
and U9103 (N_9103,N_7770,N_7752);
nand U9104 (N_9104,N_8925,N_7625);
nor U9105 (N_9105,N_7626,N_8452);
nor U9106 (N_9106,N_8278,N_8066);
and U9107 (N_9107,N_8704,N_7666);
nand U9108 (N_9108,N_8795,N_8105);
nor U9109 (N_9109,N_8522,N_7932);
nand U9110 (N_9110,N_7917,N_8056);
and U9111 (N_9111,N_8923,N_7581);
or U9112 (N_9112,N_8384,N_7853);
nand U9113 (N_9113,N_8892,N_8927);
xor U9114 (N_9114,N_7541,N_7850);
nor U9115 (N_9115,N_8459,N_7736);
nor U9116 (N_9116,N_7559,N_7904);
nand U9117 (N_9117,N_7717,N_7524);
nor U9118 (N_9118,N_8625,N_8830);
and U9119 (N_9119,N_8128,N_8499);
nand U9120 (N_9120,N_8349,N_7509);
nand U9121 (N_9121,N_7802,N_7869);
or U9122 (N_9122,N_8102,N_8694);
nand U9123 (N_9123,N_8107,N_7769);
or U9124 (N_9124,N_8358,N_8019);
and U9125 (N_9125,N_8968,N_8556);
nand U9126 (N_9126,N_8760,N_8866);
xor U9127 (N_9127,N_7539,N_7765);
or U9128 (N_9128,N_7933,N_8008);
nand U9129 (N_9129,N_8777,N_7735);
nand U9130 (N_9130,N_8013,N_8548);
nand U9131 (N_9131,N_8000,N_8964);
nor U9132 (N_9132,N_7893,N_8940);
nor U9133 (N_9133,N_8860,N_7936);
xor U9134 (N_9134,N_8362,N_7701);
nor U9135 (N_9135,N_7720,N_8494);
nand U9136 (N_9136,N_7857,N_8204);
or U9137 (N_9137,N_8862,N_8451);
or U9138 (N_9138,N_7507,N_8259);
or U9139 (N_9139,N_8205,N_8685);
xor U9140 (N_9140,N_8106,N_7879);
nor U9141 (N_9141,N_8753,N_7903);
nor U9142 (N_9142,N_8602,N_8471);
nor U9143 (N_9143,N_8502,N_8069);
xnor U9144 (N_9144,N_7827,N_8217);
nor U9145 (N_9145,N_8779,N_7510);
or U9146 (N_9146,N_8890,N_8315);
nor U9147 (N_9147,N_8719,N_8552);
nand U9148 (N_9148,N_8219,N_8254);
and U9149 (N_9149,N_8708,N_7522);
nor U9150 (N_9150,N_8767,N_8850);
or U9151 (N_9151,N_8218,N_8799);
xor U9152 (N_9152,N_8492,N_8705);
or U9153 (N_9153,N_8367,N_7836);
or U9154 (N_9154,N_8271,N_8011);
nor U9155 (N_9155,N_8449,N_7839);
or U9156 (N_9156,N_8042,N_8423);
and U9157 (N_9157,N_7943,N_8101);
nor U9158 (N_9158,N_8357,N_7881);
nor U9159 (N_9159,N_7992,N_7550);
nand U9160 (N_9160,N_8952,N_7907);
nand U9161 (N_9161,N_7826,N_8237);
nor U9162 (N_9162,N_8922,N_8354);
and U9163 (N_9163,N_7820,N_7876);
and U9164 (N_9164,N_7920,N_7797);
or U9165 (N_9165,N_8793,N_8841);
nand U9166 (N_9166,N_7645,N_8581);
nor U9167 (N_9167,N_7835,N_8856);
or U9168 (N_9168,N_7598,N_8433);
or U9169 (N_9169,N_8720,N_8699);
xnor U9170 (N_9170,N_7560,N_7815);
nand U9171 (N_9171,N_8420,N_8261);
and U9172 (N_9172,N_8672,N_8674);
or U9173 (N_9173,N_7681,N_8061);
and U9174 (N_9174,N_8709,N_7829);
nand U9175 (N_9175,N_8692,N_7587);
nand U9176 (N_9176,N_7982,N_7832);
nor U9177 (N_9177,N_7529,N_7723);
or U9178 (N_9178,N_8835,N_7856);
nand U9179 (N_9179,N_8186,N_8958);
and U9180 (N_9180,N_8122,N_7831);
nand U9181 (N_9181,N_8863,N_8136);
and U9182 (N_9182,N_7923,N_8415);
nand U9183 (N_9183,N_8604,N_8612);
nand U9184 (N_9184,N_8877,N_8734);
nand U9185 (N_9185,N_8649,N_8081);
and U9186 (N_9186,N_8053,N_7552);
and U9187 (N_9187,N_8089,N_7887);
and U9188 (N_9188,N_8335,N_7727);
and U9189 (N_9189,N_7910,N_8072);
or U9190 (N_9190,N_8093,N_7947);
xor U9191 (N_9191,N_7956,N_8025);
nand U9192 (N_9192,N_8700,N_7711);
and U9193 (N_9193,N_8112,N_8421);
nand U9194 (N_9194,N_8487,N_8479);
nand U9195 (N_9195,N_8326,N_8124);
nor U9196 (N_9196,N_8696,N_8002);
nand U9197 (N_9197,N_7571,N_8833);
and U9198 (N_9198,N_7859,N_7898);
nand U9199 (N_9199,N_8913,N_8539);
and U9200 (N_9200,N_8411,N_7551);
xor U9201 (N_9201,N_8748,N_8059);
or U9202 (N_9202,N_8414,N_7580);
or U9203 (N_9203,N_8565,N_8615);
or U9204 (N_9204,N_8328,N_8917);
xor U9205 (N_9205,N_8747,N_8214);
and U9206 (N_9206,N_8594,N_8791);
nand U9207 (N_9207,N_8230,N_8507);
nor U9208 (N_9208,N_8084,N_8686);
nor U9209 (N_9209,N_8029,N_7692);
and U9210 (N_9210,N_7716,N_8758);
and U9211 (N_9211,N_8683,N_8756);
or U9212 (N_9212,N_8316,N_8088);
and U9213 (N_9213,N_8050,N_7873);
nand U9214 (N_9214,N_8246,N_8664);
nand U9215 (N_9215,N_8839,N_8973);
or U9216 (N_9216,N_7705,N_8211);
nand U9217 (N_9217,N_8776,N_8695);
nand U9218 (N_9218,N_7937,N_8386);
and U9219 (N_9219,N_7738,N_8650);
and U9220 (N_9220,N_8157,N_8441);
or U9221 (N_9221,N_7816,N_8291);
nand U9222 (N_9222,N_8065,N_8557);
nand U9223 (N_9223,N_8546,N_8836);
or U9224 (N_9224,N_7694,N_7766);
nand U9225 (N_9225,N_8475,N_7709);
or U9226 (N_9226,N_8524,N_8823);
and U9227 (N_9227,N_8992,N_7942);
nor U9228 (N_9228,N_8681,N_8577);
or U9229 (N_9229,N_8242,N_7683);
and U9230 (N_9230,N_7792,N_8595);
nor U9231 (N_9231,N_7985,N_7525);
and U9232 (N_9232,N_8854,N_7991);
xnor U9233 (N_9233,N_8235,N_8852);
or U9234 (N_9234,N_8610,N_8653);
nor U9235 (N_9235,N_7607,N_7722);
nor U9236 (N_9236,N_8282,N_7960);
nor U9237 (N_9237,N_8169,N_8858);
nor U9238 (N_9238,N_8585,N_8810);
nand U9239 (N_9239,N_8608,N_8983);
nand U9240 (N_9240,N_7511,N_7739);
nor U9241 (N_9241,N_8279,N_8529);
or U9242 (N_9242,N_7633,N_8745);
and U9243 (N_9243,N_8885,N_7502);
and U9244 (N_9244,N_8794,N_8912);
and U9245 (N_9245,N_8934,N_7673);
nand U9246 (N_9246,N_8593,N_7562);
or U9247 (N_9247,N_8655,N_8231);
nand U9248 (N_9248,N_7854,N_7871);
xnor U9249 (N_9249,N_8307,N_8490);
nand U9250 (N_9250,N_8520,N_8652);
nor U9251 (N_9251,N_7631,N_8373);
nand U9252 (N_9252,N_8582,N_8975);
nor U9253 (N_9253,N_7546,N_7715);
or U9254 (N_9254,N_8015,N_8381);
nand U9255 (N_9255,N_8183,N_7719);
nand U9256 (N_9256,N_8044,N_8751);
or U9257 (N_9257,N_8238,N_8972);
nand U9258 (N_9258,N_7957,N_8959);
and U9259 (N_9259,N_7706,N_7671);
nand U9260 (N_9260,N_7744,N_7691);
nand U9261 (N_9261,N_8811,N_7884);
or U9262 (N_9262,N_8123,N_8871);
nor U9263 (N_9263,N_8864,N_7659);
and U9264 (N_9264,N_8097,N_8187);
or U9265 (N_9265,N_7866,N_8996);
nand U9266 (N_9266,N_7830,N_8396);
nand U9267 (N_9267,N_8372,N_8919);
nor U9268 (N_9268,N_8976,N_8142);
and U9269 (N_9269,N_8347,N_8173);
or U9270 (N_9270,N_8208,N_7808);
and U9271 (N_9271,N_7773,N_7777);
or U9272 (N_9272,N_7877,N_8970);
xor U9273 (N_9273,N_8436,N_8553);
nor U9274 (N_9274,N_8742,N_8504);
or U9275 (N_9275,N_8580,N_8609);
nand U9276 (N_9276,N_8736,N_8399);
and U9277 (N_9277,N_8550,N_8155);
and U9278 (N_9278,N_8910,N_8878);
nor U9279 (N_9279,N_7663,N_8812);
and U9280 (N_9280,N_7599,N_8829);
and U9281 (N_9281,N_8629,N_8345);
nor U9282 (N_9282,N_8394,N_7747);
xnor U9283 (N_9283,N_8137,N_7557);
nor U9284 (N_9284,N_8193,N_8990);
nor U9285 (N_9285,N_8453,N_8531);
and U9286 (N_9286,N_8009,N_7732);
nand U9287 (N_9287,N_8232,N_7864);
xor U9288 (N_9288,N_8879,N_7803);
nand U9289 (N_9289,N_8431,N_7601);
nand U9290 (N_9290,N_8070,N_7712);
and U9291 (N_9291,N_7851,N_8201);
or U9292 (N_9292,N_7868,N_7966);
and U9293 (N_9293,N_8040,N_8403);
and U9294 (N_9294,N_8073,N_8658);
nor U9295 (N_9295,N_8480,N_8196);
nand U9296 (N_9296,N_8905,N_8109);
xor U9297 (N_9297,N_8813,N_8209);
nor U9298 (N_9298,N_8549,N_8014);
nor U9299 (N_9299,N_8946,N_7883);
xor U9300 (N_9300,N_7682,N_8560);
nand U9301 (N_9301,N_8405,N_8497);
nand U9302 (N_9302,N_7624,N_7584);
or U9303 (N_9303,N_8636,N_8458);
xor U9304 (N_9304,N_8509,N_8325);
nor U9305 (N_9305,N_8306,N_8202);
and U9306 (N_9306,N_8443,N_8997);
nand U9307 (N_9307,N_8321,N_7999);
or U9308 (N_9308,N_8045,N_8590);
or U9309 (N_9309,N_7971,N_7724);
or U9310 (N_9310,N_7809,N_8739);
and U9311 (N_9311,N_8318,N_7800);
or U9312 (N_9312,N_8139,N_8016);
xnor U9313 (N_9313,N_8496,N_8574);
nand U9314 (N_9314,N_7870,N_8099);
or U9315 (N_9315,N_8998,N_7505);
xor U9316 (N_9316,N_8936,N_7979);
or U9317 (N_9317,N_8297,N_8094);
or U9318 (N_9318,N_7515,N_7726);
nor U9319 (N_9319,N_7913,N_8244);
or U9320 (N_9320,N_7635,N_8656);
or U9321 (N_9321,N_8290,N_7961);
nor U9322 (N_9322,N_7556,N_7592);
or U9323 (N_9323,N_8018,N_8544);
and U9324 (N_9324,N_8150,N_8894);
and U9325 (N_9325,N_7849,N_7647);
nor U9326 (N_9326,N_8407,N_8351);
or U9327 (N_9327,N_8374,N_8572);
nand U9328 (N_9328,N_8266,N_7713);
or U9329 (N_9329,N_8095,N_8401);
or U9330 (N_9330,N_8951,N_7642);
or U9331 (N_9331,N_8666,N_7938);
and U9332 (N_9332,N_8041,N_8597);
nand U9333 (N_9333,N_7748,N_7728);
and U9334 (N_9334,N_7861,N_8735);
or U9335 (N_9335,N_8985,N_7523);
and U9336 (N_9336,N_8966,N_8145);
xor U9337 (N_9337,N_7566,N_8076);
or U9338 (N_9338,N_8571,N_8815);
and U9339 (N_9339,N_8378,N_8530);
or U9340 (N_9340,N_8513,N_7699);
nor U9341 (N_9341,N_7997,N_7841);
or U9342 (N_9342,N_8886,N_8967);
or U9343 (N_9343,N_8662,N_7605);
nor U9344 (N_9344,N_8714,N_8828);
or U9345 (N_9345,N_8979,N_7890);
nor U9346 (N_9346,N_8224,N_8898);
nor U9347 (N_9347,N_8043,N_8797);
nand U9348 (N_9348,N_8617,N_8769);
nor U9349 (N_9349,N_8485,N_8732);
and U9350 (N_9350,N_8177,N_8086);
nand U9351 (N_9351,N_8284,N_7763);
and U9352 (N_9352,N_8605,N_8252);
nand U9353 (N_9353,N_7989,N_8439);
nor U9354 (N_9354,N_7619,N_8090);
nand U9355 (N_9355,N_8780,N_8684);
and U9356 (N_9356,N_8788,N_7731);
and U9357 (N_9357,N_8948,N_8949);
nand U9358 (N_9358,N_7964,N_8537);
nand U9359 (N_9359,N_7990,N_8820);
nor U9360 (N_9360,N_8682,N_8350);
nand U9361 (N_9361,N_8887,N_8801);
or U9362 (N_9362,N_8554,N_7949);
and U9363 (N_9363,N_8036,N_8434);
and U9364 (N_9364,N_7532,N_7780);
or U9365 (N_9365,N_7799,N_8425);
nand U9366 (N_9366,N_8771,N_8816);
and U9367 (N_9367,N_7993,N_7618);
and U9368 (N_9368,N_8118,N_8346);
or U9369 (N_9369,N_7698,N_7794);
nor U9370 (N_9370,N_8363,N_7615);
nand U9371 (N_9371,N_8868,N_8032);
and U9372 (N_9372,N_8233,N_7959);
or U9373 (N_9373,N_8115,N_8586);
xnor U9374 (N_9374,N_8368,N_7994);
nor U9375 (N_9375,N_8057,N_7512);
or U9376 (N_9376,N_7753,N_7593);
nor U9377 (N_9377,N_8891,N_8849);
nor U9378 (N_9378,N_8203,N_8762);
or U9379 (N_9379,N_8371,N_8616);
and U9380 (N_9380,N_7653,N_7656);
and U9381 (N_9381,N_8063,N_8023);
nor U9382 (N_9382,N_8098,N_8382);
xor U9383 (N_9383,N_8731,N_8077);
xnor U9384 (N_9384,N_8404,N_8566);
or U9385 (N_9385,N_8915,N_8960);
or U9386 (N_9386,N_8716,N_7782);
nand U9387 (N_9387,N_8468,N_7614);
or U9388 (N_9388,N_7958,N_8718);
nor U9389 (N_9389,N_8153,N_8024);
nor U9390 (N_9390,N_8006,N_7760);
or U9391 (N_9391,N_7843,N_8432);
and U9392 (N_9392,N_8733,N_7621);
or U9393 (N_9393,N_8725,N_8781);
nand U9394 (N_9394,N_8085,N_8635);
or U9395 (N_9395,N_8932,N_8755);
or U9396 (N_9396,N_7757,N_8324);
or U9397 (N_9397,N_8171,N_8962);
nand U9398 (N_9398,N_7838,N_8339);
or U9399 (N_9399,N_8133,N_7733);
nand U9400 (N_9400,N_7847,N_8921);
or U9401 (N_9401,N_8838,N_7880);
and U9402 (N_9402,N_7825,N_8867);
and U9403 (N_9403,N_7894,N_8379);
and U9404 (N_9404,N_8185,N_8667);
or U9405 (N_9405,N_8782,N_7922);
and U9406 (N_9406,N_8364,N_7695);
and U9407 (N_9407,N_8067,N_8149);
nand U9408 (N_9408,N_8412,N_8564);
xnor U9409 (N_9409,N_7734,N_8676);
nand U9410 (N_9410,N_8179,N_8693);
nor U9411 (N_9411,N_7745,N_8989);
nand U9412 (N_9412,N_7988,N_7863);
or U9413 (N_9413,N_7610,N_8493);
xnor U9414 (N_9414,N_8356,N_8226);
or U9415 (N_9415,N_8308,N_8803);
and U9416 (N_9416,N_7667,N_7700);
and U9417 (N_9417,N_8859,N_7558);
or U9418 (N_9418,N_8579,N_7503);
or U9419 (N_9419,N_8391,N_8677);
and U9420 (N_9420,N_8687,N_7543);
nor U9421 (N_9421,N_8909,N_8258);
nand U9422 (N_9422,N_7608,N_8535);
nand U9423 (N_9423,N_7954,N_7650);
or U9424 (N_9424,N_7740,N_8148);
and U9425 (N_9425,N_8296,N_8519);
nor U9426 (N_9426,N_8567,N_8660);
xnor U9427 (N_9427,N_8749,N_8074);
or U9428 (N_9428,N_7530,N_7902);
and U9429 (N_9429,N_7783,N_8189);
and U9430 (N_9430,N_8323,N_8447);
nand U9431 (N_9431,N_8207,N_8152);
xor U9432 (N_9432,N_8584,N_7702);
or U9433 (N_9433,N_8322,N_8457);
xor U9434 (N_9434,N_8383,N_7547);
xor U9435 (N_9435,N_8961,N_8980);
xnor U9436 (N_9436,N_8819,N_8194);
xor U9437 (N_9437,N_7500,N_8588);
and U9438 (N_9438,N_7926,N_8300);
and U9439 (N_9439,N_7590,N_7924);
nor U9440 (N_9440,N_8498,N_8551);
or U9441 (N_9441,N_8834,N_7912);
nand U9442 (N_9442,N_7929,N_8678);
and U9443 (N_9443,N_8199,N_7662);
and U9444 (N_9444,N_8790,N_8825);
and U9445 (N_9445,N_8773,N_8416);
nand U9446 (N_9446,N_8900,N_7561);
and U9447 (N_9447,N_8884,N_8775);
and U9448 (N_9448,N_8702,N_8978);
nor U9449 (N_9449,N_8589,N_8393);
and U9450 (N_9450,N_7968,N_8343);
xnor U9451 (N_9451,N_8937,N_8814);
and U9452 (N_9452,N_7921,N_8827);
nand U9453 (N_9453,N_8741,N_7897);
nor U9454 (N_9454,N_8848,N_8761);
nor U9455 (N_9455,N_7860,N_8645);
and U9456 (N_9456,N_8212,N_7995);
nor U9457 (N_9457,N_7939,N_7742);
nor U9458 (N_9458,N_8634,N_8181);
or U9459 (N_9459,N_8999,N_8846);
or U9460 (N_9460,N_7976,N_8792);
or U9461 (N_9461,N_8007,N_7822);
nand U9462 (N_9462,N_8129,N_8723);
nor U9463 (N_9463,N_8631,N_7643);
or U9464 (N_9464,N_8802,N_7909);
nor U9465 (N_9465,N_8111,N_8770);
or U9466 (N_9466,N_7652,N_8332);
or U9467 (N_9467,N_8712,N_8673);
and U9468 (N_9468,N_8166,N_8869);
and U9469 (N_9469,N_7874,N_8275);
nand U9470 (N_9470,N_8216,N_8289);
nand U9471 (N_9471,N_8172,N_8663);
nand U9472 (N_9472,N_7845,N_7882);
nor U9473 (N_9473,N_7622,N_7665);
or U9474 (N_9474,N_7875,N_8526);
nor U9475 (N_9475,N_8654,N_8243);
nor U9476 (N_9476,N_7672,N_7518);
and U9477 (N_9477,N_7594,N_7813);
nand U9478 (N_9478,N_8840,N_7603);
or U9479 (N_9479,N_8766,N_8784);
xor U9480 (N_9480,N_8798,N_8286);
and U9481 (N_9481,N_8896,N_8482);
or U9482 (N_9482,N_8375,N_8456);
and U9483 (N_9483,N_8637,N_7521);
xor U9484 (N_9484,N_8772,N_8516);
nor U9485 (N_9485,N_7600,N_8260);
or U9486 (N_9486,N_7963,N_8144);
or U9487 (N_9487,N_8428,N_7975);
nand U9488 (N_9488,N_8807,N_8703);
xnor U9489 (N_9489,N_8164,N_8888);
nand U9490 (N_9490,N_8161,N_8198);
xor U9491 (N_9491,N_7658,N_8599);
nand U9492 (N_9492,N_8119,N_7784);
nor U9493 (N_9493,N_8542,N_7846);
nand U9494 (N_9494,N_8947,N_8897);
nand U9495 (N_9495,N_8971,N_8711);
and U9496 (N_9496,N_8503,N_8474);
and U9497 (N_9497,N_8729,N_8851);
and U9498 (N_9498,N_8517,N_8287);
and U9499 (N_9499,N_8141,N_7746);
nand U9500 (N_9500,N_8470,N_7576);
or U9501 (N_9501,N_8713,N_7611);
nand U9502 (N_9502,N_7930,N_7669);
nor U9503 (N_9503,N_8532,N_7729);
and U9504 (N_9504,N_7790,N_8021);
nand U9505 (N_9505,N_7639,N_8670);
nor U9506 (N_9506,N_7689,N_8338);
nand U9507 (N_9507,N_8786,N_7758);
xor U9508 (N_9508,N_7916,N_7582);
or U9509 (N_9509,N_8249,N_7762);
and U9510 (N_9510,N_8251,N_7812);
nor U9511 (N_9511,N_7789,N_7896);
xor U9512 (N_9512,N_7657,N_7538);
or U9513 (N_9513,N_8221,N_8698);
and U9514 (N_9514,N_7889,N_8424);
and U9515 (N_9515,N_7687,N_8227);
nand U9516 (N_9516,N_8478,N_7602);
or U9517 (N_9517,N_8241,N_8309);
nand U9518 (N_9518,N_8302,N_7981);
nand U9519 (N_9519,N_7787,N_8926);
nor U9520 (N_9520,N_8484,N_7804);
nand U9521 (N_9521,N_8510,N_7842);
nand U9522 (N_9522,N_7965,N_8726);
or U9523 (N_9523,N_8525,N_8377);
nand U9524 (N_9524,N_7513,N_8256);
or U9525 (N_9525,N_7899,N_8486);
xor U9526 (N_9526,N_8872,N_7980);
nand U9527 (N_9527,N_8263,N_7872);
nor U9528 (N_9528,N_8754,N_8239);
or U9529 (N_9529,N_8646,N_7596);
nand U9530 (N_9530,N_8064,N_8644);
nand U9531 (N_9531,N_7527,N_8501);
and U9532 (N_9532,N_8659,N_8293);
and U9533 (N_9533,N_8883,N_8783);
xnor U9534 (N_9534,N_8826,N_7540);
or U9535 (N_9535,N_8472,N_7630);
and U9536 (N_9536,N_7751,N_8613);
nor U9537 (N_9537,N_8824,N_7918);
nand U9538 (N_9538,N_8170,N_8276);
nand U9539 (N_9539,N_8559,N_8387);
and U9540 (N_9540,N_8027,N_7588);
nor U9541 (N_9541,N_7984,N_8392);
and U9542 (N_9542,N_8965,N_8668);
nand U9543 (N_9543,N_8861,N_7564);
or U9544 (N_9544,N_8918,N_7572);
xnor U9545 (N_9545,N_8435,N_8465);
or U9546 (N_9546,N_7858,N_8534);
nand U9547 (N_9547,N_8563,N_8933);
or U9548 (N_9548,N_8156,N_7814);
and U9549 (N_9549,N_8508,N_8448);
nand U9550 (N_9550,N_7517,N_8722);
nand U9551 (N_9551,N_8538,N_8562);
nor U9552 (N_9552,N_8135,N_8789);
and U9553 (N_9553,N_7586,N_7516);
nor U9554 (N_9554,N_8592,N_8030);
nand U9555 (N_9555,N_7565,N_8450);
nand U9556 (N_9556,N_8623,N_7911);
nand U9557 (N_9557,N_7693,N_8247);
or U9558 (N_9558,N_8515,N_7721);
and U9559 (N_9559,N_8389,N_8624);
nor U9560 (N_9560,N_8445,N_7952);
or U9561 (N_9561,N_8234,N_7795);
nand U9562 (N_9562,N_7779,N_8518);
or U9563 (N_9563,N_8675,N_7664);
or U9564 (N_9564,N_8147,N_7567);
nand U9565 (N_9565,N_8706,N_8865);
or U9566 (N_9566,N_8265,N_7620);
nor U9567 (N_9567,N_8026,N_8028);
nand U9568 (N_9568,N_8647,N_8495);
xnor U9569 (N_9569,N_8904,N_7801);
nor U9570 (N_9570,N_8527,N_8911);
nand U9571 (N_9571,N_7834,N_7840);
nand U9572 (N_9572,N_7764,N_8461);
nand U9573 (N_9573,N_8361,N_8160);
nor U9574 (N_9574,N_8988,N_8931);
nand U9575 (N_9575,N_8336,N_8764);
or U9576 (N_9576,N_7865,N_8429);
nand U9577 (N_9577,N_7679,N_7844);
and U9578 (N_9578,N_8511,N_7928);
xnor U9579 (N_9579,N_7545,N_8151);
and U9580 (N_9580,N_7775,N_7996);
and U9581 (N_9581,N_8292,N_8938);
nor U9582 (N_9582,N_8895,N_8924);
nor U9583 (N_9583,N_7962,N_8661);
xor U9584 (N_9584,N_8195,N_8805);
nand U9585 (N_9585,N_8607,N_7519);
nand U9586 (N_9586,N_8215,N_8163);
nor U9587 (N_9587,N_8182,N_8957);
and U9588 (N_9588,N_7950,N_8080);
and U9589 (N_9589,N_8054,N_7806);
and U9590 (N_9590,N_8831,N_8818);
or U9591 (N_9591,N_8213,N_8223);
xor U9592 (N_9592,N_7796,N_8638);
and U9593 (N_9593,N_8506,N_8945);
nor U9594 (N_9594,N_8035,N_8104);
nand U9595 (N_9595,N_8409,N_8601);
nor U9596 (N_9596,N_8342,N_8628);
or U9597 (N_9597,N_8406,N_7676);
and U9598 (N_9598,N_8460,N_7948);
nor U9599 (N_9599,N_7946,N_8575);
or U9600 (N_9600,N_7817,N_8800);
nand U9601 (N_9601,N_8410,N_8092);
and U9602 (N_9602,N_8545,N_8481);
nor U9603 (N_9603,N_8333,N_7737);
nand U9604 (N_9604,N_7781,N_7791);
and U9605 (N_9605,N_8558,N_8390);
nand U9606 (N_9606,N_8398,N_8757);
or U9607 (N_9607,N_8130,N_8873);
nor U9608 (N_9608,N_8229,N_7788);
and U9609 (N_9609,N_8068,N_7617);
and U9610 (N_9610,N_8010,N_8679);
or U9611 (N_9611,N_8082,N_8707);
nand U9612 (N_9612,N_7506,N_8752);
xnor U9613 (N_9613,N_7674,N_8746);
nand U9614 (N_9614,N_8715,N_8039);
nand U9615 (N_9615,N_8078,N_8785);
nor U9616 (N_9616,N_8464,N_8874);
or U9617 (N_9617,N_8536,N_8642);
nand U9618 (N_9618,N_7563,N_7908);
xor U9619 (N_9619,N_8114,N_8768);
nand U9620 (N_9620,N_8728,N_8576);
nor U9621 (N_9621,N_8857,N_8778);
nand U9622 (N_9622,N_8245,N_7998);
and U9623 (N_9623,N_7623,N_8651);
nand U9624 (N_9624,N_7589,N_8417);
nand U9625 (N_9625,N_8730,N_7945);
nor U9626 (N_9626,N_7837,N_8491);
nor U9627 (N_9627,N_8108,N_7504);
xor U9628 (N_9628,N_8352,N_8273);
nor U9629 (N_9629,N_7867,N_8916);
xor U9630 (N_9630,N_7824,N_8626);
nand U9631 (N_9631,N_7554,N_8600);
nor U9632 (N_9632,N_8744,N_7776);
and U9633 (N_9633,N_8774,N_8533);
or U9634 (N_9634,N_8614,N_8935);
or U9635 (N_9635,N_7579,N_7595);
nor U9636 (N_9636,N_8727,N_7508);
and U9637 (N_9637,N_7730,N_7940);
nor U9638 (N_9638,N_8991,N_8426);
nand U9639 (N_9639,N_7573,N_7549);
nand U9640 (N_9640,N_8087,N_7754);
nand U9641 (N_9641,N_8353,N_7661);
nand U9642 (N_9642,N_8220,N_8176);
and U9643 (N_9643,N_8993,N_8611);
or U9644 (N_9644,N_8206,N_7953);
and U9645 (N_9645,N_8319,N_7855);
or U9646 (N_9646,N_8131,N_8606);
nor U9647 (N_9647,N_8314,N_7640);
or U9648 (N_9648,N_8005,N_8876);
and U9649 (N_9649,N_8360,N_8180);
and U9650 (N_9650,N_8903,N_7927);
xnor U9651 (N_9651,N_8413,N_8640);
xor U9652 (N_9652,N_7714,N_8473);
nand U9653 (N_9653,N_8116,N_8822);
nor U9654 (N_9654,N_8334,N_7668);
and U9655 (N_9655,N_8046,N_7680);
and U9656 (N_9656,N_8270,N_7616);
and U9657 (N_9657,N_8422,N_8902);
nor U9658 (N_9658,N_7533,N_8882);
or U9659 (N_9659,N_8939,N_8977);
xnor U9660 (N_9660,N_8031,N_8855);
and U9661 (N_9661,N_8255,N_8167);
nor U9662 (N_9662,N_7749,N_8143);
nor U9663 (N_9663,N_8853,N_8697);
and U9664 (N_9664,N_8942,N_7575);
nor U9665 (N_9665,N_7785,N_8907);
nor U9666 (N_9666,N_7649,N_8408);
and U9667 (N_9667,N_8446,N_8806);
and U9668 (N_9668,N_8737,N_7514);
nand U9669 (N_9669,N_7811,N_7553);
nor U9670 (N_9670,N_7823,N_8596);
nor U9671 (N_9671,N_8690,N_8222);
nand U9672 (N_9672,N_7678,N_8899);
nor U9673 (N_9673,N_8134,N_8083);
nand U9674 (N_9674,N_8257,N_8630);
and U9675 (N_9675,N_8743,N_7577);
nor U9676 (N_9676,N_8274,N_8165);
or U9677 (N_9677,N_8740,N_8832);
and U9678 (N_9678,N_8738,N_8310);
nand U9679 (N_9679,N_8521,N_8955);
or U9680 (N_9680,N_8796,N_8691);
or U9681 (N_9681,N_8175,N_8710);
nor U9682 (N_9682,N_8311,N_8440);
or U9683 (N_9683,N_8442,N_7597);
nor U9684 (N_9684,N_7591,N_7569);
or U9685 (N_9685,N_8430,N_8267);
nor U9686 (N_9686,N_7696,N_8022);
nor U9687 (N_9687,N_7684,N_8017);
and U9688 (N_9688,N_7609,N_8569);
xor U9689 (N_9689,N_7756,N_8669);
or U9690 (N_9690,N_8721,N_8680);
and U9691 (N_9691,N_8889,N_8305);
and U9692 (N_9692,N_8837,N_7585);
nor U9693 (N_9693,N_7604,N_8126);
and U9694 (N_9694,N_7555,N_7583);
and U9695 (N_9695,N_7951,N_8639);
and U9696 (N_9696,N_8348,N_7654);
nor U9697 (N_9697,N_7818,N_8641);
nor U9698 (N_9698,N_8982,N_7828);
nor U9699 (N_9699,N_8987,N_7710);
nand U9700 (N_9700,N_7743,N_7848);
nand U9701 (N_9701,N_8880,N_7641);
nand U9702 (N_9702,N_7570,N_8162);
nand U9703 (N_9703,N_8113,N_7697);
and U9704 (N_9704,N_7690,N_8893);
nand U9705 (N_9705,N_8984,N_7627);
or U9706 (N_9706,N_7805,N_8842);
nor U9707 (N_9707,N_8140,N_8262);
nand U9708 (N_9708,N_8340,N_7798);
nor U9709 (N_9709,N_8184,N_7977);
nor U9710 (N_9710,N_8463,N_8337);
xor U9711 (N_9711,N_8541,N_7688);
and U9712 (N_9712,N_8419,N_8941);
nand U9713 (N_9713,N_8618,N_8688);
nor U9714 (N_9714,N_8329,N_7613);
nor U9715 (N_9715,N_7895,N_8400);
or U9716 (N_9716,N_8914,N_8587);
nor U9717 (N_9717,N_8210,N_8561);
nand U9718 (N_9718,N_8048,N_7548);
xor U9719 (N_9719,N_8385,N_8366);
nor U9720 (N_9720,N_7703,N_8294);
or U9721 (N_9721,N_8462,N_7941);
xnor U9722 (N_9722,N_8944,N_8621);
and U9723 (N_9723,N_8120,N_7983);
and U9724 (N_9724,N_7646,N_8817);
nand U9725 (N_9725,N_8540,N_8071);
and U9726 (N_9726,N_7628,N_8344);
or U9727 (N_9727,N_7707,N_8103);
nand U9728 (N_9728,N_7544,N_7675);
or U9729 (N_9729,N_8047,N_8632);
nor U9730 (N_9730,N_8299,N_8001);
xnor U9731 (N_9731,N_8236,N_7768);
xor U9732 (N_9732,N_8277,N_8843);
or U9733 (N_9733,N_7636,N_8418);
or U9734 (N_9734,N_8514,N_8174);
and U9735 (N_9735,N_7612,N_8049);
or U9736 (N_9736,N_7915,N_7878);
xor U9737 (N_9737,N_8476,N_8724);
nor U9738 (N_9738,N_8248,N_7967);
and U9739 (N_9739,N_8427,N_7900);
or U9740 (N_9740,N_8370,N_8301);
and U9741 (N_9741,N_8627,N_8225);
xor U9742 (N_9742,N_8280,N_8313);
or U9743 (N_9743,N_7568,N_7578);
or U9744 (N_9744,N_8578,N_7528);
nor U9745 (N_9745,N_7644,N_7772);
nor U9746 (N_9746,N_8158,N_8454);
nor U9747 (N_9747,N_8974,N_7955);
nor U9748 (N_9748,N_8981,N_8950);
nor U9749 (N_9749,N_8620,N_8012);
or U9750 (N_9750,N_8459,N_8280);
xnor U9751 (N_9751,N_8843,N_8396);
nand U9752 (N_9752,N_8523,N_7748);
xor U9753 (N_9753,N_7864,N_8923);
or U9754 (N_9754,N_8527,N_7895);
nor U9755 (N_9755,N_8759,N_8535);
or U9756 (N_9756,N_7756,N_7528);
nor U9757 (N_9757,N_8881,N_8981);
xor U9758 (N_9758,N_8015,N_8365);
nand U9759 (N_9759,N_8289,N_8940);
nor U9760 (N_9760,N_8958,N_8405);
nor U9761 (N_9761,N_8482,N_7929);
nor U9762 (N_9762,N_8335,N_8304);
and U9763 (N_9763,N_8245,N_7700);
or U9764 (N_9764,N_8040,N_7524);
nand U9765 (N_9765,N_7612,N_7513);
and U9766 (N_9766,N_8387,N_7996);
or U9767 (N_9767,N_7742,N_8272);
or U9768 (N_9768,N_7591,N_7739);
or U9769 (N_9769,N_7681,N_7913);
nor U9770 (N_9770,N_8788,N_8552);
nand U9771 (N_9771,N_8102,N_7757);
nor U9772 (N_9772,N_8862,N_7644);
or U9773 (N_9773,N_8766,N_8991);
and U9774 (N_9774,N_8832,N_8710);
nand U9775 (N_9775,N_7686,N_8121);
nand U9776 (N_9776,N_8152,N_8347);
or U9777 (N_9777,N_8225,N_7577);
nand U9778 (N_9778,N_7860,N_7962);
nand U9779 (N_9779,N_8729,N_7987);
nand U9780 (N_9780,N_7557,N_8343);
or U9781 (N_9781,N_7936,N_8801);
nor U9782 (N_9782,N_8153,N_8124);
or U9783 (N_9783,N_8369,N_8334);
xnor U9784 (N_9784,N_7952,N_8213);
nand U9785 (N_9785,N_8658,N_8844);
xor U9786 (N_9786,N_7701,N_8990);
and U9787 (N_9787,N_8044,N_7523);
or U9788 (N_9788,N_8661,N_8201);
nor U9789 (N_9789,N_7675,N_8649);
or U9790 (N_9790,N_8145,N_7588);
or U9791 (N_9791,N_8828,N_8040);
or U9792 (N_9792,N_8945,N_7957);
nand U9793 (N_9793,N_7814,N_7592);
and U9794 (N_9794,N_8782,N_7923);
nor U9795 (N_9795,N_8725,N_8870);
nand U9796 (N_9796,N_8110,N_8182);
nand U9797 (N_9797,N_7612,N_8486);
or U9798 (N_9798,N_8967,N_7832);
and U9799 (N_9799,N_7728,N_8355);
nand U9800 (N_9800,N_8281,N_7901);
nor U9801 (N_9801,N_7964,N_8958);
or U9802 (N_9802,N_8331,N_7677);
nand U9803 (N_9803,N_8772,N_8125);
or U9804 (N_9804,N_8069,N_8476);
and U9805 (N_9805,N_8908,N_8534);
nand U9806 (N_9806,N_7506,N_7976);
or U9807 (N_9807,N_8094,N_8325);
or U9808 (N_9808,N_8496,N_7755);
and U9809 (N_9809,N_8182,N_7640);
nor U9810 (N_9810,N_7932,N_7997);
nand U9811 (N_9811,N_8669,N_8086);
or U9812 (N_9812,N_8585,N_7995);
and U9813 (N_9813,N_8702,N_7954);
nor U9814 (N_9814,N_8290,N_8790);
nand U9815 (N_9815,N_8419,N_8892);
or U9816 (N_9816,N_8032,N_8050);
nor U9817 (N_9817,N_8417,N_8839);
or U9818 (N_9818,N_8946,N_8254);
and U9819 (N_9819,N_8676,N_8401);
xnor U9820 (N_9820,N_8135,N_7526);
nor U9821 (N_9821,N_8061,N_7767);
nand U9822 (N_9822,N_7744,N_8687);
and U9823 (N_9823,N_8679,N_8375);
nand U9824 (N_9824,N_8146,N_7504);
and U9825 (N_9825,N_8678,N_7709);
nor U9826 (N_9826,N_8993,N_8790);
and U9827 (N_9827,N_8597,N_7752);
or U9828 (N_9828,N_8435,N_7555);
and U9829 (N_9829,N_8865,N_8280);
or U9830 (N_9830,N_8392,N_8212);
and U9831 (N_9831,N_7539,N_8938);
and U9832 (N_9832,N_8693,N_7832);
or U9833 (N_9833,N_7643,N_8454);
nor U9834 (N_9834,N_8281,N_7521);
and U9835 (N_9835,N_8428,N_7706);
nand U9836 (N_9836,N_7931,N_8882);
and U9837 (N_9837,N_8067,N_8827);
nand U9838 (N_9838,N_8498,N_8794);
nand U9839 (N_9839,N_8920,N_7879);
or U9840 (N_9840,N_8991,N_8763);
and U9841 (N_9841,N_8761,N_8106);
nand U9842 (N_9842,N_8435,N_8170);
or U9843 (N_9843,N_8251,N_8806);
or U9844 (N_9844,N_8384,N_8147);
nand U9845 (N_9845,N_8674,N_7695);
and U9846 (N_9846,N_8537,N_8702);
nor U9847 (N_9847,N_7777,N_8939);
nor U9848 (N_9848,N_7543,N_8215);
nand U9849 (N_9849,N_7544,N_8732);
nand U9850 (N_9850,N_8499,N_8099);
nand U9851 (N_9851,N_8932,N_8820);
or U9852 (N_9852,N_7645,N_7947);
nor U9853 (N_9853,N_8613,N_8886);
nor U9854 (N_9854,N_7753,N_8503);
and U9855 (N_9855,N_8313,N_7915);
nand U9856 (N_9856,N_8338,N_7921);
nand U9857 (N_9857,N_7987,N_7702);
nor U9858 (N_9858,N_7752,N_7906);
nor U9859 (N_9859,N_8530,N_7755);
nand U9860 (N_9860,N_8962,N_7830);
and U9861 (N_9861,N_8726,N_8498);
or U9862 (N_9862,N_7603,N_8808);
xnor U9863 (N_9863,N_8852,N_7634);
nor U9864 (N_9864,N_7636,N_7560);
nand U9865 (N_9865,N_8348,N_8600);
xnor U9866 (N_9866,N_8956,N_8148);
and U9867 (N_9867,N_8083,N_8727);
nor U9868 (N_9868,N_7795,N_7818);
nor U9869 (N_9869,N_8962,N_8892);
nand U9870 (N_9870,N_8181,N_7640);
xnor U9871 (N_9871,N_8664,N_8276);
and U9872 (N_9872,N_8208,N_8457);
or U9873 (N_9873,N_7654,N_7560);
or U9874 (N_9874,N_8092,N_7674);
nand U9875 (N_9875,N_8541,N_8783);
or U9876 (N_9876,N_8149,N_7806);
or U9877 (N_9877,N_8114,N_7522);
and U9878 (N_9878,N_8212,N_7975);
nand U9879 (N_9879,N_8316,N_8840);
or U9880 (N_9880,N_7675,N_8733);
nor U9881 (N_9881,N_8305,N_8688);
nand U9882 (N_9882,N_8272,N_7878);
or U9883 (N_9883,N_8140,N_7614);
and U9884 (N_9884,N_8518,N_8784);
and U9885 (N_9885,N_8999,N_7791);
nor U9886 (N_9886,N_8836,N_8448);
and U9887 (N_9887,N_8241,N_8064);
or U9888 (N_9888,N_7622,N_8563);
nor U9889 (N_9889,N_8080,N_8529);
and U9890 (N_9890,N_8764,N_7562);
nor U9891 (N_9891,N_8271,N_7984);
nand U9892 (N_9892,N_7573,N_8920);
or U9893 (N_9893,N_7828,N_7649);
nor U9894 (N_9894,N_7945,N_8200);
xor U9895 (N_9895,N_7934,N_8010);
nand U9896 (N_9896,N_8295,N_7691);
nor U9897 (N_9897,N_8523,N_8241);
nand U9898 (N_9898,N_8541,N_8723);
and U9899 (N_9899,N_7669,N_8044);
nor U9900 (N_9900,N_7929,N_7799);
nor U9901 (N_9901,N_8773,N_8938);
and U9902 (N_9902,N_7809,N_8389);
nor U9903 (N_9903,N_8053,N_7977);
xnor U9904 (N_9904,N_8210,N_8484);
xnor U9905 (N_9905,N_8469,N_7935);
and U9906 (N_9906,N_8387,N_8507);
nor U9907 (N_9907,N_8311,N_7811);
and U9908 (N_9908,N_8121,N_8239);
nand U9909 (N_9909,N_7725,N_8896);
nand U9910 (N_9910,N_8432,N_8493);
xor U9911 (N_9911,N_8644,N_7742);
or U9912 (N_9912,N_8868,N_7751);
and U9913 (N_9913,N_7666,N_7502);
and U9914 (N_9914,N_7649,N_8781);
or U9915 (N_9915,N_7706,N_8647);
nor U9916 (N_9916,N_8956,N_7738);
or U9917 (N_9917,N_8332,N_8680);
nor U9918 (N_9918,N_7568,N_8023);
nand U9919 (N_9919,N_8429,N_8183);
and U9920 (N_9920,N_7966,N_8033);
nor U9921 (N_9921,N_8192,N_8293);
nor U9922 (N_9922,N_7832,N_7513);
xnor U9923 (N_9923,N_8631,N_8849);
or U9924 (N_9924,N_7979,N_8078);
or U9925 (N_9925,N_8699,N_7721);
xor U9926 (N_9926,N_8865,N_8729);
nand U9927 (N_9927,N_7954,N_7517);
and U9928 (N_9928,N_7703,N_8384);
nor U9929 (N_9929,N_8320,N_7762);
and U9930 (N_9930,N_7545,N_8228);
or U9931 (N_9931,N_7591,N_8683);
xor U9932 (N_9932,N_8400,N_8937);
xor U9933 (N_9933,N_8790,N_7972);
nor U9934 (N_9934,N_7723,N_7880);
and U9935 (N_9935,N_8242,N_8943);
and U9936 (N_9936,N_8093,N_7936);
xnor U9937 (N_9937,N_7941,N_7728);
nor U9938 (N_9938,N_8738,N_8098);
or U9939 (N_9939,N_7676,N_8025);
nand U9940 (N_9940,N_8820,N_8375);
nand U9941 (N_9941,N_8818,N_8808);
nand U9942 (N_9942,N_8238,N_7704);
or U9943 (N_9943,N_8863,N_7713);
or U9944 (N_9944,N_7526,N_7523);
nor U9945 (N_9945,N_8589,N_8992);
or U9946 (N_9946,N_7536,N_7796);
and U9947 (N_9947,N_7696,N_8319);
and U9948 (N_9948,N_8908,N_8188);
nor U9949 (N_9949,N_7881,N_7652);
and U9950 (N_9950,N_8222,N_8210);
nand U9951 (N_9951,N_8225,N_7708);
and U9952 (N_9952,N_7761,N_7555);
and U9953 (N_9953,N_8366,N_7658);
or U9954 (N_9954,N_7724,N_8346);
nand U9955 (N_9955,N_7678,N_8851);
nor U9956 (N_9956,N_8955,N_8564);
and U9957 (N_9957,N_7682,N_7722);
and U9958 (N_9958,N_8467,N_8631);
nor U9959 (N_9959,N_8169,N_7588);
xor U9960 (N_9960,N_8410,N_7921);
nand U9961 (N_9961,N_8088,N_8782);
xnor U9962 (N_9962,N_7666,N_8902);
xnor U9963 (N_9963,N_8891,N_8601);
nand U9964 (N_9964,N_7688,N_7502);
nand U9965 (N_9965,N_7895,N_7606);
nor U9966 (N_9966,N_8097,N_8076);
nand U9967 (N_9967,N_8463,N_8913);
nand U9968 (N_9968,N_7687,N_8320);
nand U9969 (N_9969,N_7637,N_7943);
and U9970 (N_9970,N_8519,N_8986);
or U9971 (N_9971,N_7531,N_7885);
nor U9972 (N_9972,N_8049,N_8967);
xnor U9973 (N_9973,N_8020,N_8318);
nand U9974 (N_9974,N_8948,N_8148);
nand U9975 (N_9975,N_8689,N_7830);
nand U9976 (N_9976,N_8111,N_8558);
or U9977 (N_9977,N_8950,N_8375);
xnor U9978 (N_9978,N_7653,N_7736);
nor U9979 (N_9979,N_8652,N_8860);
nand U9980 (N_9980,N_7709,N_8068);
and U9981 (N_9981,N_8369,N_8599);
and U9982 (N_9982,N_8663,N_7972);
nor U9983 (N_9983,N_8707,N_7731);
or U9984 (N_9984,N_8429,N_8135);
nand U9985 (N_9985,N_8936,N_8731);
xnor U9986 (N_9986,N_8879,N_7774);
and U9987 (N_9987,N_8556,N_8623);
xor U9988 (N_9988,N_7875,N_8505);
nor U9989 (N_9989,N_8343,N_8188);
and U9990 (N_9990,N_8591,N_7993);
or U9991 (N_9991,N_8754,N_8749);
nor U9992 (N_9992,N_7679,N_8581);
or U9993 (N_9993,N_8007,N_8676);
nand U9994 (N_9994,N_8327,N_8087);
and U9995 (N_9995,N_7501,N_8060);
nand U9996 (N_9996,N_7611,N_7634);
nand U9997 (N_9997,N_7507,N_8749);
nor U9998 (N_9998,N_8142,N_8137);
or U9999 (N_9999,N_8244,N_7907);
nor U10000 (N_10000,N_8865,N_8285);
nor U10001 (N_10001,N_7744,N_8886);
nor U10002 (N_10002,N_7694,N_7584);
nand U10003 (N_10003,N_8691,N_7823);
nand U10004 (N_10004,N_8192,N_8308);
or U10005 (N_10005,N_8806,N_8308);
nand U10006 (N_10006,N_8646,N_7937);
nand U10007 (N_10007,N_8575,N_8722);
nor U10008 (N_10008,N_8293,N_8277);
and U10009 (N_10009,N_8656,N_8443);
and U10010 (N_10010,N_8972,N_7986);
nand U10011 (N_10011,N_8938,N_8189);
and U10012 (N_10012,N_7512,N_7795);
and U10013 (N_10013,N_7720,N_8091);
xnor U10014 (N_10014,N_8796,N_8574);
and U10015 (N_10015,N_7507,N_8566);
and U10016 (N_10016,N_8982,N_8921);
nor U10017 (N_10017,N_7766,N_8661);
nand U10018 (N_10018,N_7761,N_7739);
nor U10019 (N_10019,N_8121,N_8801);
nor U10020 (N_10020,N_8500,N_8062);
or U10021 (N_10021,N_8339,N_8295);
and U10022 (N_10022,N_7804,N_7614);
or U10023 (N_10023,N_8821,N_8388);
xor U10024 (N_10024,N_7778,N_8403);
xnor U10025 (N_10025,N_7640,N_7549);
and U10026 (N_10026,N_8137,N_7925);
nand U10027 (N_10027,N_8124,N_8202);
and U10028 (N_10028,N_8574,N_8777);
nor U10029 (N_10029,N_7830,N_8011);
nor U10030 (N_10030,N_8704,N_7935);
or U10031 (N_10031,N_8477,N_7570);
or U10032 (N_10032,N_7608,N_8301);
nor U10033 (N_10033,N_8155,N_8432);
and U10034 (N_10034,N_8007,N_7769);
or U10035 (N_10035,N_8710,N_8102);
and U10036 (N_10036,N_7801,N_8103);
xnor U10037 (N_10037,N_7893,N_8718);
nand U10038 (N_10038,N_7505,N_8609);
and U10039 (N_10039,N_7627,N_8400);
nor U10040 (N_10040,N_7745,N_8333);
xor U10041 (N_10041,N_7592,N_8493);
nor U10042 (N_10042,N_8755,N_8720);
xor U10043 (N_10043,N_7589,N_8473);
nand U10044 (N_10044,N_8438,N_7601);
nand U10045 (N_10045,N_8411,N_7623);
or U10046 (N_10046,N_8427,N_7959);
and U10047 (N_10047,N_8845,N_8978);
nor U10048 (N_10048,N_8858,N_8943);
xor U10049 (N_10049,N_8751,N_8483);
or U10050 (N_10050,N_8746,N_8891);
nand U10051 (N_10051,N_7937,N_8689);
or U10052 (N_10052,N_8935,N_8756);
nand U10053 (N_10053,N_7959,N_8676);
nand U10054 (N_10054,N_8113,N_8122);
or U10055 (N_10055,N_8792,N_7814);
nand U10056 (N_10056,N_7988,N_8095);
nor U10057 (N_10057,N_8386,N_8524);
nand U10058 (N_10058,N_8207,N_7931);
nor U10059 (N_10059,N_8848,N_8546);
nor U10060 (N_10060,N_8041,N_8244);
and U10061 (N_10061,N_8522,N_7847);
or U10062 (N_10062,N_7853,N_8979);
and U10063 (N_10063,N_8827,N_8699);
xor U10064 (N_10064,N_8281,N_7618);
and U10065 (N_10065,N_7566,N_7573);
and U10066 (N_10066,N_8571,N_8105);
xor U10067 (N_10067,N_7500,N_8583);
and U10068 (N_10068,N_7702,N_8811);
and U10069 (N_10069,N_7949,N_8473);
or U10070 (N_10070,N_7887,N_7973);
nand U10071 (N_10071,N_8925,N_8436);
and U10072 (N_10072,N_7511,N_8052);
nor U10073 (N_10073,N_8696,N_8933);
nand U10074 (N_10074,N_7697,N_7770);
nor U10075 (N_10075,N_7921,N_7772);
and U10076 (N_10076,N_8613,N_7763);
and U10077 (N_10077,N_8110,N_8221);
nor U10078 (N_10078,N_8817,N_8317);
and U10079 (N_10079,N_8561,N_8610);
nor U10080 (N_10080,N_8783,N_8069);
xnor U10081 (N_10081,N_8460,N_7846);
and U10082 (N_10082,N_7610,N_8615);
and U10083 (N_10083,N_7538,N_8680);
nand U10084 (N_10084,N_8986,N_7839);
nor U10085 (N_10085,N_8434,N_8626);
nor U10086 (N_10086,N_7664,N_8503);
or U10087 (N_10087,N_7975,N_8148);
xnor U10088 (N_10088,N_8838,N_8491);
and U10089 (N_10089,N_8170,N_8338);
xnor U10090 (N_10090,N_7780,N_8638);
nand U10091 (N_10091,N_8811,N_8262);
nor U10092 (N_10092,N_8257,N_8628);
or U10093 (N_10093,N_8194,N_8319);
nor U10094 (N_10094,N_8343,N_7660);
xor U10095 (N_10095,N_8391,N_8002);
xor U10096 (N_10096,N_7654,N_8597);
or U10097 (N_10097,N_7753,N_7794);
and U10098 (N_10098,N_7664,N_7885);
xor U10099 (N_10099,N_8326,N_7597);
and U10100 (N_10100,N_7624,N_8921);
nor U10101 (N_10101,N_8532,N_7644);
nor U10102 (N_10102,N_7868,N_8554);
nand U10103 (N_10103,N_7982,N_8574);
nor U10104 (N_10104,N_7724,N_8255);
or U10105 (N_10105,N_8475,N_8537);
and U10106 (N_10106,N_8038,N_8729);
nor U10107 (N_10107,N_8317,N_7732);
or U10108 (N_10108,N_8571,N_8022);
and U10109 (N_10109,N_8006,N_8847);
nor U10110 (N_10110,N_8535,N_7705);
nand U10111 (N_10111,N_8991,N_8191);
or U10112 (N_10112,N_7902,N_7829);
nand U10113 (N_10113,N_7552,N_8846);
and U10114 (N_10114,N_8152,N_7686);
nor U10115 (N_10115,N_7945,N_7858);
nand U10116 (N_10116,N_7649,N_8850);
or U10117 (N_10117,N_8253,N_7624);
or U10118 (N_10118,N_7906,N_8963);
nor U10119 (N_10119,N_8567,N_8659);
or U10120 (N_10120,N_8889,N_8525);
nand U10121 (N_10121,N_8932,N_8728);
nor U10122 (N_10122,N_7552,N_7917);
and U10123 (N_10123,N_8279,N_8199);
or U10124 (N_10124,N_8103,N_7911);
or U10125 (N_10125,N_8570,N_8712);
nand U10126 (N_10126,N_8676,N_8430);
nand U10127 (N_10127,N_8653,N_7789);
xnor U10128 (N_10128,N_8273,N_7587);
nand U10129 (N_10129,N_7685,N_8229);
nor U10130 (N_10130,N_8276,N_8239);
and U10131 (N_10131,N_8940,N_8958);
nand U10132 (N_10132,N_8442,N_7690);
and U10133 (N_10133,N_7559,N_8241);
and U10134 (N_10134,N_7768,N_8300);
nor U10135 (N_10135,N_7766,N_8547);
and U10136 (N_10136,N_8410,N_8732);
nand U10137 (N_10137,N_8236,N_8528);
xor U10138 (N_10138,N_8206,N_8930);
nor U10139 (N_10139,N_8945,N_7964);
xor U10140 (N_10140,N_8795,N_8787);
nor U10141 (N_10141,N_7998,N_8631);
nor U10142 (N_10142,N_8109,N_7669);
and U10143 (N_10143,N_7910,N_7750);
or U10144 (N_10144,N_8434,N_8578);
and U10145 (N_10145,N_7720,N_7990);
or U10146 (N_10146,N_8683,N_7837);
nand U10147 (N_10147,N_8161,N_8650);
xor U10148 (N_10148,N_8005,N_8980);
or U10149 (N_10149,N_8742,N_7712);
and U10150 (N_10150,N_8777,N_8717);
or U10151 (N_10151,N_8327,N_8465);
xor U10152 (N_10152,N_8792,N_7690);
or U10153 (N_10153,N_8528,N_7974);
nor U10154 (N_10154,N_7740,N_8225);
nand U10155 (N_10155,N_8441,N_8495);
xnor U10156 (N_10156,N_8554,N_7896);
or U10157 (N_10157,N_7876,N_8358);
or U10158 (N_10158,N_7817,N_8091);
or U10159 (N_10159,N_8782,N_7527);
or U10160 (N_10160,N_7515,N_8330);
or U10161 (N_10161,N_8873,N_8476);
and U10162 (N_10162,N_8793,N_8558);
nand U10163 (N_10163,N_8935,N_8167);
nor U10164 (N_10164,N_8602,N_8039);
or U10165 (N_10165,N_8709,N_7762);
nand U10166 (N_10166,N_7687,N_8867);
nand U10167 (N_10167,N_8977,N_7882);
nand U10168 (N_10168,N_8648,N_8725);
nor U10169 (N_10169,N_7849,N_8813);
nor U10170 (N_10170,N_8522,N_8403);
nor U10171 (N_10171,N_7801,N_8410);
and U10172 (N_10172,N_7913,N_8786);
and U10173 (N_10173,N_8574,N_8806);
xor U10174 (N_10174,N_8228,N_8406);
or U10175 (N_10175,N_8692,N_7503);
and U10176 (N_10176,N_7504,N_7746);
nand U10177 (N_10177,N_8059,N_8492);
nand U10178 (N_10178,N_8382,N_8903);
and U10179 (N_10179,N_8156,N_8941);
nor U10180 (N_10180,N_8366,N_7675);
or U10181 (N_10181,N_7818,N_8313);
xnor U10182 (N_10182,N_8923,N_7840);
or U10183 (N_10183,N_8897,N_8704);
nand U10184 (N_10184,N_7619,N_8924);
nor U10185 (N_10185,N_7616,N_8349);
or U10186 (N_10186,N_7578,N_8056);
or U10187 (N_10187,N_8856,N_8667);
or U10188 (N_10188,N_8455,N_8755);
and U10189 (N_10189,N_7919,N_8930);
nand U10190 (N_10190,N_7958,N_7703);
or U10191 (N_10191,N_8173,N_7687);
and U10192 (N_10192,N_8108,N_7802);
nand U10193 (N_10193,N_8648,N_8606);
or U10194 (N_10194,N_8063,N_8857);
nand U10195 (N_10195,N_8603,N_8004);
and U10196 (N_10196,N_8402,N_8914);
nand U10197 (N_10197,N_8050,N_8426);
or U10198 (N_10198,N_8674,N_7615);
nand U10199 (N_10199,N_7764,N_7824);
or U10200 (N_10200,N_8588,N_8963);
xnor U10201 (N_10201,N_8082,N_8968);
nor U10202 (N_10202,N_7965,N_8108);
nor U10203 (N_10203,N_8631,N_7731);
nor U10204 (N_10204,N_8249,N_8579);
xnor U10205 (N_10205,N_7770,N_8592);
and U10206 (N_10206,N_7993,N_8374);
or U10207 (N_10207,N_8356,N_7684);
nand U10208 (N_10208,N_7752,N_8638);
and U10209 (N_10209,N_7730,N_8862);
nand U10210 (N_10210,N_8073,N_8750);
nor U10211 (N_10211,N_8980,N_8709);
and U10212 (N_10212,N_8768,N_8847);
and U10213 (N_10213,N_7748,N_7641);
or U10214 (N_10214,N_7629,N_8380);
or U10215 (N_10215,N_8519,N_8476);
nor U10216 (N_10216,N_8249,N_8074);
nor U10217 (N_10217,N_7765,N_8790);
nand U10218 (N_10218,N_8702,N_7617);
and U10219 (N_10219,N_7856,N_8791);
or U10220 (N_10220,N_7746,N_7677);
or U10221 (N_10221,N_8291,N_8504);
xor U10222 (N_10222,N_7512,N_7601);
nand U10223 (N_10223,N_8775,N_8373);
or U10224 (N_10224,N_7895,N_7819);
and U10225 (N_10225,N_8185,N_8171);
and U10226 (N_10226,N_7648,N_8845);
nand U10227 (N_10227,N_7814,N_8536);
or U10228 (N_10228,N_8360,N_8396);
xnor U10229 (N_10229,N_7507,N_7896);
nor U10230 (N_10230,N_8351,N_7794);
and U10231 (N_10231,N_7964,N_8387);
nor U10232 (N_10232,N_7583,N_7698);
nor U10233 (N_10233,N_8227,N_7662);
nor U10234 (N_10234,N_8884,N_8572);
nor U10235 (N_10235,N_8392,N_8244);
and U10236 (N_10236,N_7827,N_8756);
nand U10237 (N_10237,N_8396,N_7665);
and U10238 (N_10238,N_8566,N_7968);
xor U10239 (N_10239,N_7802,N_8296);
and U10240 (N_10240,N_7733,N_8902);
or U10241 (N_10241,N_8176,N_7712);
or U10242 (N_10242,N_8620,N_7869);
and U10243 (N_10243,N_8765,N_8969);
or U10244 (N_10244,N_7857,N_8505);
nand U10245 (N_10245,N_7704,N_7565);
nor U10246 (N_10246,N_8039,N_8064);
and U10247 (N_10247,N_7782,N_8204);
nand U10248 (N_10248,N_8972,N_8901);
and U10249 (N_10249,N_7500,N_7702);
nand U10250 (N_10250,N_8583,N_8972);
nand U10251 (N_10251,N_8981,N_7786);
nor U10252 (N_10252,N_8851,N_8653);
or U10253 (N_10253,N_8136,N_8544);
or U10254 (N_10254,N_8275,N_7796);
nor U10255 (N_10255,N_7554,N_8231);
nand U10256 (N_10256,N_7655,N_8948);
nand U10257 (N_10257,N_8656,N_8575);
nand U10258 (N_10258,N_7925,N_8941);
xor U10259 (N_10259,N_8226,N_7685);
and U10260 (N_10260,N_7690,N_7669);
or U10261 (N_10261,N_8629,N_7901);
nand U10262 (N_10262,N_7890,N_8892);
nor U10263 (N_10263,N_8028,N_8955);
nor U10264 (N_10264,N_8512,N_8196);
and U10265 (N_10265,N_8140,N_8607);
nand U10266 (N_10266,N_8519,N_8181);
and U10267 (N_10267,N_8138,N_7742);
and U10268 (N_10268,N_8337,N_8282);
nand U10269 (N_10269,N_8012,N_8597);
and U10270 (N_10270,N_7569,N_8419);
nand U10271 (N_10271,N_7967,N_7508);
xor U10272 (N_10272,N_7645,N_8497);
nand U10273 (N_10273,N_8707,N_8048);
xor U10274 (N_10274,N_7508,N_8717);
nor U10275 (N_10275,N_8377,N_8841);
nand U10276 (N_10276,N_8255,N_8943);
or U10277 (N_10277,N_7967,N_8354);
xnor U10278 (N_10278,N_8998,N_8899);
and U10279 (N_10279,N_8993,N_7778);
nand U10280 (N_10280,N_8753,N_7577);
and U10281 (N_10281,N_8205,N_8710);
and U10282 (N_10282,N_8044,N_8331);
nor U10283 (N_10283,N_8444,N_7973);
nand U10284 (N_10284,N_8644,N_8808);
nand U10285 (N_10285,N_8225,N_8482);
or U10286 (N_10286,N_7586,N_8267);
nand U10287 (N_10287,N_8871,N_8406);
nand U10288 (N_10288,N_8266,N_7633);
nand U10289 (N_10289,N_8840,N_8209);
or U10290 (N_10290,N_7988,N_7833);
nor U10291 (N_10291,N_7660,N_8098);
and U10292 (N_10292,N_7749,N_7835);
nor U10293 (N_10293,N_8321,N_7967);
nor U10294 (N_10294,N_8392,N_8196);
nand U10295 (N_10295,N_8907,N_8183);
or U10296 (N_10296,N_7773,N_8204);
and U10297 (N_10297,N_8047,N_8132);
or U10298 (N_10298,N_7948,N_8367);
nor U10299 (N_10299,N_8386,N_8960);
and U10300 (N_10300,N_7968,N_7604);
nor U10301 (N_10301,N_7989,N_8807);
or U10302 (N_10302,N_7763,N_7995);
or U10303 (N_10303,N_8199,N_8373);
or U10304 (N_10304,N_8529,N_8422);
nand U10305 (N_10305,N_7866,N_8964);
and U10306 (N_10306,N_8185,N_8683);
or U10307 (N_10307,N_8941,N_8719);
or U10308 (N_10308,N_8733,N_8515);
and U10309 (N_10309,N_8459,N_8859);
and U10310 (N_10310,N_7933,N_8079);
nor U10311 (N_10311,N_8823,N_8119);
nor U10312 (N_10312,N_8273,N_7731);
and U10313 (N_10313,N_8296,N_8005);
or U10314 (N_10314,N_8785,N_8524);
xnor U10315 (N_10315,N_7588,N_8720);
or U10316 (N_10316,N_8684,N_8174);
or U10317 (N_10317,N_8777,N_8582);
nand U10318 (N_10318,N_8185,N_8788);
nand U10319 (N_10319,N_8361,N_7689);
or U10320 (N_10320,N_8048,N_8115);
or U10321 (N_10321,N_8135,N_8435);
or U10322 (N_10322,N_8116,N_8954);
or U10323 (N_10323,N_7729,N_8840);
and U10324 (N_10324,N_8442,N_8826);
or U10325 (N_10325,N_8679,N_8445);
nand U10326 (N_10326,N_8831,N_8545);
or U10327 (N_10327,N_8378,N_7814);
nand U10328 (N_10328,N_8466,N_8582);
nor U10329 (N_10329,N_7715,N_8729);
or U10330 (N_10330,N_7565,N_8652);
or U10331 (N_10331,N_8639,N_7551);
nor U10332 (N_10332,N_8235,N_8190);
nand U10333 (N_10333,N_8687,N_8757);
or U10334 (N_10334,N_8916,N_8566);
nor U10335 (N_10335,N_8150,N_7667);
and U10336 (N_10336,N_8486,N_8808);
or U10337 (N_10337,N_8605,N_8237);
nor U10338 (N_10338,N_8632,N_8058);
nor U10339 (N_10339,N_8282,N_8108);
and U10340 (N_10340,N_8400,N_7563);
nor U10341 (N_10341,N_7682,N_8650);
xor U10342 (N_10342,N_8672,N_8558);
or U10343 (N_10343,N_8902,N_8275);
xnor U10344 (N_10344,N_8874,N_8841);
and U10345 (N_10345,N_8496,N_7839);
or U10346 (N_10346,N_8735,N_7940);
nor U10347 (N_10347,N_7889,N_8775);
nor U10348 (N_10348,N_8144,N_8973);
nand U10349 (N_10349,N_8130,N_8916);
or U10350 (N_10350,N_8563,N_8009);
nand U10351 (N_10351,N_7617,N_8411);
or U10352 (N_10352,N_8795,N_8129);
and U10353 (N_10353,N_8976,N_8172);
nor U10354 (N_10354,N_8550,N_8776);
or U10355 (N_10355,N_7778,N_7827);
and U10356 (N_10356,N_8308,N_8360);
nand U10357 (N_10357,N_8623,N_8010);
or U10358 (N_10358,N_8469,N_8946);
or U10359 (N_10359,N_7591,N_7623);
xnor U10360 (N_10360,N_8516,N_7942);
nor U10361 (N_10361,N_7668,N_8145);
nand U10362 (N_10362,N_7897,N_8404);
and U10363 (N_10363,N_8816,N_7914);
nand U10364 (N_10364,N_7931,N_8026);
or U10365 (N_10365,N_8364,N_8242);
and U10366 (N_10366,N_7550,N_8213);
and U10367 (N_10367,N_8241,N_7805);
and U10368 (N_10368,N_7941,N_8291);
nor U10369 (N_10369,N_8394,N_7846);
or U10370 (N_10370,N_7768,N_8006);
or U10371 (N_10371,N_8417,N_7813);
nor U10372 (N_10372,N_8192,N_7692);
nor U10373 (N_10373,N_8461,N_7743);
nor U10374 (N_10374,N_8022,N_8164);
or U10375 (N_10375,N_8459,N_7935);
and U10376 (N_10376,N_7786,N_8985);
nand U10377 (N_10377,N_7528,N_7857);
nor U10378 (N_10378,N_8138,N_8491);
nand U10379 (N_10379,N_8501,N_8555);
xor U10380 (N_10380,N_8452,N_7634);
and U10381 (N_10381,N_8517,N_7575);
nand U10382 (N_10382,N_8098,N_7501);
nor U10383 (N_10383,N_8501,N_8023);
or U10384 (N_10384,N_8853,N_7697);
nor U10385 (N_10385,N_8134,N_8159);
or U10386 (N_10386,N_8704,N_8289);
nor U10387 (N_10387,N_8636,N_7740);
xnor U10388 (N_10388,N_8602,N_7839);
and U10389 (N_10389,N_7705,N_8272);
or U10390 (N_10390,N_7771,N_8663);
and U10391 (N_10391,N_8204,N_8822);
xnor U10392 (N_10392,N_7539,N_8212);
and U10393 (N_10393,N_7626,N_7974);
nand U10394 (N_10394,N_7784,N_7948);
xnor U10395 (N_10395,N_7898,N_8739);
nor U10396 (N_10396,N_8018,N_7651);
or U10397 (N_10397,N_7745,N_8629);
and U10398 (N_10398,N_8439,N_8451);
or U10399 (N_10399,N_7924,N_7823);
xor U10400 (N_10400,N_8976,N_8241);
nand U10401 (N_10401,N_7627,N_8877);
nand U10402 (N_10402,N_7753,N_8093);
nand U10403 (N_10403,N_8628,N_7823);
nand U10404 (N_10404,N_7804,N_8329);
xnor U10405 (N_10405,N_8591,N_7793);
nor U10406 (N_10406,N_8228,N_8924);
or U10407 (N_10407,N_8352,N_8027);
nand U10408 (N_10408,N_8084,N_8267);
nand U10409 (N_10409,N_8857,N_7761);
or U10410 (N_10410,N_7773,N_7620);
xnor U10411 (N_10411,N_8070,N_8506);
xor U10412 (N_10412,N_8151,N_7738);
or U10413 (N_10413,N_7814,N_8494);
nand U10414 (N_10414,N_8350,N_8684);
or U10415 (N_10415,N_8678,N_8336);
or U10416 (N_10416,N_7762,N_8825);
or U10417 (N_10417,N_7840,N_7733);
or U10418 (N_10418,N_8171,N_8542);
nor U10419 (N_10419,N_8640,N_8786);
xnor U10420 (N_10420,N_8203,N_8425);
or U10421 (N_10421,N_8450,N_7749);
nor U10422 (N_10422,N_7882,N_8533);
and U10423 (N_10423,N_7704,N_8111);
or U10424 (N_10424,N_8845,N_7600);
nand U10425 (N_10425,N_8856,N_7665);
and U10426 (N_10426,N_8178,N_8883);
or U10427 (N_10427,N_8936,N_8083);
and U10428 (N_10428,N_7665,N_8571);
nand U10429 (N_10429,N_8665,N_8138);
nor U10430 (N_10430,N_8028,N_8211);
or U10431 (N_10431,N_7504,N_8468);
nand U10432 (N_10432,N_8492,N_8314);
and U10433 (N_10433,N_8878,N_8746);
or U10434 (N_10434,N_7877,N_8018);
nand U10435 (N_10435,N_7863,N_8612);
and U10436 (N_10436,N_8967,N_8767);
nor U10437 (N_10437,N_7509,N_7517);
nor U10438 (N_10438,N_7707,N_8313);
and U10439 (N_10439,N_8940,N_7755);
nor U10440 (N_10440,N_8678,N_8594);
or U10441 (N_10441,N_7849,N_7554);
nor U10442 (N_10442,N_8935,N_8604);
nand U10443 (N_10443,N_8240,N_8345);
and U10444 (N_10444,N_7741,N_8054);
or U10445 (N_10445,N_8341,N_8919);
xor U10446 (N_10446,N_8456,N_8689);
nand U10447 (N_10447,N_8816,N_8220);
nor U10448 (N_10448,N_7631,N_8843);
and U10449 (N_10449,N_7897,N_8647);
nor U10450 (N_10450,N_8902,N_8886);
or U10451 (N_10451,N_8266,N_7908);
nor U10452 (N_10452,N_8800,N_7663);
nand U10453 (N_10453,N_7571,N_7556);
nand U10454 (N_10454,N_8117,N_8880);
or U10455 (N_10455,N_7887,N_8974);
and U10456 (N_10456,N_7884,N_8499);
nand U10457 (N_10457,N_8978,N_7550);
nor U10458 (N_10458,N_8671,N_7603);
nand U10459 (N_10459,N_8027,N_7852);
nand U10460 (N_10460,N_8285,N_7593);
or U10461 (N_10461,N_8664,N_8704);
and U10462 (N_10462,N_8244,N_8918);
xor U10463 (N_10463,N_7717,N_8014);
xor U10464 (N_10464,N_7541,N_8215);
nor U10465 (N_10465,N_8587,N_8767);
and U10466 (N_10466,N_8059,N_8692);
xnor U10467 (N_10467,N_7913,N_7888);
or U10468 (N_10468,N_8773,N_7567);
nand U10469 (N_10469,N_7836,N_7677);
and U10470 (N_10470,N_8468,N_8486);
and U10471 (N_10471,N_8761,N_8010);
and U10472 (N_10472,N_7704,N_7765);
nand U10473 (N_10473,N_8983,N_8595);
nor U10474 (N_10474,N_8350,N_8484);
and U10475 (N_10475,N_7813,N_8519);
nor U10476 (N_10476,N_7963,N_8161);
nor U10477 (N_10477,N_8119,N_8465);
xnor U10478 (N_10478,N_8745,N_7519);
or U10479 (N_10479,N_8325,N_8404);
nand U10480 (N_10480,N_8879,N_8026);
or U10481 (N_10481,N_8152,N_8917);
xor U10482 (N_10482,N_8859,N_8655);
and U10483 (N_10483,N_8482,N_7895);
nand U10484 (N_10484,N_7543,N_7614);
nor U10485 (N_10485,N_8115,N_7615);
and U10486 (N_10486,N_8466,N_8553);
or U10487 (N_10487,N_8112,N_8456);
and U10488 (N_10488,N_7836,N_8099);
nand U10489 (N_10489,N_8504,N_8571);
or U10490 (N_10490,N_7764,N_7930);
nor U10491 (N_10491,N_7632,N_7523);
nand U10492 (N_10492,N_7780,N_8218);
and U10493 (N_10493,N_8069,N_7971);
and U10494 (N_10494,N_8197,N_8378);
xnor U10495 (N_10495,N_7997,N_8296);
xnor U10496 (N_10496,N_8593,N_8415);
or U10497 (N_10497,N_8464,N_7955);
nor U10498 (N_10498,N_7903,N_8032);
nor U10499 (N_10499,N_8298,N_7679);
xor U10500 (N_10500,N_9240,N_9493);
nor U10501 (N_10501,N_10344,N_9442);
and U10502 (N_10502,N_10268,N_9817);
nor U10503 (N_10503,N_9794,N_10010);
or U10504 (N_10504,N_9754,N_9025);
or U10505 (N_10505,N_9707,N_9980);
nor U10506 (N_10506,N_10432,N_9294);
nor U10507 (N_10507,N_9168,N_9462);
or U10508 (N_10508,N_9313,N_9227);
nand U10509 (N_10509,N_9247,N_10262);
nand U10510 (N_10510,N_9795,N_9407);
and U10511 (N_10511,N_9164,N_10365);
nand U10512 (N_10512,N_10032,N_10078);
or U10513 (N_10513,N_10310,N_9360);
nor U10514 (N_10514,N_10098,N_9619);
nand U10515 (N_10515,N_9200,N_10158);
nor U10516 (N_10516,N_9455,N_9638);
or U10517 (N_10517,N_9956,N_10141);
and U10518 (N_10518,N_9554,N_9774);
nor U10519 (N_10519,N_9976,N_9665);
nand U10520 (N_10520,N_9295,N_9464);
and U10521 (N_10521,N_9426,N_9381);
nor U10522 (N_10522,N_10205,N_10222);
xor U10523 (N_10523,N_9822,N_9005);
nor U10524 (N_10524,N_10146,N_10194);
nor U10525 (N_10525,N_10248,N_9081);
or U10526 (N_10526,N_10300,N_9618);
nand U10527 (N_10527,N_9220,N_10221);
xor U10528 (N_10528,N_9978,N_9050);
and U10529 (N_10529,N_9262,N_9955);
or U10530 (N_10530,N_9226,N_9608);
nand U10531 (N_10531,N_10220,N_10293);
xnor U10532 (N_10532,N_9899,N_9655);
nand U10533 (N_10533,N_10337,N_10108);
and U10534 (N_10534,N_10465,N_9744);
or U10535 (N_10535,N_9008,N_9931);
nand U10536 (N_10536,N_9234,N_10253);
nand U10537 (N_10537,N_9031,N_10499);
xnor U10538 (N_10538,N_9743,N_9191);
nand U10539 (N_10539,N_9156,N_9596);
or U10540 (N_10540,N_10476,N_9965);
and U10541 (N_10541,N_9892,N_9528);
or U10542 (N_10542,N_9350,N_9130);
and U10543 (N_10543,N_9867,N_9022);
and U10544 (N_10544,N_9376,N_10368);
or U10545 (N_10545,N_9945,N_10087);
nand U10546 (N_10546,N_10382,N_10345);
xnor U10547 (N_10547,N_9370,N_9861);
nand U10548 (N_10548,N_9809,N_10256);
nor U10549 (N_10549,N_9369,N_9662);
nor U10550 (N_10550,N_9241,N_9679);
nand U10551 (N_10551,N_10030,N_10053);
or U10552 (N_10552,N_10112,N_9446);
nor U10553 (N_10553,N_9645,N_9209);
xor U10554 (N_10554,N_10131,N_9391);
nor U10555 (N_10555,N_10188,N_10326);
nor U10556 (N_10556,N_10213,N_9538);
xnor U10557 (N_10557,N_9524,N_9384);
and U10558 (N_10558,N_9626,N_9045);
and U10559 (N_10559,N_10464,N_9102);
xnor U10560 (N_10560,N_9534,N_9912);
or U10561 (N_10561,N_9838,N_9257);
or U10562 (N_10562,N_9552,N_9733);
and U10563 (N_10563,N_9246,N_9946);
and U10564 (N_10564,N_9006,N_9950);
or U10565 (N_10565,N_9553,N_9195);
nand U10566 (N_10566,N_9488,N_9132);
and U10567 (N_10567,N_9884,N_9482);
nand U10568 (N_10568,N_9516,N_9802);
nand U10569 (N_10569,N_9398,N_9400);
nor U10570 (N_10570,N_9985,N_10050);
nor U10571 (N_10571,N_9727,N_10116);
or U10572 (N_10572,N_9518,N_9934);
or U10573 (N_10573,N_9305,N_9916);
or U10574 (N_10574,N_10471,N_9219);
or U10575 (N_10575,N_10265,N_10289);
nor U10576 (N_10576,N_9009,N_10283);
or U10577 (N_10577,N_9770,N_9366);
or U10578 (N_10578,N_9541,N_10034);
and U10579 (N_10579,N_9768,N_9917);
nand U10580 (N_10580,N_9993,N_10057);
or U10581 (N_10581,N_9954,N_9077);
nand U10582 (N_10582,N_10139,N_10443);
nand U10583 (N_10583,N_10360,N_10343);
or U10584 (N_10584,N_10099,N_9877);
or U10585 (N_10585,N_9859,N_10356);
or U10586 (N_10586,N_9688,N_9204);
nor U10587 (N_10587,N_9601,N_9145);
and U10588 (N_10588,N_9091,N_9735);
nand U10589 (N_10589,N_9344,N_10008);
xnor U10590 (N_10590,N_9000,N_9352);
and U10591 (N_10591,N_10298,N_10025);
or U10592 (N_10592,N_10318,N_9378);
nand U10593 (N_10593,N_9717,N_9166);
or U10594 (N_10594,N_10328,N_10439);
and U10595 (N_10595,N_10269,N_9897);
or U10596 (N_10596,N_9756,N_10279);
and U10597 (N_10597,N_10460,N_9825);
and U10598 (N_10598,N_9469,N_10294);
and U10599 (N_10599,N_9926,N_9107);
and U10600 (N_10600,N_10355,N_9104);
or U10601 (N_10601,N_9289,N_9757);
nand U10602 (N_10602,N_9497,N_9372);
and U10603 (N_10603,N_9279,N_9371);
and U10604 (N_10604,N_10377,N_9751);
and U10605 (N_10605,N_9876,N_9064);
or U10606 (N_10606,N_10065,N_9712);
nor U10607 (N_10607,N_10118,N_10215);
nor U10608 (N_10608,N_9066,N_9543);
nand U10609 (N_10609,N_9745,N_9832);
nor U10610 (N_10610,N_9988,N_9141);
nor U10611 (N_10611,N_9823,N_10123);
and U10612 (N_10612,N_9821,N_9737);
xnor U10613 (N_10613,N_9715,N_9100);
xnor U10614 (N_10614,N_9728,N_9292);
and U10615 (N_10615,N_9748,N_10170);
nor U10616 (N_10616,N_10047,N_9870);
and U10617 (N_10617,N_10031,N_10081);
or U10618 (N_10618,N_9076,N_10358);
and U10619 (N_10619,N_10136,N_9167);
xor U10620 (N_10620,N_9547,N_9682);
or U10621 (N_10621,N_9374,N_9758);
and U10622 (N_10622,N_9033,N_9653);
or U10623 (N_10623,N_9694,N_9845);
nor U10624 (N_10624,N_10223,N_9478);
and U10625 (N_10625,N_10304,N_9095);
and U10626 (N_10626,N_10095,N_9385);
nand U10627 (N_10627,N_9559,N_9544);
and U10628 (N_10628,N_9625,N_10245);
and U10629 (N_10629,N_10416,N_10387);
nor U10630 (N_10630,N_9452,N_9264);
xor U10631 (N_10631,N_9448,N_10373);
xnor U10632 (N_10632,N_10378,N_10309);
and U10633 (N_10633,N_10074,N_9730);
nor U10634 (N_10634,N_9176,N_9904);
nor U10635 (N_10635,N_10453,N_9222);
or U10636 (N_10636,N_10391,N_9447);
and U10637 (N_10637,N_9738,N_10092);
nand U10638 (N_10638,N_9185,N_10012);
nand U10639 (N_10639,N_10054,N_9018);
nor U10640 (N_10640,N_10086,N_9969);
or U10641 (N_10641,N_10428,N_10437);
nor U10642 (N_10642,N_9036,N_9542);
nor U10643 (N_10643,N_9550,N_9153);
and U10644 (N_10644,N_10473,N_9392);
nor U10645 (N_10645,N_9819,N_9722);
or U10646 (N_10646,N_10442,N_10048);
nor U10647 (N_10647,N_9138,N_10462);
and U10648 (N_10648,N_9397,N_9115);
and U10649 (N_10649,N_9431,N_9129);
xnor U10650 (N_10650,N_9919,N_9517);
nand U10651 (N_10651,N_10258,N_9466);
or U10652 (N_10652,N_10291,N_10064);
or U10653 (N_10653,N_9752,N_9918);
or U10654 (N_10654,N_10470,N_9749);
or U10655 (N_10655,N_9539,N_10229);
nand U10656 (N_10656,N_9726,N_10184);
nand U10657 (N_10657,N_9231,N_9046);
or U10658 (N_10658,N_10083,N_10135);
and U10659 (N_10659,N_9967,N_10371);
and U10660 (N_10660,N_9428,N_9580);
nand U10661 (N_10661,N_9713,N_10255);
nand U10662 (N_10662,N_9984,N_9315);
nor U10663 (N_10663,N_10409,N_9327);
and U10664 (N_10664,N_9072,N_10257);
nor U10665 (N_10665,N_10426,N_9074);
nor U10666 (N_10666,N_10002,N_9276);
or U10667 (N_10667,N_9729,N_10125);
and U10668 (N_10668,N_9778,N_9406);
xor U10669 (N_10669,N_10185,N_9948);
or U10670 (N_10670,N_9113,N_9287);
xnor U10671 (N_10671,N_10142,N_10094);
and U10672 (N_10672,N_9724,N_9925);
nor U10673 (N_10673,N_9101,N_9684);
xnor U10674 (N_10674,N_10227,N_10466);
nand U10675 (N_10675,N_10488,N_10261);
xnor U10676 (N_10676,N_9924,N_10477);
nand U10677 (N_10677,N_10204,N_10237);
xor U10678 (N_10678,N_9439,N_9092);
nand U10679 (N_10679,N_10082,N_9816);
and U10680 (N_10680,N_9023,N_9930);
or U10681 (N_10681,N_9911,N_10354);
nand U10682 (N_10682,N_9964,N_10189);
and U10683 (N_10683,N_10085,N_9300);
xor U10684 (N_10684,N_9210,N_10329);
nor U10685 (N_10685,N_10070,N_10276);
or U10686 (N_10686,N_9284,N_9208);
and U10687 (N_10687,N_10015,N_9977);
nor U10688 (N_10688,N_10212,N_9927);
or U10689 (N_10689,N_9048,N_10383);
nand U10690 (N_10690,N_9971,N_9974);
and U10691 (N_10691,N_9936,N_10167);
xor U10692 (N_10692,N_9150,N_9237);
nor U10693 (N_10693,N_10376,N_9499);
xnor U10694 (N_10694,N_10180,N_9882);
nor U10695 (N_10695,N_9110,N_9806);
nor U10696 (N_10696,N_10066,N_10441);
and U10697 (N_10697,N_9913,N_10100);
xor U10698 (N_10698,N_10068,N_9419);
or U10699 (N_10699,N_9044,N_9606);
nor U10700 (N_10700,N_9531,N_9982);
nand U10701 (N_10701,N_10290,N_9014);
and U10702 (N_10702,N_9786,N_9671);
and U10703 (N_10703,N_10422,N_10270);
nor U10704 (N_10704,N_9557,N_9122);
nand U10705 (N_10705,N_9375,N_9835);
nor U10706 (N_10706,N_10132,N_9860);
nand U10707 (N_10707,N_9286,N_10021);
or U10708 (N_10708,N_10487,N_10338);
nand U10709 (N_10709,N_10312,N_9769);
and U10710 (N_10710,N_9960,N_9560);
and U10711 (N_10711,N_9124,N_10244);
nor U10712 (N_10712,N_9634,N_10127);
or U10713 (N_10713,N_9187,N_9169);
and U10714 (N_10714,N_10263,N_9864);
and U10715 (N_10715,N_9915,N_10105);
or U10716 (N_10716,N_10250,N_9624);
and U10717 (N_10717,N_9900,N_9736);
nand U10718 (N_10718,N_9181,N_10148);
nor U10719 (N_10719,N_10023,N_9088);
or U10720 (N_10720,N_9647,N_10498);
nor U10721 (N_10721,N_9432,N_9165);
and U10722 (N_10722,N_10389,N_9999);
xnor U10723 (N_10723,N_9760,N_10101);
nor U10724 (N_10724,N_10496,N_9855);
nor U10725 (N_10725,N_9986,N_10201);
and U10726 (N_10726,N_10115,N_9781);
or U10727 (N_10727,N_9693,N_10072);
nand U10728 (N_10728,N_9609,N_9274);
or U10729 (N_10729,N_10363,N_9377);
nor U10730 (N_10730,N_10140,N_9330);
and U10731 (N_10731,N_10181,N_9896);
nor U10732 (N_10732,N_10342,N_9277);
and U10733 (N_10733,N_10489,N_9603);
nand U10734 (N_10734,N_9335,N_10479);
nand U10735 (N_10735,N_9898,N_9467);
nor U10736 (N_10736,N_10417,N_9863);
or U10737 (N_10737,N_9329,N_10412);
xnor U10738 (N_10738,N_9318,N_10052);
nand U10739 (N_10739,N_10306,N_9650);
and U10740 (N_10740,N_9765,N_10176);
nand U10741 (N_10741,N_9221,N_9889);
and U10742 (N_10742,N_9687,N_9905);
nand U10743 (N_10743,N_10285,N_10120);
nand U10744 (N_10744,N_9629,N_9255);
xnor U10745 (N_10745,N_10423,N_9112);
and U10746 (N_10746,N_9854,N_10159);
nor U10747 (N_10747,N_9678,N_10339);
nor U10748 (N_10748,N_9079,N_9086);
nor U10749 (N_10749,N_10350,N_9456);
nor U10750 (N_10750,N_10286,N_9034);
and U10751 (N_10751,N_9716,N_9970);
or U10752 (N_10752,N_9062,N_10395);
nand U10753 (N_10753,N_9139,N_9013);
xnor U10754 (N_10754,N_10454,N_9811);
nor U10755 (N_10755,N_9703,N_9633);
nor U10756 (N_10756,N_9268,N_9987);
nand U10757 (N_10757,N_9979,N_9024);
nor U10758 (N_10758,N_9394,N_9672);
nor U10759 (N_10759,N_9026,N_9607);
xor U10760 (N_10760,N_10450,N_9235);
or U10761 (N_10761,N_9157,N_9324);
or U10762 (N_10762,N_9422,N_9109);
nor U10763 (N_10763,N_9353,N_10491);
xor U10764 (N_10764,N_10388,N_9020);
nand U10765 (N_10765,N_10203,N_10129);
or U10766 (N_10766,N_9218,N_10156);
nor U10767 (N_10767,N_10234,N_9496);
or U10768 (N_10768,N_9868,N_9293);
or U10769 (N_10769,N_9820,N_9498);
nor U10770 (N_10770,N_9767,N_9742);
and U10771 (N_10771,N_9399,N_9995);
xnor U10772 (N_10772,N_10169,N_9942);
nor U10773 (N_10773,N_10497,N_9520);
nand U10774 (N_10774,N_9951,N_9258);
nor U10775 (N_10775,N_9303,N_9395);
or U10776 (N_10776,N_10003,N_10027);
or U10777 (N_10777,N_9622,N_9839);
nand U10778 (N_10778,N_9105,N_10447);
nand U10779 (N_10779,N_10214,N_10469);
nand U10780 (N_10780,N_9198,N_10102);
and U10781 (N_10781,N_9908,N_9764);
nand U10782 (N_10782,N_9322,N_9089);
nand U10783 (N_10783,N_9362,N_10061);
or U10784 (N_10784,N_10278,N_9850);
or U10785 (N_10785,N_10133,N_10024);
nor U10786 (N_10786,N_9460,N_9789);
nor U10787 (N_10787,N_9163,N_10448);
and U10788 (N_10788,N_10352,N_9572);
xnor U10789 (N_10789,N_10492,N_9595);
or U10790 (N_10790,N_10226,N_9858);
nor U10791 (N_10791,N_9364,N_9762);
or U10792 (N_10792,N_10045,N_9367);
or U10793 (N_10793,N_9570,N_10224);
nand U10794 (N_10794,N_10317,N_9245);
nand U10795 (N_10795,N_9224,N_9785);
xor U10796 (N_10796,N_9127,N_10347);
nor U10797 (N_10797,N_10458,N_9578);
or U10798 (N_10798,N_9510,N_9337);
or U10799 (N_10799,N_10230,N_9990);
and U10800 (N_10800,N_10379,N_9312);
nor U10801 (N_10801,N_10266,N_10375);
or U10802 (N_10802,N_10399,N_9686);
nand U10803 (N_10803,N_9797,N_9575);
nand U10804 (N_10804,N_9963,N_10316);
nand U10805 (N_10805,N_10468,N_10006);
and U10806 (N_10806,N_9471,N_9283);
nor U10807 (N_10807,N_9067,N_9644);
or U10808 (N_10808,N_10218,N_9470);
and U10809 (N_10809,N_9847,N_10076);
and U10810 (N_10810,N_9555,N_9953);
or U10811 (N_10811,N_10461,N_9481);
or U10812 (N_10812,N_9673,N_9012);
nor U10813 (N_10813,N_9815,N_10055);
nand U10814 (N_10814,N_10071,N_9804);
and U10815 (N_10815,N_9676,N_10036);
nor U10816 (N_10816,N_9959,N_10327);
nor U10817 (N_10817,N_9415,N_9143);
and U10818 (N_10818,N_10348,N_10434);
or U10819 (N_10819,N_9389,N_9589);
and U10820 (N_10820,N_9457,N_10151);
xor U10821 (N_10821,N_10109,N_10445);
or U10822 (N_10822,N_10424,N_10037);
and U10823 (N_10823,N_10119,N_10475);
and U10824 (N_10824,N_9853,N_9007);
xor U10825 (N_10825,N_9865,N_10333);
xnor U10826 (N_10826,N_10264,N_9800);
xnor U10827 (N_10827,N_9142,N_9938);
nor U10828 (N_10828,N_9773,N_10152);
nor U10829 (N_10829,N_9306,N_10200);
nor U10830 (N_10830,N_10177,N_10367);
xor U10831 (N_10831,N_10126,N_9961);
and U10832 (N_10832,N_9051,N_10155);
nand U10833 (N_10833,N_9004,N_9373);
and U10834 (N_10834,N_9309,N_10486);
nand U10835 (N_10835,N_10208,N_9801);
xor U10836 (N_10836,N_9906,N_9252);
xor U10837 (N_10837,N_9197,N_9910);
xor U10838 (N_10838,N_10398,N_9331);
nand U10839 (N_10839,N_9347,N_9273);
nand U10840 (N_10840,N_9871,N_10251);
or U10841 (N_10841,N_10372,N_10396);
and U10842 (N_10842,N_9502,N_10104);
nor U10843 (N_10843,N_9651,N_10038);
or U10844 (N_10844,N_9849,N_10273);
xnor U10845 (N_10845,N_9179,N_9957);
and U10846 (N_10846,N_9521,N_10103);
nand U10847 (N_10847,N_9939,N_9584);
and U10848 (N_10848,N_9483,N_9424);
nand U10849 (N_10849,N_9216,N_10084);
nand U10850 (N_10850,N_9551,N_10319);
and U10851 (N_10851,N_10485,N_10259);
nor U10852 (N_10852,N_9567,N_9094);
and U10853 (N_10853,N_10191,N_10483);
or U10854 (N_10854,N_9404,N_10403);
xor U10855 (N_10855,N_10418,N_10287);
xor U10856 (N_10856,N_10435,N_10160);
nand U10857 (N_10857,N_10392,N_10178);
and U10858 (N_10858,N_10331,N_9003);
or U10859 (N_10859,N_9652,N_10157);
nor U10860 (N_10860,N_10228,N_9788);
and U10861 (N_10861,N_10444,N_9830);
and U10862 (N_10862,N_9160,N_9747);
nor U10863 (N_10863,N_9328,N_9253);
or U10864 (N_10864,N_10411,N_10239);
xor U10865 (N_10865,N_9706,N_9387);
xor U10866 (N_10866,N_10494,N_9732);
xnor U10867 (N_10867,N_9523,N_9958);
nor U10868 (N_10868,N_10039,N_9453);
nor U10869 (N_10869,N_10202,N_9581);
or U10870 (N_10870,N_9261,N_9154);
nand U10871 (N_10871,N_9791,N_9290);
nor U10872 (N_10872,N_9648,N_9405);
and U10873 (N_10873,N_9296,N_9621);
nand U10874 (N_10874,N_9674,N_10011);
nand U10875 (N_10875,N_9082,N_9841);
and U10876 (N_10876,N_9776,N_9714);
xnor U10877 (N_10877,N_10145,N_9813);
nor U10878 (N_10878,N_9075,N_9450);
nor U10879 (N_10879,N_10014,N_9338);
nand U10880 (N_10880,N_9734,N_9069);
or U10881 (N_10881,N_9172,N_9631);
nor U10882 (N_10882,N_10022,N_10236);
nor U10883 (N_10883,N_9097,N_9879);
nand U10884 (N_10884,N_9561,N_9772);
or U10885 (N_10885,N_10183,N_10190);
and U10886 (N_10886,N_9039,N_9994);
and U10887 (N_10887,N_9472,N_9001);
and U10888 (N_10888,N_10438,N_9530);
nor U10889 (N_10889,N_9015,N_10277);
nand U10890 (N_10890,N_9205,N_9212);
nand U10891 (N_10891,N_10370,N_10182);
or U10892 (N_10892,N_10400,N_10062);
or U10893 (N_10893,N_10361,N_9201);
and U10894 (N_10894,N_9443,N_9875);
xor U10895 (N_10895,N_9342,N_9620);
or U10896 (N_10896,N_10341,N_9536);
or U10897 (N_10897,N_9288,N_9746);
or U10898 (N_10898,N_9099,N_10474);
nor U10899 (N_10899,N_9623,N_9002);
and U10900 (N_10900,N_10324,N_10235);
and U10901 (N_10901,N_9412,N_9709);
and U10902 (N_10902,N_9857,N_10452);
xnor U10903 (N_10903,N_10246,N_10093);
nor U10904 (N_10904,N_10232,N_9512);
and U10905 (N_10905,N_9708,N_9040);
or U10906 (N_10906,N_9843,N_10493);
or U10907 (N_10907,N_10429,N_9435);
or U10908 (N_10908,N_10241,N_9616);
nor U10909 (N_10909,N_10330,N_9639);
xor U10910 (N_10910,N_10440,N_10134);
xor U10911 (N_10911,N_9509,N_9635);
nor U10912 (N_10912,N_10430,N_10394);
and U10913 (N_10913,N_9365,N_10254);
or U10914 (N_10914,N_9699,N_9689);
and U10915 (N_10915,N_9943,N_10427);
or U10916 (N_10916,N_9325,N_10238);
nor U10917 (N_10917,N_9149,N_9251);
nor U10918 (N_10918,N_9611,N_9041);
xnor U10919 (N_10919,N_9895,N_9304);
or U10920 (N_10920,N_9420,N_9458);
nand U10921 (N_10921,N_10097,N_9535);
nand U10922 (N_10922,N_9704,N_9133);
or U10923 (N_10923,N_10274,N_9213);
xor U10924 (N_10924,N_9571,N_9416);
nand U10925 (N_10925,N_9098,N_10449);
nand U10926 (N_10926,N_9463,N_9299);
or U10927 (N_10927,N_10280,N_9065);
nor U10928 (N_10928,N_10410,N_9361);
or U10929 (N_10929,N_9058,N_10028);
and U10930 (N_10930,N_10478,N_9232);
nand U10931 (N_10931,N_9357,N_9568);
nand U10932 (N_10932,N_9271,N_10163);
nor U10933 (N_10933,N_9604,N_9602);
or U10934 (N_10934,N_10351,N_9888);
or U10935 (N_10935,N_9011,N_10366);
nand U10936 (N_10936,N_9929,N_9920);
nand U10937 (N_10937,N_10436,N_9190);
xnor U10938 (N_10938,N_9828,N_9174);
and U10939 (N_10939,N_9390,N_9540);
nand U10940 (N_10940,N_10374,N_9940);
nor U10941 (N_10941,N_10079,N_10402);
nand U10942 (N_10942,N_10455,N_10359);
nor U10943 (N_10943,N_9787,N_9670);
nor U10944 (N_10944,N_9229,N_9627);
or U10945 (N_10945,N_9837,N_9529);
and U10946 (N_10946,N_10334,N_9332);
and U10947 (N_10947,N_9901,N_9562);
nor U10948 (N_10948,N_9675,N_9668);
nor U10949 (N_10949,N_9566,N_10346);
or U10950 (N_10950,N_9239,N_9016);
or U10951 (N_10951,N_10364,N_10325);
or U10952 (N_10952,N_9803,N_9844);
nor U10953 (N_10953,N_9848,N_9301);
nor U10954 (N_10954,N_9131,N_9386);
nand U10955 (N_10955,N_9125,N_9333);
nand U10956 (N_10956,N_9349,N_9585);
nand U10957 (N_10957,N_9574,N_10484);
nor U10958 (N_10958,N_9326,N_9495);
nand U10959 (N_10959,N_10164,N_9151);
xor U10960 (N_10960,N_10321,N_9401);
nand U10961 (N_10961,N_9739,N_9021);
nand U10962 (N_10962,N_9297,N_10490);
nand U10963 (N_10963,N_10090,N_9725);
and U10964 (N_10964,N_9032,N_9445);
nand U10965 (N_10965,N_10292,N_9383);
or U10966 (N_10966,N_10284,N_9549);
nand U10967 (N_10967,N_9840,N_10433);
xor U10968 (N_10968,N_10035,N_9178);
or U10969 (N_10969,N_10128,N_9949);
nand U10970 (N_10970,N_10405,N_9434);
nand U10971 (N_10971,N_9666,N_9577);
nand U10972 (N_10972,N_9027,N_9824);
nand U10973 (N_10973,N_9677,N_9196);
or U10974 (N_10974,N_9465,N_9272);
nand U10975 (N_10975,N_9641,N_10171);
nand U10976 (N_10976,N_10001,N_9056);
or U10977 (N_10977,N_9336,N_9880);
and U10978 (N_10978,N_9408,N_9887);
and U10979 (N_10979,N_9881,N_9720);
nor U10980 (N_10980,N_9454,N_9663);
xor U10981 (N_10981,N_9792,N_9852);
or U10982 (N_10982,N_9891,N_10275);
nor U10983 (N_10983,N_9507,N_9341);
and U10984 (N_10984,N_10089,N_9225);
or U10985 (N_10985,N_10282,N_9321);
nor U10986 (N_10986,N_9885,N_9661);
and U10987 (N_10987,N_10166,N_10174);
nand U10988 (N_10988,N_10481,N_10308);
nand U10989 (N_10989,N_9134,N_9108);
nand U10990 (N_10990,N_9238,N_10197);
nand U10991 (N_10991,N_9972,N_9159);
or U10992 (N_10992,N_10390,N_10029);
nor U10993 (N_10993,N_9563,N_9111);
and U10994 (N_10994,N_9614,N_10153);
xor U10995 (N_10995,N_9417,N_10063);
nand U10996 (N_10996,N_9490,N_10110);
or U10997 (N_10997,N_9263,N_10046);
nand U10998 (N_10998,N_10362,N_9872);
and U10999 (N_10999,N_9643,N_9579);
and U11000 (N_11000,N_9184,N_9140);
and U11001 (N_11001,N_9136,N_9669);
nand U11002 (N_11002,N_9211,N_9681);
nand U11003 (N_11003,N_9269,N_9266);
nor U11004 (N_11004,N_10196,N_9741);
nor U11005 (N_11005,N_9642,N_9701);
or U11006 (N_11006,N_9410,N_9186);
nand U11007 (N_11007,N_9937,N_9161);
xnor U11008 (N_11008,N_9117,N_9413);
xor U11009 (N_11009,N_10288,N_10480);
or U11010 (N_11010,N_9890,N_10467);
and U11011 (N_11011,N_9180,N_10172);
or U11012 (N_11012,N_10249,N_9106);
and U11013 (N_11013,N_9883,N_10240);
or U11014 (N_11014,N_10150,N_10380);
nand U11015 (N_11015,N_9846,N_9152);
nand U11016 (N_11016,N_10281,N_10207);
nor U11017 (N_11017,N_9474,N_10198);
nand U11018 (N_11018,N_9632,N_10162);
nor U11019 (N_11019,N_10143,N_10323);
and U11020 (N_11020,N_10414,N_9382);
or U11021 (N_11021,N_10311,N_9514);
nor U11022 (N_11022,N_9866,N_10091);
nand U11023 (N_11023,N_9944,N_10096);
nand U11024 (N_11024,N_10179,N_9265);
xor U11025 (N_11025,N_10017,N_10219);
nand U11026 (N_11026,N_9952,N_9340);
or U11027 (N_11027,N_10340,N_9545);
nand U11028 (N_11028,N_9418,N_9203);
and U11029 (N_11029,N_9060,N_9071);
and U11030 (N_11030,N_9148,N_9587);
nor U11031 (N_11031,N_9836,N_9719);
nand U11032 (N_11032,N_9894,N_9711);
nor U11033 (N_11033,N_10393,N_9078);
nand U11034 (N_11034,N_10385,N_10121);
and U11035 (N_11035,N_9637,N_9697);
and U11036 (N_11036,N_9975,N_9494);
nor U11037 (N_11037,N_10302,N_9981);
or U11038 (N_11038,N_9504,N_9921);
or U11039 (N_11039,N_9658,N_10408);
or U11040 (N_11040,N_9267,N_9307);
and U11041 (N_11041,N_10117,N_9194);
nand U11042 (N_11042,N_9030,N_9508);
and U11043 (N_11043,N_10124,N_9451);
nor U11044 (N_11044,N_10147,N_9433);
and U11045 (N_11045,N_9334,N_10233);
nor U11046 (N_11046,N_10168,N_10413);
nor U11047 (N_11047,N_10043,N_9615);
and U11048 (N_11048,N_10019,N_10463);
nor U11049 (N_11049,N_10080,N_9275);
nand U11050 (N_11050,N_9790,N_9317);
and U11051 (N_11051,N_9355,N_9487);
xor U11052 (N_11052,N_9636,N_9243);
or U11053 (N_11053,N_10020,N_10033);
or U11054 (N_11054,N_9548,N_9135);
nand U11055 (N_11055,N_9314,N_9522);
or U11056 (N_11056,N_9723,N_9437);
nor U11057 (N_11057,N_10457,N_10425);
and U11058 (N_11058,N_9755,N_9158);
xnor U11059 (N_11059,N_9468,N_9192);
nor U11060 (N_11060,N_9922,N_9368);
or U11061 (N_11061,N_9777,N_9348);
nor U11062 (N_11062,N_10161,N_9402);
xnor U11063 (N_11063,N_10210,N_9038);
nor U11064 (N_11064,N_9217,N_9526);
xor U11065 (N_11065,N_9799,N_9696);
xnor U11066 (N_11066,N_9775,N_10107);
nand U11067 (N_11067,N_9259,N_9617);
and U11068 (N_11068,N_10446,N_9807);
or U11069 (N_11069,N_9484,N_9783);
or U11070 (N_11070,N_9010,N_9515);
xnor U11071 (N_11071,N_9116,N_9228);
nand U11072 (N_11072,N_9233,N_9692);
or U11073 (N_11073,N_9278,N_9856);
or U11074 (N_11074,N_9147,N_9597);
nand U11075 (N_11075,N_10225,N_9533);
and U11076 (N_11076,N_9308,N_9319);
xnor U11077 (N_11077,N_9586,N_9281);
nor U11078 (N_11078,N_9793,N_10077);
xnor U11079 (N_11079,N_9182,N_9177);
nor U11080 (N_11080,N_9242,N_9998);
or U11081 (N_11081,N_9339,N_10186);
or U11082 (N_11082,N_9966,N_9814);
or U11083 (N_11083,N_10044,N_9146);
or U11084 (N_11084,N_9582,N_10459);
and U11085 (N_11085,N_9519,N_9605);
nand U11086 (N_11086,N_10252,N_10114);
or U11087 (N_11087,N_10013,N_9320);
or U11088 (N_11088,N_10336,N_10175);
and U11089 (N_11089,N_9403,N_9414);
xnor U11090 (N_11090,N_9479,N_9780);
nor U11091 (N_11091,N_9249,N_9808);
nor U11092 (N_11092,N_9096,N_9947);
nor U11093 (N_11093,N_9996,N_9396);
and U11094 (N_11094,N_10322,N_9411);
nor U11095 (N_11095,N_9093,N_10004);
and U11096 (N_11096,N_9667,N_9028);
or U11097 (N_11097,N_9311,N_9120);
xor U11098 (N_11098,N_9070,N_9763);
nor U11099 (N_11099,N_9119,N_10482);
nand U11100 (N_11100,N_9354,N_9254);
xnor U11101 (N_11101,N_9430,N_9527);
nor U11102 (N_11102,N_10067,N_9063);
and U11103 (N_11103,N_9175,N_9992);
or U11104 (N_11104,N_9649,N_10431);
or U11105 (N_11105,N_9834,N_10272);
nor U11106 (N_11106,N_9784,N_9812);
xnor U11107 (N_11107,N_9646,N_10407);
nor U11108 (N_11108,N_9680,N_9388);
or U11109 (N_11109,N_9427,N_9436);
or U11110 (N_11110,N_9236,N_9043);
and U11111 (N_11111,N_9114,N_9282);
and U11112 (N_11112,N_9591,N_10335);
and U11113 (N_11113,N_10173,N_9902);
or U11114 (N_11114,N_10267,N_9444);
nor U11115 (N_11115,N_10009,N_9590);
or U11116 (N_11116,N_10130,N_9080);
nand U11117 (N_11117,N_9761,N_10295);
and U11118 (N_11118,N_10051,N_10313);
or U11119 (N_11119,N_9423,N_9691);
or U11120 (N_11120,N_10386,N_9244);
or U11121 (N_11121,N_9962,N_9933);
or U11122 (N_11122,N_10243,N_9610);
nor U11123 (N_11123,N_9805,N_10122);
xor U11124 (N_11124,N_9084,N_10419);
xor U11125 (N_11125,N_10271,N_9476);
or U11126 (N_11126,N_9903,N_10073);
and U11127 (N_11127,N_10211,N_9118);
or U11128 (N_11128,N_9700,N_9029);
and U11129 (N_11129,N_9500,N_9505);
nor U11130 (N_11130,N_9298,N_9513);
nor U11131 (N_11131,N_9532,N_9486);
or U11132 (N_11132,N_9042,N_9057);
nor U11133 (N_11133,N_9593,N_9363);
and U11134 (N_11134,N_10192,N_10404);
nand U11135 (N_11135,N_9123,N_9558);
or U11136 (N_11136,N_9189,N_9055);
or U11137 (N_11137,N_10401,N_9656);
nor U11138 (N_11138,N_9600,N_9379);
nor U11139 (N_11139,N_9909,N_9049);
nand U11140 (N_11140,N_9260,N_9035);
or U11141 (N_11141,N_9766,N_9090);
and U11142 (N_11142,N_9199,N_9873);
and U11143 (N_11143,N_9053,N_9759);
nand U11144 (N_11144,N_9137,N_9771);
xnor U11145 (N_11145,N_9874,N_10397);
nor U11146 (N_11146,N_9556,N_9459);
xor U11147 (N_11147,N_9503,N_9842);
nand U11148 (N_11148,N_10314,N_9356);
nand U11149 (N_11149,N_10042,N_9183);
nand U11150 (N_11150,N_9907,N_9047);
nor U11151 (N_11151,N_9594,N_10420);
nor U11152 (N_11152,N_9968,N_9565);
nand U11153 (N_11153,N_10016,N_9997);
or U11154 (N_11154,N_9037,N_9475);
nor U11155 (N_11155,N_9660,N_10137);
nand U11156 (N_11156,N_10018,N_9818);
nand U11157 (N_11157,N_9973,N_9491);
and U11158 (N_11158,N_10113,N_10242);
nand U11159 (N_11159,N_9573,N_9878);
nor U11160 (N_11160,N_9473,N_10058);
or U11161 (N_11161,N_9511,N_9270);
and U11162 (N_11162,N_10421,N_9345);
and U11163 (N_11163,N_9731,N_9215);
or U11164 (N_11164,N_9054,N_9598);
nand U11165 (N_11165,N_10049,N_9128);
nor U11166 (N_11166,N_10000,N_9170);
nand U11167 (N_11167,N_9659,N_10187);
or U11168 (N_11168,N_9827,N_9438);
nor U11169 (N_11169,N_9302,N_9380);
nor U11170 (N_11170,N_10297,N_9685);
nand U11171 (N_11171,N_10056,N_9316);
xor U11172 (N_11172,N_9886,N_9346);
nand U11173 (N_11173,N_10231,N_9599);
nor U11174 (N_11174,N_10069,N_10357);
or U11175 (N_11175,N_9829,N_9343);
and U11176 (N_11176,N_10060,N_9310);
nor U11177 (N_11177,N_9059,N_9932);
xor U11178 (N_11178,N_9657,N_9941);
nor U11179 (N_11179,N_9061,N_9537);
and U11180 (N_11180,N_10216,N_10303);
or U11181 (N_11181,N_9291,N_9171);
and U11182 (N_11182,N_9230,N_9721);
xor U11183 (N_11183,N_9017,N_10059);
xor U11184 (N_11184,N_9351,N_10305);
nor U11185 (N_11185,N_10260,N_9698);
and U11186 (N_11186,N_9087,N_10349);
and U11187 (N_11187,N_9612,N_9564);
and U11188 (N_11188,N_9690,N_10451);
and U11189 (N_11189,N_9480,N_9851);
or U11190 (N_11190,N_9810,N_10320);
nand U11191 (N_11191,N_9421,N_9753);
or U11192 (N_11192,N_10353,N_9862);
xnor U11193 (N_11193,N_9358,N_9162);
nand U11194 (N_11194,N_9583,N_10040);
xnor U11195 (N_11195,N_10193,N_9193);
nand U11196 (N_11196,N_10195,N_10315);
or U11197 (N_11197,N_9214,N_10144);
and U11198 (N_11198,N_9248,N_10384);
nor U11199 (N_11199,N_9779,N_9359);
nand U11200 (N_11200,N_10301,N_9068);
xor U11201 (N_11201,N_10495,N_10106);
xnor U11202 (N_11202,N_9206,N_9576);
nor U11203 (N_11203,N_9223,N_9085);
xor U11204 (N_11204,N_10041,N_9477);
nand U11205 (N_11205,N_10369,N_9285);
or U11206 (N_11206,N_9640,N_9569);
nand U11207 (N_11207,N_10088,N_9782);
xnor U11208 (N_11208,N_9202,N_10138);
and U11209 (N_11209,N_10332,N_9664);
nor U11210 (N_11210,N_9207,N_9831);
or U11211 (N_11211,N_10381,N_10111);
or U11212 (N_11212,N_9683,N_9155);
xor U11213 (N_11213,N_9126,N_9588);
nand U11214 (N_11214,N_10199,N_9173);
nand U11215 (N_11215,N_10075,N_9323);
nor U11216 (N_11216,N_9826,N_10299);
and U11217 (N_11217,N_10217,N_10247);
nor U11218 (N_11218,N_10307,N_10472);
nand U11219 (N_11219,N_9750,N_9630);
nor U11220 (N_11220,N_9103,N_9983);
nor U11221 (N_11221,N_10209,N_9893);
nand U11222 (N_11222,N_10154,N_9695);
or U11223 (N_11223,N_9914,N_9869);
nor U11224 (N_11224,N_9256,N_10026);
nor U11225 (N_11225,N_9409,N_9506);
nor U11226 (N_11226,N_10206,N_9425);
and U11227 (N_11227,N_10149,N_9546);
nand U11228 (N_11228,N_9628,N_9019);
nor U11229 (N_11229,N_9705,N_9073);
and U11230 (N_11230,N_9280,N_9989);
and U11231 (N_11231,N_9440,N_9492);
nor U11232 (N_11232,N_9188,N_9449);
and U11233 (N_11233,N_10406,N_9121);
and U11234 (N_11234,N_9923,N_9592);
and U11235 (N_11235,N_9798,N_9654);
xnor U11236 (N_11236,N_10415,N_9393);
nand U11237 (N_11237,N_9525,N_9052);
nor U11238 (N_11238,N_9796,N_9613);
nor U11239 (N_11239,N_9702,N_9935);
xor U11240 (N_11240,N_10296,N_9928);
or U11241 (N_11241,N_9740,N_9429);
or U11242 (N_11242,N_9833,N_9441);
nor U11243 (N_11243,N_9991,N_10456);
or U11244 (N_11244,N_9485,N_9083);
and U11245 (N_11245,N_9489,N_10165);
or U11246 (N_11246,N_10007,N_10005);
xor U11247 (N_11247,N_9501,N_9461);
or U11248 (N_11248,N_9144,N_9718);
and U11249 (N_11249,N_9250,N_9710);
nor U11250 (N_11250,N_9834,N_9817);
or U11251 (N_11251,N_10255,N_9903);
or U11252 (N_11252,N_9135,N_10479);
nor U11253 (N_11253,N_9155,N_10372);
xor U11254 (N_11254,N_10477,N_9400);
and U11255 (N_11255,N_9946,N_10316);
or U11256 (N_11256,N_9957,N_9528);
nor U11257 (N_11257,N_10230,N_10465);
or U11258 (N_11258,N_9613,N_9428);
and U11259 (N_11259,N_9984,N_9459);
or U11260 (N_11260,N_9587,N_9084);
nor U11261 (N_11261,N_9661,N_9537);
xnor U11262 (N_11262,N_10142,N_9589);
xor U11263 (N_11263,N_9824,N_9631);
nand U11264 (N_11264,N_9721,N_9669);
nor U11265 (N_11265,N_9308,N_10000);
xnor U11266 (N_11266,N_10023,N_9013);
nand U11267 (N_11267,N_9967,N_9430);
or U11268 (N_11268,N_10187,N_9414);
nor U11269 (N_11269,N_9457,N_9151);
nor U11270 (N_11270,N_10011,N_10376);
and U11271 (N_11271,N_10432,N_10086);
xnor U11272 (N_11272,N_9026,N_9856);
and U11273 (N_11273,N_10164,N_9612);
nor U11274 (N_11274,N_9099,N_9175);
or U11275 (N_11275,N_9085,N_9350);
nor U11276 (N_11276,N_10454,N_9249);
or U11277 (N_11277,N_9068,N_9063);
and U11278 (N_11278,N_9745,N_9217);
xnor U11279 (N_11279,N_9044,N_9126);
and U11280 (N_11280,N_10446,N_9407);
xnor U11281 (N_11281,N_10063,N_9774);
and U11282 (N_11282,N_10483,N_10057);
nor U11283 (N_11283,N_10306,N_10449);
and U11284 (N_11284,N_10465,N_9014);
nand U11285 (N_11285,N_9845,N_9488);
and U11286 (N_11286,N_9332,N_9980);
nand U11287 (N_11287,N_9632,N_9025);
and U11288 (N_11288,N_9122,N_10388);
or U11289 (N_11289,N_10439,N_10075);
and U11290 (N_11290,N_9121,N_9028);
nand U11291 (N_11291,N_10467,N_10484);
and U11292 (N_11292,N_9512,N_10303);
nor U11293 (N_11293,N_9124,N_10082);
nor U11294 (N_11294,N_10206,N_10475);
and U11295 (N_11295,N_9397,N_9579);
nor U11296 (N_11296,N_9912,N_10492);
nor U11297 (N_11297,N_10091,N_10499);
nor U11298 (N_11298,N_9794,N_9013);
xnor U11299 (N_11299,N_9739,N_9069);
nand U11300 (N_11300,N_9992,N_10294);
nor U11301 (N_11301,N_10050,N_10208);
xnor U11302 (N_11302,N_10099,N_9942);
and U11303 (N_11303,N_9045,N_9607);
nor U11304 (N_11304,N_10033,N_9726);
xnor U11305 (N_11305,N_10253,N_9451);
xor U11306 (N_11306,N_10479,N_10105);
nand U11307 (N_11307,N_9340,N_10372);
and U11308 (N_11308,N_9290,N_9916);
nor U11309 (N_11309,N_10275,N_9709);
and U11310 (N_11310,N_9048,N_9991);
nor U11311 (N_11311,N_9185,N_10270);
nor U11312 (N_11312,N_9481,N_9529);
nor U11313 (N_11313,N_10288,N_10160);
and U11314 (N_11314,N_9516,N_10139);
nand U11315 (N_11315,N_10118,N_10044);
nor U11316 (N_11316,N_9007,N_9844);
nor U11317 (N_11317,N_9725,N_9022);
xor U11318 (N_11318,N_9190,N_10262);
or U11319 (N_11319,N_10103,N_9657);
nor U11320 (N_11320,N_9255,N_10465);
or U11321 (N_11321,N_9624,N_9971);
nand U11322 (N_11322,N_9002,N_9617);
xnor U11323 (N_11323,N_9694,N_9050);
or U11324 (N_11324,N_10406,N_9159);
nor U11325 (N_11325,N_10079,N_9286);
nor U11326 (N_11326,N_9435,N_10281);
and U11327 (N_11327,N_9083,N_9013);
and U11328 (N_11328,N_9607,N_10467);
or U11329 (N_11329,N_9471,N_10081);
nand U11330 (N_11330,N_9656,N_9331);
or U11331 (N_11331,N_9540,N_9966);
nor U11332 (N_11332,N_10199,N_10187);
nand U11333 (N_11333,N_9130,N_10452);
and U11334 (N_11334,N_9475,N_9502);
nor U11335 (N_11335,N_9245,N_10486);
nor U11336 (N_11336,N_10420,N_10203);
xor U11337 (N_11337,N_9399,N_9330);
xnor U11338 (N_11338,N_9211,N_10081);
and U11339 (N_11339,N_9831,N_9169);
nor U11340 (N_11340,N_9723,N_10135);
nor U11341 (N_11341,N_10479,N_9140);
nor U11342 (N_11342,N_9605,N_9423);
or U11343 (N_11343,N_9583,N_10093);
or U11344 (N_11344,N_9754,N_9532);
nor U11345 (N_11345,N_9072,N_10046);
nand U11346 (N_11346,N_10034,N_9387);
and U11347 (N_11347,N_10250,N_9889);
xnor U11348 (N_11348,N_10367,N_9219);
nand U11349 (N_11349,N_9758,N_9941);
nor U11350 (N_11350,N_10449,N_10007);
nand U11351 (N_11351,N_10093,N_9992);
nor U11352 (N_11352,N_9029,N_10339);
or U11353 (N_11353,N_9028,N_10365);
nor U11354 (N_11354,N_9825,N_9268);
nand U11355 (N_11355,N_9794,N_10266);
nor U11356 (N_11356,N_9160,N_9318);
nand U11357 (N_11357,N_9746,N_9994);
or U11358 (N_11358,N_9381,N_10217);
nand U11359 (N_11359,N_9114,N_10097);
nor U11360 (N_11360,N_10033,N_10268);
nand U11361 (N_11361,N_9895,N_9726);
nor U11362 (N_11362,N_9356,N_9529);
or U11363 (N_11363,N_9098,N_9832);
or U11364 (N_11364,N_9094,N_9958);
nand U11365 (N_11365,N_9121,N_9570);
nand U11366 (N_11366,N_10456,N_9027);
nand U11367 (N_11367,N_9516,N_9214);
nand U11368 (N_11368,N_9649,N_9364);
nor U11369 (N_11369,N_9055,N_9879);
nor U11370 (N_11370,N_9872,N_9061);
nand U11371 (N_11371,N_9128,N_10498);
nor U11372 (N_11372,N_9253,N_10007);
or U11373 (N_11373,N_10459,N_9484);
or U11374 (N_11374,N_10158,N_9495);
and U11375 (N_11375,N_9074,N_10309);
and U11376 (N_11376,N_10104,N_9767);
nor U11377 (N_11377,N_10222,N_9550);
nor U11378 (N_11378,N_10108,N_9121);
nor U11379 (N_11379,N_9153,N_9932);
nor U11380 (N_11380,N_10067,N_9744);
nand U11381 (N_11381,N_9101,N_9726);
nand U11382 (N_11382,N_9027,N_10151);
and U11383 (N_11383,N_10063,N_9678);
or U11384 (N_11384,N_9707,N_9576);
nand U11385 (N_11385,N_9372,N_9795);
nand U11386 (N_11386,N_10436,N_9792);
or U11387 (N_11387,N_9945,N_10006);
and U11388 (N_11388,N_10441,N_10353);
and U11389 (N_11389,N_10073,N_10094);
nand U11390 (N_11390,N_10038,N_9097);
and U11391 (N_11391,N_9604,N_9941);
or U11392 (N_11392,N_10386,N_9205);
or U11393 (N_11393,N_9387,N_9992);
xnor U11394 (N_11394,N_9567,N_9089);
and U11395 (N_11395,N_9508,N_9260);
or U11396 (N_11396,N_9670,N_9673);
nor U11397 (N_11397,N_10403,N_9571);
and U11398 (N_11398,N_9884,N_9318);
and U11399 (N_11399,N_9984,N_9701);
nand U11400 (N_11400,N_10447,N_9950);
nor U11401 (N_11401,N_10027,N_9346);
nor U11402 (N_11402,N_9758,N_9011);
nand U11403 (N_11403,N_9737,N_10051);
nor U11404 (N_11404,N_9723,N_9185);
nor U11405 (N_11405,N_9868,N_10199);
and U11406 (N_11406,N_9679,N_9298);
nand U11407 (N_11407,N_10032,N_10191);
nand U11408 (N_11408,N_9345,N_9019);
or U11409 (N_11409,N_9935,N_9746);
nand U11410 (N_11410,N_10190,N_9234);
and U11411 (N_11411,N_10175,N_10127);
nor U11412 (N_11412,N_9881,N_10051);
and U11413 (N_11413,N_9965,N_9137);
xnor U11414 (N_11414,N_9987,N_10034);
nor U11415 (N_11415,N_10467,N_10174);
and U11416 (N_11416,N_10436,N_9534);
nand U11417 (N_11417,N_10325,N_9122);
xnor U11418 (N_11418,N_9492,N_10170);
or U11419 (N_11419,N_9156,N_9647);
and U11420 (N_11420,N_9688,N_9624);
nand U11421 (N_11421,N_9276,N_9288);
or U11422 (N_11422,N_9699,N_9828);
xnor U11423 (N_11423,N_9917,N_9967);
nor U11424 (N_11424,N_9557,N_9203);
nor U11425 (N_11425,N_9027,N_9062);
or U11426 (N_11426,N_9004,N_10352);
nor U11427 (N_11427,N_9468,N_9666);
nor U11428 (N_11428,N_9710,N_10085);
and U11429 (N_11429,N_10392,N_9564);
and U11430 (N_11430,N_9222,N_10207);
nand U11431 (N_11431,N_9742,N_10279);
nor U11432 (N_11432,N_9936,N_10102);
nand U11433 (N_11433,N_10193,N_9116);
nand U11434 (N_11434,N_10002,N_9713);
or U11435 (N_11435,N_9373,N_9606);
and U11436 (N_11436,N_9890,N_9452);
nand U11437 (N_11437,N_9655,N_9076);
and U11438 (N_11438,N_9643,N_9074);
nand U11439 (N_11439,N_10059,N_10263);
and U11440 (N_11440,N_9204,N_10314);
nand U11441 (N_11441,N_9040,N_10293);
nand U11442 (N_11442,N_9787,N_10006);
nand U11443 (N_11443,N_10075,N_10256);
and U11444 (N_11444,N_9235,N_10155);
or U11445 (N_11445,N_10001,N_9388);
nand U11446 (N_11446,N_10378,N_10005);
nand U11447 (N_11447,N_10340,N_10046);
or U11448 (N_11448,N_9706,N_9243);
nor U11449 (N_11449,N_9239,N_10166);
or U11450 (N_11450,N_10122,N_9013);
or U11451 (N_11451,N_10424,N_9333);
nor U11452 (N_11452,N_10196,N_9585);
and U11453 (N_11453,N_9247,N_9347);
or U11454 (N_11454,N_9585,N_9118);
or U11455 (N_11455,N_10250,N_9928);
nand U11456 (N_11456,N_9600,N_10332);
and U11457 (N_11457,N_10385,N_9372);
xor U11458 (N_11458,N_9519,N_9524);
nand U11459 (N_11459,N_9508,N_9396);
nor U11460 (N_11460,N_9013,N_9493);
nor U11461 (N_11461,N_10348,N_10236);
nor U11462 (N_11462,N_9484,N_9138);
nand U11463 (N_11463,N_10233,N_9509);
nand U11464 (N_11464,N_10068,N_9390);
or U11465 (N_11465,N_9954,N_10304);
xnor U11466 (N_11466,N_10349,N_9104);
and U11467 (N_11467,N_9196,N_10104);
and U11468 (N_11468,N_9026,N_9769);
and U11469 (N_11469,N_10473,N_10267);
nand U11470 (N_11470,N_9306,N_9505);
and U11471 (N_11471,N_9376,N_9065);
nor U11472 (N_11472,N_9806,N_9082);
or U11473 (N_11473,N_9558,N_9432);
and U11474 (N_11474,N_10005,N_9842);
or U11475 (N_11475,N_9959,N_9424);
nand U11476 (N_11476,N_10286,N_9197);
nand U11477 (N_11477,N_9413,N_9978);
nor U11478 (N_11478,N_10258,N_9318);
nand U11479 (N_11479,N_9771,N_9572);
nor U11480 (N_11480,N_9917,N_10246);
or U11481 (N_11481,N_10301,N_10411);
nand U11482 (N_11482,N_9777,N_9397);
or U11483 (N_11483,N_10032,N_10324);
nor U11484 (N_11484,N_9963,N_10249);
and U11485 (N_11485,N_9999,N_9902);
nor U11486 (N_11486,N_10417,N_10218);
and U11487 (N_11487,N_9840,N_10064);
or U11488 (N_11488,N_9585,N_10190);
or U11489 (N_11489,N_9524,N_9807);
nand U11490 (N_11490,N_9959,N_9579);
or U11491 (N_11491,N_9631,N_9872);
or U11492 (N_11492,N_9732,N_9178);
xor U11493 (N_11493,N_9987,N_9130);
nand U11494 (N_11494,N_9366,N_9212);
xnor U11495 (N_11495,N_10000,N_9042);
or U11496 (N_11496,N_9406,N_9023);
or U11497 (N_11497,N_9002,N_9935);
xor U11498 (N_11498,N_9939,N_10368);
nand U11499 (N_11499,N_9712,N_9348);
and U11500 (N_11500,N_10321,N_10402);
or U11501 (N_11501,N_9149,N_9283);
or U11502 (N_11502,N_10088,N_9828);
or U11503 (N_11503,N_10210,N_9789);
nor U11504 (N_11504,N_10348,N_10015);
nor U11505 (N_11505,N_10123,N_9920);
nor U11506 (N_11506,N_9230,N_9284);
xnor U11507 (N_11507,N_9960,N_10100);
or U11508 (N_11508,N_10171,N_9082);
and U11509 (N_11509,N_10377,N_9477);
nor U11510 (N_11510,N_9699,N_10153);
nor U11511 (N_11511,N_10047,N_9286);
nor U11512 (N_11512,N_9608,N_9717);
or U11513 (N_11513,N_9132,N_9945);
nand U11514 (N_11514,N_10480,N_10391);
xnor U11515 (N_11515,N_10124,N_10206);
and U11516 (N_11516,N_10349,N_9026);
nand U11517 (N_11517,N_9392,N_9307);
nand U11518 (N_11518,N_9688,N_10483);
or U11519 (N_11519,N_9522,N_9931);
or U11520 (N_11520,N_9993,N_10485);
or U11521 (N_11521,N_10427,N_9883);
and U11522 (N_11522,N_9515,N_9011);
nand U11523 (N_11523,N_10033,N_10324);
nor U11524 (N_11524,N_9593,N_9995);
and U11525 (N_11525,N_9321,N_9276);
nor U11526 (N_11526,N_10292,N_9430);
and U11527 (N_11527,N_10292,N_10271);
nand U11528 (N_11528,N_9885,N_10477);
or U11529 (N_11529,N_10356,N_10495);
or U11530 (N_11530,N_9846,N_9323);
and U11531 (N_11531,N_9453,N_10220);
or U11532 (N_11532,N_9068,N_9227);
and U11533 (N_11533,N_10224,N_10468);
and U11534 (N_11534,N_9312,N_10275);
nor U11535 (N_11535,N_9557,N_9167);
or U11536 (N_11536,N_9372,N_9706);
xnor U11537 (N_11537,N_9645,N_9613);
nand U11538 (N_11538,N_9723,N_9091);
or U11539 (N_11539,N_9503,N_9476);
or U11540 (N_11540,N_9684,N_10388);
nand U11541 (N_11541,N_10294,N_10382);
nor U11542 (N_11542,N_9434,N_9477);
nand U11543 (N_11543,N_10354,N_9306);
nor U11544 (N_11544,N_10479,N_9044);
or U11545 (N_11545,N_9381,N_9869);
or U11546 (N_11546,N_10449,N_9128);
and U11547 (N_11547,N_9759,N_10078);
nor U11548 (N_11548,N_9500,N_9212);
nand U11549 (N_11549,N_10188,N_9531);
and U11550 (N_11550,N_10389,N_9970);
nor U11551 (N_11551,N_10322,N_10218);
and U11552 (N_11552,N_9856,N_9067);
and U11553 (N_11553,N_10023,N_10213);
and U11554 (N_11554,N_9078,N_9397);
nand U11555 (N_11555,N_9849,N_9634);
xnor U11556 (N_11556,N_9477,N_9514);
and U11557 (N_11557,N_10264,N_10051);
or U11558 (N_11558,N_9620,N_10084);
xnor U11559 (N_11559,N_10341,N_9742);
nand U11560 (N_11560,N_10029,N_9756);
or U11561 (N_11561,N_9755,N_9671);
nor U11562 (N_11562,N_9692,N_9010);
or U11563 (N_11563,N_9787,N_10228);
or U11564 (N_11564,N_9606,N_9881);
nor U11565 (N_11565,N_9888,N_9328);
nor U11566 (N_11566,N_9484,N_9093);
xor U11567 (N_11567,N_9707,N_10282);
and U11568 (N_11568,N_10184,N_10026);
or U11569 (N_11569,N_9548,N_9550);
nand U11570 (N_11570,N_9922,N_9311);
nand U11571 (N_11571,N_10196,N_9760);
or U11572 (N_11572,N_10038,N_9974);
or U11573 (N_11573,N_9361,N_9517);
nand U11574 (N_11574,N_9117,N_10271);
and U11575 (N_11575,N_10410,N_9497);
or U11576 (N_11576,N_9966,N_9126);
or U11577 (N_11577,N_9069,N_10234);
nor U11578 (N_11578,N_10472,N_9829);
and U11579 (N_11579,N_9079,N_9380);
or U11580 (N_11580,N_10451,N_9829);
nor U11581 (N_11581,N_10350,N_9050);
and U11582 (N_11582,N_9928,N_10225);
nor U11583 (N_11583,N_10248,N_10439);
nor U11584 (N_11584,N_9978,N_10103);
nor U11585 (N_11585,N_9849,N_10030);
nand U11586 (N_11586,N_10191,N_9178);
xor U11587 (N_11587,N_9434,N_9946);
nand U11588 (N_11588,N_9499,N_9771);
or U11589 (N_11589,N_10053,N_10497);
nand U11590 (N_11590,N_9681,N_9853);
or U11591 (N_11591,N_9695,N_9096);
nand U11592 (N_11592,N_10217,N_10409);
nand U11593 (N_11593,N_9488,N_10255);
nor U11594 (N_11594,N_9534,N_9032);
or U11595 (N_11595,N_9522,N_9853);
and U11596 (N_11596,N_9229,N_10251);
nand U11597 (N_11597,N_9776,N_9546);
or U11598 (N_11598,N_9509,N_9730);
nand U11599 (N_11599,N_9103,N_10373);
nand U11600 (N_11600,N_10056,N_9151);
and U11601 (N_11601,N_9023,N_9976);
or U11602 (N_11602,N_9500,N_10220);
xnor U11603 (N_11603,N_9997,N_9887);
or U11604 (N_11604,N_9282,N_10387);
nor U11605 (N_11605,N_9103,N_10112);
or U11606 (N_11606,N_9186,N_9077);
xnor U11607 (N_11607,N_9635,N_10226);
nor U11608 (N_11608,N_9351,N_9774);
nor U11609 (N_11609,N_9774,N_9786);
and U11610 (N_11610,N_9702,N_9666);
nand U11611 (N_11611,N_9233,N_10233);
or U11612 (N_11612,N_9413,N_10194);
nand U11613 (N_11613,N_9240,N_9801);
nor U11614 (N_11614,N_9527,N_9878);
and U11615 (N_11615,N_9912,N_9369);
nand U11616 (N_11616,N_9270,N_9356);
nand U11617 (N_11617,N_9722,N_9151);
nand U11618 (N_11618,N_9784,N_9230);
nor U11619 (N_11619,N_9387,N_9870);
and U11620 (N_11620,N_9666,N_10411);
nand U11621 (N_11621,N_9484,N_10224);
nand U11622 (N_11622,N_9373,N_10349);
and U11623 (N_11623,N_9141,N_10012);
and U11624 (N_11624,N_9595,N_9459);
or U11625 (N_11625,N_9238,N_9421);
or U11626 (N_11626,N_9588,N_9914);
nor U11627 (N_11627,N_9756,N_10383);
or U11628 (N_11628,N_9736,N_9225);
nor U11629 (N_11629,N_9912,N_9432);
or U11630 (N_11630,N_9885,N_9680);
nor U11631 (N_11631,N_9339,N_10196);
or U11632 (N_11632,N_9074,N_9335);
xnor U11633 (N_11633,N_9204,N_10358);
and U11634 (N_11634,N_9665,N_9559);
or U11635 (N_11635,N_10166,N_10224);
or U11636 (N_11636,N_10248,N_9482);
or U11637 (N_11637,N_10464,N_10357);
or U11638 (N_11638,N_9125,N_10288);
and U11639 (N_11639,N_10120,N_9458);
or U11640 (N_11640,N_10112,N_9858);
or U11641 (N_11641,N_9445,N_9204);
nand U11642 (N_11642,N_9755,N_9698);
nor U11643 (N_11643,N_10204,N_9742);
nor U11644 (N_11644,N_9265,N_9241);
and U11645 (N_11645,N_10369,N_9823);
nand U11646 (N_11646,N_10489,N_9064);
nor U11647 (N_11647,N_10359,N_9173);
nor U11648 (N_11648,N_10387,N_9497);
nand U11649 (N_11649,N_9138,N_9415);
and U11650 (N_11650,N_9054,N_9083);
nand U11651 (N_11651,N_9922,N_10214);
nor U11652 (N_11652,N_10193,N_9533);
nor U11653 (N_11653,N_10013,N_9501);
and U11654 (N_11654,N_9938,N_9399);
nand U11655 (N_11655,N_10479,N_9424);
or U11656 (N_11656,N_9360,N_9611);
nand U11657 (N_11657,N_10014,N_10027);
or U11658 (N_11658,N_10247,N_9887);
or U11659 (N_11659,N_9780,N_9909);
nor U11660 (N_11660,N_10375,N_9803);
nand U11661 (N_11661,N_9741,N_9436);
and U11662 (N_11662,N_9536,N_9071);
nor U11663 (N_11663,N_10306,N_9471);
and U11664 (N_11664,N_9999,N_9053);
and U11665 (N_11665,N_9044,N_10007);
nor U11666 (N_11666,N_10250,N_10389);
nor U11667 (N_11667,N_10341,N_9191);
nor U11668 (N_11668,N_10480,N_10024);
nor U11669 (N_11669,N_9437,N_10221);
and U11670 (N_11670,N_9534,N_9505);
nor U11671 (N_11671,N_9874,N_9000);
and U11672 (N_11672,N_10059,N_9147);
nand U11673 (N_11673,N_9292,N_9169);
nor U11674 (N_11674,N_9797,N_9555);
and U11675 (N_11675,N_9190,N_10135);
or U11676 (N_11676,N_9332,N_9258);
xnor U11677 (N_11677,N_9713,N_9015);
nor U11678 (N_11678,N_10102,N_9244);
nand U11679 (N_11679,N_9305,N_9797);
or U11680 (N_11680,N_9394,N_10421);
or U11681 (N_11681,N_10449,N_10056);
or U11682 (N_11682,N_10441,N_9777);
nand U11683 (N_11683,N_9808,N_9120);
and U11684 (N_11684,N_9035,N_9712);
nor U11685 (N_11685,N_9360,N_9496);
or U11686 (N_11686,N_10203,N_9829);
nor U11687 (N_11687,N_9705,N_9958);
or U11688 (N_11688,N_10318,N_10223);
xnor U11689 (N_11689,N_9397,N_10452);
nand U11690 (N_11690,N_9602,N_9899);
nand U11691 (N_11691,N_9261,N_9031);
or U11692 (N_11692,N_9054,N_9490);
and U11693 (N_11693,N_9474,N_9391);
and U11694 (N_11694,N_10223,N_10110);
or U11695 (N_11695,N_9188,N_9714);
and U11696 (N_11696,N_9109,N_10262);
nand U11697 (N_11697,N_9506,N_10164);
and U11698 (N_11698,N_10294,N_9192);
and U11699 (N_11699,N_9832,N_10264);
or U11700 (N_11700,N_9192,N_10209);
nor U11701 (N_11701,N_9191,N_9826);
and U11702 (N_11702,N_10256,N_9514);
nand U11703 (N_11703,N_10465,N_9541);
nor U11704 (N_11704,N_10214,N_9586);
and U11705 (N_11705,N_10208,N_10464);
nand U11706 (N_11706,N_9210,N_9383);
or U11707 (N_11707,N_10348,N_10460);
and U11708 (N_11708,N_10285,N_10129);
nor U11709 (N_11709,N_9534,N_10066);
nand U11710 (N_11710,N_9484,N_9136);
nand U11711 (N_11711,N_9372,N_9407);
or U11712 (N_11712,N_9011,N_9333);
or U11713 (N_11713,N_10294,N_9809);
and U11714 (N_11714,N_9676,N_9469);
nor U11715 (N_11715,N_9909,N_10302);
nand U11716 (N_11716,N_10056,N_9093);
and U11717 (N_11717,N_10243,N_9575);
xor U11718 (N_11718,N_9997,N_10235);
or U11719 (N_11719,N_10394,N_9931);
xor U11720 (N_11720,N_9278,N_9719);
xnor U11721 (N_11721,N_9951,N_9011);
nand U11722 (N_11722,N_10034,N_10291);
nor U11723 (N_11723,N_9512,N_9741);
or U11724 (N_11724,N_10345,N_9294);
nand U11725 (N_11725,N_9142,N_9872);
nand U11726 (N_11726,N_9897,N_9826);
or U11727 (N_11727,N_10486,N_9606);
xnor U11728 (N_11728,N_9522,N_9775);
or U11729 (N_11729,N_9475,N_9733);
or U11730 (N_11730,N_10492,N_10151);
or U11731 (N_11731,N_9595,N_9126);
nor U11732 (N_11732,N_10186,N_10029);
or U11733 (N_11733,N_10207,N_9454);
or U11734 (N_11734,N_9909,N_10050);
nor U11735 (N_11735,N_9274,N_9581);
and U11736 (N_11736,N_9637,N_9971);
nor U11737 (N_11737,N_9648,N_9187);
xor U11738 (N_11738,N_9344,N_10343);
nand U11739 (N_11739,N_10059,N_9835);
and U11740 (N_11740,N_9745,N_9537);
nor U11741 (N_11741,N_10375,N_10077);
xor U11742 (N_11742,N_9227,N_9130);
nand U11743 (N_11743,N_9359,N_10005);
xor U11744 (N_11744,N_9280,N_9233);
and U11745 (N_11745,N_9063,N_10332);
nor U11746 (N_11746,N_10369,N_10207);
and U11747 (N_11747,N_9665,N_9715);
and U11748 (N_11748,N_10018,N_9298);
or U11749 (N_11749,N_9011,N_9134);
and U11750 (N_11750,N_10119,N_9471);
and U11751 (N_11751,N_10237,N_9924);
nor U11752 (N_11752,N_9055,N_9587);
and U11753 (N_11753,N_9405,N_9233);
nor U11754 (N_11754,N_9054,N_9909);
and U11755 (N_11755,N_10499,N_9312);
or U11756 (N_11756,N_9555,N_10326);
nand U11757 (N_11757,N_9225,N_10312);
nand U11758 (N_11758,N_10277,N_10027);
and U11759 (N_11759,N_9279,N_10128);
nor U11760 (N_11760,N_10235,N_9566);
or U11761 (N_11761,N_9854,N_10355);
nor U11762 (N_11762,N_10128,N_10134);
nor U11763 (N_11763,N_10340,N_9252);
and U11764 (N_11764,N_9891,N_9794);
or U11765 (N_11765,N_10176,N_10347);
or U11766 (N_11766,N_9715,N_10159);
and U11767 (N_11767,N_10198,N_9797);
nor U11768 (N_11768,N_10385,N_9754);
nand U11769 (N_11769,N_9803,N_9937);
and U11770 (N_11770,N_10442,N_9364);
nor U11771 (N_11771,N_10182,N_10362);
nor U11772 (N_11772,N_10255,N_9848);
and U11773 (N_11773,N_10412,N_9016);
nand U11774 (N_11774,N_9334,N_10152);
or U11775 (N_11775,N_10442,N_9504);
or U11776 (N_11776,N_10359,N_9950);
and U11777 (N_11777,N_9694,N_10325);
and U11778 (N_11778,N_9404,N_10192);
nor U11779 (N_11779,N_9541,N_10438);
nor U11780 (N_11780,N_10217,N_9003);
nand U11781 (N_11781,N_10055,N_9767);
nand U11782 (N_11782,N_10293,N_10416);
nand U11783 (N_11783,N_9799,N_10422);
and U11784 (N_11784,N_9688,N_9283);
nor U11785 (N_11785,N_9064,N_9817);
and U11786 (N_11786,N_9820,N_9531);
nand U11787 (N_11787,N_10127,N_9526);
and U11788 (N_11788,N_9422,N_9015);
or U11789 (N_11789,N_9182,N_10347);
nor U11790 (N_11790,N_10223,N_9952);
and U11791 (N_11791,N_10483,N_10407);
and U11792 (N_11792,N_9708,N_9516);
nor U11793 (N_11793,N_9146,N_10428);
nand U11794 (N_11794,N_9723,N_9991);
or U11795 (N_11795,N_10391,N_10074);
or U11796 (N_11796,N_9341,N_9522);
nand U11797 (N_11797,N_10214,N_9066);
and U11798 (N_11798,N_9077,N_10266);
or U11799 (N_11799,N_9677,N_9621);
nand U11800 (N_11800,N_10291,N_10205);
xor U11801 (N_11801,N_9212,N_10111);
or U11802 (N_11802,N_9877,N_9915);
nand U11803 (N_11803,N_9005,N_10269);
nand U11804 (N_11804,N_10453,N_9678);
nand U11805 (N_11805,N_10178,N_10072);
nand U11806 (N_11806,N_9186,N_9897);
and U11807 (N_11807,N_10465,N_10467);
and U11808 (N_11808,N_9563,N_9762);
and U11809 (N_11809,N_10384,N_10294);
or U11810 (N_11810,N_9011,N_10417);
and U11811 (N_11811,N_9330,N_9133);
or U11812 (N_11812,N_10262,N_9721);
nand U11813 (N_11813,N_10043,N_9564);
nor U11814 (N_11814,N_9633,N_9664);
and U11815 (N_11815,N_9129,N_10170);
nand U11816 (N_11816,N_9017,N_9285);
and U11817 (N_11817,N_9076,N_9639);
or U11818 (N_11818,N_9627,N_9518);
nand U11819 (N_11819,N_9441,N_9890);
nor U11820 (N_11820,N_9592,N_9849);
or U11821 (N_11821,N_9333,N_9508);
nand U11822 (N_11822,N_9589,N_10165);
nor U11823 (N_11823,N_9210,N_9511);
nor U11824 (N_11824,N_9040,N_9295);
or U11825 (N_11825,N_9949,N_10134);
or U11826 (N_11826,N_9044,N_9611);
or U11827 (N_11827,N_9666,N_10455);
or U11828 (N_11828,N_9299,N_9758);
nand U11829 (N_11829,N_9405,N_9687);
nand U11830 (N_11830,N_10250,N_9969);
or U11831 (N_11831,N_9064,N_9380);
nand U11832 (N_11832,N_9407,N_10452);
and U11833 (N_11833,N_9595,N_9777);
and U11834 (N_11834,N_9025,N_9396);
nor U11835 (N_11835,N_9178,N_9021);
xnor U11836 (N_11836,N_9229,N_10317);
or U11837 (N_11837,N_9590,N_9016);
or U11838 (N_11838,N_9676,N_9208);
and U11839 (N_11839,N_9745,N_10431);
xor U11840 (N_11840,N_9925,N_9256);
and U11841 (N_11841,N_9158,N_9046);
nor U11842 (N_11842,N_9240,N_10389);
nand U11843 (N_11843,N_9185,N_9903);
nand U11844 (N_11844,N_10304,N_9753);
nor U11845 (N_11845,N_9834,N_9066);
and U11846 (N_11846,N_9454,N_9171);
xor U11847 (N_11847,N_9352,N_9518);
nand U11848 (N_11848,N_9979,N_9161);
nor U11849 (N_11849,N_9293,N_9274);
nor U11850 (N_11850,N_9265,N_9892);
and U11851 (N_11851,N_10341,N_10155);
and U11852 (N_11852,N_9469,N_9962);
or U11853 (N_11853,N_9660,N_9176);
and U11854 (N_11854,N_9884,N_10364);
nor U11855 (N_11855,N_9925,N_9792);
nor U11856 (N_11856,N_9642,N_9442);
xnor U11857 (N_11857,N_9445,N_10138);
and U11858 (N_11858,N_10068,N_10107);
nor U11859 (N_11859,N_10046,N_9868);
and U11860 (N_11860,N_9396,N_10226);
nand U11861 (N_11861,N_9017,N_10043);
xnor U11862 (N_11862,N_9669,N_10416);
nand U11863 (N_11863,N_9827,N_9535);
nor U11864 (N_11864,N_9400,N_10216);
and U11865 (N_11865,N_10031,N_9802);
and U11866 (N_11866,N_9956,N_9769);
and U11867 (N_11867,N_10158,N_9460);
and U11868 (N_11868,N_9721,N_10282);
nand U11869 (N_11869,N_9126,N_9497);
or U11870 (N_11870,N_9124,N_10473);
and U11871 (N_11871,N_9869,N_9147);
and U11872 (N_11872,N_9578,N_9626);
nor U11873 (N_11873,N_9694,N_10330);
nor U11874 (N_11874,N_9837,N_9092);
and U11875 (N_11875,N_10057,N_9795);
nor U11876 (N_11876,N_9449,N_9460);
nor U11877 (N_11877,N_9321,N_9936);
and U11878 (N_11878,N_10434,N_9555);
nor U11879 (N_11879,N_9233,N_10473);
xnor U11880 (N_11880,N_9108,N_10160);
or U11881 (N_11881,N_10479,N_9882);
and U11882 (N_11882,N_9294,N_9398);
and U11883 (N_11883,N_10276,N_9230);
nor U11884 (N_11884,N_9505,N_9602);
and U11885 (N_11885,N_9453,N_9032);
and U11886 (N_11886,N_10081,N_10381);
nor U11887 (N_11887,N_9663,N_9111);
or U11888 (N_11888,N_10404,N_9942);
or U11889 (N_11889,N_10382,N_9817);
and U11890 (N_11890,N_9831,N_10027);
or U11891 (N_11891,N_9715,N_9078);
or U11892 (N_11892,N_9552,N_10388);
and U11893 (N_11893,N_10416,N_9518);
xnor U11894 (N_11894,N_9331,N_10354);
or U11895 (N_11895,N_9350,N_10275);
or U11896 (N_11896,N_10187,N_9063);
nor U11897 (N_11897,N_9944,N_9900);
and U11898 (N_11898,N_9123,N_10496);
or U11899 (N_11899,N_9146,N_10311);
nor U11900 (N_11900,N_9325,N_9173);
nor U11901 (N_11901,N_9096,N_10189);
nand U11902 (N_11902,N_9475,N_9936);
and U11903 (N_11903,N_9666,N_9396);
nor U11904 (N_11904,N_10175,N_9837);
and U11905 (N_11905,N_9082,N_10292);
nand U11906 (N_11906,N_10402,N_10080);
and U11907 (N_11907,N_9944,N_9200);
or U11908 (N_11908,N_9406,N_9272);
nor U11909 (N_11909,N_9454,N_10256);
nor U11910 (N_11910,N_9447,N_9556);
and U11911 (N_11911,N_9749,N_9796);
nor U11912 (N_11912,N_9426,N_10161);
and U11913 (N_11913,N_9335,N_9211);
and U11914 (N_11914,N_9729,N_9831);
and U11915 (N_11915,N_9605,N_10263);
xnor U11916 (N_11916,N_10256,N_9892);
xor U11917 (N_11917,N_9926,N_9481);
and U11918 (N_11918,N_9203,N_10495);
nor U11919 (N_11919,N_9053,N_9460);
nor U11920 (N_11920,N_10465,N_9011);
or U11921 (N_11921,N_9007,N_10138);
nor U11922 (N_11922,N_9788,N_9389);
nand U11923 (N_11923,N_9230,N_10189);
nor U11924 (N_11924,N_9458,N_10312);
nor U11925 (N_11925,N_9565,N_9630);
or U11926 (N_11926,N_9829,N_10167);
nand U11927 (N_11927,N_9609,N_9597);
nor U11928 (N_11928,N_9006,N_9594);
nor U11929 (N_11929,N_9377,N_10361);
and U11930 (N_11930,N_9845,N_9964);
and U11931 (N_11931,N_9193,N_9599);
nor U11932 (N_11932,N_9611,N_9413);
and U11933 (N_11933,N_10273,N_10288);
nor U11934 (N_11934,N_9649,N_9415);
nand U11935 (N_11935,N_10489,N_10414);
or U11936 (N_11936,N_10099,N_10018);
nand U11937 (N_11937,N_10355,N_9313);
nand U11938 (N_11938,N_10421,N_9127);
and U11939 (N_11939,N_9649,N_9287);
and U11940 (N_11940,N_9143,N_9823);
or U11941 (N_11941,N_9056,N_9158);
and U11942 (N_11942,N_10017,N_10104);
or U11943 (N_11943,N_9081,N_9594);
or U11944 (N_11944,N_9302,N_10244);
or U11945 (N_11945,N_9464,N_9684);
nor U11946 (N_11946,N_10215,N_9289);
or U11947 (N_11947,N_10266,N_9201);
and U11948 (N_11948,N_9471,N_10108);
nor U11949 (N_11949,N_9862,N_10272);
and U11950 (N_11950,N_10040,N_9429);
or U11951 (N_11951,N_9221,N_10213);
nor U11952 (N_11952,N_9747,N_10018);
nand U11953 (N_11953,N_9846,N_10263);
xor U11954 (N_11954,N_9568,N_9936);
nor U11955 (N_11955,N_9773,N_10497);
nor U11956 (N_11956,N_9135,N_10488);
nand U11957 (N_11957,N_9063,N_9153);
xnor U11958 (N_11958,N_9947,N_9416);
or U11959 (N_11959,N_10049,N_9019);
and U11960 (N_11960,N_10317,N_9967);
and U11961 (N_11961,N_10004,N_9483);
or U11962 (N_11962,N_9086,N_10192);
or U11963 (N_11963,N_10344,N_10034);
nand U11964 (N_11964,N_9583,N_10218);
xnor U11965 (N_11965,N_9470,N_9703);
and U11966 (N_11966,N_10120,N_10205);
or U11967 (N_11967,N_9855,N_10004);
nand U11968 (N_11968,N_9686,N_9996);
nand U11969 (N_11969,N_9542,N_9456);
and U11970 (N_11970,N_9967,N_9918);
or U11971 (N_11971,N_9168,N_10052);
nand U11972 (N_11972,N_9941,N_9000);
nor U11973 (N_11973,N_9440,N_9740);
or U11974 (N_11974,N_9079,N_9823);
nor U11975 (N_11975,N_9119,N_10267);
and U11976 (N_11976,N_10120,N_9297);
and U11977 (N_11977,N_9874,N_9973);
nor U11978 (N_11978,N_9418,N_10221);
nor U11979 (N_11979,N_9263,N_10005);
and U11980 (N_11980,N_9838,N_9434);
xnor U11981 (N_11981,N_9904,N_10088);
and U11982 (N_11982,N_9853,N_9714);
xor U11983 (N_11983,N_9704,N_10147);
nand U11984 (N_11984,N_9097,N_10145);
and U11985 (N_11985,N_9933,N_9879);
nor U11986 (N_11986,N_9919,N_9114);
nor U11987 (N_11987,N_9735,N_9242);
nand U11988 (N_11988,N_9480,N_10409);
nor U11989 (N_11989,N_9098,N_9556);
or U11990 (N_11990,N_10002,N_10301);
or U11991 (N_11991,N_9375,N_9484);
nor U11992 (N_11992,N_9691,N_10026);
nand U11993 (N_11993,N_9563,N_9732);
or U11994 (N_11994,N_9726,N_9785);
nand U11995 (N_11995,N_9427,N_9763);
xnor U11996 (N_11996,N_10205,N_10352);
nand U11997 (N_11997,N_9866,N_9494);
nand U11998 (N_11998,N_10293,N_9100);
xnor U11999 (N_11999,N_9721,N_9117);
nor U12000 (N_12000,N_11602,N_11949);
or U12001 (N_12001,N_11335,N_11265);
nor U12002 (N_12002,N_10970,N_10894);
nand U12003 (N_12003,N_11820,N_10834);
nand U12004 (N_12004,N_11667,N_11716);
or U12005 (N_12005,N_11543,N_11337);
nor U12006 (N_12006,N_11293,N_10849);
or U12007 (N_12007,N_11141,N_10691);
nand U12008 (N_12008,N_11899,N_10687);
nor U12009 (N_12009,N_11654,N_11438);
nand U12010 (N_12010,N_10920,N_11088);
or U12011 (N_12011,N_11436,N_10637);
or U12012 (N_12012,N_11326,N_11004);
and U12013 (N_12013,N_11897,N_11706);
nand U12014 (N_12014,N_10976,N_10788);
xnor U12015 (N_12015,N_10653,N_10542);
nand U12016 (N_12016,N_11389,N_10762);
nand U12017 (N_12017,N_11940,N_11652);
and U12018 (N_12018,N_10911,N_10501);
nor U12019 (N_12019,N_11947,N_11261);
nand U12020 (N_12020,N_11833,N_10708);
or U12021 (N_12021,N_11270,N_11594);
and U12022 (N_12022,N_11924,N_10775);
nor U12023 (N_12023,N_11577,N_10870);
and U12024 (N_12024,N_11636,N_11403);
nand U12025 (N_12025,N_11761,N_10945);
xor U12026 (N_12026,N_10648,N_10810);
or U12027 (N_12027,N_11368,N_11410);
nand U12028 (N_12028,N_11343,N_11537);
and U12029 (N_12029,N_11483,N_11937);
xnor U12030 (N_12030,N_11530,N_11603);
or U12031 (N_12031,N_11830,N_11212);
or U12032 (N_12032,N_10759,N_10659);
nand U12033 (N_12033,N_11397,N_11251);
or U12034 (N_12034,N_11700,N_10909);
or U12035 (N_12035,N_10889,N_11720);
or U12036 (N_12036,N_10988,N_11339);
or U12037 (N_12037,N_11135,N_11221);
and U12038 (N_12038,N_11945,N_10580);
nor U12039 (N_12039,N_11239,N_11974);
nor U12040 (N_12040,N_10713,N_11510);
or U12041 (N_12041,N_11976,N_11964);
and U12042 (N_12042,N_11763,N_11268);
nor U12043 (N_12043,N_11573,N_11549);
nand U12044 (N_12044,N_11327,N_11130);
xnor U12045 (N_12045,N_11733,N_11844);
and U12046 (N_12046,N_11016,N_11887);
nor U12047 (N_12047,N_10673,N_11640);
nand U12048 (N_12048,N_10836,N_10609);
or U12049 (N_12049,N_11776,N_11439);
or U12050 (N_12050,N_10758,N_10838);
nor U12051 (N_12051,N_10811,N_10517);
nand U12052 (N_12052,N_11402,N_11648);
and U12053 (N_12053,N_10728,N_11091);
and U12054 (N_12054,N_11748,N_10631);
or U12055 (N_12055,N_11172,N_11298);
nand U12056 (N_12056,N_11304,N_11122);
nand U12057 (N_12057,N_11630,N_11711);
nand U12058 (N_12058,N_10956,N_10776);
or U12059 (N_12059,N_11435,N_10533);
nand U12060 (N_12060,N_11723,N_11713);
nand U12061 (N_12061,N_10915,N_11649);
nand U12062 (N_12062,N_11538,N_11236);
nor U12063 (N_12063,N_11767,N_10840);
xor U12064 (N_12064,N_11011,N_11331);
or U12065 (N_12065,N_11226,N_10558);
and U12066 (N_12066,N_10923,N_10954);
nand U12067 (N_12067,N_10783,N_11606);
nand U12068 (N_12068,N_10718,N_11854);
or U12069 (N_12069,N_11764,N_11943);
or U12070 (N_12070,N_10520,N_11249);
or U12071 (N_12071,N_11255,N_11967);
or U12072 (N_12072,N_11120,N_11469);
nand U12073 (N_12073,N_11356,N_11653);
nor U12074 (N_12074,N_10978,N_11787);
xor U12075 (N_12075,N_11592,N_11527);
and U12076 (N_12076,N_10846,N_11639);
and U12077 (N_12077,N_11168,N_11821);
nand U12078 (N_12078,N_10905,N_11097);
nor U12079 (N_12079,N_11416,N_11160);
and U12080 (N_12080,N_11053,N_10750);
or U12081 (N_12081,N_11533,N_10576);
and U12082 (N_12082,N_10716,N_10646);
or U12083 (N_12083,N_10890,N_10872);
or U12084 (N_12084,N_10722,N_11687);
and U12085 (N_12085,N_10596,N_10572);
and U12086 (N_12086,N_11825,N_11045);
or U12087 (N_12087,N_11599,N_10982);
and U12088 (N_12088,N_11256,N_11020);
nand U12089 (N_12089,N_11988,N_11994);
nand U12090 (N_12090,N_11234,N_10527);
nor U12091 (N_12091,N_11086,N_11330);
and U12092 (N_12092,N_11532,N_11412);
or U12093 (N_12093,N_11152,N_10601);
and U12094 (N_12094,N_11065,N_11344);
and U12095 (N_12095,N_11291,N_11593);
nand U12096 (N_12096,N_10743,N_11348);
and U12097 (N_12097,N_11957,N_11398);
and U12098 (N_12098,N_10627,N_11062);
nor U12099 (N_12099,N_11635,N_11218);
nand U12100 (N_12100,N_11448,N_10629);
nor U12101 (N_12101,N_11246,N_11034);
xor U12102 (N_12102,N_11401,N_10806);
or U12103 (N_12103,N_11392,N_10817);
or U12104 (N_12104,N_10655,N_11740);
nand U12105 (N_12105,N_10966,N_11774);
xor U12106 (N_12106,N_11941,N_11874);
nand U12107 (N_12107,N_11881,N_11646);
or U12108 (N_12108,N_11557,N_11801);
or U12109 (N_12109,N_10925,N_11878);
nand U12110 (N_12110,N_11560,N_11472);
or U12111 (N_12111,N_10665,N_11862);
xnor U12112 (N_12112,N_11715,N_10678);
xor U12113 (N_12113,N_11993,N_11497);
or U12114 (N_12114,N_11060,N_10560);
nor U12115 (N_12115,N_11808,N_11243);
nand U12116 (N_12116,N_11800,N_11441);
or U12117 (N_12117,N_11457,N_11111);
and U12118 (N_12118,N_11514,N_11759);
nor U12119 (N_12119,N_11099,N_10825);
nor U12120 (N_12120,N_11032,N_11487);
or U12121 (N_12121,N_10754,N_11424);
and U12122 (N_12122,N_11245,N_11340);
or U12123 (N_12123,N_11718,N_11917);
and U12124 (N_12124,N_10995,N_10525);
or U12125 (N_12125,N_11132,N_10544);
and U12126 (N_12126,N_11328,N_10635);
nor U12127 (N_12127,N_11312,N_11907);
and U12128 (N_12128,N_10599,N_10906);
nand U12129 (N_12129,N_11272,N_11822);
or U12130 (N_12130,N_10582,N_10667);
nand U12131 (N_12131,N_10530,N_11014);
nand U12132 (N_12132,N_10529,N_11714);
nor U12133 (N_12133,N_11253,N_10815);
or U12134 (N_12134,N_11936,N_11427);
and U12135 (N_12135,N_11147,N_10682);
nand U12136 (N_12136,N_10647,N_10763);
nor U12137 (N_12137,N_11562,N_11888);
or U12138 (N_12138,N_11409,N_10510);
nand U12139 (N_12139,N_10656,N_11375);
xnor U12140 (N_12140,N_10607,N_10828);
nor U12141 (N_12141,N_11224,N_11841);
and U12142 (N_12142,N_11214,N_10824);
or U12143 (N_12143,N_11669,N_11208);
nor U12144 (N_12144,N_11975,N_11737);
nand U12145 (N_12145,N_11986,N_11515);
or U12146 (N_12146,N_11999,N_10534);
xnor U12147 (N_12147,N_10803,N_11909);
nand U12148 (N_12148,N_11890,N_11710);
or U12149 (N_12149,N_11428,N_11358);
nand U12150 (N_12150,N_11210,N_11704);
and U12151 (N_12151,N_11213,N_10556);
nand U12152 (N_12152,N_10571,N_10814);
nor U12153 (N_12153,N_11492,N_10855);
xor U12154 (N_12154,N_10700,N_11100);
and U12155 (N_12155,N_10739,N_11432);
or U12156 (N_12156,N_10615,N_11217);
nor U12157 (N_12157,N_11237,N_11419);
nand U12158 (N_12158,N_11123,N_11076);
or U12159 (N_12159,N_11698,N_10674);
nand U12160 (N_12160,N_10518,N_11584);
xnor U12161 (N_12161,N_10622,N_10733);
nand U12162 (N_12162,N_11346,N_11972);
or U12163 (N_12163,N_11165,N_10785);
nand U12164 (N_12164,N_10871,N_10882);
and U12165 (N_12165,N_10774,N_11848);
and U12166 (N_12166,N_11336,N_10677);
nor U12167 (N_12167,N_11205,N_11486);
nand U12168 (N_12168,N_10848,N_11984);
and U12169 (N_12169,N_11528,N_10685);
and U12170 (N_12170,N_11240,N_10809);
or U12171 (N_12171,N_11067,N_11918);
or U12172 (N_12172,N_10614,N_10881);
nand U12173 (N_12173,N_11475,N_11181);
and U12174 (N_12174,N_11354,N_10732);
nand U12175 (N_12175,N_11028,N_10860);
or U12176 (N_12176,N_11650,N_11455);
nor U12177 (N_12177,N_11279,N_11517);
and U12178 (N_12178,N_11285,N_10726);
or U12179 (N_12179,N_11772,N_10816);
and U12180 (N_12180,N_11461,N_10551);
and U12181 (N_12181,N_10568,N_11851);
and U12182 (N_12182,N_11657,N_10742);
nor U12183 (N_12183,N_11660,N_11782);
nor U12184 (N_12184,N_10781,N_10878);
or U12185 (N_12185,N_11038,N_11857);
and U12186 (N_12186,N_10756,N_11571);
nor U12187 (N_12187,N_11842,N_11405);
nor U12188 (N_12188,N_11789,N_11333);
nand U12189 (N_12189,N_11365,N_10786);
nor U12190 (N_12190,N_11547,N_10592);
nand U12191 (N_12191,N_10874,N_10741);
or U12192 (N_12192,N_11791,N_11071);
nand U12193 (N_12193,N_11459,N_11961);
and U12194 (N_12194,N_10654,N_11553);
nor U12195 (N_12195,N_11450,N_11736);
and U12196 (N_12196,N_11509,N_10984);
nor U12197 (N_12197,N_11281,N_11741);
and U12198 (N_12198,N_11480,N_10841);
or U12199 (N_12199,N_11232,N_10536);
xnor U12200 (N_12200,N_10877,N_11896);
and U12201 (N_12201,N_11002,N_11664);
nand U12202 (N_12202,N_10903,N_11443);
nor U12203 (N_12203,N_11575,N_11886);
nand U12204 (N_12204,N_11591,N_11712);
xor U12205 (N_12205,N_11367,N_10710);
and U12206 (N_12206,N_11770,N_10548);
or U12207 (N_12207,N_11058,N_10603);
or U12208 (N_12208,N_11166,N_11678);
or U12209 (N_12209,N_11162,N_11968);
and U12210 (N_12210,N_10644,N_11834);
nand U12211 (N_12211,N_11026,N_11882);
or U12212 (N_12212,N_10546,N_10990);
xor U12213 (N_12213,N_11186,N_10594);
and U12214 (N_12214,N_11777,N_11051);
or U12215 (N_12215,N_11012,N_10935);
nand U12216 (N_12216,N_10693,N_11430);
or U12217 (N_12217,N_10565,N_11950);
nand U12218 (N_12218,N_10624,N_11811);
xor U12219 (N_12219,N_11596,N_10797);
and U12220 (N_12220,N_11452,N_10884);
and U12221 (N_12221,N_11319,N_11148);
or U12222 (N_12222,N_10616,N_10897);
and U12223 (N_12223,N_11925,N_10658);
nand U12224 (N_12224,N_11080,N_10641);
or U12225 (N_12225,N_10961,N_11728);
nand U12226 (N_12226,N_11095,N_11845);
nor U12227 (N_12227,N_11555,N_11338);
nor U12228 (N_12228,N_11534,N_10960);
nor U12229 (N_12229,N_10892,N_11381);
nand U12230 (N_12230,N_11033,N_11204);
and U12231 (N_12231,N_10524,N_11676);
and U12232 (N_12232,N_11329,N_10844);
and U12233 (N_12233,N_10714,N_11729);
or U12234 (N_12234,N_10608,N_11059);
nor U12235 (N_12235,N_11754,N_11793);
and U12236 (N_12236,N_10610,N_11101);
nor U12237 (N_12237,N_11929,N_10737);
and U12238 (N_12238,N_10612,N_11661);
nor U12239 (N_12239,N_11133,N_11695);
nand U12240 (N_12240,N_10927,N_10668);
nand U12241 (N_12241,N_11558,N_11954);
nand U12242 (N_12242,N_11134,N_10886);
nor U12243 (N_12243,N_11103,N_11703);
or U12244 (N_12244,N_11000,N_11173);
nand U12245 (N_12245,N_11373,N_10991);
nand U12246 (N_12246,N_10939,N_11536);
nor U12247 (N_12247,N_11470,N_11273);
nand U12248 (N_12248,N_10583,N_11868);
or U12249 (N_12249,N_11087,N_10839);
nand U12250 (N_12250,N_11316,N_11876);
xnor U12251 (N_12251,N_11969,N_11188);
nor U12252 (N_12252,N_11783,N_11959);
nand U12253 (N_12253,N_11699,N_11719);
nor U12254 (N_12254,N_11609,N_11295);
and U12255 (N_12255,N_11301,N_10706);
or U12256 (N_12256,N_11363,N_10914);
nor U12257 (N_12257,N_10651,N_10888);
nor U12258 (N_12258,N_11563,N_10675);
nand U12259 (N_12259,N_10799,N_11118);
nor U12260 (N_12260,N_10711,N_10953);
nand U12261 (N_12261,N_11075,N_11347);
or U12262 (N_12262,N_11131,N_11149);
nor U12263 (N_12263,N_10657,N_11803);
and U12264 (N_12264,N_11068,N_11495);
xor U12265 (N_12265,N_11275,N_11966);
nor U12266 (N_12266,N_11850,N_11965);
and U12267 (N_12267,N_10724,N_10791);
nand U12268 (N_12268,N_11771,N_10912);
or U12269 (N_12269,N_10857,N_11778);
and U12270 (N_12270,N_10908,N_10503);
and U12271 (N_12271,N_10579,N_11216);
and U12272 (N_12272,N_11855,N_10725);
and U12273 (N_12273,N_11353,N_10879);
nand U12274 (N_12274,N_11473,N_11463);
nand U12275 (N_12275,N_11914,N_11056);
or U12276 (N_12276,N_11980,N_11362);
nand U12277 (N_12277,N_10820,N_10676);
or U12278 (N_12278,N_11681,N_10819);
or U12279 (N_12279,N_11057,N_10697);
nand U12280 (N_12280,N_11502,N_11142);
nor U12281 (N_12281,N_10921,N_11422);
nor U12282 (N_12282,N_11171,N_11183);
nand U12283 (N_12283,N_10940,N_10863);
or U12284 (N_12284,N_10757,N_11048);
nor U12285 (N_12285,N_11751,N_11624);
and U12286 (N_12286,N_11137,N_10766);
or U12287 (N_12287,N_11582,N_11437);
and U12288 (N_12288,N_10620,N_11668);
nor U12289 (N_12289,N_11197,N_10867);
and U12290 (N_12290,N_11773,N_11548);
nor U12291 (N_12291,N_10919,N_11756);
nor U12292 (N_12292,N_11840,N_11616);
and U12293 (N_12293,N_10535,N_10952);
nand U12294 (N_12294,N_11228,N_11449);
nor U12295 (N_12295,N_11901,N_10744);
xnor U12296 (N_12296,N_11015,N_11580);
nor U12297 (N_12297,N_11796,N_10949);
and U12298 (N_12298,N_11146,N_11471);
nand U12299 (N_12299,N_11550,N_11102);
xor U12300 (N_12300,N_10512,N_10507);
or U12301 (N_12301,N_10618,N_11613);
xor U12302 (N_12302,N_11612,N_11190);
or U12303 (N_12303,N_10661,N_10550);
or U12304 (N_12304,N_10928,N_11590);
xor U12305 (N_12305,N_11371,N_10689);
nor U12306 (N_12306,N_11566,N_11174);
nor U12307 (N_12307,N_11317,N_11730);
and U12308 (N_12308,N_10793,N_11523);
and U12309 (N_12309,N_11926,N_11286);
and U12310 (N_12310,N_10847,N_11278);
or U12311 (N_12311,N_11179,N_11040);
nor U12312 (N_12312,N_11692,N_10532);
or U12313 (N_12313,N_10734,N_11116);
or U12314 (N_12314,N_10539,N_11884);
nand U12315 (N_12315,N_11474,N_11696);
nand U12316 (N_12316,N_11445,N_11956);
nor U12317 (N_12317,N_10736,N_11476);
nor U12318 (N_12318,N_11913,N_11078);
or U12319 (N_12319,N_10628,N_11376);
or U12320 (N_12320,N_10513,N_11390);
and U12321 (N_12321,N_11456,N_11154);
nor U12322 (N_12322,N_11288,N_11490);
or U12323 (N_12323,N_11683,N_11505);
or U12324 (N_12324,N_11911,N_11853);
or U12325 (N_12325,N_11638,N_10772);
or U12326 (N_12326,N_11079,N_10997);
nor U12327 (N_12327,N_11489,N_11063);
nor U12328 (N_12328,N_11581,N_10898);
nor U12329 (N_12329,N_11735,N_11223);
nand U12330 (N_12330,N_11423,N_11479);
nand U12331 (N_12331,N_11185,N_11037);
nand U12332 (N_12332,N_11561,N_10932);
and U12333 (N_12333,N_11644,N_11995);
or U12334 (N_12334,N_11587,N_11421);
nand U12335 (N_12335,N_11666,N_10515);
nand U12336 (N_12336,N_10778,N_10973);
nor U12337 (N_12337,N_11642,N_10942);
xor U12338 (N_12338,N_10969,N_11411);
nand U12339 (N_12339,N_10557,N_11379);
nor U12340 (N_12340,N_11151,N_10951);
or U12341 (N_12341,N_11749,N_10777);
or U12342 (N_12342,N_10831,N_11167);
nor U12343 (N_12343,N_11879,N_11585);
and U12344 (N_12344,N_10818,N_10796);
nand U12345 (N_12345,N_10703,N_11084);
and U12346 (N_12346,N_11418,N_11935);
and U12347 (N_12347,N_11110,N_11175);
or U12348 (N_12348,N_10679,N_11035);
and U12349 (N_12349,N_10975,N_11992);
nor U12350 (N_12350,N_11104,N_10562);
and U12351 (N_12351,N_11637,N_11271);
and U12352 (N_12352,N_10980,N_11209);
nand U12353 (N_12353,N_11578,N_11750);
xnor U12354 (N_12354,N_11634,N_10790);
nand U12355 (N_12355,N_10643,N_10979);
or U12356 (N_12356,N_11394,N_10729);
and U12357 (N_12357,N_11629,N_10993);
xor U12358 (N_12358,N_10563,N_11780);
nand U12359 (N_12359,N_10586,N_11541);
and U12360 (N_12360,N_11518,N_11207);
or U12361 (N_12361,N_11570,N_10701);
xor U12362 (N_12362,N_11395,N_11934);
or U12363 (N_12363,N_10985,N_11485);
nand U12364 (N_12364,N_11701,N_11478);
nand U12365 (N_12365,N_11831,N_10506);
nor U12366 (N_12366,N_11072,N_10924);
or U12367 (N_12367,N_10934,N_11039);
xor U12368 (N_12368,N_11085,N_10694);
xor U12369 (N_12369,N_11090,N_11586);
or U12370 (N_12370,N_11906,N_11551);
nor U12371 (N_12371,N_10639,N_11313);
nor U12372 (N_12372,N_10864,N_10642);
nor U12373 (N_12373,N_10917,N_10584);
or U12374 (N_12374,N_11227,N_11477);
or U12375 (N_12375,N_11184,N_10543);
nand U12376 (N_12376,N_10843,N_10595);
or U12377 (N_12377,N_11798,N_10965);
nor U12378 (N_12378,N_11302,N_11425);
nor U12379 (N_12379,N_11177,N_10523);
nor U12380 (N_12380,N_11768,N_10823);
nand U12381 (N_12381,N_10688,N_11453);
and U12382 (N_12382,N_10904,N_11804);
xnor U12383 (N_12383,N_10613,N_11875);
xnor U12384 (N_12384,N_10862,N_11196);
nand U12385 (N_12385,N_11126,N_10626);
nand U12386 (N_12386,N_11267,N_10514);
or U12387 (N_12387,N_11828,N_10946);
nand U12388 (N_12388,N_10910,N_11277);
and U12389 (N_12389,N_11870,N_11786);
nor U12390 (N_12390,N_10638,N_11195);
nand U12391 (N_12391,N_11501,N_10981);
or U12392 (N_12392,N_11274,N_11178);
and U12393 (N_12393,N_10891,N_11539);
xnor U12394 (N_12394,N_11567,N_10950);
or U12395 (N_12395,N_11109,N_10521);
xor U12396 (N_12396,N_11465,N_11601);
or U12397 (N_12397,N_11807,N_11454);
nor U12398 (N_12398,N_11632,N_11055);
nor U12399 (N_12399,N_11872,N_11694);
nor U12400 (N_12400,N_11709,N_11960);
and U12401 (N_12401,N_11050,N_10865);
or U12402 (N_12402,N_11556,N_11247);
nand U12403 (N_12403,N_11662,N_11743);
and U12404 (N_12404,N_10999,N_11838);
and U12405 (N_12405,N_11989,N_11342);
nor U12406 (N_12406,N_11607,N_11372);
or U12407 (N_12407,N_10931,N_11623);
and U12408 (N_12408,N_11380,N_10705);
nand U12409 (N_12409,N_11157,N_11987);
or U12410 (N_12410,N_10972,N_10606);
nor U12411 (N_12411,N_11521,N_11910);
nor U12412 (N_12412,N_11932,N_11355);
and U12413 (N_12413,N_11985,N_11235);
xor U12414 (N_12414,N_11615,N_11108);
or U12415 (N_12415,N_10866,N_11413);
and U12416 (N_12416,N_11017,N_10587);
and U12417 (N_12417,N_10854,N_11282);
nand U12418 (N_12418,N_11835,N_11839);
nor U12419 (N_12419,N_10761,N_11306);
nand U12420 (N_12420,N_11023,N_11025);
nor U12421 (N_12421,N_10958,N_11684);
nor U12422 (N_12422,N_11626,N_11369);
or U12423 (N_12423,N_11944,N_11263);
or U12424 (N_12424,N_11873,N_11627);
nor U12425 (N_12425,N_11797,N_11574);
nor U12426 (N_12426,N_11921,N_10663);
nor U12427 (N_12427,N_11724,N_10893);
nor U12428 (N_12428,N_11908,N_10929);
nor U12429 (N_12429,N_11462,N_10948);
or U12430 (N_12430,N_11927,N_11524);
nand U12431 (N_12431,N_11019,N_11597);
and U12432 (N_12432,N_11849,N_10549);
nor U12433 (N_12433,N_11136,N_11902);
nand U12434 (N_12434,N_11903,N_10875);
or U12435 (N_12435,N_10753,N_11589);
and U12436 (N_12436,N_11145,N_10826);
nor U12437 (N_12437,N_10787,N_10686);
and U12438 (N_12438,N_11303,N_10941);
or U12439 (N_12439,N_10770,N_10692);
nor U12440 (N_12440,N_10621,N_11052);
nand U12441 (N_12441,N_10664,N_11983);
or U12442 (N_12442,N_11760,N_11143);
nor U12443 (N_12443,N_10611,N_10504);
nand U12444 (N_12444,N_11468,N_11013);
or U12445 (N_12445,N_10570,N_11112);
or U12446 (N_12446,N_11388,N_11665);
nor U12447 (N_12447,N_10566,N_10630);
or U12448 (N_12448,N_10715,N_11264);
or U12449 (N_12449,N_11350,N_11933);
and U12450 (N_12450,N_11258,N_10943);
or U12451 (N_12451,N_11127,N_11106);
nor U12452 (N_12452,N_11257,N_10930);
nor U12453 (N_12453,N_10555,N_10869);
and U12454 (N_12454,N_10680,N_11150);
and U12455 (N_12455,N_11201,N_10760);
or U12456 (N_12456,N_11415,N_11215);
or U12457 (N_12457,N_10681,N_11442);
and U12458 (N_12458,N_10947,N_11203);
and U12459 (N_12459,N_11066,N_11098);
xnor U12460 (N_12460,N_11794,N_10649);
xor U12461 (N_12461,N_11739,N_10617);
and U12462 (N_12462,N_11507,N_10821);
or U12463 (N_12463,N_11022,N_11202);
nand U12464 (N_12464,N_11220,N_10845);
or U12465 (N_12465,N_10748,N_11323);
or U12466 (N_12466,N_11007,N_11512);
and U12467 (N_12467,N_11250,N_11813);
xor U12468 (N_12468,N_10578,N_10850);
nand U12469 (N_12469,N_11546,N_10896);
nor U12470 (N_12470,N_10807,N_11310);
xor U12471 (N_12471,N_11314,N_11341);
nor U12472 (N_12472,N_11805,N_11900);
nand U12473 (N_12473,N_10597,N_10567);
or U12474 (N_12474,N_11466,N_11345);
nand U12475 (N_12475,N_11604,N_11792);
or U12476 (N_12476,N_10669,N_11655);
nand U12477 (N_12477,N_10559,N_11672);
nor U12478 (N_12478,N_10684,N_11904);
nand U12479 (N_12479,N_11292,N_11180);
and U12480 (N_12480,N_10640,N_11554);
xnor U12481 (N_12481,N_11433,N_11970);
xor U12482 (N_12482,N_11894,N_11458);
xnor U12483 (N_12483,N_11755,N_11083);
and U12484 (N_12484,N_10625,N_10900);
nand U12485 (N_12485,N_10695,N_11565);
or U12486 (N_12486,N_10859,N_11732);
and U12487 (N_12487,N_11262,N_10650);
or U12488 (N_12488,N_10505,N_10913);
and U12489 (N_12489,N_11318,N_10690);
or U12490 (N_12490,N_11259,N_10998);
nand U12491 (N_12491,N_11817,N_10907);
nor U12492 (N_12492,N_10508,N_10589);
nor U12493 (N_12493,N_11069,N_10996);
or U12494 (N_12494,N_11816,N_11287);
nand U12495 (N_12495,N_11529,N_11193);
xnor U12496 (N_12496,N_11745,N_11544);
or U12497 (N_12497,N_10632,N_11559);
and U12498 (N_12498,N_10660,N_11349);
or U12499 (N_12499,N_11107,N_11406);
or U12500 (N_12500,N_11351,N_10957);
or U12501 (N_12501,N_11315,N_10740);
and U12502 (N_12502,N_11446,N_11895);
nand U12503 (N_12503,N_11385,N_10955);
and U12504 (N_12504,N_11790,N_11958);
and U12505 (N_12505,N_10746,N_11915);
and U12506 (N_12506,N_11981,N_10944);
nand U12507 (N_12507,N_11920,N_11496);
nand U12508 (N_12508,N_10738,N_10830);
and U12509 (N_12509,N_11440,N_11753);
xor U12510 (N_12510,N_11189,N_11155);
and U12511 (N_12511,N_11404,N_10699);
nor U12512 (N_12512,N_11407,N_11863);
or U12513 (N_12513,N_11871,N_11861);
nand U12514 (N_12514,N_10901,N_11742);
or U12515 (N_12515,N_10696,N_11620);
nor U12516 (N_12516,N_11552,N_11765);
nor U12517 (N_12517,N_10794,N_10749);
nor U12518 (N_12518,N_11880,N_11621);
and U12519 (N_12519,N_11885,N_11625);
or U12520 (N_12520,N_11889,N_11766);
nor U12521 (N_12521,N_11384,N_10540);
or U12522 (N_12522,N_10755,N_11856);
nor U12523 (N_12523,N_11916,N_10538);
nor U12524 (N_12524,N_11296,N_11628);
and U12525 (N_12525,N_11826,N_11818);
and U12526 (N_12526,N_10994,N_11260);
nand U12527 (N_12527,N_10519,N_11008);
xor U12528 (N_12528,N_10500,N_11357);
nand U12529 (N_12529,N_11891,N_11311);
nor U12530 (N_12530,N_11633,N_11158);
nand U12531 (N_12531,N_11883,N_11568);
xor U12532 (N_12532,N_11081,N_10709);
and U12533 (N_12533,N_10902,N_10581);
nand U12534 (N_12534,N_11722,N_11061);
nor U12535 (N_12535,N_11417,N_10832);
or U12536 (N_12536,N_11866,N_11192);
nand U12537 (N_12537,N_11758,N_10598);
nand U12538 (N_12538,N_11041,N_11673);
xor U12539 (N_12539,N_11810,N_10789);
nand U12540 (N_12540,N_10856,N_10842);
or U12541 (N_12541,N_11182,N_11785);
or U12542 (N_12542,N_11491,N_11674);
and U12543 (N_12543,N_11645,N_11161);
and U12544 (N_12544,N_11252,N_10666);
nand U12545 (N_12545,N_11860,N_11289);
nand U12546 (N_12546,N_11176,N_10735);
or U12547 (N_12547,N_11093,N_10619);
nor U12548 (N_12548,N_10683,N_11996);
xnor U12549 (N_12549,N_11688,N_11070);
nor U12550 (N_12550,N_11869,N_10767);
nor U12551 (N_12551,N_11955,N_11690);
or U12552 (N_12552,N_10959,N_11641);
nand U12553 (N_12553,N_11089,N_11024);
or U12554 (N_12554,N_11129,N_11321);
nand U12555 (N_12555,N_10717,N_11299);
and U12556 (N_12556,N_11018,N_11021);
nor U12557 (N_12557,N_11843,N_10773);
and U12558 (N_12558,N_10916,N_11781);
nand U12559 (N_12559,N_11977,N_11656);
nor U12560 (N_12560,N_11734,N_10964);
or U12561 (N_12561,N_11663,N_10808);
and U12562 (N_12562,N_11611,N_11386);
nand U12563 (N_12563,N_11322,N_11504);
and U12564 (N_12564,N_11159,N_10764);
nor U12565 (N_12565,N_11588,N_10782);
or U12566 (N_12566,N_11036,N_10765);
nand U12567 (N_12567,N_11671,N_11324);
nand U12568 (N_12568,N_10822,N_10798);
nand U12569 (N_12569,N_11200,N_11429);
or U12570 (N_12570,N_11717,N_11010);
and U12571 (N_12571,N_11511,N_10604);
xnor U12572 (N_12572,N_10779,N_10813);
xnor U12573 (N_12573,N_10593,N_11516);
nand U12574 (N_12574,N_11608,N_11928);
and U12575 (N_12575,N_11500,N_11484);
nand U12576 (N_12576,N_11211,N_11689);
xor U12577 (N_12577,N_10992,N_11997);
nor U12578 (N_12578,N_10805,N_11451);
and U12579 (N_12579,N_11283,N_11998);
nor U12580 (N_12580,N_10868,N_11726);
or U12581 (N_12581,N_11991,N_10747);
or U12582 (N_12582,N_11266,N_10623);
and U12583 (N_12583,N_11962,N_11113);
and U12584 (N_12584,N_11074,N_11003);
nand U12585 (N_12585,N_11948,N_10745);
and U12586 (N_12586,N_11332,N_10633);
nand U12587 (N_12587,N_10983,N_11054);
nor U12588 (N_12588,N_10835,N_11795);
or U12589 (N_12589,N_10752,N_11679);
nand U12590 (N_12590,N_11513,N_11115);
and U12591 (N_12591,N_11614,N_11752);
xnor U12592 (N_12592,N_10707,N_11946);
or U12593 (N_12593,N_11520,N_10522);
and U12594 (N_12594,N_10968,N_11309);
nand U12595 (N_12595,N_11930,N_11400);
nand U12596 (N_12596,N_11610,N_11697);
nand U12597 (N_12597,N_10883,N_11294);
nand U12598 (N_12598,N_10802,N_11721);
or U12599 (N_12599,N_11824,N_11702);
nand U12600 (N_12600,N_10564,N_11675);
nand U12601 (N_12601,N_10989,N_11467);
nor U12602 (N_12602,N_11494,N_11815);
and U12603 (N_12603,N_10730,N_11762);
nand U12604 (N_12604,N_11535,N_10895);
or U12605 (N_12605,N_10552,N_11374);
and U12606 (N_12606,N_10918,N_11540);
or U12607 (N_12607,N_11393,N_11414);
or U12608 (N_12608,N_11125,N_10926);
and U12609 (N_12609,N_11979,N_11242);
nor U12610 (N_12610,N_10780,N_10547);
or U12611 (N_12611,N_10670,N_11049);
or U12612 (N_12612,N_10858,N_11460);
or U12613 (N_12613,N_10880,N_11498);
nor U12614 (N_12614,N_11042,N_11846);
nor U12615 (N_12615,N_11757,N_10569);
nor U12616 (N_12616,N_11044,N_10727);
nand U12617 (N_12617,N_11128,N_10971);
nor U12618 (N_12618,N_10590,N_11297);
or U12619 (N_12619,N_11230,N_11583);
nor U12620 (N_12620,N_11938,N_11680);
nand U12621 (N_12621,N_11809,N_11659);
nor U12622 (N_12622,N_10634,N_10833);
nor U12623 (N_12623,N_11225,N_11576);
nor U12624 (N_12624,N_10537,N_11140);
and U12625 (N_12625,N_10645,N_11092);
and U12626 (N_12626,N_11788,N_11525);
and U12627 (N_12627,N_11852,N_10731);
nor U12628 (N_12628,N_11094,N_11170);
xnor U12629 (N_12629,N_10652,N_11931);
and U12630 (N_12630,N_11579,N_11799);
and U12631 (N_12631,N_11290,N_10804);
or U12632 (N_12632,N_11307,N_11686);
and U12633 (N_12633,N_10575,N_11163);
nor U12634 (N_12634,N_11951,N_11522);
and U12635 (N_12635,N_11334,N_11647);
xnor U12636 (N_12636,N_11222,N_11464);
nand U12637 (N_12637,N_11391,N_10636);
nor U12638 (N_12638,N_11806,N_11031);
nand U12639 (N_12639,N_11677,N_11444);
and U12640 (N_12640,N_10977,N_11238);
and U12641 (N_12641,N_11707,N_11631);
and U12642 (N_12642,N_10986,N_10936);
nor U12643 (N_12643,N_11731,N_10800);
nor U12644 (N_12644,N_11519,N_10937);
or U12645 (N_12645,N_11194,N_11531);
nor U12646 (N_12646,N_11827,N_10554);
nor U12647 (N_12647,N_11506,N_11124);
or U12648 (N_12648,N_11206,N_11378);
nor U12649 (N_12649,N_10829,N_11847);
nor U12650 (N_12650,N_11138,N_11325);
nor U12651 (N_12651,N_11953,N_11396);
nand U12652 (N_12652,N_11082,N_11682);
or U12653 (N_12653,N_10887,N_11744);
and U12654 (N_12654,N_11139,N_11865);
or U12655 (N_12655,N_11233,N_11364);
nor U12656 (N_12656,N_10577,N_11705);
and U12657 (N_12657,N_10852,N_11829);
nand U12658 (N_12658,N_11658,N_11605);
nor U12659 (N_12659,N_11982,N_11426);
or U12660 (N_12660,N_11009,N_11978);
xor U12661 (N_12661,N_10720,N_11905);
nand U12662 (N_12662,N_11499,N_11867);
or U12663 (N_12663,N_11893,N_10795);
xnor U12664 (N_12664,N_11963,N_11858);
and U12665 (N_12665,N_11305,N_11359);
nor U12666 (N_12666,N_11229,N_11030);
or U12667 (N_12667,N_11725,N_11399);
nor U12668 (N_12668,N_11670,N_11244);
xor U12669 (N_12669,N_11187,N_11027);
nor U12670 (N_12670,N_11096,N_10509);
nand U12671 (N_12671,N_11361,N_11814);
nand U12672 (N_12672,N_10792,N_11117);
or U12673 (N_12673,N_10502,N_10974);
nor U12674 (N_12674,N_11043,N_10531);
xor U12675 (N_12675,N_11819,N_11542);
or U12676 (N_12676,N_11493,N_11382);
or U12677 (N_12677,N_11990,N_11370);
nand U12678 (N_12678,N_11005,N_11508);
nand U12679 (N_12679,N_11064,N_11923);
or U12680 (N_12680,N_11300,N_10873);
and U12681 (N_12681,N_10561,N_11939);
nor U12682 (N_12682,N_11823,N_10702);
xor U12683 (N_12683,N_11617,N_10837);
nand U12684 (N_12684,N_10541,N_10511);
nor U12685 (N_12685,N_11779,N_11942);
nand U12686 (N_12686,N_11526,N_11892);
nor U12687 (N_12687,N_11600,N_11708);
nand U12688 (N_12688,N_11691,N_11366);
nor U12689 (N_12689,N_11481,N_11775);
nor U12690 (N_12690,N_11269,N_10933);
or U12691 (N_12691,N_11029,N_10526);
nor U12692 (N_12692,N_11727,N_10602);
and U12693 (N_12693,N_10719,N_11219);
nand U12694 (N_12694,N_10922,N_11308);
nand U12695 (N_12695,N_10885,N_11564);
and U12696 (N_12696,N_11859,N_11121);
nor U12697 (N_12697,N_11352,N_10812);
nand U12698 (N_12698,N_11280,N_11420);
nor U12699 (N_12699,N_10528,N_10698);
or U12700 (N_12700,N_11431,N_10962);
nor U12701 (N_12701,N_10938,N_11073);
xnor U12702 (N_12702,N_11198,N_11254);
nor U12703 (N_12703,N_10827,N_11952);
or U12704 (N_12704,N_11387,N_11545);
xor U12705 (N_12705,N_10967,N_11482);
nand U12706 (N_12706,N_11276,N_11919);
nor U12707 (N_12707,N_11746,N_11769);
xor U12708 (N_12708,N_10899,N_11832);
nand U12709 (N_12709,N_11408,N_11119);
nor U12710 (N_12710,N_11284,N_11738);
xnor U12711 (N_12711,N_11144,N_10861);
xor U12712 (N_12712,N_11572,N_10801);
or U12713 (N_12713,N_11877,N_10784);
or U12714 (N_12714,N_11434,N_11047);
nor U12715 (N_12715,N_11837,N_11377);
or U12716 (N_12716,N_10721,N_11488);
and U12717 (N_12717,N_10769,N_11618);
nand U12718 (N_12718,N_11651,N_11802);
nor U12719 (N_12719,N_10771,N_11973);
and U12720 (N_12720,N_10662,N_11169);
or U12721 (N_12721,N_11320,N_10516);
and U12722 (N_12722,N_11114,N_10704);
nor U12723 (N_12723,N_11619,N_10600);
and U12724 (N_12724,N_10573,N_11812);
nor U12725 (N_12725,N_11191,N_11164);
or U12726 (N_12726,N_10768,N_11685);
and U12727 (N_12727,N_11383,N_11077);
xnor U12728 (N_12728,N_11864,N_11248);
nor U12729 (N_12729,N_10671,N_10712);
and U12730 (N_12730,N_10751,N_10545);
xor U12731 (N_12731,N_11447,N_10853);
or U12732 (N_12732,N_11971,N_11622);
and U12733 (N_12733,N_11598,N_11001);
nand U12734 (N_12734,N_11898,N_11231);
nor U12735 (N_12735,N_11006,N_10553);
or U12736 (N_12736,N_11503,N_10591);
or U12737 (N_12737,N_10605,N_11784);
or U12738 (N_12738,N_10574,N_10588);
nand U12739 (N_12739,N_11595,N_11199);
and U12740 (N_12740,N_11569,N_10723);
nand U12741 (N_12741,N_11241,N_11912);
nand U12742 (N_12742,N_11922,N_11360);
and U12743 (N_12743,N_11046,N_10672);
or U12744 (N_12744,N_11693,N_10876);
or U12745 (N_12745,N_11643,N_11747);
and U12746 (N_12746,N_11105,N_10585);
or U12747 (N_12747,N_10963,N_11156);
xnor U12748 (N_12748,N_11836,N_11153);
nand U12749 (N_12749,N_10851,N_10987);
xor U12750 (N_12750,N_11227,N_10538);
xor U12751 (N_12751,N_11327,N_10839);
and U12752 (N_12752,N_11485,N_10891);
nand U12753 (N_12753,N_10622,N_11191);
and U12754 (N_12754,N_11645,N_11274);
or U12755 (N_12755,N_11126,N_11496);
and U12756 (N_12756,N_10813,N_11637);
nor U12757 (N_12757,N_10654,N_11594);
nor U12758 (N_12758,N_11486,N_11467);
or U12759 (N_12759,N_10590,N_10971);
nor U12760 (N_12760,N_11862,N_10644);
and U12761 (N_12761,N_10907,N_10839);
nor U12762 (N_12762,N_11853,N_11770);
nand U12763 (N_12763,N_11786,N_11468);
or U12764 (N_12764,N_11650,N_11121);
nor U12765 (N_12765,N_10937,N_10806);
nand U12766 (N_12766,N_10965,N_11098);
and U12767 (N_12767,N_10789,N_10769);
nand U12768 (N_12768,N_11500,N_11872);
nor U12769 (N_12769,N_11382,N_11199);
xnor U12770 (N_12770,N_10548,N_11554);
and U12771 (N_12771,N_10791,N_10932);
or U12772 (N_12772,N_11829,N_11959);
nand U12773 (N_12773,N_11239,N_11576);
and U12774 (N_12774,N_11363,N_11831);
nor U12775 (N_12775,N_11935,N_11433);
nor U12776 (N_12776,N_11136,N_11452);
or U12777 (N_12777,N_11482,N_11532);
nand U12778 (N_12778,N_10707,N_10879);
nor U12779 (N_12779,N_11153,N_10923);
or U12780 (N_12780,N_10827,N_11611);
nand U12781 (N_12781,N_11037,N_11169);
and U12782 (N_12782,N_11985,N_11391);
or U12783 (N_12783,N_10558,N_11571);
nand U12784 (N_12784,N_10526,N_11799);
or U12785 (N_12785,N_11640,N_11667);
nand U12786 (N_12786,N_11442,N_11907);
or U12787 (N_12787,N_11634,N_11418);
and U12788 (N_12788,N_10730,N_10757);
or U12789 (N_12789,N_11082,N_11484);
nand U12790 (N_12790,N_11266,N_11454);
and U12791 (N_12791,N_10931,N_10880);
and U12792 (N_12792,N_11021,N_11721);
and U12793 (N_12793,N_11798,N_11390);
nor U12794 (N_12794,N_10726,N_11587);
and U12795 (N_12795,N_10657,N_11764);
nor U12796 (N_12796,N_11899,N_11651);
xor U12797 (N_12797,N_11592,N_11292);
or U12798 (N_12798,N_10626,N_11726);
nand U12799 (N_12799,N_11683,N_10924);
nor U12800 (N_12800,N_11003,N_11469);
nor U12801 (N_12801,N_11586,N_11870);
xnor U12802 (N_12802,N_11842,N_11312);
nor U12803 (N_12803,N_11018,N_11134);
nand U12804 (N_12804,N_11175,N_11995);
nor U12805 (N_12805,N_10967,N_11677);
or U12806 (N_12806,N_10858,N_11559);
or U12807 (N_12807,N_11173,N_11145);
nor U12808 (N_12808,N_10992,N_11655);
nand U12809 (N_12809,N_11048,N_10546);
nor U12810 (N_12810,N_10689,N_10730);
nand U12811 (N_12811,N_11737,N_11773);
nor U12812 (N_12812,N_11506,N_11030);
nand U12813 (N_12813,N_11514,N_11096);
xor U12814 (N_12814,N_10561,N_11953);
nand U12815 (N_12815,N_10789,N_10528);
and U12816 (N_12816,N_11196,N_11246);
nand U12817 (N_12817,N_10881,N_11692);
and U12818 (N_12818,N_11515,N_10650);
or U12819 (N_12819,N_10684,N_11049);
and U12820 (N_12820,N_11680,N_10731);
and U12821 (N_12821,N_11458,N_11469);
nand U12822 (N_12822,N_11869,N_11723);
nor U12823 (N_12823,N_10929,N_11631);
and U12824 (N_12824,N_11668,N_10934);
or U12825 (N_12825,N_10715,N_10723);
xor U12826 (N_12826,N_11018,N_11226);
nand U12827 (N_12827,N_11377,N_10601);
xor U12828 (N_12828,N_11355,N_11918);
nand U12829 (N_12829,N_11900,N_11014);
xor U12830 (N_12830,N_10714,N_10927);
xnor U12831 (N_12831,N_10593,N_11025);
or U12832 (N_12832,N_11290,N_11190);
and U12833 (N_12833,N_11341,N_11305);
and U12834 (N_12834,N_11794,N_10846);
nor U12835 (N_12835,N_11684,N_11362);
or U12836 (N_12836,N_10845,N_11138);
nor U12837 (N_12837,N_10983,N_11903);
nand U12838 (N_12838,N_10533,N_11165);
and U12839 (N_12839,N_11389,N_11085);
xor U12840 (N_12840,N_10578,N_10800);
nand U12841 (N_12841,N_11528,N_11103);
nand U12842 (N_12842,N_10598,N_11986);
nor U12843 (N_12843,N_11675,N_10782);
xor U12844 (N_12844,N_10658,N_10652);
nor U12845 (N_12845,N_11843,N_11919);
nand U12846 (N_12846,N_11521,N_11786);
or U12847 (N_12847,N_11773,N_11188);
nand U12848 (N_12848,N_10578,N_11860);
nor U12849 (N_12849,N_10644,N_11521);
or U12850 (N_12850,N_11366,N_11540);
nand U12851 (N_12851,N_11322,N_11370);
and U12852 (N_12852,N_11603,N_10866);
nor U12853 (N_12853,N_11784,N_11221);
nand U12854 (N_12854,N_11970,N_10571);
and U12855 (N_12855,N_11441,N_11435);
or U12856 (N_12856,N_10781,N_11722);
nand U12857 (N_12857,N_10811,N_10701);
and U12858 (N_12858,N_11815,N_11140);
nand U12859 (N_12859,N_11200,N_10708);
nor U12860 (N_12860,N_11271,N_11200);
nand U12861 (N_12861,N_11041,N_11955);
xor U12862 (N_12862,N_11595,N_10782);
xnor U12863 (N_12863,N_11538,N_10884);
nor U12864 (N_12864,N_10605,N_11440);
xor U12865 (N_12865,N_10844,N_11514);
nor U12866 (N_12866,N_11463,N_11914);
and U12867 (N_12867,N_11242,N_11901);
xor U12868 (N_12868,N_11411,N_11233);
xor U12869 (N_12869,N_11393,N_10850);
xnor U12870 (N_12870,N_10637,N_11607);
nand U12871 (N_12871,N_11362,N_11199);
or U12872 (N_12872,N_11148,N_11592);
nand U12873 (N_12873,N_10905,N_11242);
or U12874 (N_12874,N_10630,N_11672);
or U12875 (N_12875,N_11711,N_10506);
nand U12876 (N_12876,N_11226,N_10873);
and U12877 (N_12877,N_10628,N_11171);
nor U12878 (N_12878,N_11250,N_11873);
nand U12879 (N_12879,N_11804,N_11280);
xnor U12880 (N_12880,N_10636,N_11740);
and U12881 (N_12881,N_11231,N_11317);
nand U12882 (N_12882,N_11063,N_11065);
or U12883 (N_12883,N_11630,N_10776);
or U12884 (N_12884,N_10991,N_11464);
nand U12885 (N_12885,N_11681,N_11506);
nor U12886 (N_12886,N_11101,N_10981);
and U12887 (N_12887,N_11768,N_11776);
and U12888 (N_12888,N_11522,N_11240);
xnor U12889 (N_12889,N_10935,N_11169);
or U12890 (N_12890,N_11232,N_11948);
xnor U12891 (N_12891,N_10992,N_11982);
and U12892 (N_12892,N_11405,N_11374);
or U12893 (N_12893,N_11612,N_10835);
and U12894 (N_12894,N_10971,N_11467);
nand U12895 (N_12895,N_11863,N_11749);
xor U12896 (N_12896,N_10623,N_11138);
nand U12897 (N_12897,N_10974,N_11642);
and U12898 (N_12898,N_11152,N_11632);
nand U12899 (N_12899,N_10951,N_10534);
nand U12900 (N_12900,N_11405,N_11838);
nand U12901 (N_12901,N_11635,N_11787);
nor U12902 (N_12902,N_10725,N_11584);
nor U12903 (N_12903,N_11323,N_11026);
or U12904 (N_12904,N_10890,N_11211);
nor U12905 (N_12905,N_11936,N_10953);
or U12906 (N_12906,N_11371,N_11921);
or U12907 (N_12907,N_11788,N_10514);
nand U12908 (N_12908,N_10569,N_11405);
or U12909 (N_12909,N_10688,N_11583);
nor U12910 (N_12910,N_11664,N_11356);
and U12911 (N_12911,N_11225,N_10886);
and U12912 (N_12912,N_11942,N_10773);
and U12913 (N_12913,N_11331,N_11363);
nand U12914 (N_12914,N_11891,N_11700);
and U12915 (N_12915,N_11505,N_11829);
or U12916 (N_12916,N_11797,N_11072);
or U12917 (N_12917,N_10914,N_11483);
nand U12918 (N_12918,N_10806,N_11802);
or U12919 (N_12919,N_11617,N_11616);
xor U12920 (N_12920,N_10797,N_10678);
and U12921 (N_12921,N_11041,N_10586);
or U12922 (N_12922,N_11080,N_11861);
or U12923 (N_12923,N_11254,N_10787);
nor U12924 (N_12924,N_10847,N_11122);
or U12925 (N_12925,N_11867,N_10893);
and U12926 (N_12926,N_11913,N_11874);
and U12927 (N_12927,N_10609,N_11690);
or U12928 (N_12928,N_11368,N_11241);
and U12929 (N_12929,N_11319,N_10513);
nand U12930 (N_12930,N_11590,N_11535);
xnor U12931 (N_12931,N_11677,N_11749);
nand U12932 (N_12932,N_11091,N_11683);
nor U12933 (N_12933,N_11140,N_10820);
nor U12934 (N_12934,N_10760,N_10559);
and U12935 (N_12935,N_11900,N_11020);
nor U12936 (N_12936,N_11740,N_11173);
and U12937 (N_12937,N_11456,N_10993);
or U12938 (N_12938,N_11469,N_11892);
or U12939 (N_12939,N_11584,N_11580);
nand U12940 (N_12940,N_11052,N_11668);
xnor U12941 (N_12941,N_11754,N_11410);
and U12942 (N_12942,N_11252,N_10543);
xor U12943 (N_12943,N_11084,N_11941);
nor U12944 (N_12944,N_11990,N_11419);
and U12945 (N_12945,N_11443,N_11560);
or U12946 (N_12946,N_11336,N_11294);
or U12947 (N_12947,N_11612,N_11698);
nand U12948 (N_12948,N_11327,N_10979);
or U12949 (N_12949,N_11517,N_11425);
nor U12950 (N_12950,N_11704,N_11339);
or U12951 (N_12951,N_11284,N_10907);
and U12952 (N_12952,N_10979,N_11250);
nor U12953 (N_12953,N_11541,N_11571);
nor U12954 (N_12954,N_10562,N_10603);
and U12955 (N_12955,N_10581,N_11742);
xnor U12956 (N_12956,N_10660,N_11709);
and U12957 (N_12957,N_11442,N_11305);
or U12958 (N_12958,N_11047,N_11722);
nand U12959 (N_12959,N_10657,N_11361);
nand U12960 (N_12960,N_11824,N_11120);
nor U12961 (N_12961,N_11020,N_11622);
nor U12962 (N_12962,N_11923,N_10715);
nor U12963 (N_12963,N_10998,N_11205);
nand U12964 (N_12964,N_11994,N_11083);
nor U12965 (N_12965,N_10648,N_10598);
nor U12966 (N_12966,N_11987,N_11747);
and U12967 (N_12967,N_10580,N_11443);
and U12968 (N_12968,N_11203,N_10533);
and U12969 (N_12969,N_11683,N_11048);
and U12970 (N_12970,N_11134,N_11062);
or U12971 (N_12971,N_11375,N_11527);
nand U12972 (N_12972,N_11577,N_10681);
and U12973 (N_12973,N_11625,N_11445);
or U12974 (N_12974,N_11657,N_11028);
nand U12975 (N_12975,N_10620,N_11321);
xor U12976 (N_12976,N_11756,N_10825);
nand U12977 (N_12977,N_11438,N_10700);
and U12978 (N_12978,N_11736,N_11367);
nand U12979 (N_12979,N_11765,N_11767);
xnor U12980 (N_12980,N_11185,N_10771);
or U12981 (N_12981,N_11143,N_11497);
and U12982 (N_12982,N_11443,N_11887);
xnor U12983 (N_12983,N_10932,N_11348);
nand U12984 (N_12984,N_11585,N_11815);
nor U12985 (N_12985,N_10781,N_11612);
nand U12986 (N_12986,N_11434,N_11288);
or U12987 (N_12987,N_11811,N_11416);
xor U12988 (N_12988,N_11822,N_10921);
nor U12989 (N_12989,N_11698,N_11503);
and U12990 (N_12990,N_11514,N_11094);
nor U12991 (N_12991,N_11966,N_11300);
or U12992 (N_12992,N_11291,N_11715);
and U12993 (N_12993,N_11202,N_11981);
xnor U12994 (N_12994,N_11137,N_11763);
nand U12995 (N_12995,N_11068,N_11739);
or U12996 (N_12996,N_10884,N_11687);
nand U12997 (N_12997,N_10849,N_11051);
nor U12998 (N_12998,N_10866,N_10981);
nand U12999 (N_12999,N_11422,N_10908);
and U13000 (N_13000,N_10857,N_11497);
xnor U13001 (N_13001,N_10527,N_10730);
and U13002 (N_13002,N_10904,N_11481);
or U13003 (N_13003,N_11605,N_11237);
nand U13004 (N_13004,N_11194,N_10615);
nor U13005 (N_13005,N_11030,N_10795);
nand U13006 (N_13006,N_11535,N_11540);
and U13007 (N_13007,N_10566,N_11043);
and U13008 (N_13008,N_10947,N_10710);
nor U13009 (N_13009,N_11625,N_10739);
nand U13010 (N_13010,N_10753,N_10731);
and U13011 (N_13011,N_10775,N_11036);
nand U13012 (N_13012,N_11674,N_11652);
xor U13013 (N_13013,N_10530,N_10619);
or U13014 (N_13014,N_10542,N_10971);
nand U13015 (N_13015,N_10852,N_11027);
nor U13016 (N_13016,N_10526,N_11084);
nor U13017 (N_13017,N_10794,N_11474);
nand U13018 (N_13018,N_11207,N_11686);
nand U13019 (N_13019,N_10514,N_10715);
and U13020 (N_13020,N_10950,N_10694);
or U13021 (N_13021,N_10925,N_11848);
and U13022 (N_13022,N_11505,N_10865);
nor U13023 (N_13023,N_11130,N_11073);
and U13024 (N_13024,N_11049,N_10560);
xor U13025 (N_13025,N_10892,N_10904);
nand U13026 (N_13026,N_11142,N_10910);
nand U13027 (N_13027,N_11695,N_10703);
and U13028 (N_13028,N_10637,N_11849);
nor U13029 (N_13029,N_11288,N_10936);
xor U13030 (N_13030,N_11992,N_11467);
nand U13031 (N_13031,N_11679,N_11467);
or U13032 (N_13032,N_10698,N_11386);
nor U13033 (N_13033,N_11017,N_11926);
nand U13034 (N_13034,N_11254,N_11876);
nand U13035 (N_13035,N_10857,N_10927);
or U13036 (N_13036,N_11238,N_11066);
and U13037 (N_13037,N_11055,N_11945);
xor U13038 (N_13038,N_11237,N_11119);
and U13039 (N_13039,N_10964,N_11474);
nor U13040 (N_13040,N_10551,N_10537);
nor U13041 (N_13041,N_11250,N_10976);
nor U13042 (N_13042,N_11307,N_10574);
xor U13043 (N_13043,N_11257,N_11861);
or U13044 (N_13044,N_10636,N_11666);
nand U13045 (N_13045,N_11594,N_11389);
nor U13046 (N_13046,N_11268,N_10633);
xor U13047 (N_13047,N_11725,N_11493);
xor U13048 (N_13048,N_10505,N_11830);
nor U13049 (N_13049,N_11366,N_11061);
and U13050 (N_13050,N_11531,N_10695);
nand U13051 (N_13051,N_11040,N_11212);
nand U13052 (N_13052,N_11585,N_11435);
nor U13053 (N_13053,N_10878,N_11133);
nor U13054 (N_13054,N_11844,N_10547);
xor U13055 (N_13055,N_11849,N_11505);
nor U13056 (N_13056,N_11718,N_10778);
and U13057 (N_13057,N_11668,N_11024);
nor U13058 (N_13058,N_11856,N_11818);
nand U13059 (N_13059,N_11434,N_10626);
nor U13060 (N_13060,N_11327,N_10710);
nand U13061 (N_13061,N_11925,N_10939);
and U13062 (N_13062,N_10945,N_11010);
nand U13063 (N_13063,N_10815,N_11358);
nand U13064 (N_13064,N_11684,N_10833);
nor U13065 (N_13065,N_11663,N_11354);
or U13066 (N_13066,N_10816,N_10834);
and U13067 (N_13067,N_11417,N_11459);
or U13068 (N_13068,N_11051,N_11382);
xor U13069 (N_13069,N_11015,N_11507);
nand U13070 (N_13070,N_11471,N_11216);
nor U13071 (N_13071,N_10625,N_10727);
xnor U13072 (N_13072,N_10880,N_10928);
nand U13073 (N_13073,N_11747,N_11437);
and U13074 (N_13074,N_11365,N_10847);
or U13075 (N_13075,N_11157,N_11036);
nand U13076 (N_13076,N_11513,N_11319);
and U13077 (N_13077,N_10918,N_11887);
nor U13078 (N_13078,N_10971,N_11824);
nand U13079 (N_13079,N_11917,N_11334);
nor U13080 (N_13080,N_11696,N_11273);
nand U13081 (N_13081,N_11625,N_11923);
and U13082 (N_13082,N_11499,N_11406);
or U13083 (N_13083,N_11877,N_10805);
nand U13084 (N_13084,N_10999,N_11049);
nor U13085 (N_13085,N_11271,N_10779);
nand U13086 (N_13086,N_10906,N_11729);
nand U13087 (N_13087,N_11612,N_11330);
nand U13088 (N_13088,N_11962,N_11760);
nor U13089 (N_13089,N_10952,N_11486);
and U13090 (N_13090,N_11123,N_10856);
nand U13091 (N_13091,N_11546,N_11673);
and U13092 (N_13092,N_10803,N_11603);
or U13093 (N_13093,N_11710,N_11592);
and U13094 (N_13094,N_11943,N_11682);
and U13095 (N_13095,N_10656,N_11355);
or U13096 (N_13096,N_10931,N_11591);
nand U13097 (N_13097,N_11562,N_11907);
nor U13098 (N_13098,N_11661,N_11602);
nor U13099 (N_13099,N_10778,N_11826);
nand U13100 (N_13100,N_10811,N_11032);
or U13101 (N_13101,N_10962,N_11268);
nor U13102 (N_13102,N_11943,N_11966);
nor U13103 (N_13103,N_10654,N_11533);
or U13104 (N_13104,N_11779,N_11049);
and U13105 (N_13105,N_11598,N_11192);
and U13106 (N_13106,N_11035,N_11206);
xnor U13107 (N_13107,N_11866,N_10582);
or U13108 (N_13108,N_10980,N_11820);
nand U13109 (N_13109,N_11175,N_10935);
nand U13110 (N_13110,N_10913,N_11042);
nor U13111 (N_13111,N_10681,N_11866);
nand U13112 (N_13112,N_11615,N_10565);
or U13113 (N_13113,N_11180,N_11143);
nor U13114 (N_13114,N_11556,N_10701);
and U13115 (N_13115,N_11780,N_10511);
nor U13116 (N_13116,N_11632,N_11972);
or U13117 (N_13117,N_11542,N_11145);
nand U13118 (N_13118,N_11365,N_11940);
nand U13119 (N_13119,N_11079,N_11781);
nand U13120 (N_13120,N_11751,N_11957);
or U13121 (N_13121,N_10816,N_10792);
nand U13122 (N_13122,N_10967,N_10635);
or U13123 (N_13123,N_11498,N_11202);
nor U13124 (N_13124,N_11149,N_11058);
nor U13125 (N_13125,N_11217,N_11032);
or U13126 (N_13126,N_11326,N_11305);
nand U13127 (N_13127,N_11492,N_11899);
or U13128 (N_13128,N_11459,N_10805);
and U13129 (N_13129,N_10993,N_11149);
nor U13130 (N_13130,N_11965,N_11173);
and U13131 (N_13131,N_11733,N_10525);
or U13132 (N_13132,N_11034,N_11260);
or U13133 (N_13133,N_11385,N_11912);
xor U13134 (N_13134,N_11289,N_10561);
nand U13135 (N_13135,N_10611,N_10771);
nand U13136 (N_13136,N_11581,N_11814);
nor U13137 (N_13137,N_11302,N_11318);
nand U13138 (N_13138,N_11387,N_10625);
nand U13139 (N_13139,N_11425,N_11391);
or U13140 (N_13140,N_11724,N_11639);
nand U13141 (N_13141,N_10948,N_11559);
and U13142 (N_13142,N_10957,N_11414);
nand U13143 (N_13143,N_10879,N_11036);
or U13144 (N_13144,N_11580,N_11974);
nand U13145 (N_13145,N_10513,N_10941);
nor U13146 (N_13146,N_11684,N_11903);
nor U13147 (N_13147,N_11990,N_10892);
and U13148 (N_13148,N_11837,N_11755);
or U13149 (N_13149,N_11450,N_10711);
or U13150 (N_13150,N_11056,N_10548);
nor U13151 (N_13151,N_11572,N_10746);
xor U13152 (N_13152,N_10600,N_11898);
nor U13153 (N_13153,N_11853,N_10882);
or U13154 (N_13154,N_11678,N_11457);
or U13155 (N_13155,N_11477,N_11643);
and U13156 (N_13156,N_11141,N_11701);
xor U13157 (N_13157,N_11758,N_11255);
or U13158 (N_13158,N_11784,N_10575);
or U13159 (N_13159,N_11479,N_11901);
or U13160 (N_13160,N_10745,N_11617);
nor U13161 (N_13161,N_10594,N_11925);
nand U13162 (N_13162,N_10573,N_10993);
or U13163 (N_13163,N_11814,N_10846);
nor U13164 (N_13164,N_11063,N_11130);
and U13165 (N_13165,N_10851,N_11190);
and U13166 (N_13166,N_10776,N_11509);
or U13167 (N_13167,N_11318,N_10713);
or U13168 (N_13168,N_11866,N_11409);
xnor U13169 (N_13169,N_10507,N_11412);
and U13170 (N_13170,N_10744,N_11656);
or U13171 (N_13171,N_10952,N_10949);
xor U13172 (N_13172,N_10740,N_11167);
and U13173 (N_13173,N_11490,N_11966);
and U13174 (N_13174,N_11024,N_10810);
and U13175 (N_13175,N_11088,N_11756);
nor U13176 (N_13176,N_10639,N_11982);
and U13177 (N_13177,N_10665,N_11428);
or U13178 (N_13178,N_11626,N_11947);
nand U13179 (N_13179,N_11757,N_11748);
nand U13180 (N_13180,N_10769,N_10524);
xnor U13181 (N_13181,N_11250,N_11947);
nor U13182 (N_13182,N_10692,N_11922);
nor U13183 (N_13183,N_11544,N_11142);
and U13184 (N_13184,N_11147,N_10740);
and U13185 (N_13185,N_10839,N_10625);
xor U13186 (N_13186,N_11473,N_10565);
and U13187 (N_13187,N_11714,N_11855);
and U13188 (N_13188,N_10727,N_11285);
nor U13189 (N_13189,N_10942,N_10891);
and U13190 (N_13190,N_11155,N_11110);
nor U13191 (N_13191,N_11974,N_11922);
nor U13192 (N_13192,N_10646,N_11336);
xnor U13193 (N_13193,N_11587,N_10932);
nand U13194 (N_13194,N_10899,N_10884);
or U13195 (N_13195,N_11959,N_11567);
or U13196 (N_13196,N_11693,N_10640);
nand U13197 (N_13197,N_10578,N_11515);
and U13198 (N_13198,N_11118,N_11364);
or U13199 (N_13199,N_10809,N_10951);
and U13200 (N_13200,N_11900,N_10993);
xor U13201 (N_13201,N_11793,N_11735);
nand U13202 (N_13202,N_11142,N_10613);
nand U13203 (N_13203,N_11394,N_11564);
nand U13204 (N_13204,N_11162,N_10951);
xor U13205 (N_13205,N_11551,N_10661);
and U13206 (N_13206,N_10673,N_11397);
xor U13207 (N_13207,N_10515,N_10585);
or U13208 (N_13208,N_10971,N_11704);
nor U13209 (N_13209,N_11146,N_10585);
nor U13210 (N_13210,N_10562,N_11197);
nand U13211 (N_13211,N_11180,N_11917);
and U13212 (N_13212,N_11864,N_11083);
or U13213 (N_13213,N_11977,N_11007);
nand U13214 (N_13214,N_11328,N_11087);
xor U13215 (N_13215,N_11856,N_10648);
or U13216 (N_13216,N_11763,N_11397);
nand U13217 (N_13217,N_11113,N_11643);
xor U13218 (N_13218,N_11021,N_10944);
nand U13219 (N_13219,N_11065,N_11935);
or U13220 (N_13220,N_11801,N_11176);
or U13221 (N_13221,N_11482,N_11554);
xnor U13222 (N_13222,N_10836,N_11480);
and U13223 (N_13223,N_10730,N_11551);
nor U13224 (N_13224,N_11834,N_11347);
and U13225 (N_13225,N_11076,N_10912);
or U13226 (N_13226,N_10812,N_11702);
or U13227 (N_13227,N_11221,N_10817);
nor U13228 (N_13228,N_11440,N_11327);
nand U13229 (N_13229,N_11545,N_11735);
nand U13230 (N_13230,N_11449,N_11989);
or U13231 (N_13231,N_10529,N_11068);
and U13232 (N_13232,N_11867,N_11729);
nor U13233 (N_13233,N_11063,N_10964);
or U13234 (N_13234,N_11773,N_11323);
and U13235 (N_13235,N_10793,N_11537);
nand U13236 (N_13236,N_11790,N_11967);
nor U13237 (N_13237,N_10663,N_11144);
or U13238 (N_13238,N_10844,N_11773);
xnor U13239 (N_13239,N_11284,N_11217);
xor U13240 (N_13240,N_11473,N_11174);
nor U13241 (N_13241,N_11951,N_10904);
or U13242 (N_13242,N_10534,N_11821);
or U13243 (N_13243,N_11955,N_11290);
xor U13244 (N_13244,N_11665,N_10553);
or U13245 (N_13245,N_11803,N_11062);
xnor U13246 (N_13246,N_11695,N_11495);
nor U13247 (N_13247,N_11697,N_11641);
xor U13248 (N_13248,N_11557,N_11876);
or U13249 (N_13249,N_11053,N_10739);
or U13250 (N_13250,N_10784,N_10718);
nor U13251 (N_13251,N_11557,N_11643);
nand U13252 (N_13252,N_11679,N_11600);
or U13253 (N_13253,N_10895,N_11258);
nand U13254 (N_13254,N_11163,N_11210);
nand U13255 (N_13255,N_11850,N_11004);
xor U13256 (N_13256,N_11438,N_11058);
and U13257 (N_13257,N_11340,N_10922);
nand U13258 (N_13258,N_11128,N_11816);
nand U13259 (N_13259,N_11242,N_11424);
nor U13260 (N_13260,N_11428,N_10595);
and U13261 (N_13261,N_11187,N_10508);
or U13262 (N_13262,N_11610,N_11246);
or U13263 (N_13263,N_11441,N_11124);
and U13264 (N_13264,N_10559,N_11431);
nand U13265 (N_13265,N_11953,N_11982);
nor U13266 (N_13266,N_11051,N_11247);
and U13267 (N_13267,N_11421,N_10646);
nand U13268 (N_13268,N_11819,N_10712);
nand U13269 (N_13269,N_10604,N_11830);
nand U13270 (N_13270,N_11036,N_10610);
xnor U13271 (N_13271,N_11149,N_10756);
and U13272 (N_13272,N_10991,N_11881);
or U13273 (N_13273,N_11833,N_11553);
nand U13274 (N_13274,N_11445,N_11283);
nor U13275 (N_13275,N_11512,N_10630);
xor U13276 (N_13276,N_10524,N_11944);
or U13277 (N_13277,N_10982,N_11543);
nor U13278 (N_13278,N_11290,N_10902);
and U13279 (N_13279,N_11826,N_10927);
or U13280 (N_13280,N_10882,N_11448);
nand U13281 (N_13281,N_11854,N_11414);
nor U13282 (N_13282,N_10970,N_11997);
nand U13283 (N_13283,N_11488,N_11087);
nand U13284 (N_13284,N_11293,N_11682);
and U13285 (N_13285,N_11212,N_11955);
nand U13286 (N_13286,N_11534,N_11535);
or U13287 (N_13287,N_10953,N_11278);
or U13288 (N_13288,N_11891,N_11598);
or U13289 (N_13289,N_11142,N_11492);
nor U13290 (N_13290,N_11144,N_11087);
nor U13291 (N_13291,N_11494,N_11589);
and U13292 (N_13292,N_11163,N_11825);
nor U13293 (N_13293,N_11365,N_11396);
or U13294 (N_13294,N_11969,N_11823);
nor U13295 (N_13295,N_10979,N_11037);
or U13296 (N_13296,N_10596,N_10551);
and U13297 (N_13297,N_11322,N_11354);
nor U13298 (N_13298,N_10633,N_11639);
or U13299 (N_13299,N_11832,N_11611);
nor U13300 (N_13300,N_10935,N_11364);
nor U13301 (N_13301,N_11575,N_11195);
or U13302 (N_13302,N_10841,N_11149);
nor U13303 (N_13303,N_11301,N_10744);
nor U13304 (N_13304,N_11262,N_10838);
or U13305 (N_13305,N_10635,N_11487);
or U13306 (N_13306,N_11490,N_10721);
xnor U13307 (N_13307,N_10513,N_11823);
nor U13308 (N_13308,N_11128,N_11015);
nor U13309 (N_13309,N_11222,N_10787);
nor U13310 (N_13310,N_11777,N_11928);
nor U13311 (N_13311,N_11716,N_10919);
nor U13312 (N_13312,N_11220,N_10668);
xnor U13313 (N_13313,N_11369,N_11410);
nand U13314 (N_13314,N_11285,N_10693);
nand U13315 (N_13315,N_11256,N_10626);
nor U13316 (N_13316,N_11782,N_11615);
and U13317 (N_13317,N_11436,N_11245);
and U13318 (N_13318,N_11231,N_11597);
nand U13319 (N_13319,N_11176,N_11370);
xnor U13320 (N_13320,N_11804,N_10760);
nand U13321 (N_13321,N_10864,N_11792);
and U13322 (N_13322,N_11548,N_11375);
nand U13323 (N_13323,N_11940,N_10995);
nor U13324 (N_13324,N_11706,N_10951);
or U13325 (N_13325,N_10881,N_11357);
or U13326 (N_13326,N_11538,N_11657);
and U13327 (N_13327,N_11711,N_11463);
nor U13328 (N_13328,N_11392,N_11408);
nor U13329 (N_13329,N_11843,N_11000);
nand U13330 (N_13330,N_11626,N_10803);
or U13331 (N_13331,N_10962,N_11884);
nand U13332 (N_13332,N_11241,N_11316);
nand U13333 (N_13333,N_10734,N_11746);
or U13334 (N_13334,N_10676,N_10753);
xor U13335 (N_13335,N_11550,N_10623);
nand U13336 (N_13336,N_10565,N_11004);
nand U13337 (N_13337,N_11012,N_11768);
nand U13338 (N_13338,N_11469,N_11784);
or U13339 (N_13339,N_11564,N_10583);
or U13340 (N_13340,N_11437,N_11450);
xnor U13341 (N_13341,N_11036,N_11895);
nor U13342 (N_13342,N_11835,N_11210);
nor U13343 (N_13343,N_10884,N_11105);
nand U13344 (N_13344,N_10898,N_11286);
nor U13345 (N_13345,N_11447,N_11497);
and U13346 (N_13346,N_11130,N_11865);
nand U13347 (N_13347,N_11206,N_11768);
or U13348 (N_13348,N_11047,N_10708);
and U13349 (N_13349,N_10838,N_10836);
nor U13350 (N_13350,N_11868,N_11727);
nand U13351 (N_13351,N_11641,N_11300);
nand U13352 (N_13352,N_11087,N_11299);
and U13353 (N_13353,N_10555,N_11347);
and U13354 (N_13354,N_11487,N_11734);
and U13355 (N_13355,N_11802,N_11637);
and U13356 (N_13356,N_11311,N_11873);
nor U13357 (N_13357,N_11174,N_10852);
nor U13358 (N_13358,N_11330,N_11710);
nor U13359 (N_13359,N_11716,N_11101);
and U13360 (N_13360,N_11945,N_11303);
and U13361 (N_13361,N_10911,N_10926);
or U13362 (N_13362,N_10874,N_11107);
and U13363 (N_13363,N_10560,N_10647);
nor U13364 (N_13364,N_11212,N_11487);
nor U13365 (N_13365,N_10860,N_11012);
or U13366 (N_13366,N_11726,N_11735);
nor U13367 (N_13367,N_11830,N_11868);
xor U13368 (N_13368,N_10732,N_10843);
and U13369 (N_13369,N_11093,N_11428);
and U13370 (N_13370,N_11053,N_10610);
nand U13371 (N_13371,N_11736,N_11507);
and U13372 (N_13372,N_10984,N_11085);
and U13373 (N_13373,N_10843,N_11918);
nand U13374 (N_13374,N_10890,N_11238);
and U13375 (N_13375,N_11436,N_11012);
nand U13376 (N_13376,N_10847,N_11568);
nand U13377 (N_13377,N_11371,N_11920);
xnor U13378 (N_13378,N_11760,N_10853);
or U13379 (N_13379,N_11862,N_10696);
and U13380 (N_13380,N_11205,N_11526);
and U13381 (N_13381,N_10831,N_11736);
or U13382 (N_13382,N_10844,N_11031);
or U13383 (N_13383,N_11089,N_10845);
or U13384 (N_13384,N_10821,N_11567);
or U13385 (N_13385,N_11829,N_10960);
nor U13386 (N_13386,N_11148,N_11276);
nor U13387 (N_13387,N_11793,N_11774);
or U13388 (N_13388,N_10577,N_10697);
xnor U13389 (N_13389,N_11135,N_11157);
nor U13390 (N_13390,N_11356,N_11160);
or U13391 (N_13391,N_11029,N_11962);
and U13392 (N_13392,N_11661,N_10954);
nor U13393 (N_13393,N_11414,N_11729);
or U13394 (N_13394,N_10507,N_11798);
or U13395 (N_13395,N_11886,N_11654);
nor U13396 (N_13396,N_11104,N_11931);
nor U13397 (N_13397,N_11320,N_11211);
nand U13398 (N_13398,N_10613,N_11050);
nand U13399 (N_13399,N_11845,N_10789);
nand U13400 (N_13400,N_10715,N_10911);
nor U13401 (N_13401,N_10510,N_11686);
nand U13402 (N_13402,N_10817,N_11109);
and U13403 (N_13403,N_10552,N_11401);
nor U13404 (N_13404,N_10671,N_10664);
nand U13405 (N_13405,N_11844,N_11947);
and U13406 (N_13406,N_10770,N_11540);
or U13407 (N_13407,N_11280,N_10960);
nor U13408 (N_13408,N_11346,N_10651);
and U13409 (N_13409,N_11032,N_11682);
and U13410 (N_13410,N_11638,N_10895);
nand U13411 (N_13411,N_11950,N_11589);
and U13412 (N_13412,N_11109,N_11761);
xor U13413 (N_13413,N_11418,N_11593);
or U13414 (N_13414,N_10737,N_11335);
or U13415 (N_13415,N_11970,N_11122);
and U13416 (N_13416,N_11583,N_11270);
and U13417 (N_13417,N_11964,N_11624);
and U13418 (N_13418,N_11692,N_10976);
nor U13419 (N_13419,N_11558,N_11397);
nand U13420 (N_13420,N_10798,N_11708);
xor U13421 (N_13421,N_11276,N_11540);
nand U13422 (N_13422,N_11893,N_11140);
or U13423 (N_13423,N_11499,N_11236);
and U13424 (N_13424,N_11456,N_11800);
or U13425 (N_13425,N_11413,N_11945);
nand U13426 (N_13426,N_11260,N_10560);
nor U13427 (N_13427,N_11662,N_10800);
and U13428 (N_13428,N_11553,N_10535);
and U13429 (N_13429,N_10557,N_10725);
nor U13430 (N_13430,N_11177,N_11332);
nand U13431 (N_13431,N_10635,N_11812);
and U13432 (N_13432,N_10840,N_10978);
nor U13433 (N_13433,N_10547,N_11806);
nor U13434 (N_13434,N_11300,N_11201);
and U13435 (N_13435,N_10826,N_11854);
or U13436 (N_13436,N_11131,N_11482);
nor U13437 (N_13437,N_11733,N_11132);
nand U13438 (N_13438,N_11121,N_11350);
and U13439 (N_13439,N_11943,N_11766);
and U13440 (N_13440,N_11889,N_10706);
nand U13441 (N_13441,N_11872,N_11107);
nor U13442 (N_13442,N_11369,N_10764);
and U13443 (N_13443,N_11173,N_10738);
or U13444 (N_13444,N_11000,N_11160);
xnor U13445 (N_13445,N_10894,N_11142);
or U13446 (N_13446,N_10679,N_10709);
or U13447 (N_13447,N_11162,N_11686);
nand U13448 (N_13448,N_11806,N_11103);
or U13449 (N_13449,N_10718,N_10833);
nand U13450 (N_13450,N_11553,N_11360);
nand U13451 (N_13451,N_10654,N_11659);
and U13452 (N_13452,N_11987,N_11040);
and U13453 (N_13453,N_11621,N_11541);
or U13454 (N_13454,N_11989,N_10603);
or U13455 (N_13455,N_11499,N_11534);
nand U13456 (N_13456,N_10615,N_11614);
or U13457 (N_13457,N_11312,N_11567);
and U13458 (N_13458,N_11439,N_10941);
or U13459 (N_13459,N_10889,N_11387);
and U13460 (N_13460,N_11973,N_11143);
and U13461 (N_13461,N_10958,N_11249);
or U13462 (N_13462,N_11762,N_11405);
and U13463 (N_13463,N_11979,N_11354);
or U13464 (N_13464,N_11195,N_10884);
nand U13465 (N_13465,N_11536,N_11751);
nor U13466 (N_13466,N_10996,N_11307);
nor U13467 (N_13467,N_10542,N_11148);
nor U13468 (N_13468,N_11429,N_10616);
or U13469 (N_13469,N_11782,N_11365);
nand U13470 (N_13470,N_10984,N_10667);
or U13471 (N_13471,N_11155,N_11623);
and U13472 (N_13472,N_10624,N_11631);
or U13473 (N_13473,N_11270,N_10823);
nor U13474 (N_13474,N_10891,N_11669);
nor U13475 (N_13475,N_11928,N_10566);
xor U13476 (N_13476,N_11253,N_11755);
or U13477 (N_13477,N_10864,N_10504);
and U13478 (N_13478,N_11838,N_11136);
nand U13479 (N_13479,N_11070,N_11858);
or U13480 (N_13480,N_10720,N_11504);
or U13481 (N_13481,N_11539,N_10523);
and U13482 (N_13482,N_11037,N_10921);
nand U13483 (N_13483,N_11336,N_11146);
xnor U13484 (N_13484,N_11402,N_11513);
nand U13485 (N_13485,N_10888,N_11038);
or U13486 (N_13486,N_11825,N_11452);
and U13487 (N_13487,N_11559,N_10551);
nor U13488 (N_13488,N_11328,N_11640);
or U13489 (N_13489,N_11444,N_11514);
and U13490 (N_13490,N_11259,N_10540);
nand U13491 (N_13491,N_11093,N_10727);
xnor U13492 (N_13492,N_11465,N_11112);
nand U13493 (N_13493,N_11196,N_10752);
or U13494 (N_13494,N_11686,N_11620);
nor U13495 (N_13495,N_11060,N_10830);
xor U13496 (N_13496,N_10634,N_10706);
and U13497 (N_13497,N_11847,N_11503);
nor U13498 (N_13498,N_11139,N_11756);
or U13499 (N_13499,N_10509,N_11764);
and U13500 (N_13500,N_12591,N_12589);
nand U13501 (N_13501,N_13075,N_13152);
nor U13502 (N_13502,N_12736,N_13114);
and U13503 (N_13503,N_12770,N_13094);
nand U13504 (N_13504,N_12944,N_12050);
nor U13505 (N_13505,N_12037,N_12728);
xor U13506 (N_13506,N_12376,N_13345);
and U13507 (N_13507,N_13007,N_12653);
nor U13508 (N_13508,N_13387,N_12695);
and U13509 (N_13509,N_13100,N_12140);
or U13510 (N_13510,N_12069,N_13462);
nand U13511 (N_13511,N_12823,N_13312);
and U13512 (N_13512,N_13081,N_12664);
nand U13513 (N_13513,N_12675,N_12532);
nand U13514 (N_13514,N_12021,N_12084);
nand U13515 (N_13515,N_12253,N_12072);
nand U13516 (N_13516,N_12788,N_12649);
xnor U13517 (N_13517,N_12509,N_13493);
nand U13518 (N_13518,N_12264,N_13218);
or U13519 (N_13519,N_13121,N_12075);
nor U13520 (N_13520,N_13402,N_12131);
or U13521 (N_13521,N_13316,N_13353);
and U13522 (N_13522,N_12166,N_12560);
xor U13523 (N_13523,N_12053,N_13141);
and U13524 (N_13524,N_12153,N_13056);
nand U13525 (N_13525,N_12401,N_13236);
or U13526 (N_13526,N_12135,N_12827);
nor U13527 (N_13527,N_13201,N_12546);
nand U13528 (N_13528,N_13290,N_12298);
or U13529 (N_13529,N_12446,N_13054);
nand U13530 (N_13530,N_13012,N_12779);
nand U13531 (N_13531,N_12909,N_12385);
nor U13532 (N_13532,N_12711,N_13017);
nor U13533 (N_13533,N_12801,N_13037);
and U13534 (N_13534,N_13004,N_13317);
or U13535 (N_13535,N_13257,N_12608);
xnor U13536 (N_13536,N_13367,N_12771);
nor U13537 (N_13537,N_13458,N_13372);
nand U13538 (N_13538,N_12793,N_13259);
or U13539 (N_13539,N_12420,N_12899);
nand U13540 (N_13540,N_13178,N_12838);
nor U13541 (N_13541,N_12055,N_12088);
nand U13542 (N_13542,N_12470,N_12937);
and U13543 (N_13543,N_12698,N_12928);
nand U13544 (N_13544,N_12662,N_13237);
xor U13545 (N_13545,N_12670,N_12477);
nor U13546 (N_13546,N_13242,N_12611);
or U13547 (N_13547,N_13092,N_12355);
xnor U13548 (N_13548,N_13277,N_12442);
nor U13549 (N_13549,N_13072,N_13483);
nand U13550 (N_13550,N_13003,N_13404);
xnor U13551 (N_13551,N_12438,N_12757);
or U13552 (N_13552,N_13410,N_13263);
nor U13553 (N_13553,N_12969,N_12331);
nor U13554 (N_13554,N_12782,N_12350);
or U13555 (N_13555,N_13133,N_12354);
nand U13556 (N_13556,N_13479,N_13232);
nor U13557 (N_13557,N_13470,N_12745);
or U13558 (N_13558,N_13348,N_13226);
nor U13559 (N_13559,N_12747,N_13030);
nand U13560 (N_13560,N_13328,N_12179);
nor U13561 (N_13561,N_13352,N_12289);
nand U13562 (N_13562,N_13274,N_13199);
nor U13563 (N_13563,N_12254,N_13040);
nor U13564 (N_13564,N_12461,N_12258);
xnor U13565 (N_13565,N_12555,N_12154);
nand U13566 (N_13566,N_12231,N_12042);
and U13567 (N_13567,N_12839,N_12162);
and U13568 (N_13568,N_12735,N_12222);
nand U13569 (N_13569,N_12357,N_12661);
nand U13570 (N_13570,N_12898,N_12250);
nand U13571 (N_13571,N_12404,N_12007);
nand U13572 (N_13572,N_12144,N_12557);
nor U13573 (N_13573,N_13216,N_12086);
nand U13574 (N_13574,N_13371,N_13467);
nor U13575 (N_13575,N_12766,N_13091);
nand U13576 (N_13576,N_12062,N_13433);
or U13577 (N_13577,N_12709,N_12468);
and U13578 (N_13578,N_12837,N_13489);
nand U13579 (N_13579,N_12332,N_12262);
and U13580 (N_13580,N_12568,N_13424);
nor U13581 (N_13581,N_12267,N_12876);
and U13582 (N_13582,N_12241,N_13456);
nand U13583 (N_13583,N_12505,N_12345);
nand U13584 (N_13584,N_12526,N_12829);
and U13585 (N_13585,N_12469,N_13304);
nor U13586 (N_13586,N_12121,N_13373);
nand U13587 (N_13587,N_12058,N_13022);
xor U13588 (N_13588,N_12979,N_13480);
and U13589 (N_13589,N_13397,N_12986);
or U13590 (N_13590,N_13231,N_13418);
nand U13591 (N_13591,N_12506,N_13109);
and U13592 (N_13592,N_12160,N_12825);
and U13593 (N_13593,N_12377,N_13084);
xor U13594 (N_13594,N_13358,N_12559);
and U13595 (N_13595,N_12847,N_13378);
and U13596 (N_13596,N_12205,N_12798);
and U13597 (N_13597,N_12739,N_12614);
nand U13598 (N_13598,N_13093,N_12775);
nand U13599 (N_13599,N_12027,N_12636);
and U13600 (N_13600,N_13087,N_12048);
and U13601 (N_13601,N_13491,N_12361);
nand U13602 (N_13602,N_13339,N_12529);
nand U13603 (N_13603,N_12374,N_13130);
xor U13604 (N_13604,N_13222,N_13076);
nand U13605 (N_13605,N_13357,N_12269);
or U13606 (N_13606,N_12044,N_12031);
and U13607 (N_13607,N_12233,N_13207);
nand U13608 (N_13608,N_12105,N_12943);
and U13609 (N_13609,N_13211,N_12811);
and U13610 (N_13610,N_12046,N_12902);
xnor U13611 (N_13611,N_12753,N_12752);
nor U13612 (N_13612,N_12984,N_13015);
nand U13613 (N_13613,N_12921,N_12858);
nor U13614 (N_13614,N_13191,N_12817);
and U13615 (N_13615,N_12276,N_12466);
or U13616 (N_13616,N_12464,N_12625);
nor U13617 (N_13617,N_12449,N_13240);
and U13618 (N_13618,N_12663,N_12497);
or U13619 (N_13619,N_12888,N_12440);
nand U13620 (N_13620,N_12147,N_12132);
nor U13621 (N_13621,N_12606,N_12599);
nor U13622 (N_13622,N_12039,N_12856);
and U13623 (N_13623,N_12704,N_12408);
nor U13624 (N_13624,N_13276,N_13202);
nand U13625 (N_13625,N_12875,N_13171);
and U13626 (N_13626,N_13213,N_12453);
nor U13627 (N_13627,N_12930,N_12809);
and U13628 (N_13628,N_12997,N_12656);
nand U13629 (N_13629,N_12009,N_13282);
nor U13630 (N_13630,N_12304,N_12645);
and U13631 (N_13631,N_12395,N_13436);
or U13632 (N_13632,N_12683,N_13457);
and U13633 (N_13633,N_12761,N_13058);
and U13634 (N_13634,N_12962,N_13374);
nand U13635 (N_13635,N_12203,N_13098);
nor U13636 (N_13636,N_12278,N_12201);
and U13637 (N_13637,N_12508,N_13368);
or U13638 (N_13638,N_12318,N_12637);
nor U13639 (N_13639,N_12422,N_12521);
or U13640 (N_13640,N_12392,N_12286);
nand U13641 (N_13641,N_12441,N_12623);
or U13642 (N_13642,N_12041,N_13338);
nor U13643 (N_13643,N_13495,N_13044);
nand U13644 (N_13644,N_12033,N_13016);
or U13645 (N_13645,N_12128,N_13010);
nor U13646 (N_13646,N_12814,N_12681);
or U13647 (N_13647,N_12896,N_13468);
nand U13648 (N_13648,N_13145,N_12587);
and U13649 (N_13649,N_12878,N_13175);
nor U13650 (N_13650,N_12467,N_13041);
and U13651 (N_13651,N_13370,N_13297);
xor U13652 (N_13652,N_12202,N_12139);
or U13653 (N_13653,N_12530,N_13448);
nor U13654 (N_13654,N_12429,N_12200);
nor U13655 (N_13655,N_13050,N_12189);
nand U13656 (N_13656,N_12904,N_12717);
or U13657 (N_13657,N_12789,N_13454);
nand U13658 (N_13658,N_12305,N_13005);
nand U13659 (N_13659,N_12593,N_12538);
and U13660 (N_13660,N_12638,N_12475);
nand U13661 (N_13661,N_13413,N_12018);
nor U13662 (N_13662,N_13067,N_12812);
nor U13663 (N_13663,N_12598,N_12540);
nor U13664 (N_13664,N_12684,N_12686);
and U13665 (N_13665,N_13105,N_12485);
or U13666 (N_13666,N_12976,N_13026);
nor U13667 (N_13667,N_13278,N_12874);
nand U13668 (N_13668,N_13013,N_12352);
nor U13669 (N_13669,N_12666,N_13296);
and U13670 (N_13670,N_12630,N_12524);
or U13671 (N_13671,N_13382,N_12767);
or U13672 (N_13672,N_12407,N_12006);
nand U13673 (N_13673,N_13332,N_13138);
nand U13674 (N_13674,N_13329,N_12690);
nor U13675 (N_13675,N_12556,N_12870);
and U13676 (N_13676,N_12426,N_12585);
nand U13677 (N_13677,N_12841,N_13180);
and U13678 (N_13678,N_12784,N_13172);
nor U13679 (N_13679,N_12078,N_12119);
nor U13680 (N_13680,N_12196,N_12403);
or U13681 (N_13681,N_12609,N_12057);
nand U13682 (N_13682,N_12191,N_12641);
or U13683 (N_13683,N_12565,N_12881);
nor U13684 (N_13684,N_13399,N_13002);
nor U13685 (N_13685,N_12954,N_12073);
or U13686 (N_13686,N_12941,N_13389);
and U13687 (N_13687,N_12145,N_13181);
nor U13688 (N_13688,N_12503,N_12300);
nor U13689 (N_13689,N_12288,N_12938);
nand U13690 (N_13690,N_12873,N_12601);
nor U13691 (N_13691,N_12240,N_12038);
or U13692 (N_13692,N_12400,N_12834);
and U13693 (N_13693,N_13187,N_13273);
nand U13694 (N_13694,N_13365,N_12756);
and U13695 (N_13695,N_12992,N_12014);
xnor U13696 (N_13696,N_13082,N_12257);
and U13697 (N_13697,N_12256,N_13465);
xor U13698 (N_13698,N_12894,N_13193);
and U13699 (N_13699,N_12916,N_12184);
nand U13700 (N_13700,N_12323,N_13243);
and U13701 (N_13701,N_12799,N_12434);
xor U13702 (N_13702,N_12292,N_13225);
xor U13703 (N_13703,N_12547,N_12927);
nor U13704 (N_13704,N_12171,N_12488);
and U13705 (N_13705,N_12622,N_13043);
nand U13706 (N_13706,N_12772,N_12708);
or U13707 (N_13707,N_12730,N_12134);
or U13708 (N_13708,N_12012,N_12610);
or U13709 (N_13709,N_12691,N_13061);
nor U13710 (N_13710,N_12657,N_12685);
xnor U13711 (N_13711,N_12741,N_12965);
nor U13712 (N_13712,N_12866,N_12225);
or U13713 (N_13713,N_12764,N_12915);
and U13714 (N_13714,N_12689,N_13059);
or U13715 (N_13715,N_13233,N_13071);
nand U13716 (N_13716,N_12310,N_12268);
nand U13717 (N_13717,N_12650,N_12312);
nor U13718 (N_13718,N_12060,N_12759);
and U13719 (N_13719,N_12848,N_12076);
nor U13720 (N_13720,N_12971,N_12541);
nand U13721 (N_13721,N_13350,N_13264);
nor U13722 (N_13722,N_12877,N_12341);
nand U13723 (N_13723,N_13272,N_13356);
and U13724 (N_13724,N_13239,N_13147);
nand U13725 (N_13725,N_13112,N_12390);
and U13726 (N_13726,N_13011,N_12970);
or U13727 (N_13727,N_12066,N_12074);
nand U13728 (N_13728,N_12324,N_12972);
nor U13729 (N_13729,N_12826,N_12284);
xnor U13730 (N_13730,N_12148,N_13166);
xnor U13731 (N_13731,N_13205,N_12755);
and U13732 (N_13732,N_13336,N_12835);
nor U13733 (N_13733,N_12845,N_12079);
or U13734 (N_13734,N_13452,N_13461);
and U13735 (N_13735,N_12862,N_13453);
nand U13736 (N_13736,N_12161,N_12627);
or U13737 (N_13737,N_13140,N_12010);
nand U13738 (N_13738,N_12552,N_12581);
and U13739 (N_13739,N_12099,N_13032);
nand U13740 (N_13740,N_13146,N_12431);
and U13741 (N_13741,N_13409,N_13220);
nand U13742 (N_13742,N_12116,N_12476);
xnor U13743 (N_13743,N_12537,N_12337);
or U13744 (N_13744,N_13113,N_12901);
and U13745 (N_13745,N_13354,N_12749);
nor U13746 (N_13746,N_13421,N_13128);
nor U13747 (N_13747,N_12563,N_12209);
and U13748 (N_13748,N_12492,N_12781);
or U13749 (N_13749,N_12214,N_13307);
and U13750 (N_13750,N_13131,N_12586);
nand U13751 (N_13751,N_12785,N_13362);
and U13752 (N_13752,N_12558,N_12696);
or U13753 (N_13753,N_12229,N_12525);
xor U13754 (N_13754,N_12487,N_13322);
nand U13755 (N_13755,N_12989,N_12644);
or U13756 (N_13756,N_13208,N_12141);
nand U13757 (N_13757,N_13115,N_13223);
and U13758 (N_13758,N_12742,N_12237);
nand U13759 (N_13759,N_13301,N_13124);
and U13760 (N_13760,N_12479,N_12564);
or U13761 (N_13761,N_12633,N_12803);
nand U13762 (N_13762,N_13442,N_12607);
xnor U13763 (N_13763,N_12882,N_12891);
and U13764 (N_13764,N_13441,N_13311);
nor U13765 (N_13765,N_12085,N_12910);
nand U13766 (N_13766,N_12528,N_12832);
nor U13767 (N_13767,N_12617,N_12316);
nand U13768 (N_13768,N_12673,N_12999);
nor U13769 (N_13769,N_13288,N_12892);
nor U13770 (N_13770,N_12493,N_12167);
and U13771 (N_13771,N_12271,N_12378);
or U13772 (N_13772,N_13077,N_12418);
nor U13773 (N_13773,N_13349,N_12536);
and U13774 (N_13774,N_12239,N_13034);
and U13775 (N_13775,N_12996,N_13425);
nor U13776 (N_13776,N_12983,N_13283);
nor U13777 (N_13777,N_13401,N_12880);
nor U13778 (N_13778,N_13340,N_13136);
nand U13779 (N_13779,N_13396,N_12389);
nor U13780 (N_13780,N_12707,N_12313);
xor U13781 (N_13781,N_13342,N_12867);
nor U13782 (N_13782,N_13038,N_12406);
and U13783 (N_13783,N_12995,N_13089);
and U13784 (N_13784,N_13066,N_12512);
nand U13785 (N_13785,N_12156,N_12501);
nor U13786 (N_13786,N_12384,N_12919);
or U13787 (N_13787,N_12967,N_12150);
or U13788 (N_13788,N_12631,N_12329);
or U13789 (N_13789,N_12101,N_13334);
nor U13790 (N_13790,N_13251,N_12405);
nor U13791 (N_13791,N_12857,N_13486);
and U13792 (N_13792,N_12399,N_12106);
nand U13793 (N_13793,N_13435,N_12291);
nor U13794 (N_13794,N_13247,N_13057);
and U13795 (N_13795,N_12490,N_12259);
or U13796 (N_13796,N_13069,N_12905);
nor U13797 (N_13797,N_12906,N_12486);
or U13798 (N_13798,N_13381,N_13174);
and U13799 (N_13799,N_12951,N_12806);
xor U13800 (N_13800,N_12594,N_13460);
xor U13801 (N_13801,N_12471,N_12504);
nor U13802 (N_13802,N_13132,N_12173);
nor U13803 (N_13803,N_12227,N_12124);
or U13804 (N_13804,N_13028,N_12914);
nor U13805 (N_13805,N_13169,N_13035);
or U13806 (N_13806,N_12815,N_12566);
and U13807 (N_13807,N_12562,N_13021);
or U13808 (N_13808,N_13118,N_13001);
or U13809 (N_13809,N_13472,N_12480);
nand U13810 (N_13810,N_12948,N_12248);
nor U13811 (N_13811,N_13437,N_12722);
nand U13812 (N_13812,N_12998,N_12713);
nand U13813 (N_13813,N_13229,N_12776);
and U13814 (N_13814,N_13106,N_12281);
nand U13815 (N_13815,N_12172,N_12448);
xor U13816 (N_13816,N_12953,N_12265);
nand U13817 (N_13817,N_12247,N_13320);
nor U13818 (N_13818,N_12249,N_12109);
nand U13819 (N_13819,N_13164,N_13039);
or U13820 (N_13820,N_12977,N_13475);
xor U13821 (N_13821,N_12648,N_13159);
nand U13822 (N_13822,N_12758,N_13499);
and U13823 (N_13823,N_12011,N_12301);
xnor U13824 (N_13824,N_12561,N_13405);
and U13825 (N_13825,N_12430,N_13110);
nand U13826 (N_13826,N_12342,N_12714);
nor U13827 (N_13827,N_12534,N_13268);
or U13828 (N_13828,N_12388,N_13255);
nand U13829 (N_13829,N_12445,N_12181);
and U13830 (N_13830,N_13261,N_12700);
nand U13831 (N_13831,N_12932,N_12296);
nand U13832 (N_13832,N_13170,N_12182);
or U13833 (N_13833,N_13079,N_12804);
or U13834 (N_13834,N_12744,N_12907);
xor U13835 (N_13835,N_12596,N_12942);
nand U13836 (N_13836,N_12208,N_13315);
nor U13837 (N_13837,N_12386,N_12550);
or U13838 (N_13838,N_13244,N_12152);
nor U13839 (N_13839,N_12082,N_12340);
nand U13840 (N_13840,N_12516,N_12917);
or U13841 (N_13841,N_13107,N_12195);
nand U13842 (N_13842,N_12754,N_13139);
xnor U13843 (N_13843,N_12737,N_12863);
nor U13844 (N_13844,N_13376,N_12155);
nand U13845 (N_13845,N_12658,N_13151);
nor U13846 (N_13846,N_13380,N_13434);
nand U13847 (N_13847,N_13427,N_13129);
nand U13848 (N_13848,N_13347,N_12339);
and U13849 (N_13849,N_12308,N_12454);
and U13850 (N_13850,N_13463,N_12865);
nand U13851 (N_13851,N_12729,N_12277);
and U13852 (N_13852,N_12008,N_12047);
nand U13853 (N_13853,N_13143,N_13333);
and U13854 (N_13854,N_12647,N_12897);
or U13855 (N_13855,N_12146,N_13033);
nor U13856 (N_13856,N_12213,N_12346);
nor U13857 (N_13857,N_12040,N_12368);
nor U13858 (N_13858,N_13125,N_13149);
or U13859 (N_13859,N_12245,N_12107);
nand U13860 (N_13860,N_12303,N_13269);
nor U13861 (N_13861,N_12026,N_12900);
and U13862 (N_13862,N_12978,N_12723);
nand U13863 (N_13863,N_12787,N_13246);
nand U13864 (N_13864,N_13300,N_12706);
nor U13865 (N_13865,N_12478,N_13490);
nor U13866 (N_13866,N_12242,N_12083);
or U13867 (N_13867,N_12913,N_12760);
xor U13868 (N_13868,N_13428,N_13161);
nand U13869 (N_13869,N_12846,N_13209);
and U13870 (N_13870,N_13024,N_12104);
nand U13871 (N_13871,N_13471,N_12103);
or U13872 (N_13872,N_13275,N_12024);
nand U13873 (N_13873,N_12791,N_12013);
nand U13874 (N_13874,N_12016,N_13250);
or U13875 (N_13875,N_12223,N_13403);
or U13876 (N_13876,N_13398,N_13214);
and U13877 (N_13877,N_12371,N_13422);
nor U13878 (N_13878,N_13327,N_12108);
xor U13879 (N_13879,N_13488,N_12272);
nor U13880 (N_13880,N_13271,N_12718);
or U13881 (N_13881,N_12294,N_13411);
nand U13882 (N_13882,N_12879,N_12703);
nor U13883 (N_13883,N_13451,N_13383);
nand U13884 (N_13884,N_12235,N_13321);
nor U13885 (N_13885,N_13230,N_12660);
xnor U13886 (N_13886,N_12514,N_12260);
and U13887 (N_13887,N_12343,N_12626);
or U13888 (N_13888,N_13198,N_13306);
nor U13889 (N_13889,N_12192,N_12005);
and U13890 (N_13890,N_12003,N_12499);
nand U13891 (N_13891,N_12089,N_12813);
nor U13892 (N_13892,N_12110,N_12618);
xnor U13893 (N_13893,N_13314,N_12251);
nor U13894 (N_13894,N_13265,N_13086);
and U13895 (N_13895,N_13027,N_12774);
nand U13896 (N_13896,N_12212,N_13256);
or U13897 (N_13897,N_12777,N_13310);
or U13898 (N_13898,N_13155,N_13280);
nand U13899 (N_13899,N_12415,N_13364);
and U13900 (N_13900,N_12483,N_12895);
or U13901 (N_13901,N_12705,N_13194);
nand U13902 (N_13902,N_12314,N_13279);
and U13903 (N_13903,N_12176,N_12988);
nor U13904 (N_13904,N_13177,N_13459);
and U13905 (N_13905,N_12436,N_12952);
or U13906 (N_13906,N_12659,N_12669);
and U13907 (N_13907,N_13388,N_12455);
nor U13908 (N_13908,N_12692,N_12411);
or U13909 (N_13909,N_12980,N_12322);
nor U13910 (N_13910,N_13189,N_13386);
nand U13911 (N_13911,N_12890,N_12080);
and U13912 (N_13912,N_13473,N_12973);
nand U13913 (N_13913,N_12679,N_12054);
nand U13914 (N_13914,N_13186,N_13192);
nor U13915 (N_13915,N_12137,N_13184);
and U13916 (N_13916,N_12710,N_12924);
and U13917 (N_13917,N_12765,N_13221);
nor U13918 (N_13918,N_12731,N_12215);
xor U13919 (N_13919,N_13065,N_13391);
and U13920 (N_13920,N_12678,N_13219);
nor U13921 (N_13921,N_12567,N_13469);
or U13922 (N_13922,N_13165,N_12338);
nand U13923 (N_13923,N_12369,N_13379);
xnor U13924 (N_13924,N_12893,N_12359);
nor U13925 (N_13925,N_12790,N_12800);
xor U13926 (N_13926,N_12335,N_12419);
and U13927 (N_13927,N_12396,N_12416);
or U13928 (N_13928,N_13298,N_13062);
nand U13929 (N_13929,N_12373,N_12402);
nand U13930 (N_13930,N_12712,N_12808);
or U13931 (N_13931,N_12883,N_12619);
and U13932 (N_13932,N_12138,N_13200);
nand U13933 (N_13933,N_13481,N_12588);
nand U13934 (N_13934,N_13014,N_12939);
or U13935 (N_13935,N_13484,N_12067);
xor U13936 (N_13936,N_12961,N_12615);
and U13937 (N_13937,N_13366,N_13415);
or U13938 (N_13938,N_12077,N_13009);
nor U13939 (N_13939,N_12802,N_12494);
nor U13940 (N_13940,N_13337,N_12836);
xor U13941 (N_13941,N_13137,N_12945);
and U13942 (N_13942,N_12168,N_12315);
and U13943 (N_13943,N_13235,N_12535);
xor U13944 (N_13944,N_12417,N_12629);
nand U13945 (N_13945,N_13440,N_12348);
nand U13946 (N_13946,N_12719,N_12549);
or U13947 (N_13947,N_12502,N_13053);
nor U13948 (N_13948,N_13390,N_12425);
or U13949 (N_13949,N_12092,N_12960);
nand U13950 (N_13950,N_12035,N_13095);
xor U13951 (N_13951,N_12726,N_12093);
and U13952 (N_13952,N_13070,N_12853);
or U13953 (N_13953,N_12194,N_12363);
and U13954 (N_13954,N_13217,N_12577);
nand U13955 (N_13955,N_12981,N_12274);
nor U13956 (N_13956,N_13210,N_12792);
nand U13957 (N_13957,N_12740,N_12394);
nand U13958 (N_13958,N_12409,N_13190);
or U13959 (N_13959,N_12533,N_13134);
and U13960 (N_13960,N_12634,N_12545);
or U13961 (N_13961,N_12061,N_13258);
nand U13962 (N_13962,N_12868,N_13392);
or U13963 (N_13963,N_12571,N_12570);
nor U13964 (N_13964,N_13309,N_13074);
nor U13965 (N_13965,N_13455,N_12911);
and U13966 (N_13966,N_12190,N_12423);
or U13967 (N_13967,N_12472,N_12025);
xor U13968 (N_13968,N_12398,N_12118);
or U13969 (N_13969,N_13203,N_12720);
nand U13970 (N_13970,N_13295,N_12844);
xnor U13971 (N_13971,N_12531,N_12946);
nor U13972 (N_13972,N_12188,N_12052);
nor U13973 (N_13973,N_12603,N_12743);
nand U13974 (N_13974,N_12697,N_13485);
or U13975 (N_13975,N_13104,N_12850);
nand U13976 (N_13976,N_12127,N_12266);
nor U13977 (N_13977,N_13360,N_12548);
xnor U13978 (N_13978,N_13045,N_12518);
nand U13979 (N_13979,N_13393,N_12095);
and U13980 (N_13980,N_12520,N_12958);
xor U13981 (N_13981,N_13179,N_13308);
nor U13982 (N_13982,N_12206,N_13299);
nor U13983 (N_13983,N_12238,N_13412);
nand U13984 (N_13984,N_13144,N_12087);
nand U13985 (N_13985,N_12451,N_13414);
nand U13986 (N_13986,N_12985,N_12903);
and U13987 (N_13987,N_12498,N_12624);
nand U13988 (N_13988,N_12435,N_12462);
and U13989 (N_13989,N_13182,N_12126);
and U13990 (N_13990,N_12612,N_13088);
and U13991 (N_13991,N_12081,N_12311);
xor U13992 (N_13992,N_12143,N_12828);
nand U13993 (N_13993,N_13023,N_12326);
and U13994 (N_13994,N_13188,N_13051);
or U13995 (N_13995,N_12515,N_12920);
xor U13996 (N_13996,N_12872,N_13423);
nand U13997 (N_13997,N_13083,N_13055);
and U13998 (N_13998,N_12198,N_12680);
xnor U13999 (N_13999,N_12064,N_12360);
nor U14000 (N_14000,N_12218,N_12507);
xnor U14001 (N_14001,N_12115,N_13117);
nor U14002 (N_14002,N_12620,N_12665);
and U14003 (N_14003,N_13343,N_12600);
nand U14004 (N_14004,N_13326,N_13123);
nor U14005 (N_14005,N_13122,N_12869);
or U14006 (N_14006,N_12157,N_12643);
xnor U14007 (N_14007,N_12397,N_13487);
nor U14008 (N_14008,N_12321,N_12187);
and U14009 (N_14009,N_13270,N_12317);
nor U14010 (N_14010,N_12358,N_12063);
and U14011 (N_14011,N_12583,N_12170);
nor U14012 (N_14012,N_12830,N_12849);
nor U14013 (N_14013,N_13443,N_12216);
xor U14014 (N_14014,N_12676,N_13498);
and U14015 (N_14015,N_12575,N_12595);
xor U14016 (N_14016,N_12183,N_13173);
and U14017 (N_14017,N_12030,N_12908);
or U14018 (N_14018,N_13068,N_12651);
nand U14019 (N_14019,N_12750,N_13154);
or U14020 (N_14020,N_12129,N_12519);
and U14021 (N_14021,N_13085,N_13000);
xor U14022 (N_14022,N_12023,N_12275);
nor U14023 (N_14023,N_13325,N_13319);
and U14024 (N_14024,N_12287,N_13416);
or U14025 (N_14025,N_13266,N_12574);
xnor U14026 (N_14026,N_12362,N_12036);
nand U14027 (N_14027,N_12217,N_12458);
or U14028 (N_14028,N_12957,N_12821);
xnor U14029 (N_14029,N_12372,N_12819);
nor U14030 (N_14030,N_13163,N_13431);
and U14031 (N_14031,N_12456,N_13176);
nor U14032 (N_14032,N_12211,N_12632);
and U14033 (N_14033,N_13286,N_13408);
nor U14034 (N_14034,N_12186,N_13432);
or U14035 (N_14035,N_13227,N_12474);
and U14036 (N_14036,N_12097,N_12822);
nor U14037 (N_14037,N_12513,N_12482);
and U14038 (N_14038,N_12319,N_13073);
nor U14039 (N_14039,N_12022,N_12439);
nand U14040 (N_14040,N_13063,N_13096);
xnor U14041 (N_14041,N_12654,N_12029);
nor U14042 (N_14042,N_12860,N_12810);
xnor U14043 (N_14043,N_12232,N_13385);
nor U14044 (N_14044,N_12113,N_12746);
or U14045 (N_14045,N_13291,N_12255);
nand U14046 (N_14046,N_12299,N_12114);
nand U14047 (N_14047,N_12886,N_12783);
and U14048 (N_14048,N_12734,N_13395);
nand U14049 (N_14049,N_13494,N_12721);
xor U14050 (N_14050,N_13020,N_12169);
xor U14051 (N_14051,N_13351,N_13430);
and U14052 (N_14052,N_12762,N_12220);
nor U14053 (N_14053,N_13482,N_12344);
or U14054 (N_14054,N_13445,N_12751);
nor U14055 (N_14055,N_12621,N_13429);
xnor U14056 (N_14056,N_13305,N_13162);
nor U14057 (N_14057,N_12383,N_12929);
and U14058 (N_14058,N_12185,N_12270);
and U14059 (N_14059,N_13284,N_12796);
nor U14060 (N_14060,N_13294,N_12017);
xor U14061 (N_14061,N_12991,N_12120);
and U14062 (N_14062,N_12934,N_13206);
nand U14063 (N_14063,N_13363,N_13245);
nor U14064 (N_14064,N_12032,N_12094);
and U14065 (N_14065,N_12221,N_12333);
and U14066 (N_14066,N_12573,N_12347);
or U14067 (N_14067,N_12059,N_13450);
and U14068 (N_14068,N_12460,N_12261);
nand U14069 (N_14069,N_12602,N_12306);
xor U14070 (N_14070,N_12912,N_12543);
and U14071 (N_14071,N_12780,N_13267);
or U14072 (N_14072,N_13042,N_12786);
or U14073 (N_14073,N_12163,N_12671);
nor U14074 (N_14074,N_12702,N_12956);
nor U14075 (N_14075,N_12457,N_12178);
xnor U14076 (N_14076,N_13111,N_13359);
or U14077 (N_14077,N_12578,N_13406);
nor U14078 (N_14078,N_12635,N_12646);
nand U14079 (N_14079,N_12580,N_12071);
or U14080 (N_14080,N_12100,N_12351);
nor U14081 (N_14081,N_13474,N_12175);
xnor U14082 (N_14082,N_12732,N_12642);
and U14083 (N_14083,N_12197,N_13344);
xnor U14084 (N_14084,N_12413,N_12366);
nand U14085 (N_14085,N_12820,N_12285);
nor U14086 (N_14086,N_13446,N_13419);
nand U14087 (N_14087,N_12283,N_12947);
and U14088 (N_14088,N_13102,N_12993);
and U14089 (N_14089,N_12230,N_12884);
nand U14090 (N_14090,N_12159,N_12051);
or U14091 (N_14091,N_12773,N_12701);
xor U14092 (N_14092,N_12843,N_12738);
and U14093 (N_14093,N_12795,N_12177);
nor U14094 (N_14094,N_13127,N_12336);
and U14095 (N_14095,N_12500,N_12797);
and U14096 (N_14096,N_12699,N_13049);
nand U14097 (N_14097,N_13323,N_12495);
xnor U14098 (N_14098,N_12854,N_12065);
or U14099 (N_14099,N_12667,N_13097);
or U14100 (N_14100,N_12391,N_12356);
and U14101 (N_14101,N_12484,N_12859);
or U14102 (N_14102,N_13253,N_13215);
xnor U14103 (N_14103,N_12925,N_12070);
and U14104 (N_14104,N_13120,N_13148);
or U14105 (N_14105,N_13346,N_12955);
xnor U14106 (N_14106,N_12807,N_12443);
xor U14107 (N_14107,N_12102,N_12375);
or U14108 (N_14108,N_12282,N_13116);
or U14109 (N_14109,N_12174,N_12885);
nor U14110 (N_14110,N_13156,N_13108);
nand U14111 (N_14111,N_12437,N_12694);
nor U14112 (N_14112,N_12043,N_12049);
nand U14113 (N_14113,N_12542,N_12640);
or U14114 (N_14114,N_12004,N_13047);
nand U14115 (N_14115,N_12414,N_12001);
xor U14116 (N_14116,N_13006,N_12523);
or U14117 (N_14117,N_12481,N_12364);
nand U14118 (N_14118,N_12551,N_12450);
or U14119 (N_14119,N_13355,N_12715);
nor U14120 (N_14120,N_12297,N_13289);
nor U14121 (N_14121,N_12940,N_12544);
nand U14122 (N_14122,N_12410,N_12693);
xor U14123 (N_14123,N_13018,N_12327);
xor U14124 (N_14124,N_12778,N_12130);
or U14125 (N_14125,N_12252,N_12123);
and U14126 (N_14126,N_13361,N_12968);
and U14127 (N_14127,N_13318,N_12539);
and U14128 (N_14128,N_12840,N_12056);
nor U14129 (N_14129,N_12725,N_13126);
and U14130 (N_14130,N_12496,N_12511);
or U14131 (N_14131,N_12831,N_12923);
or U14132 (N_14132,N_12463,N_12975);
or U14133 (N_14133,N_13330,N_13407);
nor U14134 (N_14134,N_13099,N_12861);
nor U14135 (N_14135,N_12228,N_13497);
and U14136 (N_14136,N_12922,N_12091);
nand U14137 (N_14137,N_12244,N_12164);
or U14138 (N_14138,N_12987,N_12125);
nor U14139 (N_14139,N_13167,N_12687);
xnor U14140 (N_14140,N_13197,N_13036);
nand U14141 (N_14141,N_12045,N_12672);
and U14142 (N_14142,N_12427,N_13394);
and U14143 (N_14143,N_12180,N_12465);
and U14144 (N_14144,N_13228,N_12432);
nand U14145 (N_14145,N_13029,N_13234);
or U14146 (N_14146,N_13254,N_13052);
xnor U14147 (N_14147,N_13195,N_12768);
nand U14148 (N_14148,N_12887,N_12020);
and U14149 (N_14149,N_12553,N_12605);
xnor U14150 (N_14150,N_12349,N_12489);
or U14151 (N_14151,N_12219,N_13331);
nor U14152 (N_14152,N_12982,N_12290);
or U14153 (N_14153,N_13335,N_12334);
and U14154 (N_14154,N_12851,N_13341);
nor U14155 (N_14155,N_12428,N_12974);
or U14156 (N_14156,N_12616,N_13262);
and U14157 (N_14157,N_12748,N_13400);
nor U14158 (N_14158,N_12864,N_12224);
nor U14159 (N_14159,N_12330,N_13377);
nor U14160 (N_14160,N_13168,N_12949);
nor U14161 (N_14161,N_12933,N_12682);
and U14162 (N_14162,N_13238,N_13153);
and U14163 (N_14163,N_13160,N_12613);
nand U14164 (N_14164,N_12353,N_12424);
and U14165 (N_14165,N_12674,N_13060);
nand U14166 (N_14166,N_12433,N_13449);
or U14167 (N_14167,N_12295,N_13185);
xnor U14168 (N_14168,N_12320,N_12459);
nor U14169 (N_14169,N_12234,N_12510);
and U14170 (N_14170,N_12590,N_12226);
xor U14171 (N_14171,N_13281,N_13426);
nand U14172 (N_14172,N_13438,N_13303);
nor U14173 (N_14173,N_13078,N_13048);
xnor U14174 (N_14174,N_12473,N_12959);
and U14175 (N_14175,N_13183,N_12365);
xnor U14176 (N_14176,N_12133,N_12628);
nand U14177 (N_14177,N_12569,N_13375);
or U14178 (N_14178,N_12019,N_12117);
or U14179 (N_14179,N_12302,N_12028);
nor U14180 (N_14180,N_12572,N_13090);
or U14181 (N_14181,N_12688,N_12279);
nor U14182 (N_14182,N_13031,N_12246);
xor U14183 (N_14183,N_12964,N_13466);
nor U14184 (N_14184,N_13101,N_12149);
and U14185 (N_14185,N_13252,N_12852);
nand U14186 (N_14186,N_13324,N_12136);
nand U14187 (N_14187,N_12210,N_12096);
or U14188 (N_14188,N_13204,N_12412);
nor U14189 (N_14189,N_12652,N_12015);
and U14190 (N_14190,N_12769,N_13196);
and U14191 (N_14191,N_12936,N_12527);
or U14192 (N_14192,N_12733,N_12855);
or U14193 (N_14193,N_12090,N_12990);
nand U14194 (N_14194,N_12452,N_12236);
and U14195 (N_14195,N_12307,N_12491);
xor U14196 (N_14196,N_12668,N_13249);
nor U14197 (N_14197,N_13384,N_12576);
or U14198 (N_14198,N_13224,N_12367);
and U14199 (N_14199,N_12677,N_13212);
nor U14200 (N_14200,N_13287,N_13439);
and U14201 (N_14201,N_12380,N_12963);
and U14202 (N_14202,N_13158,N_12517);
nand U14203 (N_14203,N_12582,N_12716);
nand U14204 (N_14204,N_12918,N_12655);
and U14205 (N_14205,N_12122,N_12387);
nand U14206 (N_14206,N_12328,N_13119);
nor U14207 (N_14207,N_12597,N_12034);
and U14208 (N_14208,N_12098,N_12966);
nand U14209 (N_14209,N_12889,N_13420);
and U14210 (N_14210,N_12263,N_12604);
nor U14211 (N_14211,N_12151,N_13302);
or U14212 (N_14212,N_13492,N_12000);
nor U14213 (N_14213,N_13417,N_12370);
nand U14214 (N_14214,N_12724,N_13241);
xor U14215 (N_14215,N_12931,N_12950);
xor U14216 (N_14216,N_13150,N_13447);
or U14217 (N_14217,N_13313,N_12158);
nand U14218 (N_14218,N_12193,N_12421);
or U14219 (N_14219,N_13135,N_13248);
xnor U14220 (N_14220,N_13476,N_13260);
nand U14221 (N_14221,N_12325,N_13478);
nand U14222 (N_14222,N_13477,N_12871);
nand U14223 (N_14223,N_12805,N_13369);
xnor U14224 (N_14224,N_12816,N_12142);
and U14225 (N_14225,N_13444,N_12447);
and U14226 (N_14226,N_12824,N_12794);
or U14227 (N_14227,N_12727,N_12381);
nor U14228 (N_14228,N_12935,N_13008);
and U14229 (N_14229,N_12584,N_12002);
or U14230 (N_14230,N_12763,N_12379);
and U14231 (N_14231,N_13103,N_12554);
and U14232 (N_14232,N_13019,N_12068);
xor U14233 (N_14233,N_12112,N_12280);
and U14234 (N_14234,N_13025,N_13285);
nand U14235 (N_14235,N_12309,N_13157);
or U14236 (N_14236,N_12818,N_12842);
nor U14237 (N_14237,N_12165,N_12273);
xnor U14238 (N_14238,N_12293,N_13064);
xor U14239 (N_14239,N_13496,N_13080);
and U14240 (N_14240,N_13046,N_12204);
nor U14241 (N_14241,N_12382,N_12393);
or U14242 (N_14242,N_12111,N_12994);
or U14243 (N_14243,N_12207,N_13464);
nor U14244 (N_14244,N_12926,N_12579);
and U14245 (N_14245,N_12199,N_12592);
nor U14246 (N_14246,N_13293,N_12833);
or U14247 (N_14247,N_12444,N_12243);
nor U14248 (N_14248,N_13292,N_13142);
and U14249 (N_14249,N_12639,N_12522);
nor U14250 (N_14250,N_13128,N_12678);
and U14251 (N_14251,N_12406,N_13138);
nand U14252 (N_14252,N_12977,N_12593);
and U14253 (N_14253,N_13029,N_12275);
xnor U14254 (N_14254,N_13089,N_12115);
nor U14255 (N_14255,N_12599,N_12149);
nand U14256 (N_14256,N_13228,N_12489);
and U14257 (N_14257,N_13257,N_12737);
and U14258 (N_14258,N_12184,N_12955);
and U14259 (N_14259,N_12879,N_12267);
or U14260 (N_14260,N_12212,N_12009);
and U14261 (N_14261,N_12570,N_13082);
or U14262 (N_14262,N_13443,N_12011);
or U14263 (N_14263,N_13093,N_12106);
nor U14264 (N_14264,N_12587,N_13313);
nor U14265 (N_14265,N_12935,N_12297);
nand U14266 (N_14266,N_12911,N_13486);
and U14267 (N_14267,N_12399,N_12566);
xnor U14268 (N_14268,N_12981,N_12228);
or U14269 (N_14269,N_12161,N_13217);
or U14270 (N_14270,N_12236,N_12780);
nor U14271 (N_14271,N_12035,N_12079);
nor U14272 (N_14272,N_13140,N_13208);
or U14273 (N_14273,N_12933,N_12937);
or U14274 (N_14274,N_12603,N_12896);
and U14275 (N_14275,N_12957,N_12321);
and U14276 (N_14276,N_12144,N_13256);
or U14277 (N_14277,N_12465,N_12234);
nor U14278 (N_14278,N_13000,N_13163);
nor U14279 (N_14279,N_12738,N_12022);
and U14280 (N_14280,N_12835,N_13492);
and U14281 (N_14281,N_12026,N_13129);
nor U14282 (N_14282,N_12389,N_12084);
nor U14283 (N_14283,N_13277,N_13057);
or U14284 (N_14284,N_12862,N_12321);
and U14285 (N_14285,N_12542,N_12862);
xnor U14286 (N_14286,N_12506,N_12175);
nand U14287 (N_14287,N_12822,N_12342);
or U14288 (N_14288,N_12152,N_13256);
nor U14289 (N_14289,N_12369,N_13306);
nand U14290 (N_14290,N_12060,N_13401);
and U14291 (N_14291,N_12780,N_12782);
nand U14292 (N_14292,N_12795,N_12186);
or U14293 (N_14293,N_12209,N_13003);
and U14294 (N_14294,N_12942,N_12340);
nand U14295 (N_14295,N_13235,N_12991);
and U14296 (N_14296,N_13064,N_12238);
nor U14297 (N_14297,N_13414,N_12768);
nand U14298 (N_14298,N_12934,N_12014);
or U14299 (N_14299,N_12615,N_12231);
nor U14300 (N_14300,N_12899,N_12472);
or U14301 (N_14301,N_13180,N_13115);
nor U14302 (N_14302,N_13059,N_12987);
nor U14303 (N_14303,N_12807,N_13206);
xor U14304 (N_14304,N_13016,N_12362);
nor U14305 (N_14305,N_12537,N_12707);
and U14306 (N_14306,N_12025,N_12665);
nand U14307 (N_14307,N_12431,N_12710);
and U14308 (N_14308,N_13139,N_12452);
and U14309 (N_14309,N_12635,N_12985);
and U14310 (N_14310,N_12536,N_13310);
nor U14311 (N_14311,N_12118,N_12614);
xnor U14312 (N_14312,N_13182,N_12857);
nor U14313 (N_14313,N_13201,N_12907);
and U14314 (N_14314,N_12988,N_12386);
or U14315 (N_14315,N_12094,N_12596);
or U14316 (N_14316,N_12723,N_12886);
nand U14317 (N_14317,N_12484,N_12348);
nand U14318 (N_14318,N_13141,N_13186);
and U14319 (N_14319,N_12644,N_12196);
or U14320 (N_14320,N_12959,N_12603);
and U14321 (N_14321,N_12377,N_12444);
nand U14322 (N_14322,N_12297,N_13458);
nand U14323 (N_14323,N_13389,N_12242);
nand U14324 (N_14324,N_13183,N_12897);
or U14325 (N_14325,N_12269,N_13208);
nor U14326 (N_14326,N_12643,N_12860);
nand U14327 (N_14327,N_12974,N_13182);
xor U14328 (N_14328,N_13418,N_12045);
nand U14329 (N_14329,N_12173,N_13314);
nand U14330 (N_14330,N_12653,N_12335);
xnor U14331 (N_14331,N_13305,N_13026);
or U14332 (N_14332,N_12196,N_12558);
and U14333 (N_14333,N_12348,N_12994);
xnor U14334 (N_14334,N_12356,N_12887);
nand U14335 (N_14335,N_12880,N_12095);
nand U14336 (N_14336,N_12359,N_12955);
and U14337 (N_14337,N_12447,N_13390);
nand U14338 (N_14338,N_12471,N_13474);
and U14339 (N_14339,N_12118,N_12089);
or U14340 (N_14340,N_12886,N_12359);
or U14341 (N_14341,N_12866,N_12746);
nor U14342 (N_14342,N_12640,N_12712);
nor U14343 (N_14343,N_13057,N_12482);
xnor U14344 (N_14344,N_12266,N_12920);
nor U14345 (N_14345,N_12770,N_12649);
nor U14346 (N_14346,N_12679,N_12292);
xnor U14347 (N_14347,N_12265,N_12432);
nor U14348 (N_14348,N_12749,N_12129);
nand U14349 (N_14349,N_12399,N_13138);
nor U14350 (N_14350,N_12532,N_13001);
or U14351 (N_14351,N_12524,N_13351);
or U14352 (N_14352,N_12902,N_12468);
xor U14353 (N_14353,N_13151,N_13493);
nand U14354 (N_14354,N_12601,N_12507);
nand U14355 (N_14355,N_12834,N_12448);
or U14356 (N_14356,N_13342,N_12811);
nor U14357 (N_14357,N_13147,N_13490);
nor U14358 (N_14358,N_12372,N_12412);
or U14359 (N_14359,N_12677,N_12849);
or U14360 (N_14360,N_12488,N_12309);
nand U14361 (N_14361,N_12844,N_13256);
nor U14362 (N_14362,N_12042,N_13098);
and U14363 (N_14363,N_12539,N_13151);
xnor U14364 (N_14364,N_13368,N_12200);
nand U14365 (N_14365,N_12815,N_13430);
and U14366 (N_14366,N_13474,N_12519);
or U14367 (N_14367,N_12849,N_12569);
xnor U14368 (N_14368,N_12453,N_13299);
xor U14369 (N_14369,N_12314,N_12248);
nor U14370 (N_14370,N_12588,N_13267);
nand U14371 (N_14371,N_12078,N_13250);
nor U14372 (N_14372,N_13262,N_12089);
or U14373 (N_14373,N_12866,N_13114);
or U14374 (N_14374,N_13468,N_12085);
nor U14375 (N_14375,N_13420,N_12008);
and U14376 (N_14376,N_13233,N_12600);
or U14377 (N_14377,N_12975,N_12907);
nand U14378 (N_14378,N_12056,N_12260);
nand U14379 (N_14379,N_12267,N_12624);
xor U14380 (N_14380,N_13121,N_12860);
or U14381 (N_14381,N_12039,N_13319);
nor U14382 (N_14382,N_12168,N_13025);
nand U14383 (N_14383,N_12391,N_13106);
or U14384 (N_14384,N_12521,N_12031);
nand U14385 (N_14385,N_12593,N_12539);
or U14386 (N_14386,N_12643,N_13186);
nand U14387 (N_14387,N_12622,N_12265);
or U14388 (N_14388,N_13018,N_12126);
and U14389 (N_14389,N_13111,N_13243);
nand U14390 (N_14390,N_12640,N_12441);
nor U14391 (N_14391,N_12415,N_12044);
nor U14392 (N_14392,N_12163,N_12929);
nor U14393 (N_14393,N_13115,N_12043);
nand U14394 (N_14394,N_12365,N_13376);
nand U14395 (N_14395,N_12474,N_12097);
and U14396 (N_14396,N_13197,N_13072);
xor U14397 (N_14397,N_12923,N_12139);
nor U14398 (N_14398,N_12458,N_12193);
or U14399 (N_14399,N_12496,N_13470);
nand U14400 (N_14400,N_13148,N_12231);
nand U14401 (N_14401,N_13430,N_13170);
nand U14402 (N_14402,N_13454,N_13054);
xnor U14403 (N_14403,N_12890,N_13109);
and U14404 (N_14404,N_13097,N_12415);
nand U14405 (N_14405,N_12121,N_12027);
and U14406 (N_14406,N_13315,N_13198);
nor U14407 (N_14407,N_13432,N_13233);
and U14408 (N_14408,N_12664,N_12304);
and U14409 (N_14409,N_13355,N_12539);
nor U14410 (N_14410,N_13249,N_12984);
and U14411 (N_14411,N_12388,N_12599);
and U14412 (N_14412,N_12859,N_12605);
and U14413 (N_14413,N_12121,N_13335);
nor U14414 (N_14414,N_12657,N_13006);
nand U14415 (N_14415,N_12487,N_12059);
and U14416 (N_14416,N_12946,N_12156);
or U14417 (N_14417,N_12785,N_12754);
nand U14418 (N_14418,N_12533,N_12521);
and U14419 (N_14419,N_12952,N_12049);
or U14420 (N_14420,N_12335,N_13400);
and U14421 (N_14421,N_12603,N_12888);
xor U14422 (N_14422,N_13367,N_12263);
or U14423 (N_14423,N_12821,N_12302);
nand U14424 (N_14424,N_12052,N_13490);
xor U14425 (N_14425,N_13415,N_12900);
nand U14426 (N_14426,N_12026,N_12597);
or U14427 (N_14427,N_12064,N_12658);
and U14428 (N_14428,N_12234,N_13342);
or U14429 (N_14429,N_12180,N_12678);
nand U14430 (N_14430,N_12152,N_12401);
nand U14431 (N_14431,N_13355,N_13430);
xnor U14432 (N_14432,N_12016,N_12456);
nand U14433 (N_14433,N_12947,N_12413);
and U14434 (N_14434,N_13465,N_12838);
and U14435 (N_14435,N_12864,N_12045);
xor U14436 (N_14436,N_13205,N_12792);
nand U14437 (N_14437,N_13387,N_12527);
xnor U14438 (N_14438,N_12870,N_13460);
nor U14439 (N_14439,N_13338,N_12956);
nor U14440 (N_14440,N_12119,N_12144);
nor U14441 (N_14441,N_12300,N_12418);
nor U14442 (N_14442,N_12548,N_12420);
and U14443 (N_14443,N_12544,N_12874);
or U14444 (N_14444,N_12763,N_13391);
and U14445 (N_14445,N_13221,N_12577);
and U14446 (N_14446,N_12051,N_12133);
xor U14447 (N_14447,N_12203,N_12208);
and U14448 (N_14448,N_13248,N_12258);
or U14449 (N_14449,N_13092,N_12619);
xor U14450 (N_14450,N_12900,N_12165);
and U14451 (N_14451,N_12088,N_12887);
nor U14452 (N_14452,N_12173,N_13436);
xor U14453 (N_14453,N_12227,N_12436);
xor U14454 (N_14454,N_13136,N_12010);
nand U14455 (N_14455,N_12326,N_13093);
and U14456 (N_14456,N_13061,N_12851);
nand U14457 (N_14457,N_13185,N_13221);
or U14458 (N_14458,N_12434,N_12531);
or U14459 (N_14459,N_12341,N_13304);
or U14460 (N_14460,N_13242,N_12752);
nor U14461 (N_14461,N_12275,N_12598);
nor U14462 (N_14462,N_12493,N_13170);
nand U14463 (N_14463,N_13377,N_13173);
and U14464 (N_14464,N_12535,N_12260);
nor U14465 (N_14465,N_13492,N_13222);
nor U14466 (N_14466,N_13274,N_12466);
nand U14467 (N_14467,N_12256,N_12871);
or U14468 (N_14468,N_12551,N_12543);
and U14469 (N_14469,N_12736,N_12984);
or U14470 (N_14470,N_13177,N_12551);
xnor U14471 (N_14471,N_13364,N_12012);
or U14472 (N_14472,N_13237,N_12234);
or U14473 (N_14473,N_12527,N_12636);
nor U14474 (N_14474,N_13005,N_12584);
and U14475 (N_14475,N_13065,N_13026);
or U14476 (N_14476,N_12454,N_12477);
nor U14477 (N_14477,N_12073,N_12837);
nor U14478 (N_14478,N_13018,N_13182);
nor U14479 (N_14479,N_12445,N_13356);
or U14480 (N_14480,N_12771,N_12150);
xnor U14481 (N_14481,N_12976,N_12994);
nand U14482 (N_14482,N_12754,N_12649);
nand U14483 (N_14483,N_12973,N_13398);
xnor U14484 (N_14484,N_13259,N_12747);
nand U14485 (N_14485,N_12948,N_12697);
nand U14486 (N_14486,N_13331,N_13247);
and U14487 (N_14487,N_12373,N_12148);
xor U14488 (N_14488,N_12568,N_12732);
or U14489 (N_14489,N_13122,N_12596);
or U14490 (N_14490,N_13239,N_13006);
nand U14491 (N_14491,N_13104,N_12475);
nor U14492 (N_14492,N_12649,N_13248);
nor U14493 (N_14493,N_13113,N_12459);
nor U14494 (N_14494,N_13425,N_12906);
nor U14495 (N_14495,N_13425,N_12617);
nor U14496 (N_14496,N_12228,N_12827);
nand U14497 (N_14497,N_12062,N_13472);
and U14498 (N_14498,N_12095,N_12413);
or U14499 (N_14499,N_12220,N_12717);
or U14500 (N_14500,N_12616,N_12650);
xnor U14501 (N_14501,N_12646,N_13075);
xor U14502 (N_14502,N_12818,N_12123);
or U14503 (N_14503,N_13326,N_13126);
and U14504 (N_14504,N_12410,N_13222);
nand U14505 (N_14505,N_12113,N_12389);
and U14506 (N_14506,N_12631,N_13471);
or U14507 (N_14507,N_12308,N_13372);
or U14508 (N_14508,N_12599,N_12671);
and U14509 (N_14509,N_13352,N_12746);
or U14510 (N_14510,N_12708,N_13281);
nand U14511 (N_14511,N_12640,N_12808);
xor U14512 (N_14512,N_12815,N_12847);
and U14513 (N_14513,N_12381,N_13422);
or U14514 (N_14514,N_12803,N_13163);
nor U14515 (N_14515,N_13324,N_12033);
and U14516 (N_14516,N_12307,N_13162);
or U14517 (N_14517,N_12277,N_12409);
nand U14518 (N_14518,N_12183,N_12961);
nor U14519 (N_14519,N_12034,N_12282);
nand U14520 (N_14520,N_13253,N_12321);
or U14521 (N_14521,N_12386,N_13416);
xnor U14522 (N_14522,N_12453,N_12031);
or U14523 (N_14523,N_13263,N_12592);
xor U14524 (N_14524,N_13399,N_13147);
xor U14525 (N_14525,N_12668,N_12157);
nand U14526 (N_14526,N_12458,N_13370);
and U14527 (N_14527,N_12728,N_12356);
nand U14528 (N_14528,N_12266,N_12008);
or U14529 (N_14529,N_13427,N_12452);
nor U14530 (N_14530,N_12294,N_12730);
and U14531 (N_14531,N_12729,N_12527);
nand U14532 (N_14532,N_12946,N_13135);
nor U14533 (N_14533,N_12294,N_12743);
nor U14534 (N_14534,N_13410,N_12667);
nor U14535 (N_14535,N_12180,N_12076);
and U14536 (N_14536,N_12782,N_12204);
and U14537 (N_14537,N_13128,N_13031);
or U14538 (N_14538,N_12106,N_12491);
nand U14539 (N_14539,N_12287,N_12213);
nor U14540 (N_14540,N_12229,N_13299);
and U14541 (N_14541,N_13479,N_12466);
nand U14542 (N_14542,N_12678,N_12931);
nor U14543 (N_14543,N_12028,N_12452);
and U14544 (N_14544,N_12621,N_13107);
or U14545 (N_14545,N_13458,N_12609);
nand U14546 (N_14546,N_13231,N_12173);
xnor U14547 (N_14547,N_12843,N_13190);
nor U14548 (N_14548,N_12171,N_12057);
nand U14549 (N_14549,N_12686,N_12140);
nor U14550 (N_14550,N_12460,N_13318);
nand U14551 (N_14551,N_13101,N_12422);
or U14552 (N_14552,N_12543,N_13072);
nor U14553 (N_14553,N_12596,N_12340);
nor U14554 (N_14554,N_13061,N_12044);
and U14555 (N_14555,N_12453,N_12778);
or U14556 (N_14556,N_12695,N_12397);
and U14557 (N_14557,N_13473,N_12637);
nor U14558 (N_14558,N_13279,N_13217);
nand U14559 (N_14559,N_12444,N_12981);
nor U14560 (N_14560,N_13458,N_12698);
xnor U14561 (N_14561,N_12847,N_13459);
and U14562 (N_14562,N_12559,N_12027);
and U14563 (N_14563,N_13366,N_12855);
nand U14564 (N_14564,N_12711,N_12845);
nand U14565 (N_14565,N_12429,N_13318);
nand U14566 (N_14566,N_12233,N_13092);
nor U14567 (N_14567,N_13486,N_13266);
or U14568 (N_14568,N_12651,N_12988);
nand U14569 (N_14569,N_12518,N_12445);
nor U14570 (N_14570,N_12362,N_13278);
or U14571 (N_14571,N_12644,N_12075);
or U14572 (N_14572,N_12290,N_12292);
nand U14573 (N_14573,N_12210,N_12078);
nor U14574 (N_14574,N_13271,N_12003);
and U14575 (N_14575,N_12216,N_13400);
and U14576 (N_14576,N_12080,N_12434);
and U14577 (N_14577,N_13435,N_12621);
and U14578 (N_14578,N_12869,N_12764);
nor U14579 (N_14579,N_12114,N_13287);
and U14580 (N_14580,N_12308,N_12775);
and U14581 (N_14581,N_12915,N_12835);
nand U14582 (N_14582,N_12977,N_12745);
nand U14583 (N_14583,N_12413,N_12379);
nor U14584 (N_14584,N_12764,N_13418);
nor U14585 (N_14585,N_12206,N_12120);
nand U14586 (N_14586,N_12419,N_12333);
nand U14587 (N_14587,N_13110,N_12537);
and U14588 (N_14588,N_13240,N_12158);
or U14589 (N_14589,N_13396,N_12116);
nand U14590 (N_14590,N_12247,N_12600);
nor U14591 (N_14591,N_12498,N_12536);
xnor U14592 (N_14592,N_13084,N_12275);
xor U14593 (N_14593,N_12773,N_12153);
or U14594 (N_14594,N_13189,N_13428);
and U14595 (N_14595,N_13040,N_12651);
or U14596 (N_14596,N_12840,N_12741);
nor U14597 (N_14597,N_13362,N_13382);
or U14598 (N_14598,N_13023,N_12353);
and U14599 (N_14599,N_12612,N_12487);
nand U14600 (N_14600,N_12752,N_12171);
and U14601 (N_14601,N_13408,N_12020);
and U14602 (N_14602,N_12064,N_12969);
and U14603 (N_14603,N_12685,N_12811);
nand U14604 (N_14604,N_12020,N_12142);
xor U14605 (N_14605,N_12190,N_12879);
nor U14606 (N_14606,N_13151,N_12237);
or U14607 (N_14607,N_12301,N_12387);
or U14608 (N_14608,N_12704,N_12354);
or U14609 (N_14609,N_13384,N_12551);
nand U14610 (N_14610,N_12621,N_12464);
and U14611 (N_14611,N_12975,N_12785);
or U14612 (N_14612,N_12157,N_12745);
xor U14613 (N_14613,N_12926,N_12551);
nor U14614 (N_14614,N_13374,N_12445);
nor U14615 (N_14615,N_13142,N_12341);
and U14616 (N_14616,N_12844,N_12328);
and U14617 (N_14617,N_12187,N_12312);
nor U14618 (N_14618,N_12130,N_12480);
and U14619 (N_14619,N_13304,N_13298);
nor U14620 (N_14620,N_12594,N_12187);
nand U14621 (N_14621,N_13222,N_13410);
nor U14622 (N_14622,N_13242,N_12077);
or U14623 (N_14623,N_13017,N_13060);
and U14624 (N_14624,N_12651,N_12767);
nor U14625 (N_14625,N_13480,N_13483);
nand U14626 (N_14626,N_12689,N_12211);
or U14627 (N_14627,N_12697,N_13253);
nor U14628 (N_14628,N_12485,N_12429);
xnor U14629 (N_14629,N_13206,N_12688);
xnor U14630 (N_14630,N_12493,N_13084);
nor U14631 (N_14631,N_13486,N_13027);
or U14632 (N_14632,N_13133,N_12695);
and U14633 (N_14633,N_12792,N_12350);
and U14634 (N_14634,N_13458,N_12397);
and U14635 (N_14635,N_12428,N_12363);
xnor U14636 (N_14636,N_13360,N_12966);
and U14637 (N_14637,N_12234,N_12914);
nor U14638 (N_14638,N_12749,N_12198);
nand U14639 (N_14639,N_12780,N_12600);
and U14640 (N_14640,N_12447,N_12401);
nor U14641 (N_14641,N_12581,N_13066);
xnor U14642 (N_14642,N_12119,N_12768);
or U14643 (N_14643,N_13329,N_13010);
or U14644 (N_14644,N_13435,N_12685);
nor U14645 (N_14645,N_12630,N_13072);
nor U14646 (N_14646,N_13346,N_12343);
xor U14647 (N_14647,N_13291,N_12783);
or U14648 (N_14648,N_13039,N_13295);
xor U14649 (N_14649,N_12437,N_12115);
nand U14650 (N_14650,N_12793,N_12282);
or U14651 (N_14651,N_12066,N_13106);
nor U14652 (N_14652,N_13476,N_12017);
nand U14653 (N_14653,N_12626,N_13448);
xnor U14654 (N_14654,N_12298,N_12694);
nor U14655 (N_14655,N_13239,N_13012);
or U14656 (N_14656,N_12978,N_13447);
xnor U14657 (N_14657,N_12901,N_13024);
xnor U14658 (N_14658,N_13260,N_12686);
nand U14659 (N_14659,N_12685,N_12092);
nor U14660 (N_14660,N_13335,N_12764);
nor U14661 (N_14661,N_12879,N_12915);
and U14662 (N_14662,N_12258,N_12984);
or U14663 (N_14663,N_12680,N_12556);
nor U14664 (N_14664,N_12527,N_12824);
nand U14665 (N_14665,N_12358,N_12761);
and U14666 (N_14666,N_13300,N_12124);
nor U14667 (N_14667,N_12483,N_13058);
nand U14668 (N_14668,N_12834,N_12805);
and U14669 (N_14669,N_12864,N_12445);
nor U14670 (N_14670,N_12909,N_12048);
nor U14671 (N_14671,N_13348,N_13046);
or U14672 (N_14672,N_12926,N_13196);
xnor U14673 (N_14673,N_12708,N_13168);
nor U14674 (N_14674,N_13294,N_12987);
or U14675 (N_14675,N_12431,N_12060);
and U14676 (N_14676,N_12972,N_12894);
nand U14677 (N_14677,N_13483,N_12265);
and U14678 (N_14678,N_12538,N_13151);
or U14679 (N_14679,N_13272,N_13126);
nand U14680 (N_14680,N_12239,N_12053);
or U14681 (N_14681,N_13031,N_12616);
nand U14682 (N_14682,N_12171,N_12071);
nor U14683 (N_14683,N_12315,N_12870);
and U14684 (N_14684,N_12975,N_12281);
nor U14685 (N_14685,N_13008,N_12496);
or U14686 (N_14686,N_12082,N_12554);
nand U14687 (N_14687,N_12685,N_12181);
xnor U14688 (N_14688,N_12579,N_12769);
or U14689 (N_14689,N_12460,N_12912);
or U14690 (N_14690,N_13372,N_13090);
nor U14691 (N_14691,N_12898,N_12281);
nand U14692 (N_14692,N_12671,N_12921);
or U14693 (N_14693,N_12536,N_12665);
and U14694 (N_14694,N_12571,N_12763);
nand U14695 (N_14695,N_13401,N_13022);
or U14696 (N_14696,N_12977,N_12317);
nand U14697 (N_14697,N_13257,N_12653);
and U14698 (N_14698,N_12906,N_12382);
nor U14699 (N_14699,N_12106,N_12149);
or U14700 (N_14700,N_12504,N_12814);
nand U14701 (N_14701,N_12443,N_12098);
and U14702 (N_14702,N_12953,N_12003);
nor U14703 (N_14703,N_12197,N_13398);
nand U14704 (N_14704,N_13244,N_13258);
nand U14705 (N_14705,N_13103,N_13141);
nand U14706 (N_14706,N_13404,N_13295);
nor U14707 (N_14707,N_12250,N_12023);
nor U14708 (N_14708,N_12854,N_12873);
and U14709 (N_14709,N_12715,N_12060);
nor U14710 (N_14710,N_12142,N_12428);
nand U14711 (N_14711,N_12566,N_12809);
nand U14712 (N_14712,N_12441,N_12134);
or U14713 (N_14713,N_12103,N_12940);
and U14714 (N_14714,N_13240,N_13118);
xnor U14715 (N_14715,N_13193,N_12814);
or U14716 (N_14716,N_13209,N_13138);
and U14717 (N_14717,N_12467,N_13414);
nand U14718 (N_14718,N_12113,N_12392);
nand U14719 (N_14719,N_12008,N_13345);
or U14720 (N_14720,N_12958,N_13145);
or U14721 (N_14721,N_12421,N_13403);
and U14722 (N_14722,N_12329,N_13376);
nor U14723 (N_14723,N_13018,N_12279);
and U14724 (N_14724,N_12651,N_13258);
nand U14725 (N_14725,N_13498,N_12627);
nand U14726 (N_14726,N_12600,N_13440);
xnor U14727 (N_14727,N_13349,N_12210);
nor U14728 (N_14728,N_13385,N_12448);
and U14729 (N_14729,N_13147,N_12391);
nor U14730 (N_14730,N_13442,N_12472);
nor U14731 (N_14731,N_12988,N_12251);
nor U14732 (N_14732,N_13046,N_13313);
nor U14733 (N_14733,N_12773,N_12053);
nand U14734 (N_14734,N_12943,N_13436);
and U14735 (N_14735,N_12732,N_12219);
and U14736 (N_14736,N_12931,N_12276);
nand U14737 (N_14737,N_12240,N_13308);
and U14738 (N_14738,N_13285,N_12611);
nand U14739 (N_14739,N_12686,N_13210);
or U14740 (N_14740,N_12418,N_12209);
nand U14741 (N_14741,N_12408,N_12139);
nand U14742 (N_14742,N_12194,N_12916);
xnor U14743 (N_14743,N_13036,N_12290);
nand U14744 (N_14744,N_12463,N_12785);
nand U14745 (N_14745,N_13436,N_12839);
nand U14746 (N_14746,N_13476,N_12913);
and U14747 (N_14747,N_12506,N_12518);
xnor U14748 (N_14748,N_12514,N_12714);
or U14749 (N_14749,N_13179,N_12566);
nor U14750 (N_14750,N_12207,N_13111);
or U14751 (N_14751,N_13127,N_12490);
nand U14752 (N_14752,N_12270,N_13071);
nand U14753 (N_14753,N_13336,N_13444);
and U14754 (N_14754,N_13491,N_12992);
and U14755 (N_14755,N_13226,N_12825);
nand U14756 (N_14756,N_12186,N_12984);
nand U14757 (N_14757,N_13479,N_12929);
nand U14758 (N_14758,N_12847,N_12999);
and U14759 (N_14759,N_13372,N_13126);
xor U14760 (N_14760,N_12732,N_13354);
or U14761 (N_14761,N_13129,N_13195);
nor U14762 (N_14762,N_13494,N_12446);
nor U14763 (N_14763,N_12224,N_12388);
and U14764 (N_14764,N_12253,N_12017);
or U14765 (N_14765,N_13252,N_13312);
and U14766 (N_14766,N_13396,N_12955);
nand U14767 (N_14767,N_12040,N_12716);
or U14768 (N_14768,N_12932,N_12818);
and U14769 (N_14769,N_12280,N_12936);
xnor U14770 (N_14770,N_12061,N_12380);
and U14771 (N_14771,N_12426,N_12670);
xnor U14772 (N_14772,N_13063,N_12636);
nand U14773 (N_14773,N_12713,N_13443);
or U14774 (N_14774,N_12924,N_12119);
nand U14775 (N_14775,N_12625,N_12405);
nor U14776 (N_14776,N_12688,N_13216);
xor U14777 (N_14777,N_13313,N_12272);
or U14778 (N_14778,N_12507,N_12809);
or U14779 (N_14779,N_12266,N_12438);
or U14780 (N_14780,N_13052,N_13243);
and U14781 (N_14781,N_12623,N_12978);
or U14782 (N_14782,N_12209,N_13481);
nor U14783 (N_14783,N_12148,N_12529);
nand U14784 (N_14784,N_13438,N_12974);
nor U14785 (N_14785,N_12708,N_13316);
or U14786 (N_14786,N_13323,N_12344);
nand U14787 (N_14787,N_13468,N_12515);
nand U14788 (N_14788,N_13169,N_12437);
nor U14789 (N_14789,N_12767,N_12175);
and U14790 (N_14790,N_12762,N_12548);
or U14791 (N_14791,N_13433,N_12970);
nand U14792 (N_14792,N_12644,N_12338);
or U14793 (N_14793,N_13068,N_12943);
nand U14794 (N_14794,N_13423,N_12588);
and U14795 (N_14795,N_13001,N_12925);
nand U14796 (N_14796,N_12076,N_13085);
or U14797 (N_14797,N_12241,N_13343);
nor U14798 (N_14798,N_12836,N_12235);
nand U14799 (N_14799,N_12928,N_13226);
nor U14800 (N_14800,N_12627,N_12559);
nor U14801 (N_14801,N_12451,N_12763);
nand U14802 (N_14802,N_12642,N_12739);
nand U14803 (N_14803,N_12056,N_12169);
xnor U14804 (N_14804,N_12361,N_12682);
xor U14805 (N_14805,N_13161,N_13072);
or U14806 (N_14806,N_13074,N_12983);
and U14807 (N_14807,N_13490,N_12014);
nor U14808 (N_14808,N_13322,N_12799);
nand U14809 (N_14809,N_12445,N_13422);
and U14810 (N_14810,N_12204,N_12964);
nand U14811 (N_14811,N_13298,N_12322);
xor U14812 (N_14812,N_12081,N_12199);
or U14813 (N_14813,N_12357,N_13423);
nor U14814 (N_14814,N_13049,N_13487);
nand U14815 (N_14815,N_12601,N_13203);
nor U14816 (N_14816,N_13460,N_13182);
nand U14817 (N_14817,N_13071,N_13169);
and U14818 (N_14818,N_12423,N_12273);
or U14819 (N_14819,N_13454,N_12689);
nand U14820 (N_14820,N_12613,N_13269);
nor U14821 (N_14821,N_12773,N_12631);
xor U14822 (N_14822,N_12834,N_13188);
nand U14823 (N_14823,N_12769,N_12587);
nor U14824 (N_14824,N_12588,N_12767);
nor U14825 (N_14825,N_13301,N_12579);
or U14826 (N_14826,N_12185,N_12126);
nand U14827 (N_14827,N_12729,N_13334);
nand U14828 (N_14828,N_12276,N_13166);
nand U14829 (N_14829,N_12204,N_12540);
nor U14830 (N_14830,N_12528,N_12030);
nand U14831 (N_14831,N_12439,N_12940);
xor U14832 (N_14832,N_13469,N_13147);
nand U14833 (N_14833,N_12378,N_12742);
nand U14834 (N_14834,N_12960,N_13428);
nand U14835 (N_14835,N_12433,N_12654);
or U14836 (N_14836,N_12949,N_12280);
nand U14837 (N_14837,N_12781,N_12682);
and U14838 (N_14838,N_12204,N_12226);
xor U14839 (N_14839,N_13428,N_12362);
and U14840 (N_14840,N_13464,N_12603);
xnor U14841 (N_14841,N_12666,N_12243);
nor U14842 (N_14842,N_13289,N_12472);
nand U14843 (N_14843,N_12234,N_12209);
xnor U14844 (N_14844,N_13261,N_13058);
and U14845 (N_14845,N_12842,N_12073);
nor U14846 (N_14846,N_13064,N_12797);
or U14847 (N_14847,N_12215,N_12338);
xnor U14848 (N_14848,N_12467,N_13309);
nor U14849 (N_14849,N_12079,N_12014);
nand U14850 (N_14850,N_12198,N_12216);
xor U14851 (N_14851,N_13036,N_12129);
nor U14852 (N_14852,N_13150,N_12699);
and U14853 (N_14853,N_12956,N_12169);
xnor U14854 (N_14854,N_12987,N_13141);
nand U14855 (N_14855,N_13249,N_13183);
and U14856 (N_14856,N_12452,N_12895);
xnor U14857 (N_14857,N_12823,N_12312);
nor U14858 (N_14858,N_12407,N_12257);
nand U14859 (N_14859,N_12723,N_13091);
or U14860 (N_14860,N_13127,N_12759);
or U14861 (N_14861,N_12172,N_13115);
nand U14862 (N_14862,N_12006,N_12660);
nand U14863 (N_14863,N_13355,N_13387);
nand U14864 (N_14864,N_13363,N_12713);
and U14865 (N_14865,N_12033,N_12123);
or U14866 (N_14866,N_12809,N_12685);
or U14867 (N_14867,N_13315,N_12403);
nor U14868 (N_14868,N_13343,N_13197);
nand U14869 (N_14869,N_12078,N_13455);
and U14870 (N_14870,N_13262,N_13481);
or U14871 (N_14871,N_13479,N_13224);
nor U14872 (N_14872,N_13499,N_12336);
or U14873 (N_14873,N_12914,N_13040);
nor U14874 (N_14874,N_12482,N_13139);
or U14875 (N_14875,N_13025,N_12730);
and U14876 (N_14876,N_12030,N_13199);
or U14877 (N_14877,N_12318,N_13274);
or U14878 (N_14878,N_13096,N_13072);
or U14879 (N_14879,N_12431,N_12169);
or U14880 (N_14880,N_13270,N_13466);
nand U14881 (N_14881,N_12149,N_12417);
or U14882 (N_14882,N_12450,N_12126);
nor U14883 (N_14883,N_12883,N_12227);
nand U14884 (N_14884,N_13362,N_13219);
nor U14885 (N_14885,N_12132,N_13207);
nor U14886 (N_14886,N_12335,N_12205);
or U14887 (N_14887,N_13470,N_12844);
or U14888 (N_14888,N_12430,N_12216);
nor U14889 (N_14889,N_12004,N_13114);
nor U14890 (N_14890,N_12190,N_13272);
or U14891 (N_14891,N_13273,N_13032);
or U14892 (N_14892,N_12822,N_13239);
xnor U14893 (N_14893,N_12370,N_12702);
and U14894 (N_14894,N_12759,N_12521);
nand U14895 (N_14895,N_12626,N_12474);
nor U14896 (N_14896,N_12412,N_13137);
nand U14897 (N_14897,N_13469,N_12191);
nand U14898 (N_14898,N_13457,N_12601);
nand U14899 (N_14899,N_13086,N_12515);
and U14900 (N_14900,N_12490,N_12985);
or U14901 (N_14901,N_12338,N_13210);
nor U14902 (N_14902,N_12710,N_12070);
nand U14903 (N_14903,N_12971,N_12784);
nand U14904 (N_14904,N_13468,N_12280);
nor U14905 (N_14905,N_12537,N_13400);
nor U14906 (N_14906,N_12615,N_12620);
and U14907 (N_14907,N_12096,N_12080);
xnor U14908 (N_14908,N_12150,N_13010);
nand U14909 (N_14909,N_12821,N_12434);
nand U14910 (N_14910,N_12846,N_12563);
or U14911 (N_14911,N_12677,N_13039);
or U14912 (N_14912,N_13382,N_12636);
xor U14913 (N_14913,N_13111,N_13370);
or U14914 (N_14914,N_12560,N_13292);
xnor U14915 (N_14915,N_13023,N_12869);
xor U14916 (N_14916,N_12677,N_12908);
nand U14917 (N_14917,N_13263,N_12921);
nor U14918 (N_14918,N_12949,N_12274);
or U14919 (N_14919,N_13334,N_13131);
nand U14920 (N_14920,N_12534,N_13477);
nand U14921 (N_14921,N_13367,N_12847);
nand U14922 (N_14922,N_12947,N_12313);
nor U14923 (N_14923,N_13307,N_12249);
or U14924 (N_14924,N_12832,N_12789);
and U14925 (N_14925,N_13107,N_12409);
nor U14926 (N_14926,N_13051,N_13385);
or U14927 (N_14927,N_12846,N_12151);
nor U14928 (N_14928,N_12019,N_13067);
xor U14929 (N_14929,N_13265,N_12871);
or U14930 (N_14930,N_12776,N_13358);
or U14931 (N_14931,N_13288,N_13329);
or U14932 (N_14932,N_12364,N_13488);
or U14933 (N_14933,N_12445,N_13451);
and U14934 (N_14934,N_12995,N_12340);
nor U14935 (N_14935,N_13041,N_13382);
nand U14936 (N_14936,N_12317,N_13430);
and U14937 (N_14937,N_12112,N_12171);
nor U14938 (N_14938,N_12646,N_12415);
and U14939 (N_14939,N_12136,N_12869);
and U14940 (N_14940,N_12290,N_12828);
nor U14941 (N_14941,N_12897,N_12353);
and U14942 (N_14942,N_13476,N_12807);
nand U14943 (N_14943,N_12778,N_12309);
and U14944 (N_14944,N_12519,N_13487);
or U14945 (N_14945,N_12124,N_13206);
nand U14946 (N_14946,N_13373,N_12878);
nand U14947 (N_14947,N_12188,N_12673);
or U14948 (N_14948,N_12652,N_13095);
nor U14949 (N_14949,N_13205,N_13376);
and U14950 (N_14950,N_13131,N_12171);
and U14951 (N_14951,N_13445,N_12377);
nor U14952 (N_14952,N_12230,N_12182);
nand U14953 (N_14953,N_12146,N_13286);
nor U14954 (N_14954,N_12741,N_12596);
or U14955 (N_14955,N_12359,N_12075);
and U14956 (N_14956,N_13293,N_13230);
nand U14957 (N_14957,N_12981,N_13074);
or U14958 (N_14958,N_13429,N_12824);
xor U14959 (N_14959,N_12050,N_13164);
nand U14960 (N_14960,N_12767,N_13026);
and U14961 (N_14961,N_12920,N_12763);
nand U14962 (N_14962,N_12482,N_12346);
or U14963 (N_14963,N_12123,N_13485);
or U14964 (N_14964,N_12333,N_13135);
and U14965 (N_14965,N_12128,N_13109);
xor U14966 (N_14966,N_13088,N_12484);
nor U14967 (N_14967,N_13455,N_12420);
nand U14968 (N_14968,N_13215,N_12100);
and U14969 (N_14969,N_12492,N_13407);
or U14970 (N_14970,N_13018,N_12105);
xor U14971 (N_14971,N_12764,N_12007);
and U14972 (N_14972,N_12896,N_12125);
and U14973 (N_14973,N_12040,N_12106);
or U14974 (N_14974,N_12093,N_12360);
xor U14975 (N_14975,N_12839,N_12003);
and U14976 (N_14976,N_12469,N_12671);
and U14977 (N_14977,N_12664,N_12566);
nor U14978 (N_14978,N_12206,N_13427);
nand U14979 (N_14979,N_12555,N_12198);
and U14980 (N_14980,N_12821,N_12829);
or U14981 (N_14981,N_12725,N_12913);
nand U14982 (N_14982,N_12902,N_13496);
nand U14983 (N_14983,N_13404,N_12349);
nor U14984 (N_14984,N_13271,N_12889);
and U14985 (N_14985,N_12861,N_13380);
or U14986 (N_14986,N_12067,N_12041);
nor U14987 (N_14987,N_12417,N_12532);
or U14988 (N_14988,N_13452,N_13038);
or U14989 (N_14989,N_13329,N_13468);
nor U14990 (N_14990,N_12297,N_12416);
and U14991 (N_14991,N_12428,N_12380);
and U14992 (N_14992,N_13048,N_12934);
nand U14993 (N_14993,N_12832,N_12483);
nor U14994 (N_14994,N_12323,N_12622);
nor U14995 (N_14995,N_12454,N_12705);
or U14996 (N_14996,N_13385,N_12111);
or U14997 (N_14997,N_13069,N_12344);
nor U14998 (N_14998,N_13261,N_12075);
nand U14999 (N_14999,N_12749,N_12224);
and UO_0 (O_0,N_13696,N_14401);
nor UO_1 (O_1,N_13766,N_14686);
or UO_2 (O_2,N_14273,N_14144);
xor UO_3 (O_3,N_13582,N_13682);
or UO_4 (O_4,N_14634,N_14675);
nor UO_5 (O_5,N_13756,N_14498);
nand UO_6 (O_6,N_14674,N_14856);
or UO_7 (O_7,N_14578,N_14229);
nor UO_8 (O_8,N_14691,N_14302);
nor UO_9 (O_9,N_14966,N_14372);
nand UO_10 (O_10,N_13914,N_14268);
or UO_11 (O_11,N_14140,N_14960);
nand UO_12 (O_12,N_13524,N_14033);
nor UO_13 (O_13,N_14280,N_14105);
and UO_14 (O_14,N_14985,N_14010);
xor UO_15 (O_15,N_14221,N_14698);
and UO_16 (O_16,N_13509,N_13936);
or UO_17 (O_17,N_14684,N_14837);
nand UO_18 (O_18,N_14619,N_13703);
nor UO_19 (O_19,N_14715,N_14690);
or UO_20 (O_20,N_13721,N_14679);
nand UO_21 (O_21,N_14238,N_14877);
and UO_22 (O_22,N_14834,N_13955);
nand UO_23 (O_23,N_13709,N_14699);
or UO_24 (O_24,N_14972,N_14883);
nand UO_25 (O_25,N_14112,N_13840);
and UO_26 (O_26,N_14599,N_14850);
nand UO_27 (O_27,N_13844,N_14571);
and UO_28 (O_28,N_14831,N_14631);
nand UO_29 (O_29,N_14037,N_14050);
and UO_30 (O_30,N_14941,N_14067);
nand UO_31 (O_31,N_13549,N_14129);
or UO_32 (O_32,N_14641,N_13934);
and UO_33 (O_33,N_14847,N_13853);
or UO_34 (O_34,N_14270,N_14006);
xnor UO_35 (O_35,N_14753,N_14740);
and UO_36 (O_36,N_14255,N_14083);
nor UO_37 (O_37,N_14978,N_14988);
nand UO_38 (O_38,N_14253,N_13856);
nand UO_39 (O_39,N_14477,N_13841);
or UO_40 (O_40,N_14704,N_14009);
or UO_41 (O_41,N_14812,N_13565);
and UO_42 (O_42,N_13802,N_14373);
or UO_43 (O_43,N_14975,N_13546);
xor UO_44 (O_44,N_14165,N_13718);
and UO_45 (O_45,N_14421,N_14882);
nand UO_46 (O_46,N_14977,N_13662);
nand UO_47 (O_47,N_14863,N_13601);
nand UO_48 (O_48,N_14974,N_14888);
and UO_49 (O_49,N_13708,N_14916);
or UO_50 (O_50,N_14569,N_14597);
nand UO_51 (O_51,N_14038,N_14355);
nor UO_52 (O_52,N_14514,N_13882);
and UO_53 (O_53,N_13630,N_13704);
and UO_54 (O_54,N_14091,N_14832);
nor UO_55 (O_55,N_14558,N_14130);
or UO_56 (O_56,N_13566,N_13655);
or UO_57 (O_57,N_14555,N_14608);
nor UO_58 (O_58,N_14466,N_13780);
xnor UO_59 (O_59,N_14456,N_14262);
nand UO_60 (O_60,N_13518,N_14939);
and UO_61 (O_61,N_14470,N_14746);
xnor UO_62 (O_62,N_14322,N_14900);
nor UO_63 (O_63,N_14334,N_13647);
nand UO_64 (O_64,N_14611,N_13644);
and UO_65 (O_65,N_14428,N_14046);
xor UO_66 (O_66,N_13563,N_13595);
or UO_67 (O_67,N_13817,N_13801);
nor UO_68 (O_68,N_14156,N_13998);
nand UO_69 (O_69,N_14486,N_14458);
and UO_70 (O_70,N_14271,N_14598);
nor UO_71 (O_71,N_13541,N_14707);
or UO_72 (O_72,N_13847,N_14892);
or UO_73 (O_73,N_14057,N_14248);
and UO_74 (O_74,N_14749,N_14809);
nand UO_75 (O_75,N_14092,N_14729);
nor UO_76 (O_76,N_13665,N_14683);
or UO_77 (O_77,N_13827,N_14895);
xnor UO_78 (O_78,N_14234,N_14744);
nor UO_79 (O_79,N_13962,N_14907);
nand UO_80 (O_80,N_14543,N_13553);
nand UO_81 (O_81,N_14663,N_14074);
nand UO_82 (O_82,N_14220,N_14371);
xnor UO_83 (O_83,N_14168,N_13559);
and UO_84 (O_84,N_14068,N_13578);
and UO_85 (O_85,N_14993,N_14910);
nand UO_86 (O_86,N_14361,N_14040);
or UO_87 (O_87,N_14306,N_14648);
nor UO_88 (O_88,N_14760,N_13821);
or UO_89 (O_89,N_13651,N_13814);
nor UO_90 (O_90,N_14885,N_13738);
nand UO_91 (O_91,N_13669,N_14471);
nor UO_92 (O_92,N_13577,N_13830);
or UO_93 (O_93,N_14433,N_14169);
xor UO_94 (O_94,N_13616,N_13674);
or UO_95 (O_95,N_14383,N_14246);
nand UO_96 (O_96,N_14504,N_14703);
nor UO_97 (O_97,N_14199,N_14560);
nor UO_98 (O_98,N_14030,N_14182);
and UO_99 (O_99,N_14152,N_13656);
and UO_100 (O_100,N_13520,N_14376);
and UO_101 (O_101,N_14327,N_13728);
nor UO_102 (O_102,N_14184,N_14000);
and UO_103 (O_103,N_14844,N_13660);
nand UO_104 (O_104,N_14084,N_14438);
xor UO_105 (O_105,N_14922,N_14748);
nor UO_106 (O_106,N_14469,N_13504);
or UO_107 (O_107,N_14515,N_14434);
or UO_108 (O_108,N_14319,N_14287);
nor UO_109 (O_109,N_14020,N_14128);
nor UO_110 (O_110,N_14120,N_14418);
nor UO_111 (O_111,N_14100,N_13762);
xnor UO_112 (O_112,N_14940,N_14285);
or UO_113 (O_113,N_13768,N_14846);
nor UO_114 (O_114,N_13554,N_13899);
or UO_115 (O_115,N_14687,N_13938);
or UO_116 (O_116,N_14449,N_14823);
nand UO_117 (O_117,N_14118,N_13981);
nand UO_118 (O_118,N_13940,N_13650);
or UO_119 (O_119,N_14399,N_14995);
nor UO_120 (O_120,N_14138,N_13871);
and UO_121 (O_121,N_14398,N_14170);
or UO_122 (O_122,N_13888,N_14113);
xor UO_123 (O_123,N_13972,N_13673);
nand UO_124 (O_124,N_14713,N_13985);
and UO_125 (O_125,N_13736,N_13956);
or UO_126 (O_126,N_13843,N_13773);
or UO_127 (O_127,N_13706,N_14981);
nor UO_128 (O_128,N_13959,N_14700);
nor UO_129 (O_129,N_14017,N_13711);
nand UO_130 (O_130,N_13842,N_14768);
nor UO_131 (O_131,N_14938,N_13992);
or UO_132 (O_132,N_13685,N_14076);
and UO_133 (O_133,N_13661,N_14624);
and UO_134 (O_134,N_13627,N_13807);
nand UO_135 (O_135,N_14780,N_14147);
xnor UO_136 (O_136,N_13606,N_13621);
nand UO_137 (O_137,N_13838,N_14388);
nand UO_138 (O_138,N_13924,N_14717);
or UO_139 (O_139,N_13548,N_14407);
nand UO_140 (O_140,N_14468,N_14781);
nor UO_141 (O_141,N_14189,N_14123);
and UO_142 (O_142,N_13539,N_14653);
or UO_143 (O_143,N_13832,N_13982);
nor UO_144 (O_144,N_14521,N_14096);
nand UO_145 (O_145,N_14166,N_14720);
and UO_146 (O_146,N_14927,N_14164);
nor UO_147 (O_147,N_14392,N_14216);
or UO_148 (O_148,N_14251,N_14053);
and UO_149 (O_149,N_14175,N_13861);
xor UO_150 (O_150,N_14036,N_13749);
nor UO_151 (O_151,N_14906,N_14437);
or UO_152 (O_152,N_14934,N_13759);
nor UO_153 (O_153,N_14650,N_14816);
and UO_154 (O_154,N_13592,N_13624);
and UO_155 (O_155,N_14902,N_13689);
or UO_156 (O_156,N_14143,N_14158);
or UO_157 (O_157,N_14627,N_14594);
or UO_158 (O_158,N_14602,N_14921);
xor UO_159 (O_159,N_14820,N_13954);
nor UO_160 (O_160,N_14549,N_13907);
and UO_161 (O_161,N_14357,N_14931);
nor UO_162 (O_162,N_14511,N_13866);
nand UO_163 (O_163,N_14080,N_13725);
xor UO_164 (O_164,N_14177,N_14427);
and UO_165 (O_165,N_14461,N_14948);
nor UO_166 (O_166,N_14654,N_14374);
and UO_167 (O_167,N_14580,N_14148);
nand UO_168 (O_168,N_14465,N_13911);
nand UO_169 (O_169,N_14708,N_14971);
nor UO_170 (O_170,N_14440,N_14911);
and UO_171 (O_171,N_14097,N_13737);
nand UO_172 (O_172,N_14423,N_13868);
nand UO_173 (O_173,N_14267,N_13675);
and UO_174 (O_174,N_13776,N_13699);
or UO_175 (O_175,N_14194,N_13839);
nor UO_176 (O_176,N_13625,N_13700);
nor UO_177 (O_177,N_14467,N_13600);
nor UO_178 (O_178,N_14843,N_14070);
nor UO_179 (O_179,N_14394,N_13555);
nand UO_180 (O_180,N_14970,N_14786);
or UO_181 (O_181,N_14642,N_14799);
nor UO_182 (O_182,N_14378,N_14808);
or UO_183 (O_183,N_14716,N_14485);
or UO_184 (O_184,N_14052,N_14114);
and UO_185 (O_185,N_14409,N_14345);
and UO_186 (O_186,N_13785,N_14542);
nand UO_187 (O_187,N_14866,N_14051);
nor UO_188 (O_188,N_14257,N_14730);
nand UO_189 (O_189,N_14884,N_13734);
or UO_190 (O_190,N_14572,N_14904);
or UO_191 (O_191,N_14630,N_14081);
nor UO_192 (O_192,N_13564,N_14575);
and UO_193 (O_193,N_14775,N_13730);
and UO_194 (O_194,N_13623,N_14849);
or UO_195 (O_195,N_13834,N_13926);
nand UO_196 (O_196,N_14665,N_14230);
nand UO_197 (O_197,N_14794,N_14926);
or UO_198 (O_198,N_14079,N_14737);
or UO_199 (O_199,N_13905,N_14860);
or UO_200 (O_200,N_13690,N_13583);
and UO_201 (O_201,N_14875,N_14281);
and UO_202 (O_202,N_13790,N_13750);
or UO_203 (O_203,N_14098,N_13976);
or UO_204 (O_204,N_14620,N_13714);
nor UO_205 (O_205,N_14451,N_14623);
and UO_206 (O_206,N_13800,N_14589);
nand UO_207 (O_207,N_14763,N_14329);
and UO_208 (O_208,N_14499,N_14830);
nor UO_209 (O_209,N_14350,N_14532);
nand UO_210 (O_210,N_13540,N_14154);
nor UO_211 (O_211,N_13603,N_14478);
xnor UO_212 (O_212,N_13501,N_14901);
nand UO_213 (O_213,N_13960,N_14232);
nor UO_214 (O_214,N_14402,N_13598);
xnor UO_215 (O_215,N_14537,N_13778);
and UO_216 (O_216,N_13631,N_13788);
nor UO_217 (O_217,N_13909,N_13671);
or UO_218 (O_218,N_14366,N_13813);
nor UO_219 (O_219,N_14325,N_14864);
or UO_220 (O_220,N_13668,N_14520);
nor UO_221 (O_221,N_13898,N_14672);
nor UO_222 (O_222,N_13724,N_14593);
or UO_223 (O_223,N_13921,N_13617);
or UO_224 (O_224,N_13642,N_13543);
nor UO_225 (O_225,N_13740,N_13816);
and UO_226 (O_226,N_13747,N_14206);
nand UO_227 (O_227,N_14964,N_13993);
nor UO_228 (O_228,N_13729,N_14913);
or UO_229 (O_229,N_14344,N_13772);
xor UO_230 (O_230,N_14807,N_13987);
xor UO_231 (O_231,N_14836,N_14301);
and UO_232 (O_232,N_14303,N_13915);
nor UO_233 (O_233,N_14342,N_14568);
nand UO_234 (O_234,N_13752,N_14377);
and UO_235 (O_235,N_13628,N_14996);
xor UO_236 (O_236,N_13533,N_13530);
or UO_237 (O_237,N_14738,N_13798);
nor UO_238 (O_238,N_14591,N_13535);
nand UO_239 (O_239,N_14969,N_13964);
xor UO_240 (O_240,N_14311,N_13684);
nand UO_241 (O_241,N_14493,N_14497);
and UO_242 (O_242,N_14207,N_14517);
or UO_243 (O_243,N_14029,N_13626);
and UO_244 (O_244,N_13692,N_14370);
and UO_245 (O_245,N_14735,N_14722);
nor UO_246 (O_246,N_14309,N_14436);
and UO_247 (O_247,N_13681,N_13596);
or UO_248 (O_248,N_14805,N_13670);
or UO_249 (O_249,N_14439,N_14828);
or UO_250 (O_250,N_13851,N_14929);
or UO_251 (O_251,N_14474,N_14386);
nand UO_252 (O_252,N_13903,N_14065);
or UO_253 (O_253,N_14610,N_13619);
and UO_254 (O_254,N_14779,N_14064);
and UO_255 (O_255,N_14073,N_13883);
nand UO_256 (O_256,N_14833,N_14857);
or UO_257 (O_257,N_13585,N_13507);
nand UO_258 (O_258,N_14404,N_14173);
nor UO_259 (O_259,N_14039,N_14237);
and UO_260 (O_260,N_14526,N_14576);
nand UO_261 (O_261,N_14317,N_14706);
nor UO_262 (O_262,N_14088,N_13570);
nand UO_263 (O_263,N_14852,N_13679);
nor UO_264 (O_264,N_14546,N_14818);
and UO_265 (O_265,N_13567,N_14601);
and UO_266 (O_266,N_14007,N_14759);
and UO_267 (O_267,N_14106,N_14695);
nor UO_268 (O_268,N_14688,N_14562);
nand UO_269 (O_269,N_14798,N_14227);
nor UO_270 (O_270,N_13867,N_14936);
nor UO_271 (O_271,N_13769,N_13743);
nor UO_272 (O_272,N_14283,N_14349);
or UO_273 (O_273,N_13948,N_13608);
or UO_274 (O_274,N_14797,N_14115);
or UO_275 (O_275,N_14473,N_13855);
and UO_276 (O_276,N_13633,N_13805);
nor UO_277 (O_277,N_13913,N_14489);
xnor UO_278 (O_278,N_13719,N_14644);
xnor UO_279 (O_279,N_14587,N_14914);
nor UO_280 (O_280,N_14258,N_14032);
or UO_281 (O_281,N_14762,N_14297);
nand UO_282 (O_282,N_14200,N_13602);
nor UO_283 (O_283,N_13562,N_14416);
or UO_284 (O_284,N_14890,N_14354);
or UO_285 (O_285,N_14536,N_13968);
or UO_286 (O_286,N_14802,N_14321);
nor UO_287 (O_287,N_14932,N_14647);
nand UO_288 (O_288,N_14307,N_14259);
nand UO_289 (O_289,N_13591,N_14444);
nand UO_290 (O_290,N_13865,N_13939);
and UO_291 (O_291,N_13605,N_14494);
xnor UO_292 (O_292,N_14390,N_14765);
or UO_293 (O_293,N_14887,N_13612);
xor UO_294 (O_294,N_13947,N_14294);
nor UO_295 (O_295,N_13922,N_14353);
nand UO_296 (O_296,N_14968,N_14646);
and UO_297 (O_297,N_14803,N_13536);
nor UO_298 (O_298,N_14111,N_13761);
nand UO_299 (O_299,N_13731,N_14909);
and UO_300 (O_300,N_13765,N_14382);
nor UO_301 (O_301,N_14956,N_13910);
nand UO_302 (O_302,N_14893,N_14450);
nand UO_303 (O_303,N_13908,N_13710);
xnor UO_304 (O_304,N_14413,N_13500);
nand UO_305 (O_305,N_13818,N_13568);
nor UO_306 (O_306,N_13763,N_14275);
nor UO_307 (O_307,N_13950,N_13594);
or UO_308 (O_308,N_14241,N_14157);
nand UO_309 (O_309,N_14905,N_13806);
nor UO_310 (O_310,N_13529,N_13989);
and UO_311 (O_311,N_13957,N_14240);
or UO_312 (O_312,N_14785,N_13923);
or UO_313 (O_313,N_13918,N_14919);
nor UO_314 (O_314,N_14346,N_14894);
or UO_315 (O_315,N_13688,N_13521);
and UO_316 (O_316,N_14718,N_13808);
nand UO_317 (O_317,N_14615,N_14659);
and UO_318 (O_318,N_13809,N_13537);
and UO_319 (O_319,N_14197,N_14314);
nor UO_320 (O_320,N_13774,N_14279);
xnor UO_321 (O_321,N_14223,N_13912);
or UO_322 (O_322,N_14186,N_14595);
nor UO_323 (O_323,N_14481,N_13561);
xor UO_324 (O_324,N_14313,N_14570);
nand UO_325 (O_325,N_14645,N_13760);
or UO_326 (O_326,N_14668,N_14187);
and UO_327 (O_327,N_14245,N_14455);
nor UO_328 (O_328,N_14089,N_14400);
and UO_329 (O_329,N_14935,N_14483);
nor UO_330 (O_330,N_13787,N_14772);
nand UO_331 (O_331,N_13904,N_13837);
nor UO_332 (O_332,N_13797,N_14869);
xor UO_333 (O_333,N_14649,N_14214);
nor UO_334 (O_334,N_13860,N_14202);
and UO_335 (O_335,N_13715,N_14351);
nor UO_336 (O_336,N_13513,N_14358);
xor UO_337 (O_337,N_14621,N_13525);
xnor UO_338 (O_338,N_14278,N_13900);
and UO_339 (O_339,N_13825,N_14132);
or UO_340 (O_340,N_13512,N_14584);
nor UO_341 (O_341,N_14190,N_14639);
xor UO_342 (O_342,N_13686,N_14326);
nand UO_343 (O_343,N_14291,N_14491);
and UO_344 (O_344,N_13781,N_14581);
xor UO_345 (O_345,N_14419,N_13945);
nand UO_346 (O_346,N_14447,N_14626);
or UO_347 (O_347,N_14586,N_14841);
nor UO_348 (O_348,N_14825,N_14651);
and UO_349 (O_349,N_14523,N_14629);
or UO_350 (O_350,N_13735,N_14443);
or UO_351 (O_351,N_14774,N_14918);
xnor UO_352 (O_352,N_14209,N_13589);
or UO_353 (O_353,N_14003,N_14756);
or UO_354 (O_354,N_14728,N_14026);
or UO_355 (O_355,N_14012,N_14806);
xor UO_356 (O_356,N_13978,N_14415);
nor UO_357 (O_357,N_14529,N_14263);
nand UO_358 (O_358,N_14178,N_14035);
nand UO_359 (O_359,N_13753,N_13942);
nor UO_360 (O_360,N_14984,N_14613);
nor UO_361 (O_361,N_14333,N_14561);
nor UO_362 (O_362,N_14340,N_13580);
nor UO_363 (O_363,N_14702,N_13849);
nor UO_364 (O_364,N_13927,N_14947);
or UO_365 (O_365,N_14955,N_13952);
and UO_366 (O_366,N_13744,N_14638);
nor UO_367 (O_367,N_14060,N_14673);
and UO_368 (O_368,N_13872,N_13572);
or UO_369 (O_369,N_14410,N_14146);
and UO_370 (O_370,N_14566,N_13694);
nor UO_371 (O_371,N_13786,N_14607);
or UO_372 (O_372,N_14535,N_14463);
xnor UO_373 (O_373,N_14369,N_14272);
nor UO_374 (O_374,N_14550,N_13599);
xnor UO_375 (O_375,N_14777,N_14133);
nand UO_376 (O_376,N_14235,N_14305);
xor UO_377 (O_377,N_14677,N_13538);
nand UO_378 (O_378,N_14711,N_14195);
and UO_379 (O_379,N_14556,N_14876);
or UO_380 (O_380,N_13820,N_14185);
nand UO_381 (O_381,N_14264,N_14331);
or UO_382 (O_382,N_14403,N_14171);
or UO_383 (O_383,N_13779,N_13733);
or UO_384 (O_384,N_13556,N_14878);
nor UO_385 (O_385,N_14145,N_14490);
or UO_386 (O_386,N_14192,N_13590);
or UO_387 (O_387,N_14530,N_13946);
nor UO_388 (O_388,N_13857,N_14149);
nor UO_389 (O_389,N_14903,N_14509);
and UO_390 (O_390,N_13534,N_14920);
nand UO_391 (O_391,N_14609,N_14819);
xnor UO_392 (O_392,N_14573,N_14590);
or UO_393 (O_393,N_13963,N_13720);
or UO_394 (O_394,N_13526,N_13611);
nor UO_395 (O_395,N_14360,N_14821);
xnor UO_396 (O_396,N_13819,N_14338);
nand UO_397 (O_397,N_14827,N_14337);
and UO_398 (O_398,N_14225,N_14244);
and UO_399 (O_399,N_14767,N_14747);
nand UO_400 (O_400,N_14539,N_14332);
nor UO_401 (O_401,N_14180,N_14845);
or UO_402 (O_402,N_14290,N_14405);
or UO_403 (O_403,N_14506,N_13949);
xnor UO_404 (O_404,N_13510,N_14066);
nor UO_405 (O_405,N_13574,N_13648);
or UO_406 (O_406,N_14525,N_14752);
nor UO_407 (O_407,N_13880,N_14395);
nand UO_408 (O_408,N_13705,N_14151);
and UO_409 (O_409,N_14848,N_14365);
nor UO_410 (O_410,N_14736,N_14320);
nand UO_411 (O_411,N_14953,N_14356);
nand UO_412 (O_412,N_13979,N_14260);
nor UO_413 (O_413,N_14824,N_14082);
or UO_414 (O_414,N_14897,N_14343);
xnor UO_415 (O_415,N_14750,N_14588);
nor UO_416 (O_416,N_14804,N_13875);
nor UO_417 (O_417,N_14480,N_13547);
nor UO_418 (O_418,N_14336,N_14662);
or UO_419 (O_419,N_14276,N_13726);
nor UO_420 (O_420,N_13902,N_14999);
or UO_421 (O_421,N_14505,N_13693);
nand UO_422 (O_422,N_13917,N_14963);
xnor UO_423 (O_423,N_14121,N_14422);
nor UO_424 (O_424,N_14109,N_14381);
nand UO_425 (O_425,N_13852,N_14384);
nor UO_426 (O_426,N_14754,N_14364);
and UO_427 (O_427,N_14072,N_14231);
nor UO_428 (O_428,N_14296,N_14873);
or UO_429 (O_429,N_13944,N_14101);
xor UO_430 (O_430,N_13973,N_13584);
or UO_431 (O_431,N_14766,N_14393);
or UO_432 (O_432,N_13609,N_14513);
nand UO_433 (O_433,N_14379,N_14742);
or UO_434 (O_434,N_13943,N_14842);
nand UO_435 (O_435,N_13919,N_14563);
nor UO_436 (O_436,N_14656,N_14104);
and UO_437 (O_437,N_14965,N_14693);
xor UO_438 (O_438,N_14637,N_14583);
xor UO_439 (O_439,N_13984,N_14254);
nand UO_440 (O_440,N_14475,N_13523);
or UO_441 (O_441,N_14669,N_14817);
or UO_442 (O_442,N_14603,N_14508);
or UO_443 (O_443,N_13892,N_13643);
nor UO_444 (O_444,N_14099,N_14982);
xnor UO_445 (O_445,N_14951,N_13508);
and UO_446 (O_446,N_14219,N_14042);
nand UO_447 (O_447,N_13638,N_14242);
nand UO_448 (O_448,N_14605,N_14274);
nand UO_449 (O_449,N_13845,N_13522);
nand UO_450 (O_450,N_14600,N_14923);
and UO_451 (O_451,N_14269,N_14552);
nand UO_452 (O_452,N_14987,N_14176);
nor UO_453 (O_453,N_13629,N_13712);
nor UO_454 (O_454,N_13732,N_14950);
or UO_455 (O_455,N_14479,N_14359);
and UO_456 (O_456,N_13649,N_14541);
xnor UO_457 (O_457,N_13754,N_14212);
nand UO_458 (O_458,N_14617,N_14862);
or UO_459 (O_459,N_14266,N_14967);
nand UO_460 (O_460,N_14952,N_14424);
nand UO_461 (O_461,N_13824,N_14949);
nor UO_462 (O_462,N_14492,N_13552);
or UO_463 (O_463,N_14660,N_14770);
and UO_464 (O_464,N_14406,N_14090);
nor UO_465 (O_465,N_13727,N_13558);
nand UO_466 (O_466,N_14606,N_14814);
or UO_467 (O_467,N_14874,N_13739);
nand UO_468 (O_468,N_13971,N_14487);
or UO_469 (O_469,N_14701,N_14328);
xor UO_470 (O_470,N_13874,N_14635);
xor UO_471 (O_471,N_14041,N_14915);
and UO_472 (O_472,N_14942,N_14618);
nand UO_473 (O_473,N_13610,N_13767);
nand UO_474 (O_474,N_14252,N_13977);
nor UO_475 (O_475,N_13618,N_14757);
and UO_476 (O_476,N_13697,N_14697);
and UO_477 (O_477,N_14095,N_13931);
nand UO_478 (O_478,N_13983,N_13937);
nor UO_479 (O_479,N_14045,N_14933);
xor UO_480 (O_480,N_14201,N_13879);
nand UO_481 (O_481,N_14516,N_13683);
nor UO_482 (O_482,N_13862,N_14135);
nand UO_483 (O_483,N_14024,N_13966);
nor UO_484 (O_484,N_13550,N_14043);
nand UO_485 (O_485,N_14502,N_13901);
nor UO_486 (O_486,N_13873,N_14891);
or UO_487 (O_487,N_14671,N_13782);
and UO_488 (O_488,N_14063,N_13593);
nand UO_489 (O_489,N_14930,N_14997);
or UO_490 (O_490,N_13634,N_14107);
nand UO_491 (O_491,N_14983,N_14004);
and UO_492 (O_492,N_14181,N_14002);
nand UO_493 (O_493,N_13758,N_14957);
and UO_494 (O_494,N_13723,N_14131);
nor UO_495 (O_495,N_14476,N_14265);
nor UO_496 (O_496,N_14464,N_14822);
xor UO_497 (O_497,N_13799,N_13614);
xor UO_498 (O_498,N_14008,N_13579);
and UO_499 (O_499,N_14791,N_13951);
or UO_500 (O_500,N_13958,N_14636);
nor UO_501 (O_501,N_14658,N_14094);
or UO_502 (O_502,N_14160,N_14183);
nor UO_503 (O_503,N_13869,N_14134);
nor UO_504 (O_504,N_14868,N_14937);
nand UO_505 (O_505,N_14973,N_14155);
nor UO_506 (O_506,N_14292,N_13932);
xor UO_507 (O_507,N_13916,N_14069);
xor UO_508 (O_508,N_13935,N_14655);
xor UO_509 (O_509,N_13505,N_14375);
nor UO_510 (O_510,N_14025,N_14524);
nor UO_511 (O_511,N_14554,N_13557);
and UO_512 (O_512,N_14495,N_14122);
or UO_513 (O_513,N_13795,N_14858);
xnor UO_514 (O_514,N_14034,N_14330);
nand UO_515 (O_515,N_13659,N_13794);
nor UO_516 (O_516,N_14193,N_14719);
or UO_517 (O_517,N_14815,N_14943);
nand UO_518 (O_518,N_13641,N_13953);
or UO_519 (O_519,N_13637,N_14510);
nand UO_520 (O_520,N_14559,N_14908);
or UO_521 (O_521,N_14612,N_14676);
nand UO_522 (O_522,N_13576,N_13986);
or UO_523 (O_523,N_13755,N_13991);
nand UO_524 (O_524,N_13680,N_13859);
nand UO_525 (O_525,N_13974,N_14826);
or UO_526 (O_526,N_13925,N_14783);
nor UO_527 (O_527,N_14103,N_14778);
or UO_528 (O_528,N_14881,N_14564);
and UO_529 (O_529,N_14397,N_13545);
xor UO_530 (O_530,N_13663,N_13995);
and UO_531 (O_531,N_14055,N_14385);
nor UO_532 (O_532,N_14986,N_13695);
nor UO_533 (O_533,N_14776,N_14380);
or UO_534 (O_534,N_13858,N_14712);
and UO_535 (O_535,N_14093,N_14013);
nand UO_536 (O_536,N_14734,N_14445);
nor UO_537 (O_537,N_13928,N_13676);
xnor UO_538 (O_538,N_14462,N_14389);
or UO_539 (O_539,N_14980,N_13897);
or UO_540 (O_540,N_13691,N_14496);
nand UO_541 (O_541,N_13597,N_13775);
or UO_542 (O_542,N_14298,N_13771);
nand UO_543 (O_543,N_13864,N_13996);
nor UO_544 (O_544,N_14622,N_14126);
and UO_545 (O_545,N_14284,N_14429);
nor UO_546 (O_546,N_13742,N_13620);
or UO_547 (O_547,N_13586,N_14457);
nand UO_548 (O_548,N_13503,N_13639);
and UO_549 (O_549,N_13672,N_14861);
or UO_550 (O_550,N_14188,N_13920);
and UO_551 (O_551,N_13894,N_13646);
or UO_552 (O_552,N_13878,N_14512);
nand UO_553 (O_553,N_14835,N_14945);
and UO_554 (O_554,N_14696,N_14153);
xnor UO_555 (O_555,N_14839,N_14579);
xor UO_556 (O_556,N_14482,N_14217);
and UO_557 (O_557,N_13622,N_14640);
xnor UO_558 (O_558,N_14813,N_13516);
and UO_559 (O_559,N_14518,N_13653);
or UO_560 (O_560,N_14218,N_14019);
nor UO_561 (O_561,N_14414,N_13891);
xnor UO_562 (O_562,N_14059,N_14886);
or UO_563 (O_563,N_13890,N_14990);
and UO_564 (O_564,N_13511,N_14247);
or UO_565 (O_565,N_14787,N_14507);
nand UO_566 (O_566,N_13804,N_13929);
nand UO_567 (O_567,N_13887,N_14299);
xor UO_568 (O_568,N_14840,N_13707);
or UO_569 (O_569,N_14664,N_13783);
and UO_570 (O_570,N_14117,N_14871);
nor UO_571 (O_571,N_14723,N_13810);
and UO_572 (O_572,N_13965,N_13573);
nand UO_573 (O_573,N_14522,N_14408);
xor UO_574 (O_574,N_13811,N_14204);
nor UO_575 (O_575,N_13698,N_13635);
and UO_576 (O_576,N_13886,N_14137);
nand UO_577 (O_577,N_13741,N_14989);
or UO_578 (O_578,N_14745,N_13517);
nor UO_579 (O_579,N_14367,N_14547);
nand UO_580 (O_580,N_13652,N_14021);
or UO_581 (O_581,N_13746,N_14396);
or UO_582 (O_582,N_14682,N_13836);
nand UO_583 (O_583,N_14224,N_13613);
nand UO_584 (O_584,N_14454,N_13664);
xor UO_585 (O_585,N_14503,N_14310);
and UO_586 (O_586,N_14233,N_14758);
xnor UO_587 (O_587,N_14442,N_14453);
and UO_588 (O_588,N_14167,N_14896);
and UO_589 (O_589,N_14567,N_14574);
nand UO_590 (O_590,N_14859,N_13969);
or UO_591 (O_591,N_13658,N_14341);
nand UO_592 (O_592,N_14282,N_13975);
and UO_593 (O_593,N_13997,N_13588);
nor UO_594 (O_594,N_13702,N_14743);
nand UO_595 (O_595,N_14533,N_14727);
and UO_596 (O_596,N_13528,N_13777);
or UO_597 (O_597,N_14139,N_14633);
nand UO_598 (O_598,N_14992,N_14110);
nand UO_599 (O_599,N_14300,N_14213);
and UO_600 (O_600,N_14058,N_13826);
nor UO_601 (O_601,N_14604,N_14085);
or UO_602 (O_602,N_13560,N_14174);
and UO_603 (O_603,N_14548,N_14652);
or UO_604 (O_604,N_13716,N_14685);
and UO_605 (O_605,N_14018,N_14016);
and UO_606 (O_606,N_14448,N_14994);
nor UO_607 (O_607,N_14005,N_14557);
nor UO_608 (O_608,N_14838,N_13713);
xor UO_609 (O_609,N_14141,N_14391);
nand UO_610 (O_610,N_14553,N_13994);
or UO_611 (O_611,N_14261,N_13569);
nand UO_612 (O_612,N_13889,N_14771);
and UO_613 (O_613,N_14077,N_14751);
nor UO_614 (O_614,N_14670,N_14725);
nand UO_615 (O_615,N_14432,N_14724);
nor UO_616 (O_616,N_14339,N_14527);
nand UO_617 (O_617,N_14228,N_14540);
nand UO_618 (O_618,N_13657,N_13515);
nand UO_619 (O_619,N_14577,N_13514);
and UO_620 (O_620,N_13575,N_14958);
nor UO_621 (O_621,N_14796,N_14027);
nor UO_622 (O_622,N_14028,N_14198);
and UO_623 (O_623,N_13757,N_13846);
or UO_624 (O_624,N_14425,N_14054);
or UO_625 (O_625,N_13793,N_14801);
nor UO_626 (O_626,N_14222,N_14348);
and UO_627 (O_627,N_14741,N_13863);
nand UO_628 (O_628,N_14739,N_14001);
and UO_629 (O_629,N_14792,N_13701);
and UO_630 (O_630,N_14534,N_13796);
and UO_631 (O_631,N_13615,N_13848);
nand UO_632 (O_632,N_14944,N_14087);
nand UO_633 (O_633,N_14015,N_13967);
nand UO_634 (O_634,N_14721,N_14898);
nor UO_635 (O_635,N_13751,N_14061);
xnor UO_636 (O_636,N_14323,N_13870);
or UO_637 (O_637,N_13893,N_13835);
xnor UO_638 (O_638,N_14071,N_13789);
and UO_639 (O_639,N_13667,N_14048);
nor UO_640 (O_640,N_14011,N_13678);
nor UO_641 (O_641,N_14179,N_13792);
or UO_642 (O_642,N_14312,N_13531);
xor UO_643 (O_643,N_14161,N_14962);
nor UO_644 (O_644,N_13666,N_14899);
or UO_645 (O_645,N_14643,N_14733);
xnor UO_646 (O_646,N_14924,N_14681);
and UO_647 (O_647,N_14710,N_14782);
nand UO_648 (O_648,N_13896,N_13812);
or UO_649 (O_649,N_14979,N_14854);
or UO_650 (O_650,N_14912,N_14142);
nand UO_651 (O_651,N_14308,N_13876);
or UO_652 (O_652,N_14667,N_14800);
and UO_653 (O_653,N_14998,N_14692);
nor UO_654 (O_654,N_14203,N_13988);
nand UO_655 (O_655,N_14755,N_14441);
or UO_656 (O_656,N_14277,N_13506);
or UO_657 (O_657,N_14196,N_13542);
xor UO_658 (O_658,N_13632,N_13748);
or UO_659 (O_659,N_14022,N_14872);
nor UO_660 (O_660,N_14023,N_14324);
nor UO_661 (O_661,N_14208,N_13831);
nand UO_662 (O_662,N_13581,N_14784);
and UO_663 (O_663,N_14236,N_14411);
or UO_664 (O_664,N_14592,N_14865);
nand UO_665 (O_665,N_13815,N_14732);
nor UO_666 (O_666,N_13877,N_13722);
and UO_667 (O_667,N_13551,N_14125);
and UO_668 (O_668,N_14239,N_13527);
nor UO_669 (O_669,N_14709,N_14031);
and UO_670 (O_670,N_14582,N_14347);
or UO_671 (O_671,N_14250,N_14689);
or UO_672 (O_672,N_14431,N_13895);
nand UO_673 (O_673,N_14211,N_14976);
nand UO_674 (O_674,N_14056,N_13640);
and UO_675 (O_675,N_14215,N_13519);
and UO_676 (O_676,N_14769,N_14628);
nor UO_677 (O_677,N_14210,N_14531);
or UO_678 (O_678,N_14426,N_13571);
and UO_679 (O_679,N_14078,N_14538);
nand UO_680 (O_680,N_14044,N_14108);
nor UO_681 (O_681,N_13829,N_14810);
or UO_682 (O_682,N_14764,N_14086);
and UO_683 (O_683,N_14205,N_13532);
nand UO_684 (O_684,N_13884,N_14501);
nor UO_685 (O_685,N_14289,N_14075);
nor UO_686 (O_686,N_13654,N_14295);
xnor UO_687 (O_687,N_14565,N_14127);
nand UO_688 (O_688,N_14119,N_14293);
nor UO_689 (O_689,N_14315,N_14867);
and UO_690 (O_690,N_13999,N_14102);
and UO_691 (O_691,N_13930,N_14335);
nand UO_692 (O_692,N_14773,N_14991);
or UO_693 (O_693,N_14430,N_14853);
and UO_694 (O_694,N_13854,N_13803);
and UO_695 (O_695,N_14925,N_14363);
and UO_696 (O_696,N_14726,N_14666);
nor UO_697 (O_697,N_14116,N_14946);
or UO_698 (O_698,N_14829,N_13823);
nor UO_699 (O_699,N_14452,N_13502);
nor UO_700 (O_700,N_14368,N_14256);
or UO_701 (O_701,N_14544,N_14625);
or UO_702 (O_702,N_14484,N_14678);
or UO_703 (O_703,N_14417,N_14616);
or UO_704 (O_704,N_14163,N_14062);
or UO_705 (O_705,N_14661,N_14446);
and UO_706 (O_706,N_14545,N_14136);
and UO_707 (O_707,N_14889,N_13906);
nor UO_708 (O_708,N_13636,N_14049);
xnor UO_709 (O_709,N_13764,N_14788);
nor UO_710 (O_710,N_14761,N_13604);
nand UO_711 (O_711,N_13881,N_14870);
or UO_712 (O_712,N_14614,N_14162);
or UO_713 (O_713,N_14632,N_13933);
nor UO_714 (O_714,N_14795,N_13885);
and UO_715 (O_715,N_13833,N_14172);
nand UO_716 (O_716,N_14124,N_13587);
and UO_717 (O_717,N_14657,N_14047);
nand UO_718 (O_718,N_14851,N_14460);
nand UO_719 (O_719,N_14412,N_14705);
or UO_720 (O_720,N_13770,N_13677);
or UO_721 (O_721,N_13745,N_13687);
nor UO_722 (O_722,N_14855,N_14226);
nand UO_723 (O_723,N_14585,N_14304);
xor UO_724 (O_724,N_13544,N_14959);
and UO_725 (O_725,N_14435,N_13717);
or UO_726 (O_726,N_14150,N_13980);
or UO_727 (O_727,N_13645,N_14288);
nor UO_728 (O_728,N_14472,N_14387);
or UO_729 (O_729,N_13970,N_14318);
or UO_730 (O_730,N_14694,N_14680);
or UO_731 (O_731,N_14014,N_14249);
and UO_732 (O_732,N_14362,N_14789);
nor UO_733 (O_733,N_13961,N_13791);
or UO_734 (O_734,N_14961,N_13784);
or UO_735 (O_735,N_13990,N_14500);
nor UO_736 (O_736,N_13607,N_14928);
nand UO_737 (O_737,N_13822,N_14528);
and UO_738 (O_738,N_13850,N_14459);
nor UO_739 (O_739,N_14551,N_14352);
and UO_740 (O_740,N_14316,N_14159);
or UO_741 (O_741,N_14488,N_14714);
nor UO_742 (O_742,N_14596,N_14879);
or UO_743 (O_743,N_14191,N_14917);
xor UO_744 (O_744,N_14793,N_14243);
and UO_745 (O_745,N_14286,N_13828);
nor UO_746 (O_746,N_14731,N_13941);
xor UO_747 (O_747,N_14790,N_14420);
nand UO_748 (O_748,N_14519,N_14880);
and UO_749 (O_749,N_14811,N_14954);
nand UO_750 (O_750,N_14635,N_13595);
nand UO_751 (O_751,N_13920,N_14480);
and UO_752 (O_752,N_13879,N_13571);
xnor UO_753 (O_753,N_13903,N_14996);
or UO_754 (O_754,N_14502,N_14087);
xor UO_755 (O_755,N_14486,N_13575);
and UO_756 (O_756,N_14172,N_13724);
nand UO_757 (O_757,N_14632,N_13763);
nor UO_758 (O_758,N_14514,N_13501);
or UO_759 (O_759,N_14521,N_13731);
nor UO_760 (O_760,N_14975,N_14450);
and UO_761 (O_761,N_13670,N_14073);
and UO_762 (O_762,N_13548,N_14479);
or UO_763 (O_763,N_14353,N_14292);
and UO_764 (O_764,N_14288,N_13607);
and UO_765 (O_765,N_14622,N_14739);
nand UO_766 (O_766,N_14183,N_13864);
nand UO_767 (O_767,N_13907,N_13738);
nand UO_768 (O_768,N_14151,N_13501);
xnor UO_769 (O_769,N_13954,N_13590);
xnor UO_770 (O_770,N_14212,N_14348);
or UO_771 (O_771,N_13646,N_13509);
nand UO_772 (O_772,N_13976,N_13993);
or UO_773 (O_773,N_13651,N_13985);
nand UO_774 (O_774,N_13865,N_13762);
and UO_775 (O_775,N_14758,N_14549);
xnor UO_776 (O_776,N_14961,N_14072);
and UO_777 (O_777,N_14102,N_14504);
or UO_778 (O_778,N_14608,N_14752);
xor UO_779 (O_779,N_14422,N_13791);
nor UO_780 (O_780,N_14489,N_14230);
nand UO_781 (O_781,N_14461,N_14712);
xnor UO_782 (O_782,N_14022,N_14524);
and UO_783 (O_783,N_13801,N_14278);
and UO_784 (O_784,N_14938,N_14421);
and UO_785 (O_785,N_13782,N_14417);
nor UO_786 (O_786,N_14082,N_13621);
xor UO_787 (O_787,N_14573,N_14031);
xor UO_788 (O_788,N_14451,N_14396);
nor UO_789 (O_789,N_14220,N_14914);
nand UO_790 (O_790,N_13678,N_14722);
or UO_791 (O_791,N_14486,N_14509);
xnor UO_792 (O_792,N_14788,N_14379);
and UO_793 (O_793,N_14603,N_14090);
nor UO_794 (O_794,N_14062,N_13902);
nor UO_795 (O_795,N_14440,N_13589);
or UO_796 (O_796,N_13849,N_14317);
or UO_797 (O_797,N_13647,N_13928);
or UO_798 (O_798,N_13767,N_13807);
nor UO_799 (O_799,N_14473,N_13935);
and UO_800 (O_800,N_14558,N_13749);
nor UO_801 (O_801,N_14780,N_14282);
nand UO_802 (O_802,N_14250,N_14352);
and UO_803 (O_803,N_13530,N_14960);
xnor UO_804 (O_804,N_13977,N_14896);
or UO_805 (O_805,N_13834,N_13999);
or UO_806 (O_806,N_14502,N_13925);
nor UO_807 (O_807,N_14136,N_14911);
nand UO_808 (O_808,N_14221,N_13757);
nor UO_809 (O_809,N_14512,N_13853);
and UO_810 (O_810,N_14912,N_13871);
and UO_811 (O_811,N_14514,N_13704);
or UO_812 (O_812,N_14690,N_14287);
nand UO_813 (O_813,N_14793,N_13844);
xor UO_814 (O_814,N_13678,N_14336);
or UO_815 (O_815,N_14291,N_14699);
and UO_816 (O_816,N_13522,N_14867);
and UO_817 (O_817,N_14764,N_14971);
and UO_818 (O_818,N_14201,N_14953);
xnor UO_819 (O_819,N_14969,N_14496);
or UO_820 (O_820,N_14183,N_14257);
and UO_821 (O_821,N_14390,N_13809);
nor UO_822 (O_822,N_13527,N_14997);
nand UO_823 (O_823,N_14783,N_14793);
nand UO_824 (O_824,N_13628,N_13745);
nand UO_825 (O_825,N_14152,N_14149);
and UO_826 (O_826,N_14897,N_14362);
nand UO_827 (O_827,N_13981,N_13864);
nand UO_828 (O_828,N_14875,N_14323);
or UO_829 (O_829,N_14850,N_14683);
nand UO_830 (O_830,N_14976,N_14434);
and UO_831 (O_831,N_14645,N_14784);
or UO_832 (O_832,N_14439,N_13764);
xnor UO_833 (O_833,N_13745,N_13610);
or UO_834 (O_834,N_14664,N_13538);
nand UO_835 (O_835,N_14879,N_13611);
xor UO_836 (O_836,N_13670,N_14178);
xor UO_837 (O_837,N_13524,N_13846);
nand UO_838 (O_838,N_14741,N_14929);
xor UO_839 (O_839,N_13594,N_14976);
nor UO_840 (O_840,N_13920,N_13968);
or UO_841 (O_841,N_14199,N_14107);
nor UO_842 (O_842,N_14399,N_13763);
or UO_843 (O_843,N_14572,N_13632);
and UO_844 (O_844,N_14287,N_14536);
nand UO_845 (O_845,N_14569,N_14769);
nor UO_846 (O_846,N_14831,N_14176);
and UO_847 (O_847,N_14848,N_13908);
or UO_848 (O_848,N_14300,N_14454);
or UO_849 (O_849,N_14351,N_13901);
nand UO_850 (O_850,N_14949,N_14179);
and UO_851 (O_851,N_14085,N_14296);
nor UO_852 (O_852,N_14977,N_13836);
nand UO_853 (O_853,N_14268,N_13545);
or UO_854 (O_854,N_14421,N_14720);
nor UO_855 (O_855,N_13615,N_14009);
xor UO_856 (O_856,N_14858,N_14410);
and UO_857 (O_857,N_14704,N_13676);
and UO_858 (O_858,N_14023,N_14876);
nor UO_859 (O_859,N_14213,N_14651);
nand UO_860 (O_860,N_13672,N_14701);
and UO_861 (O_861,N_14907,N_14980);
nand UO_862 (O_862,N_14361,N_13702);
nand UO_863 (O_863,N_14708,N_14070);
nor UO_864 (O_864,N_14233,N_13659);
or UO_865 (O_865,N_13897,N_13835);
xnor UO_866 (O_866,N_14416,N_13651);
or UO_867 (O_867,N_14090,N_14982);
xor UO_868 (O_868,N_14824,N_14907);
nor UO_869 (O_869,N_14992,N_13576);
nand UO_870 (O_870,N_14285,N_14299);
and UO_871 (O_871,N_14690,N_13552);
or UO_872 (O_872,N_14527,N_14249);
and UO_873 (O_873,N_14722,N_14899);
nor UO_874 (O_874,N_14036,N_14835);
nand UO_875 (O_875,N_14555,N_14955);
xor UO_876 (O_876,N_14665,N_14914);
and UO_877 (O_877,N_13653,N_14708);
or UO_878 (O_878,N_13921,N_14057);
nand UO_879 (O_879,N_14100,N_13953);
xnor UO_880 (O_880,N_13531,N_14090);
nand UO_881 (O_881,N_14704,N_14494);
or UO_882 (O_882,N_13744,N_14220);
or UO_883 (O_883,N_13515,N_13813);
nor UO_884 (O_884,N_14432,N_13595);
nor UO_885 (O_885,N_14377,N_14068);
nor UO_886 (O_886,N_13582,N_13783);
nor UO_887 (O_887,N_13562,N_13855);
or UO_888 (O_888,N_13970,N_14464);
or UO_889 (O_889,N_13885,N_13695);
and UO_890 (O_890,N_13711,N_13566);
nor UO_891 (O_891,N_14836,N_13935);
and UO_892 (O_892,N_13901,N_14126);
nand UO_893 (O_893,N_14678,N_14626);
or UO_894 (O_894,N_13760,N_14253);
and UO_895 (O_895,N_14036,N_14259);
or UO_896 (O_896,N_13586,N_14913);
nor UO_897 (O_897,N_13812,N_13790);
nor UO_898 (O_898,N_13982,N_14666);
or UO_899 (O_899,N_14331,N_14507);
nor UO_900 (O_900,N_14764,N_13830);
nand UO_901 (O_901,N_14909,N_13684);
nand UO_902 (O_902,N_13528,N_14672);
xor UO_903 (O_903,N_13753,N_14677);
and UO_904 (O_904,N_14786,N_14398);
nand UO_905 (O_905,N_14979,N_14035);
nor UO_906 (O_906,N_14378,N_14446);
and UO_907 (O_907,N_14916,N_14766);
and UO_908 (O_908,N_14629,N_13679);
or UO_909 (O_909,N_14367,N_14875);
nand UO_910 (O_910,N_13741,N_14015);
or UO_911 (O_911,N_14303,N_13797);
or UO_912 (O_912,N_14543,N_14885);
and UO_913 (O_913,N_14786,N_14108);
nor UO_914 (O_914,N_14242,N_14043);
and UO_915 (O_915,N_13956,N_14327);
nor UO_916 (O_916,N_14754,N_14517);
and UO_917 (O_917,N_14865,N_13589);
and UO_918 (O_918,N_14305,N_13865);
nor UO_919 (O_919,N_14287,N_14797);
and UO_920 (O_920,N_14854,N_13638);
or UO_921 (O_921,N_13605,N_13517);
nand UO_922 (O_922,N_14268,N_14823);
and UO_923 (O_923,N_13662,N_13975);
and UO_924 (O_924,N_13870,N_14022);
nand UO_925 (O_925,N_13519,N_13532);
or UO_926 (O_926,N_14163,N_14613);
nand UO_927 (O_927,N_13739,N_14080);
nand UO_928 (O_928,N_14586,N_13549);
or UO_929 (O_929,N_14799,N_14726);
or UO_930 (O_930,N_13878,N_14470);
or UO_931 (O_931,N_14949,N_13937);
and UO_932 (O_932,N_14634,N_14877);
nor UO_933 (O_933,N_14160,N_14978);
and UO_934 (O_934,N_14057,N_13902);
and UO_935 (O_935,N_14282,N_14197);
or UO_936 (O_936,N_14753,N_14256);
nor UO_937 (O_937,N_14003,N_13504);
and UO_938 (O_938,N_14040,N_14958);
and UO_939 (O_939,N_14938,N_13957);
nor UO_940 (O_940,N_14620,N_14585);
nor UO_941 (O_941,N_14852,N_13678);
nor UO_942 (O_942,N_13902,N_13728);
nor UO_943 (O_943,N_14031,N_14710);
nor UO_944 (O_944,N_14791,N_14049);
or UO_945 (O_945,N_14528,N_14028);
nor UO_946 (O_946,N_13943,N_14185);
nor UO_947 (O_947,N_14320,N_13776);
xnor UO_948 (O_948,N_14569,N_14564);
or UO_949 (O_949,N_14838,N_14232);
or UO_950 (O_950,N_13764,N_14345);
nand UO_951 (O_951,N_14412,N_14041);
xnor UO_952 (O_952,N_14028,N_14184);
nand UO_953 (O_953,N_13625,N_14077);
and UO_954 (O_954,N_14765,N_14443);
nand UO_955 (O_955,N_14480,N_13661);
xnor UO_956 (O_956,N_14520,N_14485);
nor UO_957 (O_957,N_14901,N_14450);
or UO_958 (O_958,N_14422,N_13611);
or UO_959 (O_959,N_14378,N_14586);
or UO_960 (O_960,N_14514,N_14847);
or UO_961 (O_961,N_13972,N_14317);
nand UO_962 (O_962,N_14128,N_13897);
nand UO_963 (O_963,N_14396,N_14768);
nand UO_964 (O_964,N_14367,N_13843);
and UO_965 (O_965,N_13949,N_13816);
nand UO_966 (O_966,N_14088,N_14618);
or UO_967 (O_967,N_13525,N_14232);
or UO_968 (O_968,N_14165,N_14824);
or UO_969 (O_969,N_14183,N_14771);
and UO_970 (O_970,N_13819,N_14280);
nand UO_971 (O_971,N_14268,N_14721);
and UO_972 (O_972,N_14168,N_13939);
nor UO_973 (O_973,N_14021,N_14383);
or UO_974 (O_974,N_14761,N_13553);
or UO_975 (O_975,N_14699,N_13598);
nor UO_976 (O_976,N_13713,N_14203);
or UO_977 (O_977,N_13839,N_13898);
or UO_978 (O_978,N_13786,N_13774);
nor UO_979 (O_979,N_14561,N_14106);
or UO_980 (O_980,N_13745,N_13685);
nor UO_981 (O_981,N_14788,N_13982);
nand UO_982 (O_982,N_14990,N_13927);
nor UO_983 (O_983,N_13747,N_13877);
nand UO_984 (O_984,N_14214,N_13728);
and UO_985 (O_985,N_14852,N_14499);
or UO_986 (O_986,N_13661,N_14071);
and UO_987 (O_987,N_14586,N_14438);
nand UO_988 (O_988,N_13702,N_14638);
nor UO_989 (O_989,N_13718,N_13568);
nor UO_990 (O_990,N_14459,N_14079);
nand UO_991 (O_991,N_14212,N_14817);
nor UO_992 (O_992,N_13839,N_13941);
nand UO_993 (O_993,N_14212,N_14542);
and UO_994 (O_994,N_13664,N_14308);
nand UO_995 (O_995,N_14591,N_14837);
nor UO_996 (O_996,N_14545,N_14401);
and UO_997 (O_997,N_14676,N_14120);
nor UO_998 (O_998,N_14284,N_14508);
nor UO_999 (O_999,N_14653,N_13981);
xnor UO_1000 (O_1000,N_14002,N_14046);
or UO_1001 (O_1001,N_14039,N_13886);
or UO_1002 (O_1002,N_14538,N_14822);
and UO_1003 (O_1003,N_14515,N_13501);
or UO_1004 (O_1004,N_14156,N_14589);
nand UO_1005 (O_1005,N_14891,N_14060);
nand UO_1006 (O_1006,N_14538,N_14409);
xor UO_1007 (O_1007,N_13677,N_14233);
nor UO_1008 (O_1008,N_13787,N_13698);
nor UO_1009 (O_1009,N_13710,N_14465);
nor UO_1010 (O_1010,N_14732,N_13790);
nor UO_1011 (O_1011,N_14943,N_13934);
nor UO_1012 (O_1012,N_14496,N_14744);
nor UO_1013 (O_1013,N_14697,N_13856);
xnor UO_1014 (O_1014,N_14283,N_14197);
or UO_1015 (O_1015,N_13505,N_14747);
xnor UO_1016 (O_1016,N_14361,N_14155);
nand UO_1017 (O_1017,N_14514,N_14369);
nor UO_1018 (O_1018,N_14196,N_13850);
or UO_1019 (O_1019,N_14611,N_14366);
nand UO_1020 (O_1020,N_14277,N_14522);
and UO_1021 (O_1021,N_13996,N_13662);
nand UO_1022 (O_1022,N_14258,N_14276);
and UO_1023 (O_1023,N_14371,N_14886);
nor UO_1024 (O_1024,N_14938,N_14490);
nor UO_1025 (O_1025,N_14437,N_14198);
nor UO_1026 (O_1026,N_14220,N_14401);
nand UO_1027 (O_1027,N_14858,N_14744);
or UO_1028 (O_1028,N_13828,N_14187);
nand UO_1029 (O_1029,N_13797,N_14510);
or UO_1030 (O_1030,N_14816,N_13693);
nor UO_1031 (O_1031,N_13807,N_14963);
and UO_1032 (O_1032,N_14653,N_13592);
nor UO_1033 (O_1033,N_13651,N_14164);
and UO_1034 (O_1034,N_14163,N_14409);
nor UO_1035 (O_1035,N_13953,N_13780);
or UO_1036 (O_1036,N_13562,N_13530);
or UO_1037 (O_1037,N_14720,N_13573);
nor UO_1038 (O_1038,N_14945,N_13680);
or UO_1039 (O_1039,N_14112,N_14471);
nor UO_1040 (O_1040,N_14583,N_14522);
nor UO_1041 (O_1041,N_13570,N_13576);
xnor UO_1042 (O_1042,N_13678,N_14905);
or UO_1043 (O_1043,N_13706,N_13629);
nand UO_1044 (O_1044,N_14482,N_14166);
nand UO_1045 (O_1045,N_14181,N_14335);
nand UO_1046 (O_1046,N_14426,N_14856);
nand UO_1047 (O_1047,N_13555,N_14305);
xor UO_1048 (O_1048,N_14879,N_14672);
xnor UO_1049 (O_1049,N_14934,N_13682);
and UO_1050 (O_1050,N_14559,N_14634);
nor UO_1051 (O_1051,N_14980,N_14915);
and UO_1052 (O_1052,N_13560,N_14458);
nand UO_1053 (O_1053,N_14310,N_14282);
or UO_1054 (O_1054,N_13868,N_14868);
or UO_1055 (O_1055,N_14217,N_14013);
xnor UO_1056 (O_1056,N_14150,N_13820);
and UO_1057 (O_1057,N_13668,N_13965);
nand UO_1058 (O_1058,N_13581,N_14588);
or UO_1059 (O_1059,N_14681,N_13745);
or UO_1060 (O_1060,N_14444,N_14040);
nor UO_1061 (O_1061,N_13814,N_14067);
nand UO_1062 (O_1062,N_14518,N_14423);
or UO_1063 (O_1063,N_13955,N_13634);
nor UO_1064 (O_1064,N_14687,N_14068);
nor UO_1065 (O_1065,N_14188,N_13546);
nor UO_1066 (O_1066,N_13830,N_13844);
nor UO_1067 (O_1067,N_13807,N_14905);
xor UO_1068 (O_1068,N_13868,N_14095);
or UO_1069 (O_1069,N_13619,N_13559);
nand UO_1070 (O_1070,N_13614,N_13516);
nor UO_1071 (O_1071,N_13859,N_14406);
or UO_1072 (O_1072,N_14281,N_14596);
or UO_1073 (O_1073,N_14180,N_14889);
or UO_1074 (O_1074,N_13744,N_14519);
or UO_1075 (O_1075,N_13790,N_14897);
and UO_1076 (O_1076,N_14459,N_14094);
xnor UO_1077 (O_1077,N_13899,N_13865);
nand UO_1078 (O_1078,N_14350,N_13859);
nor UO_1079 (O_1079,N_13610,N_14209);
xor UO_1080 (O_1080,N_14110,N_14348);
and UO_1081 (O_1081,N_14880,N_14944);
nand UO_1082 (O_1082,N_14956,N_14247);
or UO_1083 (O_1083,N_13998,N_14475);
and UO_1084 (O_1084,N_14897,N_14034);
or UO_1085 (O_1085,N_14771,N_14342);
nand UO_1086 (O_1086,N_14886,N_13659);
nor UO_1087 (O_1087,N_14752,N_14477);
and UO_1088 (O_1088,N_13885,N_14200);
or UO_1089 (O_1089,N_14430,N_13780);
or UO_1090 (O_1090,N_13576,N_14209);
nor UO_1091 (O_1091,N_13750,N_14372);
nor UO_1092 (O_1092,N_14635,N_14142);
or UO_1093 (O_1093,N_14805,N_14191);
xnor UO_1094 (O_1094,N_14997,N_13863);
and UO_1095 (O_1095,N_14451,N_14681);
and UO_1096 (O_1096,N_13735,N_13567);
or UO_1097 (O_1097,N_14278,N_14531);
nor UO_1098 (O_1098,N_14899,N_14322);
xnor UO_1099 (O_1099,N_13567,N_14936);
and UO_1100 (O_1100,N_14326,N_14809);
nand UO_1101 (O_1101,N_13955,N_14548);
and UO_1102 (O_1102,N_13921,N_14076);
or UO_1103 (O_1103,N_14056,N_14266);
nor UO_1104 (O_1104,N_14359,N_13511);
or UO_1105 (O_1105,N_14433,N_14694);
and UO_1106 (O_1106,N_14952,N_14912);
nor UO_1107 (O_1107,N_14541,N_14497);
and UO_1108 (O_1108,N_13893,N_13551);
nor UO_1109 (O_1109,N_13532,N_14220);
and UO_1110 (O_1110,N_13610,N_13921);
nand UO_1111 (O_1111,N_13934,N_13869);
nor UO_1112 (O_1112,N_14921,N_14624);
nand UO_1113 (O_1113,N_13512,N_14686);
nand UO_1114 (O_1114,N_13599,N_14967);
xor UO_1115 (O_1115,N_14251,N_14476);
xnor UO_1116 (O_1116,N_14796,N_14736);
or UO_1117 (O_1117,N_14679,N_14169);
nor UO_1118 (O_1118,N_14675,N_13952);
nand UO_1119 (O_1119,N_13684,N_14966);
nand UO_1120 (O_1120,N_14037,N_13976);
xnor UO_1121 (O_1121,N_14781,N_13863);
nor UO_1122 (O_1122,N_14795,N_14781);
nand UO_1123 (O_1123,N_13885,N_13582);
and UO_1124 (O_1124,N_14023,N_14657);
nand UO_1125 (O_1125,N_13847,N_13812);
nor UO_1126 (O_1126,N_14505,N_14304);
nor UO_1127 (O_1127,N_13787,N_14999);
and UO_1128 (O_1128,N_14575,N_14038);
nand UO_1129 (O_1129,N_14660,N_14067);
nand UO_1130 (O_1130,N_14835,N_14890);
nor UO_1131 (O_1131,N_14298,N_14907);
or UO_1132 (O_1132,N_13752,N_14479);
or UO_1133 (O_1133,N_14609,N_14209);
nor UO_1134 (O_1134,N_14233,N_14155);
xnor UO_1135 (O_1135,N_13694,N_14049);
nand UO_1136 (O_1136,N_14090,N_13721);
or UO_1137 (O_1137,N_14248,N_14751);
nand UO_1138 (O_1138,N_14349,N_14588);
nand UO_1139 (O_1139,N_14682,N_13563);
and UO_1140 (O_1140,N_14489,N_13970);
nor UO_1141 (O_1141,N_14764,N_13967);
and UO_1142 (O_1142,N_14909,N_14465);
nor UO_1143 (O_1143,N_13817,N_13834);
or UO_1144 (O_1144,N_14218,N_14774);
or UO_1145 (O_1145,N_14383,N_14509);
or UO_1146 (O_1146,N_14003,N_14370);
and UO_1147 (O_1147,N_14396,N_14603);
nor UO_1148 (O_1148,N_14833,N_14491);
nor UO_1149 (O_1149,N_14463,N_13647);
xnor UO_1150 (O_1150,N_13835,N_13747);
nand UO_1151 (O_1151,N_14017,N_14168);
or UO_1152 (O_1152,N_14415,N_14379);
nor UO_1153 (O_1153,N_13957,N_13742);
and UO_1154 (O_1154,N_14249,N_14402);
and UO_1155 (O_1155,N_14234,N_14325);
nand UO_1156 (O_1156,N_14142,N_14616);
nor UO_1157 (O_1157,N_13924,N_14167);
or UO_1158 (O_1158,N_14178,N_14308);
nor UO_1159 (O_1159,N_14263,N_14670);
nand UO_1160 (O_1160,N_14509,N_14817);
or UO_1161 (O_1161,N_14949,N_13724);
nor UO_1162 (O_1162,N_14192,N_13749);
or UO_1163 (O_1163,N_13978,N_14864);
nor UO_1164 (O_1164,N_14842,N_14582);
or UO_1165 (O_1165,N_14492,N_14413);
nor UO_1166 (O_1166,N_13857,N_14667);
nor UO_1167 (O_1167,N_14979,N_14209);
xnor UO_1168 (O_1168,N_13541,N_14354);
nand UO_1169 (O_1169,N_14759,N_13795);
or UO_1170 (O_1170,N_14769,N_14982);
nor UO_1171 (O_1171,N_13736,N_14609);
nand UO_1172 (O_1172,N_14567,N_14051);
or UO_1173 (O_1173,N_13532,N_14766);
nor UO_1174 (O_1174,N_13908,N_14334);
or UO_1175 (O_1175,N_14667,N_14886);
nor UO_1176 (O_1176,N_14370,N_14983);
xnor UO_1177 (O_1177,N_14890,N_14360);
xnor UO_1178 (O_1178,N_14515,N_13793);
or UO_1179 (O_1179,N_14977,N_14456);
xnor UO_1180 (O_1180,N_14021,N_14052);
nand UO_1181 (O_1181,N_13682,N_14900);
and UO_1182 (O_1182,N_13670,N_14983);
nand UO_1183 (O_1183,N_14638,N_13782);
and UO_1184 (O_1184,N_14539,N_13546);
xor UO_1185 (O_1185,N_14520,N_13638);
nor UO_1186 (O_1186,N_14581,N_14155);
and UO_1187 (O_1187,N_13510,N_14713);
and UO_1188 (O_1188,N_14796,N_13646);
xor UO_1189 (O_1189,N_13593,N_13977);
and UO_1190 (O_1190,N_14243,N_13713);
and UO_1191 (O_1191,N_14912,N_14816);
xor UO_1192 (O_1192,N_14079,N_14444);
nand UO_1193 (O_1193,N_13700,N_13647);
nor UO_1194 (O_1194,N_13856,N_14417);
nor UO_1195 (O_1195,N_13790,N_13648);
nand UO_1196 (O_1196,N_13583,N_13970);
nor UO_1197 (O_1197,N_14888,N_13859);
nor UO_1198 (O_1198,N_14851,N_13657);
xor UO_1199 (O_1199,N_14381,N_14562);
nand UO_1200 (O_1200,N_14464,N_13705);
nor UO_1201 (O_1201,N_13843,N_13859);
nor UO_1202 (O_1202,N_14479,N_14181);
or UO_1203 (O_1203,N_14425,N_14281);
nand UO_1204 (O_1204,N_13689,N_14746);
nor UO_1205 (O_1205,N_14101,N_13565);
and UO_1206 (O_1206,N_13665,N_14833);
and UO_1207 (O_1207,N_14996,N_13650);
nand UO_1208 (O_1208,N_14744,N_14868);
xor UO_1209 (O_1209,N_13555,N_14118);
nor UO_1210 (O_1210,N_14147,N_14418);
nand UO_1211 (O_1211,N_14586,N_14934);
xor UO_1212 (O_1212,N_14110,N_14557);
or UO_1213 (O_1213,N_14575,N_14822);
nor UO_1214 (O_1214,N_14031,N_14726);
nand UO_1215 (O_1215,N_13895,N_13763);
or UO_1216 (O_1216,N_13614,N_14756);
and UO_1217 (O_1217,N_14999,N_14485);
and UO_1218 (O_1218,N_13782,N_14051);
nand UO_1219 (O_1219,N_14667,N_13912);
or UO_1220 (O_1220,N_14603,N_13501);
or UO_1221 (O_1221,N_14815,N_13819);
or UO_1222 (O_1222,N_13936,N_14404);
xor UO_1223 (O_1223,N_13663,N_14216);
nand UO_1224 (O_1224,N_14703,N_14243);
and UO_1225 (O_1225,N_14880,N_13911);
nor UO_1226 (O_1226,N_13832,N_14803);
nand UO_1227 (O_1227,N_14482,N_13622);
or UO_1228 (O_1228,N_14214,N_14065);
nor UO_1229 (O_1229,N_14194,N_14191);
or UO_1230 (O_1230,N_13545,N_14769);
or UO_1231 (O_1231,N_13586,N_14073);
or UO_1232 (O_1232,N_14255,N_14471);
nor UO_1233 (O_1233,N_14197,N_14229);
and UO_1234 (O_1234,N_14569,N_14755);
nor UO_1235 (O_1235,N_14701,N_14825);
xnor UO_1236 (O_1236,N_14905,N_14352);
nand UO_1237 (O_1237,N_14608,N_13616);
and UO_1238 (O_1238,N_14189,N_14143);
or UO_1239 (O_1239,N_13677,N_13705);
nand UO_1240 (O_1240,N_14026,N_14499);
and UO_1241 (O_1241,N_14144,N_13764);
and UO_1242 (O_1242,N_14389,N_14260);
nor UO_1243 (O_1243,N_14943,N_13755);
or UO_1244 (O_1244,N_13613,N_13751);
nor UO_1245 (O_1245,N_14301,N_14645);
nor UO_1246 (O_1246,N_14196,N_14914);
nand UO_1247 (O_1247,N_13922,N_14098);
and UO_1248 (O_1248,N_14746,N_13536);
and UO_1249 (O_1249,N_14382,N_14233);
or UO_1250 (O_1250,N_14901,N_14772);
nand UO_1251 (O_1251,N_13960,N_14940);
or UO_1252 (O_1252,N_14939,N_13754);
and UO_1253 (O_1253,N_14622,N_14951);
nor UO_1254 (O_1254,N_14549,N_13628);
nand UO_1255 (O_1255,N_13682,N_14309);
or UO_1256 (O_1256,N_13558,N_14005);
and UO_1257 (O_1257,N_14410,N_13850);
or UO_1258 (O_1258,N_13639,N_14757);
nor UO_1259 (O_1259,N_14195,N_14959);
nand UO_1260 (O_1260,N_14298,N_14285);
nor UO_1261 (O_1261,N_13885,N_13893);
nor UO_1262 (O_1262,N_13822,N_14862);
or UO_1263 (O_1263,N_13831,N_13687);
nor UO_1264 (O_1264,N_13684,N_13705);
nor UO_1265 (O_1265,N_14526,N_13610);
nor UO_1266 (O_1266,N_14360,N_14799);
xor UO_1267 (O_1267,N_13797,N_14377);
and UO_1268 (O_1268,N_13642,N_14477);
xor UO_1269 (O_1269,N_14471,N_13511);
and UO_1270 (O_1270,N_14785,N_13700);
or UO_1271 (O_1271,N_14937,N_13774);
or UO_1272 (O_1272,N_13936,N_14705);
nand UO_1273 (O_1273,N_13921,N_14480);
nand UO_1274 (O_1274,N_14892,N_14851);
nand UO_1275 (O_1275,N_14586,N_13991);
or UO_1276 (O_1276,N_13898,N_13526);
nor UO_1277 (O_1277,N_13959,N_14161);
or UO_1278 (O_1278,N_13994,N_14191);
or UO_1279 (O_1279,N_14670,N_13695);
nor UO_1280 (O_1280,N_14790,N_13967);
and UO_1281 (O_1281,N_14327,N_14346);
nor UO_1282 (O_1282,N_13725,N_14805);
and UO_1283 (O_1283,N_13560,N_14951);
and UO_1284 (O_1284,N_14458,N_14723);
and UO_1285 (O_1285,N_13981,N_14411);
nor UO_1286 (O_1286,N_14257,N_14080);
and UO_1287 (O_1287,N_13987,N_14887);
or UO_1288 (O_1288,N_13921,N_14374);
nor UO_1289 (O_1289,N_14473,N_14720);
nor UO_1290 (O_1290,N_13983,N_13788);
nand UO_1291 (O_1291,N_13945,N_14067);
or UO_1292 (O_1292,N_13728,N_14171);
and UO_1293 (O_1293,N_13552,N_13736);
nor UO_1294 (O_1294,N_14315,N_14885);
and UO_1295 (O_1295,N_14905,N_14193);
xor UO_1296 (O_1296,N_14058,N_13768);
nor UO_1297 (O_1297,N_13808,N_14774);
nor UO_1298 (O_1298,N_14376,N_14910);
and UO_1299 (O_1299,N_14498,N_14691);
nand UO_1300 (O_1300,N_14259,N_14200);
or UO_1301 (O_1301,N_13871,N_14703);
or UO_1302 (O_1302,N_14285,N_13587);
nor UO_1303 (O_1303,N_14581,N_14721);
xnor UO_1304 (O_1304,N_14606,N_14223);
xnor UO_1305 (O_1305,N_14028,N_14190);
and UO_1306 (O_1306,N_14460,N_13859);
nand UO_1307 (O_1307,N_14104,N_14914);
nand UO_1308 (O_1308,N_14891,N_13758);
nand UO_1309 (O_1309,N_13597,N_13974);
nor UO_1310 (O_1310,N_14005,N_14990);
nor UO_1311 (O_1311,N_14428,N_13557);
or UO_1312 (O_1312,N_14027,N_14029);
xnor UO_1313 (O_1313,N_13679,N_13572);
xnor UO_1314 (O_1314,N_14074,N_13734);
nand UO_1315 (O_1315,N_13615,N_13754);
or UO_1316 (O_1316,N_14790,N_14040);
nor UO_1317 (O_1317,N_14447,N_13899);
nand UO_1318 (O_1318,N_14097,N_13819);
nor UO_1319 (O_1319,N_13553,N_14712);
or UO_1320 (O_1320,N_13500,N_14993);
xor UO_1321 (O_1321,N_13693,N_13771);
nand UO_1322 (O_1322,N_13582,N_14505);
nor UO_1323 (O_1323,N_14423,N_13598);
nand UO_1324 (O_1324,N_14966,N_14462);
or UO_1325 (O_1325,N_14694,N_14570);
xor UO_1326 (O_1326,N_14779,N_13995);
or UO_1327 (O_1327,N_13648,N_14806);
nor UO_1328 (O_1328,N_13943,N_13844);
nand UO_1329 (O_1329,N_13555,N_13574);
nor UO_1330 (O_1330,N_14700,N_13891);
nand UO_1331 (O_1331,N_14416,N_13633);
and UO_1332 (O_1332,N_14928,N_13984);
nor UO_1333 (O_1333,N_14697,N_13524);
and UO_1334 (O_1334,N_14948,N_13530);
nand UO_1335 (O_1335,N_14218,N_13721);
nor UO_1336 (O_1336,N_14224,N_14229);
and UO_1337 (O_1337,N_13949,N_13856);
nor UO_1338 (O_1338,N_13513,N_13880);
or UO_1339 (O_1339,N_14099,N_13601);
and UO_1340 (O_1340,N_14933,N_14875);
xnor UO_1341 (O_1341,N_14280,N_14300);
nand UO_1342 (O_1342,N_13699,N_13873);
or UO_1343 (O_1343,N_14611,N_13987);
or UO_1344 (O_1344,N_14335,N_14113);
xnor UO_1345 (O_1345,N_14074,N_13997);
nand UO_1346 (O_1346,N_14745,N_14151);
nand UO_1347 (O_1347,N_14500,N_14240);
and UO_1348 (O_1348,N_13622,N_14581);
nor UO_1349 (O_1349,N_14579,N_13660);
and UO_1350 (O_1350,N_14041,N_13913);
or UO_1351 (O_1351,N_14140,N_14209);
or UO_1352 (O_1352,N_14287,N_14334);
and UO_1353 (O_1353,N_13875,N_14710);
nor UO_1354 (O_1354,N_14207,N_14182);
and UO_1355 (O_1355,N_13934,N_14479);
nand UO_1356 (O_1356,N_14320,N_14005);
xnor UO_1357 (O_1357,N_13749,N_14175);
nand UO_1358 (O_1358,N_14299,N_14307);
or UO_1359 (O_1359,N_14940,N_14659);
nor UO_1360 (O_1360,N_13548,N_13944);
nor UO_1361 (O_1361,N_14584,N_14360);
xor UO_1362 (O_1362,N_14109,N_14092);
xor UO_1363 (O_1363,N_14047,N_14136);
nor UO_1364 (O_1364,N_13618,N_13988);
and UO_1365 (O_1365,N_13603,N_13844);
and UO_1366 (O_1366,N_14752,N_13657);
and UO_1367 (O_1367,N_14966,N_13862);
nor UO_1368 (O_1368,N_14744,N_14296);
nand UO_1369 (O_1369,N_14841,N_14880);
nor UO_1370 (O_1370,N_14825,N_14910);
nor UO_1371 (O_1371,N_14519,N_14321);
nor UO_1372 (O_1372,N_13889,N_13617);
nor UO_1373 (O_1373,N_13960,N_14130);
and UO_1374 (O_1374,N_13791,N_14003);
nand UO_1375 (O_1375,N_14079,N_13915);
nand UO_1376 (O_1376,N_14690,N_14145);
or UO_1377 (O_1377,N_14007,N_14733);
nand UO_1378 (O_1378,N_14304,N_13701);
nand UO_1379 (O_1379,N_14779,N_14870);
or UO_1380 (O_1380,N_14997,N_14189);
or UO_1381 (O_1381,N_14326,N_13574);
xor UO_1382 (O_1382,N_14608,N_14794);
or UO_1383 (O_1383,N_14801,N_13904);
and UO_1384 (O_1384,N_13657,N_14666);
and UO_1385 (O_1385,N_14191,N_13881);
nand UO_1386 (O_1386,N_13860,N_14421);
or UO_1387 (O_1387,N_14510,N_14827);
and UO_1388 (O_1388,N_14540,N_13865);
nand UO_1389 (O_1389,N_14486,N_13715);
xor UO_1390 (O_1390,N_14024,N_14899);
and UO_1391 (O_1391,N_14592,N_14910);
or UO_1392 (O_1392,N_14519,N_14439);
nor UO_1393 (O_1393,N_14796,N_14051);
or UO_1394 (O_1394,N_13600,N_14320);
nand UO_1395 (O_1395,N_14140,N_13985);
and UO_1396 (O_1396,N_13633,N_14861);
nand UO_1397 (O_1397,N_14721,N_14872);
and UO_1398 (O_1398,N_13950,N_13800);
nand UO_1399 (O_1399,N_14830,N_14953);
xor UO_1400 (O_1400,N_14438,N_14642);
or UO_1401 (O_1401,N_14706,N_13678);
or UO_1402 (O_1402,N_14922,N_13771);
nand UO_1403 (O_1403,N_13796,N_13708);
xor UO_1404 (O_1404,N_13517,N_14505);
nor UO_1405 (O_1405,N_13799,N_14134);
nand UO_1406 (O_1406,N_14153,N_14220);
nor UO_1407 (O_1407,N_14364,N_14804);
and UO_1408 (O_1408,N_13770,N_14618);
and UO_1409 (O_1409,N_14664,N_14618);
and UO_1410 (O_1410,N_14117,N_14529);
and UO_1411 (O_1411,N_14270,N_14595);
nor UO_1412 (O_1412,N_13755,N_14634);
xor UO_1413 (O_1413,N_13761,N_14360);
nor UO_1414 (O_1414,N_14621,N_14594);
nor UO_1415 (O_1415,N_14135,N_14810);
nand UO_1416 (O_1416,N_13534,N_14342);
and UO_1417 (O_1417,N_13663,N_13979);
nor UO_1418 (O_1418,N_14105,N_13511);
and UO_1419 (O_1419,N_13667,N_13873);
and UO_1420 (O_1420,N_14283,N_14567);
nand UO_1421 (O_1421,N_14222,N_14211);
nor UO_1422 (O_1422,N_14553,N_14315);
and UO_1423 (O_1423,N_13689,N_14734);
nand UO_1424 (O_1424,N_13735,N_14472);
and UO_1425 (O_1425,N_14705,N_14873);
or UO_1426 (O_1426,N_14432,N_14588);
and UO_1427 (O_1427,N_13521,N_14970);
and UO_1428 (O_1428,N_14637,N_13727);
nand UO_1429 (O_1429,N_14029,N_13985);
nor UO_1430 (O_1430,N_14630,N_14931);
nor UO_1431 (O_1431,N_14762,N_14861);
nand UO_1432 (O_1432,N_14866,N_14662);
and UO_1433 (O_1433,N_13763,N_14686);
and UO_1434 (O_1434,N_14202,N_14098);
or UO_1435 (O_1435,N_14967,N_14516);
nand UO_1436 (O_1436,N_14287,N_13629);
nor UO_1437 (O_1437,N_14961,N_14673);
xor UO_1438 (O_1438,N_14433,N_14414);
nand UO_1439 (O_1439,N_14431,N_14138);
nand UO_1440 (O_1440,N_14056,N_14090);
xnor UO_1441 (O_1441,N_14459,N_14444);
or UO_1442 (O_1442,N_14354,N_14274);
xor UO_1443 (O_1443,N_14502,N_13847);
xnor UO_1444 (O_1444,N_14809,N_13988);
nand UO_1445 (O_1445,N_14176,N_14646);
or UO_1446 (O_1446,N_14045,N_13932);
or UO_1447 (O_1447,N_13662,N_13575);
nor UO_1448 (O_1448,N_14180,N_14676);
or UO_1449 (O_1449,N_14173,N_13652);
nand UO_1450 (O_1450,N_14140,N_14752);
and UO_1451 (O_1451,N_14699,N_14177);
nor UO_1452 (O_1452,N_13685,N_14592);
and UO_1453 (O_1453,N_14900,N_14767);
and UO_1454 (O_1454,N_13609,N_14118);
or UO_1455 (O_1455,N_14494,N_13903);
or UO_1456 (O_1456,N_14562,N_13741);
xor UO_1457 (O_1457,N_13778,N_14607);
nand UO_1458 (O_1458,N_14339,N_14220);
nor UO_1459 (O_1459,N_14538,N_13823);
or UO_1460 (O_1460,N_14652,N_13978);
and UO_1461 (O_1461,N_13988,N_14694);
or UO_1462 (O_1462,N_14798,N_14042);
nand UO_1463 (O_1463,N_14482,N_14206);
or UO_1464 (O_1464,N_14033,N_13546);
nor UO_1465 (O_1465,N_13829,N_13926);
or UO_1466 (O_1466,N_14820,N_13927);
or UO_1467 (O_1467,N_14876,N_14724);
nor UO_1468 (O_1468,N_13626,N_13761);
or UO_1469 (O_1469,N_14677,N_13645);
or UO_1470 (O_1470,N_14082,N_14174);
nor UO_1471 (O_1471,N_13955,N_14378);
nand UO_1472 (O_1472,N_14675,N_14359);
nor UO_1473 (O_1473,N_13928,N_14913);
or UO_1474 (O_1474,N_13644,N_14080);
and UO_1475 (O_1475,N_13655,N_14363);
or UO_1476 (O_1476,N_13812,N_14454);
nand UO_1477 (O_1477,N_13785,N_13941);
nor UO_1478 (O_1478,N_14174,N_13722);
nor UO_1479 (O_1479,N_14857,N_14738);
or UO_1480 (O_1480,N_14073,N_14561);
xor UO_1481 (O_1481,N_13907,N_13783);
nor UO_1482 (O_1482,N_14247,N_14466);
and UO_1483 (O_1483,N_14822,N_14015);
nand UO_1484 (O_1484,N_13796,N_14285);
xnor UO_1485 (O_1485,N_13621,N_13793);
nand UO_1486 (O_1486,N_14108,N_14152);
and UO_1487 (O_1487,N_13654,N_14743);
and UO_1488 (O_1488,N_14688,N_14454);
nand UO_1489 (O_1489,N_14693,N_13719);
or UO_1490 (O_1490,N_14442,N_13714);
nor UO_1491 (O_1491,N_13704,N_13601);
and UO_1492 (O_1492,N_14983,N_14619);
or UO_1493 (O_1493,N_13720,N_13618);
or UO_1494 (O_1494,N_14408,N_13672);
xnor UO_1495 (O_1495,N_14777,N_13579);
or UO_1496 (O_1496,N_13829,N_14977);
or UO_1497 (O_1497,N_14735,N_14740);
and UO_1498 (O_1498,N_14431,N_14698);
nor UO_1499 (O_1499,N_14777,N_14890);
nand UO_1500 (O_1500,N_13885,N_14454);
or UO_1501 (O_1501,N_13733,N_14874);
xor UO_1502 (O_1502,N_14089,N_14829);
nand UO_1503 (O_1503,N_14090,N_14962);
nor UO_1504 (O_1504,N_13951,N_13870);
nor UO_1505 (O_1505,N_14850,N_14869);
and UO_1506 (O_1506,N_14565,N_14997);
xor UO_1507 (O_1507,N_14337,N_13973);
and UO_1508 (O_1508,N_14776,N_14643);
nand UO_1509 (O_1509,N_13525,N_14099);
nand UO_1510 (O_1510,N_13724,N_13765);
or UO_1511 (O_1511,N_14873,N_13911);
and UO_1512 (O_1512,N_14522,N_14926);
nor UO_1513 (O_1513,N_14336,N_13772);
nand UO_1514 (O_1514,N_14930,N_14019);
nor UO_1515 (O_1515,N_14395,N_14723);
nand UO_1516 (O_1516,N_13823,N_14864);
xor UO_1517 (O_1517,N_13678,N_14053);
and UO_1518 (O_1518,N_14217,N_14410);
and UO_1519 (O_1519,N_14909,N_14771);
and UO_1520 (O_1520,N_14371,N_14229);
or UO_1521 (O_1521,N_13893,N_13675);
xor UO_1522 (O_1522,N_13579,N_14334);
or UO_1523 (O_1523,N_14473,N_13823);
nor UO_1524 (O_1524,N_14309,N_13615);
nand UO_1525 (O_1525,N_14045,N_13966);
xnor UO_1526 (O_1526,N_13665,N_14654);
and UO_1527 (O_1527,N_14530,N_13901);
or UO_1528 (O_1528,N_14096,N_14586);
nor UO_1529 (O_1529,N_14640,N_13982);
or UO_1530 (O_1530,N_13564,N_13953);
and UO_1531 (O_1531,N_14088,N_14772);
or UO_1532 (O_1532,N_13949,N_13995);
and UO_1533 (O_1533,N_14434,N_13675);
nand UO_1534 (O_1534,N_13667,N_14959);
nand UO_1535 (O_1535,N_14243,N_14614);
or UO_1536 (O_1536,N_14513,N_14204);
xor UO_1537 (O_1537,N_14593,N_14363);
and UO_1538 (O_1538,N_13558,N_14836);
or UO_1539 (O_1539,N_13786,N_13535);
nor UO_1540 (O_1540,N_14146,N_14768);
nor UO_1541 (O_1541,N_14491,N_14226);
or UO_1542 (O_1542,N_14164,N_14631);
nor UO_1543 (O_1543,N_14640,N_14148);
or UO_1544 (O_1544,N_14395,N_14716);
and UO_1545 (O_1545,N_14364,N_13765);
nand UO_1546 (O_1546,N_14838,N_14776);
nor UO_1547 (O_1547,N_14281,N_14684);
or UO_1548 (O_1548,N_14330,N_14394);
and UO_1549 (O_1549,N_14135,N_13736);
xnor UO_1550 (O_1550,N_14820,N_14427);
nor UO_1551 (O_1551,N_14719,N_13881);
nor UO_1552 (O_1552,N_13668,N_14481);
nand UO_1553 (O_1553,N_14634,N_13861);
nand UO_1554 (O_1554,N_14049,N_14340);
and UO_1555 (O_1555,N_14945,N_13653);
nand UO_1556 (O_1556,N_14997,N_14801);
nand UO_1557 (O_1557,N_13565,N_14960);
xnor UO_1558 (O_1558,N_13859,N_13573);
nand UO_1559 (O_1559,N_14378,N_14249);
and UO_1560 (O_1560,N_13610,N_13637);
and UO_1561 (O_1561,N_14239,N_14522);
nand UO_1562 (O_1562,N_13611,N_14380);
or UO_1563 (O_1563,N_14708,N_14218);
nand UO_1564 (O_1564,N_13635,N_14252);
nor UO_1565 (O_1565,N_14502,N_13521);
or UO_1566 (O_1566,N_14269,N_14754);
xor UO_1567 (O_1567,N_14234,N_14761);
or UO_1568 (O_1568,N_14585,N_14280);
and UO_1569 (O_1569,N_14430,N_13559);
nor UO_1570 (O_1570,N_14113,N_14048);
nor UO_1571 (O_1571,N_13545,N_13582);
or UO_1572 (O_1572,N_14294,N_13740);
nand UO_1573 (O_1573,N_14712,N_14214);
nand UO_1574 (O_1574,N_13533,N_13808);
and UO_1575 (O_1575,N_14095,N_13781);
nand UO_1576 (O_1576,N_13596,N_14471);
nor UO_1577 (O_1577,N_13607,N_14015);
nor UO_1578 (O_1578,N_14577,N_14415);
or UO_1579 (O_1579,N_13764,N_13836);
or UO_1580 (O_1580,N_14511,N_13569);
nand UO_1581 (O_1581,N_13820,N_13770);
xor UO_1582 (O_1582,N_14040,N_14602);
and UO_1583 (O_1583,N_13654,N_14537);
and UO_1584 (O_1584,N_14390,N_14095);
or UO_1585 (O_1585,N_14368,N_14505);
nand UO_1586 (O_1586,N_14233,N_14402);
nand UO_1587 (O_1587,N_13509,N_14744);
or UO_1588 (O_1588,N_13699,N_14247);
nand UO_1589 (O_1589,N_14204,N_13620);
nor UO_1590 (O_1590,N_13856,N_14804);
or UO_1591 (O_1591,N_13844,N_14683);
nand UO_1592 (O_1592,N_13905,N_14208);
nor UO_1593 (O_1593,N_13846,N_14007);
nor UO_1594 (O_1594,N_14831,N_14379);
nand UO_1595 (O_1595,N_13740,N_13671);
and UO_1596 (O_1596,N_14316,N_14623);
xor UO_1597 (O_1597,N_14065,N_13736);
and UO_1598 (O_1598,N_14136,N_13749);
nand UO_1599 (O_1599,N_14794,N_14988);
nand UO_1600 (O_1600,N_14340,N_14809);
nor UO_1601 (O_1601,N_13533,N_14323);
or UO_1602 (O_1602,N_14882,N_13970);
nor UO_1603 (O_1603,N_13514,N_14155);
nor UO_1604 (O_1604,N_13924,N_14020);
and UO_1605 (O_1605,N_14839,N_14285);
xor UO_1606 (O_1606,N_14068,N_13568);
nor UO_1607 (O_1607,N_14962,N_14433);
or UO_1608 (O_1608,N_14300,N_14796);
or UO_1609 (O_1609,N_14482,N_13888);
nand UO_1610 (O_1610,N_13946,N_14392);
and UO_1611 (O_1611,N_14381,N_14944);
nor UO_1612 (O_1612,N_14975,N_13842);
xor UO_1613 (O_1613,N_14612,N_14169);
nand UO_1614 (O_1614,N_14040,N_13863);
nor UO_1615 (O_1615,N_14429,N_13699);
nor UO_1616 (O_1616,N_14817,N_13794);
and UO_1617 (O_1617,N_14682,N_13607);
nand UO_1618 (O_1618,N_14024,N_13817);
nor UO_1619 (O_1619,N_14679,N_13833);
nor UO_1620 (O_1620,N_14946,N_14097);
nor UO_1621 (O_1621,N_14146,N_14197);
nor UO_1622 (O_1622,N_13778,N_14327);
and UO_1623 (O_1623,N_14629,N_14484);
nand UO_1624 (O_1624,N_14142,N_14092);
and UO_1625 (O_1625,N_14152,N_14847);
and UO_1626 (O_1626,N_13878,N_14473);
or UO_1627 (O_1627,N_14273,N_14113);
nand UO_1628 (O_1628,N_13903,N_13968);
and UO_1629 (O_1629,N_13553,N_13746);
and UO_1630 (O_1630,N_14596,N_14454);
nor UO_1631 (O_1631,N_13869,N_13801);
and UO_1632 (O_1632,N_14699,N_14020);
and UO_1633 (O_1633,N_14128,N_14905);
nand UO_1634 (O_1634,N_14655,N_14469);
or UO_1635 (O_1635,N_14917,N_13521);
or UO_1636 (O_1636,N_13834,N_13564);
or UO_1637 (O_1637,N_14569,N_13635);
or UO_1638 (O_1638,N_14592,N_14161);
nor UO_1639 (O_1639,N_14132,N_14498);
nor UO_1640 (O_1640,N_14217,N_13915);
xor UO_1641 (O_1641,N_14491,N_13500);
nand UO_1642 (O_1642,N_14852,N_13501);
nand UO_1643 (O_1643,N_14156,N_14249);
xor UO_1644 (O_1644,N_13891,N_14995);
or UO_1645 (O_1645,N_13999,N_14747);
nor UO_1646 (O_1646,N_14529,N_14956);
and UO_1647 (O_1647,N_14913,N_14882);
nand UO_1648 (O_1648,N_14717,N_13792);
and UO_1649 (O_1649,N_13987,N_14287);
or UO_1650 (O_1650,N_14000,N_13613);
or UO_1651 (O_1651,N_13515,N_14323);
nor UO_1652 (O_1652,N_14939,N_14749);
nand UO_1653 (O_1653,N_14647,N_13845);
nand UO_1654 (O_1654,N_14716,N_13819);
xnor UO_1655 (O_1655,N_14448,N_14410);
nand UO_1656 (O_1656,N_13888,N_13675);
and UO_1657 (O_1657,N_13609,N_13893);
and UO_1658 (O_1658,N_14910,N_14712);
nor UO_1659 (O_1659,N_13568,N_13958);
or UO_1660 (O_1660,N_14524,N_13539);
nand UO_1661 (O_1661,N_13830,N_13637);
or UO_1662 (O_1662,N_14923,N_14681);
and UO_1663 (O_1663,N_14004,N_14722);
or UO_1664 (O_1664,N_13911,N_14421);
and UO_1665 (O_1665,N_14361,N_14820);
or UO_1666 (O_1666,N_14075,N_13809);
nand UO_1667 (O_1667,N_14178,N_14677);
or UO_1668 (O_1668,N_14917,N_14948);
xor UO_1669 (O_1669,N_13541,N_13993);
nor UO_1670 (O_1670,N_13934,N_14113);
nor UO_1671 (O_1671,N_13862,N_13898);
nor UO_1672 (O_1672,N_14110,N_14788);
nand UO_1673 (O_1673,N_13671,N_14199);
nand UO_1674 (O_1674,N_13755,N_14007);
or UO_1675 (O_1675,N_13765,N_13503);
nand UO_1676 (O_1676,N_14888,N_14532);
nand UO_1677 (O_1677,N_14367,N_13543);
nor UO_1678 (O_1678,N_14620,N_14066);
and UO_1679 (O_1679,N_14879,N_14883);
nand UO_1680 (O_1680,N_14622,N_13762);
nand UO_1681 (O_1681,N_13879,N_14496);
nor UO_1682 (O_1682,N_14555,N_14634);
and UO_1683 (O_1683,N_13970,N_14707);
xor UO_1684 (O_1684,N_14662,N_13985);
and UO_1685 (O_1685,N_14313,N_14597);
and UO_1686 (O_1686,N_14146,N_14491);
or UO_1687 (O_1687,N_14442,N_14865);
xnor UO_1688 (O_1688,N_13817,N_13823);
or UO_1689 (O_1689,N_14838,N_14238);
nor UO_1690 (O_1690,N_14517,N_13695);
or UO_1691 (O_1691,N_14338,N_13997);
nor UO_1692 (O_1692,N_14569,N_13963);
nand UO_1693 (O_1693,N_13608,N_14336);
nand UO_1694 (O_1694,N_13924,N_14511);
or UO_1695 (O_1695,N_14631,N_14893);
nor UO_1696 (O_1696,N_13731,N_14250);
and UO_1697 (O_1697,N_13977,N_14615);
nor UO_1698 (O_1698,N_14646,N_13968);
nand UO_1699 (O_1699,N_13996,N_14587);
nor UO_1700 (O_1700,N_14839,N_14985);
and UO_1701 (O_1701,N_14330,N_13509);
nand UO_1702 (O_1702,N_14335,N_14411);
xor UO_1703 (O_1703,N_13611,N_14135);
nor UO_1704 (O_1704,N_14341,N_14519);
and UO_1705 (O_1705,N_14984,N_14555);
nor UO_1706 (O_1706,N_14489,N_14460);
nor UO_1707 (O_1707,N_14847,N_14222);
and UO_1708 (O_1708,N_14898,N_13660);
nand UO_1709 (O_1709,N_14733,N_14055);
and UO_1710 (O_1710,N_14267,N_14674);
or UO_1711 (O_1711,N_14264,N_14631);
xnor UO_1712 (O_1712,N_14868,N_14644);
and UO_1713 (O_1713,N_14562,N_13627);
nand UO_1714 (O_1714,N_14380,N_14428);
nor UO_1715 (O_1715,N_14377,N_13709);
or UO_1716 (O_1716,N_13900,N_14709);
nand UO_1717 (O_1717,N_14707,N_13607);
and UO_1718 (O_1718,N_13669,N_13868);
nand UO_1719 (O_1719,N_13968,N_14237);
nand UO_1720 (O_1720,N_14825,N_14064);
nand UO_1721 (O_1721,N_14636,N_14677);
nor UO_1722 (O_1722,N_14966,N_14890);
nand UO_1723 (O_1723,N_13986,N_14578);
nor UO_1724 (O_1724,N_14950,N_13867);
nand UO_1725 (O_1725,N_13983,N_14443);
and UO_1726 (O_1726,N_14881,N_13910);
nand UO_1727 (O_1727,N_13888,N_14370);
or UO_1728 (O_1728,N_14607,N_14062);
and UO_1729 (O_1729,N_14497,N_14870);
nor UO_1730 (O_1730,N_13850,N_14775);
and UO_1731 (O_1731,N_14754,N_13715);
or UO_1732 (O_1732,N_14531,N_14826);
nand UO_1733 (O_1733,N_13880,N_14063);
nor UO_1734 (O_1734,N_14200,N_14092);
and UO_1735 (O_1735,N_14539,N_13894);
nor UO_1736 (O_1736,N_14975,N_14419);
nor UO_1737 (O_1737,N_14938,N_13651);
and UO_1738 (O_1738,N_13564,N_14951);
nand UO_1739 (O_1739,N_13742,N_14040);
xor UO_1740 (O_1740,N_14102,N_13777);
or UO_1741 (O_1741,N_14569,N_14510);
nor UO_1742 (O_1742,N_13792,N_14698);
nand UO_1743 (O_1743,N_14700,N_13802);
or UO_1744 (O_1744,N_14183,N_14343);
xor UO_1745 (O_1745,N_13791,N_14211);
nor UO_1746 (O_1746,N_13922,N_13662);
or UO_1747 (O_1747,N_14649,N_14999);
nor UO_1748 (O_1748,N_14462,N_14178);
nor UO_1749 (O_1749,N_14485,N_14513);
nor UO_1750 (O_1750,N_14648,N_14351);
nor UO_1751 (O_1751,N_14842,N_14008);
nor UO_1752 (O_1752,N_14478,N_13541);
nand UO_1753 (O_1753,N_14220,N_14383);
or UO_1754 (O_1754,N_14672,N_14286);
nor UO_1755 (O_1755,N_13964,N_14934);
or UO_1756 (O_1756,N_14562,N_13898);
nor UO_1757 (O_1757,N_14444,N_14155);
nor UO_1758 (O_1758,N_14098,N_14732);
nand UO_1759 (O_1759,N_14467,N_14399);
nor UO_1760 (O_1760,N_13782,N_13666);
and UO_1761 (O_1761,N_14012,N_13693);
nand UO_1762 (O_1762,N_14128,N_13756);
nor UO_1763 (O_1763,N_13825,N_13855);
nand UO_1764 (O_1764,N_13904,N_14525);
and UO_1765 (O_1765,N_14526,N_14229);
nor UO_1766 (O_1766,N_14292,N_13985);
or UO_1767 (O_1767,N_13765,N_14493);
nor UO_1768 (O_1768,N_14716,N_14145);
or UO_1769 (O_1769,N_14687,N_14992);
or UO_1770 (O_1770,N_14216,N_13897);
nand UO_1771 (O_1771,N_14256,N_14628);
or UO_1772 (O_1772,N_14983,N_14544);
nor UO_1773 (O_1773,N_13829,N_13939);
nand UO_1774 (O_1774,N_14020,N_13598);
or UO_1775 (O_1775,N_13701,N_14570);
and UO_1776 (O_1776,N_13885,N_14477);
and UO_1777 (O_1777,N_13654,N_13710);
xor UO_1778 (O_1778,N_14693,N_14979);
nand UO_1779 (O_1779,N_14601,N_14833);
or UO_1780 (O_1780,N_14081,N_14073);
or UO_1781 (O_1781,N_14877,N_14204);
nor UO_1782 (O_1782,N_14500,N_13914);
xnor UO_1783 (O_1783,N_14443,N_14979);
nor UO_1784 (O_1784,N_13778,N_14804);
or UO_1785 (O_1785,N_14415,N_14422);
nand UO_1786 (O_1786,N_13573,N_14359);
or UO_1787 (O_1787,N_14276,N_14616);
and UO_1788 (O_1788,N_14004,N_13912);
and UO_1789 (O_1789,N_13657,N_13735);
nor UO_1790 (O_1790,N_14904,N_13997);
xor UO_1791 (O_1791,N_13619,N_14524);
nand UO_1792 (O_1792,N_13909,N_14809);
and UO_1793 (O_1793,N_13966,N_13761);
nand UO_1794 (O_1794,N_14668,N_13660);
nor UO_1795 (O_1795,N_13893,N_13928);
nand UO_1796 (O_1796,N_13563,N_14754);
or UO_1797 (O_1797,N_14345,N_13628);
nor UO_1798 (O_1798,N_14139,N_14834);
nand UO_1799 (O_1799,N_13662,N_13884);
and UO_1800 (O_1800,N_14018,N_13910);
nand UO_1801 (O_1801,N_14799,N_13801);
or UO_1802 (O_1802,N_14289,N_14412);
or UO_1803 (O_1803,N_13905,N_14261);
xnor UO_1804 (O_1804,N_13942,N_14817);
nand UO_1805 (O_1805,N_14209,N_14494);
xor UO_1806 (O_1806,N_14613,N_13548);
or UO_1807 (O_1807,N_14068,N_14471);
or UO_1808 (O_1808,N_14146,N_14821);
nand UO_1809 (O_1809,N_14399,N_14637);
and UO_1810 (O_1810,N_13991,N_14078);
nand UO_1811 (O_1811,N_14485,N_13685);
or UO_1812 (O_1812,N_13777,N_14457);
and UO_1813 (O_1813,N_13609,N_14436);
or UO_1814 (O_1814,N_14484,N_14320);
or UO_1815 (O_1815,N_14099,N_14321);
nand UO_1816 (O_1816,N_14992,N_14237);
or UO_1817 (O_1817,N_14983,N_14382);
xor UO_1818 (O_1818,N_14909,N_13529);
nor UO_1819 (O_1819,N_14250,N_13646);
and UO_1820 (O_1820,N_14708,N_14701);
nor UO_1821 (O_1821,N_14317,N_14259);
nor UO_1822 (O_1822,N_14463,N_14469);
nor UO_1823 (O_1823,N_14531,N_14180);
or UO_1824 (O_1824,N_14374,N_14239);
nand UO_1825 (O_1825,N_14679,N_13815);
and UO_1826 (O_1826,N_14986,N_13794);
nor UO_1827 (O_1827,N_14280,N_14784);
and UO_1828 (O_1828,N_13637,N_13982);
or UO_1829 (O_1829,N_14133,N_14952);
and UO_1830 (O_1830,N_14538,N_14903);
and UO_1831 (O_1831,N_14573,N_13981);
nor UO_1832 (O_1832,N_14261,N_14305);
and UO_1833 (O_1833,N_14912,N_13951);
nor UO_1834 (O_1834,N_13654,N_14491);
nor UO_1835 (O_1835,N_14112,N_14564);
and UO_1836 (O_1836,N_13725,N_14091);
nand UO_1837 (O_1837,N_14503,N_14775);
or UO_1838 (O_1838,N_14377,N_13539);
and UO_1839 (O_1839,N_14554,N_14669);
or UO_1840 (O_1840,N_13961,N_13962);
nand UO_1841 (O_1841,N_14068,N_14221);
nor UO_1842 (O_1842,N_14536,N_14172);
and UO_1843 (O_1843,N_14108,N_14192);
nor UO_1844 (O_1844,N_13881,N_14678);
nand UO_1845 (O_1845,N_14364,N_14463);
and UO_1846 (O_1846,N_14898,N_14400);
xnor UO_1847 (O_1847,N_13665,N_14140);
nand UO_1848 (O_1848,N_14734,N_13773);
nand UO_1849 (O_1849,N_13794,N_13563);
xor UO_1850 (O_1850,N_13886,N_14835);
or UO_1851 (O_1851,N_14943,N_14313);
nand UO_1852 (O_1852,N_14557,N_14595);
nor UO_1853 (O_1853,N_14936,N_13806);
and UO_1854 (O_1854,N_13679,N_14236);
nand UO_1855 (O_1855,N_14657,N_14036);
or UO_1856 (O_1856,N_14358,N_14767);
nand UO_1857 (O_1857,N_14079,N_13838);
and UO_1858 (O_1858,N_14220,N_14006);
and UO_1859 (O_1859,N_14745,N_14103);
nor UO_1860 (O_1860,N_13676,N_14145);
and UO_1861 (O_1861,N_13523,N_14099);
nor UO_1862 (O_1862,N_13675,N_14641);
xnor UO_1863 (O_1863,N_14637,N_13827);
and UO_1864 (O_1864,N_14066,N_13942);
or UO_1865 (O_1865,N_14651,N_14882);
xnor UO_1866 (O_1866,N_13665,N_13976);
nand UO_1867 (O_1867,N_14064,N_14475);
nor UO_1868 (O_1868,N_14345,N_13742);
xor UO_1869 (O_1869,N_13669,N_14798);
xnor UO_1870 (O_1870,N_14898,N_13928);
and UO_1871 (O_1871,N_14191,N_14537);
and UO_1872 (O_1872,N_14891,N_14530);
nor UO_1873 (O_1873,N_14665,N_13533);
or UO_1874 (O_1874,N_13859,N_13835);
xor UO_1875 (O_1875,N_14004,N_13531);
and UO_1876 (O_1876,N_14388,N_13505);
nand UO_1877 (O_1877,N_14779,N_14767);
nor UO_1878 (O_1878,N_13967,N_13786);
xnor UO_1879 (O_1879,N_13626,N_14493);
nor UO_1880 (O_1880,N_14649,N_13570);
nor UO_1881 (O_1881,N_13588,N_13536);
nor UO_1882 (O_1882,N_14457,N_13605);
and UO_1883 (O_1883,N_14285,N_14250);
nor UO_1884 (O_1884,N_14003,N_13635);
nor UO_1885 (O_1885,N_13774,N_14141);
and UO_1886 (O_1886,N_14213,N_13667);
and UO_1887 (O_1887,N_13586,N_14745);
and UO_1888 (O_1888,N_13527,N_14850);
nand UO_1889 (O_1889,N_14545,N_14280);
xnor UO_1890 (O_1890,N_13823,N_14649);
and UO_1891 (O_1891,N_14531,N_14070);
or UO_1892 (O_1892,N_13580,N_13786);
xnor UO_1893 (O_1893,N_14484,N_14341);
and UO_1894 (O_1894,N_14925,N_14253);
and UO_1895 (O_1895,N_13805,N_14632);
and UO_1896 (O_1896,N_14865,N_13793);
nand UO_1897 (O_1897,N_14577,N_14204);
and UO_1898 (O_1898,N_14937,N_14108);
nand UO_1899 (O_1899,N_14501,N_14866);
nor UO_1900 (O_1900,N_14407,N_13920);
or UO_1901 (O_1901,N_14999,N_14006);
nand UO_1902 (O_1902,N_14280,N_14094);
nand UO_1903 (O_1903,N_13863,N_14277);
and UO_1904 (O_1904,N_14490,N_13996);
or UO_1905 (O_1905,N_14468,N_14581);
nor UO_1906 (O_1906,N_14276,N_13834);
nor UO_1907 (O_1907,N_14712,N_14555);
and UO_1908 (O_1908,N_14582,N_14854);
nand UO_1909 (O_1909,N_14913,N_14189);
nor UO_1910 (O_1910,N_13726,N_14439);
and UO_1911 (O_1911,N_14361,N_14314);
and UO_1912 (O_1912,N_14651,N_13935);
nand UO_1913 (O_1913,N_14460,N_14470);
nand UO_1914 (O_1914,N_14886,N_14151);
xor UO_1915 (O_1915,N_14313,N_13753);
nor UO_1916 (O_1916,N_14769,N_14792);
nand UO_1917 (O_1917,N_14678,N_13561);
nand UO_1918 (O_1918,N_14866,N_14068);
nor UO_1919 (O_1919,N_14852,N_13865);
nor UO_1920 (O_1920,N_14877,N_13777);
and UO_1921 (O_1921,N_14657,N_13983);
or UO_1922 (O_1922,N_13991,N_13909);
nor UO_1923 (O_1923,N_13963,N_13651);
nand UO_1924 (O_1924,N_13655,N_14428);
nand UO_1925 (O_1925,N_14480,N_14769);
or UO_1926 (O_1926,N_14095,N_14574);
or UO_1927 (O_1927,N_13875,N_14919);
xnor UO_1928 (O_1928,N_13945,N_14003);
nor UO_1929 (O_1929,N_14588,N_14554);
xor UO_1930 (O_1930,N_14454,N_14341);
or UO_1931 (O_1931,N_14711,N_14197);
nor UO_1932 (O_1932,N_13715,N_13837);
xnor UO_1933 (O_1933,N_14597,N_14492);
nand UO_1934 (O_1934,N_14133,N_13605);
or UO_1935 (O_1935,N_13793,N_14433);
nand UO_1936 (O_1936,N_14083,N_14177);
or UO_1937 (O_1937,N_14067,N_14805);
or UO_1938 (O_1938,N_14042,N_14966);
nor UO_1939 (O_1939,N_14266,N_14539);
or UO_1940 (O_1940,N_14070,N_14609);
nand UO_1941 (O_1941,N_14709,N_14044);
and UO_1942 (O_1942,N_13980,N_14139);
xor UO_1943 (O_1943,N_14882,N_14415);
or UO_1944 (O_1944,N_14859,N_14028);
nand UO_1945 (O_1945,N_14190,N_13584);
and UO_1946 (O_1946,N_14047,N_14126);
or UO_1947 (O_1947,N_13659,N_13744);
xnor UO_1948 (O_1948,N_14893,N_13905);
and UO_1949 (O_1949,N_14695,N_14991);
nand UO_1950 (O_1950,N_14232,N_13808);
or UO_1951 (O_1951,N_14960,N_14082);
nor UO_1952 (O_1952,N_14015,N_14164);
or UO_1953 (O_1953,N_13803,N_14321);
nand UO_1954 (O_1954,N_14810,N_14953);
nand UO_1955 (O_1955,N_13603,N_13548);
nand UO_1956 (O_1956,N_14127,N_14656);
and UO_1957 (O_1957,N_14315,N_13989);
xor UO_1958 (O_1958,N_14888,N_14925);
nor UO_1959 (O_1959,N_13876,N_14120);
and UO_1960 (O_1960,N_14832,N_13850);
nand UO_1961 (O_1961,N_14796,N_14188);
nor UO_1962 (O_1962,N_13628,N_13632);
and UO_1963 (O_1963,N_14015,N_14718);
or UO_1964 (O_1964,N_14754,N_13893);
and UO_1965 (O_1965,N_14433,N_13884);
nand UO_1966 (O_1966,N_14689,N_14920);
nand UO_1967 (O_1967,N_14172,N_13549);
and UO_1968 (O_1968,N_14687,N_13686);
nand UO_1969 (O_1969,N_14416,N_13753);
nor UO_1970 (O_1970,N_14775,N_14595);
nor UO_1971 (O_1971,N_14570,N_14539);
nand UO_1972 (O_1972,N_14323,N_13611);
nand UO_1973 (O_1973,N_14795,N_14385);
and UO_1974 (O_1974,N_14387,N_14655);
nand UO_1975 (O_1975,N_13836,N_14538);
and UO_1976 (O_1976,N_14517,N_13861);
nor UO_1977 (O_1977,N_13854,N_14741);
xnor UO_1978 (O_1978,N_14461,N_13680);
nor UO_1979 (O_1979,N_14987,N_14886);
nor UO_1980 (O_1980,N_14737,N_13607);
nand UO_1981 (O_1981,N_13987,N_14746);
or UO_1982 (O_1982,N_14183,N_13881);
nor UO_1983 (O_1983,N_13863,N_14133);
nand UO_1984 (O_1984,N_14453,N_14540);
nand UO_1985 (O_1985,N_13641,N_14388);
nor UO_1986 (O_1986,N_14538,N_13674);
or UO_1987 (O_1987,N_14826,N_14782);
nor UO_1988 (O_1988,N_14108,N_14896);
nand UO_1989 (O_1989,N_14456,N_14449);
or UO_1990 (O_1990,N_14029,N_14013);
nor UO_1991 (O_1991,N_14005,N_14406);
or UO_1992 (O_1992,N_14889,N_13914);
or UO_1993 (O_1993,N_14417,N_14807);
and UO_1994 (O_1994,N_14521,N_14614);
xor UO_1995 (O_1995,N_14915,N_14242);
and UO_1996 (O_1996,N_14816,N_14824);
nor UO_1997 (O_1997,N_13585,N_14192);
or UO_1998 (O_1998,N_14400,N_14497);
nor UO_1999 (O_1999,N_14724,N_13769);
endmodule